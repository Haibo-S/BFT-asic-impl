module pi_switch (ce,
    clk,
    done,
    l_i_bp,
    l_i_v,
    l_o_bp,
    l_o_v,
    r_i_bp,
    r_i_v,
    r_o_bp,
    r_o_v,
    rst,
    u0_i_bp,
    u0_i_v,
    u0_o_bp,
    u0_o_v,
    u1_i_bp,
    u1_i_v,
    u1_o_bp,
    u1_o_v,
    l_i,
    l_o,
    r_i,
    r_o,
    u0_i,
    u0_o,
    u1_i,
    u1_o);
 input ce;
 input clk;
 output done;
 output l_i_bp;
 input l_i_v;
 input l_o_bp;
 output l_o_v;
 output r_i_bp;
 input r_i_v;
 input r_o_bp;
 output r_o_v;
 input rst;
 output u0_i_bp;
 input u0_i_v;
 input u0_o_bp;
 output u0_o_v;
 output u1_i_bp;
 input u1_i_v;
 input u1_o_bp;
 output u1_o_v;
 input [35:0] l_i;
 output [35:0] l_o;
 input [35:0] r_i;
 output [35:0] r_o;
 input [35:0] u0_i;
 output [35:0] u0_o;
 input [35:0] u1_i;
 output [35:0] u1_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire clknet_0_clk;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net303;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 OA21x2_ASAP7_75t_R _0767_ (.A1(net65),
    .A2(net64),
    .B(net150),
    .Y(_0564_));
 INVx2_ASAP7_75t_R _0768_ (.A(_0115_),
    .Y(_0565_));
 AND2x4_ASAP7_75t_R _0769_ (.A(_0153_),
    .B(_0155_),
    .Y(_0566_));
 INVx2_ASAP7_75t_R _0770_ (.A(net138),
    .Y(_0567_));
 OA211x2_ASAP7_75t_R _0771_ (.A1(_0565_),
    .A2(_0566_),
    .B(net149),
    .C(_0567_),
    .Y(_0568_));
 BUFx6f_ASAP7_75t_R _0772_ (.A(u0_i_v),
    .Y(_0569_));
 INVx2_ASAP7_75t_R _0773_ (.A(net101),
    .Y(_0570_));
 AND2x4_ASAP7_75t_R _0774_ (.A(_0115_),
    .B(_0155_),
    .Y(_0571_));
 BUFx6f_ASAP7_75t_R _0775_ (.A(l_o_bp),
    .Y(_0572_));
 AO31x2_ASAP7_75t_R _0776_ (.A1(_0569_),
    .A2(_0570_),
    .A3(_0571_),
    .B(_0572_),
    .Y(_0573_));
 INVx1_ASAP7_75t_R _0777_ (.A(net63),
    .Y(_0574_));
 NOR2x1_ASAP7_75t_R _0778_ (.A(net65),
    .B(net64),
    .Y(_0575_));
 OA211x2_ASAP7_75t_R _0779_ (.A1(_0568_),
    .A2(_0573_),
    .B(_0574_),
    .C(_0575_),
    .Y(_0576_));
 OAI21x1_ASAP7_75t_R _0780_ (.A1(_0564_),
    .A2(_0576_),
    .B(net74),
    .Y(_0577_));
 INVx1_ASAP7_75t_R _0781_ (.A(_0577_),
    .Y(net189));
 INVx2_ASAP7_75t_R _0782_ (.A(_0154_),
    .Y(_0578_));
 AND2x6_ASAP7_75t_R _0783_ (.A(_0569_),
    .B(net101),
    .Y(_0579_));
 OA21x2_ASAP7_75t_R _0784_ (.A1(_0578_),
    .A2(_0566_),
    .B(_0579_),
    .Y(_0580_));
 AND2x2_ASAP7_75t_R _0785_ (.A(_0153_),
    .B(_0154_),
    .Y(_0581_));
 AND2x4_ASAP7_75t_R _0786_ (.A(net149),
    .B(net138),
    .Y(_0582_));
 AO21x1_ASAP7_75t_R _0787_ (.A1(_0581_),
    .A2(_0582_),
    .B(net75),
    .Y(_0583_));
 OR2x6_ASAP7_75t_R _0788_ (.A(_0580_),
    .B(_0583_),
    .Y(_0584_));
 NOR2x2_ASAP7_75t_R _0789_ (.A(net28),
    .B(net27),
    .Y(_0585_));
 AND2x6_ASAP7_75t_R _0790_ (.A(net37),
    .B(net26),
    .Y(_0586_));
 AND2x2_ASAP7_75t_R _0791_ (.A(_0585_),
    .B(_0586_),
    .Y(_0587_));
 OR2x2_ASAP7_75t_R _0792_ (.A(net28),
    .B(net27),
    .Y(_0588_));
 AND3x1_ASAP7_75t_R _0793_ (.A(net37),
    .B(net112),
    .C(_0588_),
    .Y(_0589_));
 AOI21x1_ASAP7_75t_R _0794_ (.A1(_0584_),
    .A2(_0587_),
    .B(_0589_),
    .Y(_0590_));
 INVx2_ASAP7_75t_R _0795_ (.A(_0590_),
    .Y(net151));
 INVx1_ASAP7_75t_R _0796_ (.A(net74),
    .Y(_0591_));
 OR5x1_ASAP7_75t_R _0797_ (.A(_0591_),
    .B(net63),
    .C(net65),
    .D(net64),
    .E(_0155_),
    .Y(_0592_));
 BUFx6f_ASAP7_75t_R _0798_ (.A(_0592_),
    .Y(_0593_));
 INVx2_ASAP7_75t_R _0799_ (.A(net75),
    .Y(_0594_));
 NAND2x2_ASAP7_75t_R _0800_ (.A(_0115_),
    .B(_0155_),
    .Y(_0595_));
 AND2x2_ASAP7_75t_R _0801_ (.A(_0594_),
    .B(_0595_),
    .Y(_0596_));
 NAND2x2_ASAP7_75t_R _0802_ (.A(_0569_),
    .B(net101),
    .Y(_0597_));
 AND2x2_ASAP7_75t_R _0803_ (.A(_0594_),
    .B(_0597_),
    .Y(_0598_));
 NAND2x2_ASAP7_75t_R _0804_ (.A(_0585_),
    .B(_0586_),
    .Y(_0599_));
 NAND2x1_ASAP7_75t_R _0805_ (.A(net149),
    .B(net138),
    .Y(_0600_));
 AO221x1_ASAP7_75t_R _0806_ (.A1(_0593_),
    .A2(_0596_),
    .B1(_0598_),
    .B2(_0599_),
    .C(_0600_),
    .Y(_0601_));
 NOR2x1_ASAP7_75t_R _0807_ (.A(_0572_),
    .B(_0571_),
    .Y(_0602_));
 AOI21x1_ASAP7_75t_R _0808_ (.A1(_0569_),
    .A2(_0570_),
    .B(_0572_),
    .Y(_0603_));
 OR4x1_ASAP7_75t_R _0809_ (.A(_0591_),
    .B(net63),
    .C(net65),
    .D(net64),
    .Y(_0604_));
 NAND2x1_ASAP7_75t_R _0810_ (.A(net149),
    .B(_0567_),
    .Y(_0605_));
 AO221x1_ASAP7_75t_R _0811_ (.A1(_0593_),
    .A2(_0602_),
    .B1(_0603_),
    .B2(_0604_),
    .C(_0605_),
    .Y(_0606_));
 AND2x4_ASAP7_75t_R _0812_ (.A(_0601_),
    .B(_0606_),
    .Y(_0607_));
 INVx1_ASAP7_75t_R _0813_ (.A(_0607_),
    .Y(net265));
 AND2x2_ASAP7_75t_R _0814_ (.A(_0569_),
    .B(_0570_),
    .Y(_0608_));
 INVx2_ASAP7_75t_R _0815_ (.A(_0153_),
    .Y(_0609_));
 AO31x2_ASAP7_75t_R _0816_ (.A1(_0609_),
    .A2(_0585_),
    .A3(_0586_),
    .B(_0581_),
    .Y(_0610_));
 AO32x1_ASAP7_75t_R _0817_ (.A1(net74),
    .A2(_0574_),
    .A3(_0575_),
    .B1(_0567_),
    .B2(net149),
    .Y(_0611_));
 AO21x1_ASAP7_75t_R _0818_ (.A1(_0610_),
    .A2(_0611_),
    .B(_0572_),
    .Y(_0612_));
 AO21x1_ASAP7_75t_R _0819_ (.A1(_0585_),
    .A2(_0586_),
    .B(_0582_),
    .Y(_0613_));
 AO21x1_ASAP7_75t_R _0820_ (.A1(_0610_),
    .A2(_0613_),
    .B(net75),
    .Y(_0614_));
 AOI22x1_ASAP7_75t_R _0821_ (.A1(_0608_),
    .A2(_0612_),
    .B1(_0614_),
    .B2(_0579_),
    .Y(_0615_));
 INVx1_ASAP7_75t_R _0822_ (.A(_0615_),
    .Y(net227));
 INVx2_ASAP7_75t_R _0823_ (.A(_0155_),
    .Y(_0616_));
 AND4x1_ASAP7_75t_R _0824_ (.A(_0616_),
    .B(_0590_),
    .C(_0607_),
    .D(_0615_),
    .Y(_0617_));
 AO31x2_ASAP7_75t_R _0825_ (.A1(_0578_),
    .A2(_0601_),
    .A3(_0606_),
    .B(_0565_),
    .Y(_0618_));
 AND3x1_ASAP7_75t_R _0826_ (.A(net189),
    .B(_0590_),
    .C(_0618_),
    .Y(_0619_));
 AND2x2_ASAP7_75t_R _0827_ (.A(_0609_),
    .B(net189),
    .Y(_0620_));
 BUFx6f_ASAP7_75t_R _0828_ (.A(rst),
    .Y(_0621_));
 INVx5_ASAP7_75t_R _0829_ (.A(_0621_),
    .Y(_0622_));
 BUFx12f_ASAP7_75t_R _0830_ (.A(_0622_),
    .Y(_0623_));
 BUFx6f_ASAP7_75t_R _0831_ (.A(_0623_),
    .Y(_0624_));
 OA31x2_ASAP7_75t_R _0832_ (.A1(_0617_),
    .A2(_0619_),
    .A3(_0620_),
    .B1(_0624_),
    .Y(_0002_));
 OAI21x1_ASAP7_75t_R _0833_ (.A1(_0115_),
    .A2(net151),
    .B(_0566_),
    .Y(_0625_));
 BUFx6f_ASAP7_75t_R _0834_ (.A(_0622_),
    .Y(_0626_));
 OA211x2_ASAP7_75t_R _0835_ (.A1(_0616_),
    .A2(_0577_),
    .B(net227),
    .C(_0626_),
    .Y(_0627_));
 AND5x1_ASAP7_75t_R _0836_ (.A(_0626_),
    .B(_0578_),
    .C(_0577_),
    .D(_0590_),
    .E(_0607_),
    .Y(_0628_));
 AO21x1_ASAP7_75t_R _0837_ (.A1(_0625_),
    .A2(_0627_),
    .B(_0628_),
    .Y(_0001_));
 AO31x2_ASAP7_75t_R _0838_ (.A1(_0616_),
    .A2(_0607_),
    .A3(_0615_),
    .B(_0618_),
    .Y(_0629_));
 AND4x1_ASAP7_75t_R _0839_ (.A(_0609_),
    .B(_0577_),
    .C(_0607_),
    .D(_0615_),
    .Y(_0630_));
 BUFx12f_ASAP7_75t_R _0840_ (.A(_0621_),
    .Y(_0631_));
 AO211x2_ASAP7_75t_R _0841_ (.A1(net151),
    .A2(_0629_),
    .B(_0630_),
    .C(_0631_),
    .Y(_0000_));
 AND2x2_ASAP7_75t_R _0842_ (.A(_0626_),
    .B(net265),
    .Y(_0632_));
 AO21x1_ASAP7_75t_R _0843_ (.A1(_0609_),
    .A2(_0577_),
    .B(_0616_),
    .Y(_0633_));
 AND3x1_ASAP7_75t_R _0844_ (.A(_0626_),
    .B(net265),
    .C(_0615_),
    .Y(_0634_));
 AND5x1_ASAP7_75t_R _0845_ (.A(_0623_),
    .B(_0565_),
    .C(_0577_),
    .D(_0590_),
    .E(_0615_),
    .Y(_0635_));
 AO221x1_ASAP7_75t_R _0846_ (.A1(_0578_),
    .A2(_0632_),
    .B1(_0633_),
    .B2(_0634_),
    .C(_0635_),
    .Y(_0003_));
 INVx1_ASAP7_75t_R _0847_ (.A(_0004_),
    .Y(net302));
 INVx1_ASAP7_75t_R _0848_ (.A(_0005_),
    .Y(net301));
 INVx1_ASAP7_75t_R _0849_ (.A(_0006_),
    .Y(net300));
 INVx1_ASAP7_75t_R _0850_ (.A(_0007_),
    .Y(net299));
 INVx1_ASAP7_75t_R _0851_ (.A(_0008_),
    .Y(net298));
 INVx1_ASAP7_75t_R _0852_ (.A(_0009_),
    .Y(net297));
 INVx1_ASAP7_75t_R _0853_ (.A(_0010_),
    .Y(net296));
 INVx1_ASAP7_75t_R _0854_ (.A(_0011_),
    .Y(net295));
 INVx1_ASAP7_75t_R _0855_ (.A(_0012_),
    .Y(net294));
 INVx1_ASAP7_75t_R _0856_ (.A(_0013_),
    .Y(net293));
 INVx1_ASAP7_75t_R _0857_ (.A(_0014_),
    .Y(net292));
 INVx1_ASAP7_75t_R _0858_ (.A(_0015_),
    .Y(net291));
 INVx1_ASAP7_75t_R _0859_ (.A(_0016_),
    .Y(net290));
 INVx1_ASAP7_75t_R _0860_ (.A(_0017_),
    .Y(net289));
 INVx1_ASAP7_75t_R _0861_ (.A(_0018_),
    .Y(net288));
 INVx1_ASAP7_75t_R _0862_ (.A(_0019_),
    .Y(net287));
 INVx1_ASAP7_75t_R _0863_ (.A(_0020_),
    .Y(net286));
 INVx1_ASAP7_75t_R _0864_ (.A(_0021_),
    .Y(net285));
 INVx1_ASAP7_75t_R _0865_ (.A(_0022_),
    .Y(net284));
 INVx1_ASAP7_75t_R _0866_ (.A(_0023_),
    .Y(net283));
 INVx1_ASAP7_75t_R _0867_ (.A(_0024_),
    .Y(net282));
 INVx1_ASAP7_75t_R _0868_ (.A(_0025_),
    .Y(net281));
 INVx1_ASAP7_75t_R _0869_ (.A(_0026_),
    .Y(net280));
 INVx1_ASAP7_75t_R _0870_ (.A(_0027_),
    .Y(net279));
 INVx1_ASAP7_75t_R _0871_ (.A(_0028_),
    .Y(net278));
 INVx1_ASAP7_75t_R _0872_ (.A(_0029_),
    .Y(net277));
 INVx1_ASAP7_75t_R _0873_ (.A(_0030_),
    .Y(net276));
 INVx1_ASAP7_75t_R _0874_ (.A(_0031_),
    .Y(net275));
 INVx1_ASAP7_75t_R _0875_ (.A(_0032_),
    .Y(net274));
 INVx1_ASAP7_75t_R _0876_ (.A(_0033_),
    .Y(net273));
 INVx1_ASAP7_75t_R _0877_ (.A(_0034_),
    .Y(net272));
 INVx1_ASAP7_75t_R _0878_ (.A(_0035_),
    .Y(net271));
 INVx1_ASAP7_75t_R _0879_ (.A(_0036_),
    .Y(net270));
 INVx1_ASAP7_75t_R _0880_ (.A(_0037_),
    .Y(net269));
 INVx1_ASAP7_75t_R _0881_ (.A(_0038_),
    .Y(net268));
 INVx1_ASAP7_75t_R _0882_ (.A(_0039_),
    .Y(net267));
 INVx1_ASAP7_75t_R _0883_ (.A(_0040_),
    .Y(net266));
 INVx1_ASAP7_75t_R _0884_ (.A(_0041_),
    .Y(net264));
 INVx1_ASAP7_75t_R _0885_ (.A(_0042_),
    .Y(net263));
 INVx1_ASAP7_75t_R _0886_ (.A(_0043_),
    .Y(net262));
 INVx1_ASAP7_75t_R _0887_ (.A(_0044_),
    .Y(net261));
 INVx1_ASAP7_75t_R _0888_ (.A(_0045_),
    .Y(net260));
 INVx1_ASAP7_75t_R _0889_ (.A(_0046_),
    .Y(net259));
 INVx1_ASAP7_75t_R _0890_ (.A(_0047_),
    .Y(net258));
 INVx1_ASAP7_75t_R _0891_ (.A(_0048_),
    .Y(net257));
 INVx1_ASAP7_75t_R _0892_ (.A(_0049_),
    .Y(net256));
 INVx1_ASAP7_75t_R _0893_ (.A(_0050_),
    .Y(net255));
 INVx1_ASAP7_75t_R _0894_ (.A(_0051_),
    .Y(net254));
 INVx1_ASAP7_75t_R _0895_ (.A(_0052_),
    .Y(net253));
 INVx1_ASAP7_75t_R _0896_ (.A(_0053_),
    .Y(net252));
 INVx1_ASAP7_75t_R _0897_ (.A(_0054_),
    .Y(net251));
 INVx1_ASAP7_75t_R _0898_ (.A(_0055_),
    .Y(net250));
 INVx1_ASAP7_75t_R _0899_ (.A(_0056_),
    .Y(net249));
 INVx1_ASAP7_75t_R _0900_ (.A(_0057_),
    .Y(net248));
 INVx1_ASAP7_75t_R _0901_ (.A(_0058_),
    .Y(net247));
 INVx1_ASAP7_75t_R _0902_ (.A(_0059_),
    .Y(net246));
 INVx1_ASAP7_75t_R _0903_ (.A(_0060_),
    .Y(net245));
 INVx1_ASAP7_75t_R _0904_ (.A(_0061_),
    .Y(net244));
 INVx1_ASAP7_75t_R _0905_ (.A(_0062_),
    .Y(net243));
 INVx1_ASAP7_75t_R _0906_ (.A(_0063_),
    .Y(net242));
 INVx1_ASAP7_75t_R _0907_ (.A(_0064_),
    .Y(net241));
 INVx1_ASAP7_75t_R _0908_ (.A(_0065_),
    .Y(net240));
 INVx1_ASAP7_75t_R _0909_ (.A(_0066_),
    .Y(net239));
 INVx1_ASAP7_75t_R _0910_ (.A(_0067_),
    .Y(net238));
 INVx1_ASAP7_75t_R _0911_ (.A(_0068_),
    .Y(net237));
 INVx1_ASAP7_75t_R _0912_ (.A(_0069_),
    .Y(net236));
 INVx1_ASAP7_75t_R _0913_ (.A(_0070_),
    .Y(net235));
 INVx1_ASAP7_75t_R _0914_ (.A(_0071_),
    .Y(net234));
 INVx1_ASAP7_75t_R _0915_ (.A(_0072_),
    .Y(net233));
 INVx1_ASAP7_75t_R _0916_ (.A(_0073_),
    .Y(net232));
 INVx1_ASAP7_75t_R _0917_ (.A(_0074_),
    .Y(net231));
 INVx1_ASAP7_75t_R _0918_ (.A(_0075_),
    .Y(net230));
 INVx1_ASAP7_75t_R _0919_ (.A(_0076_),
    .Y(net229));
 INVx1_ASAP7_75t_R _0920_ (.A(_0077_),
    .Y(net228));
 INVx1_ASAP7_75t_R _0921_ (.A(_0078_),
    .Y(net226));
 INVx1_ASAP7_75t_R _0922_ (.A(_0079_),
    .Y(net225));
 INVx1_ASAP7_75t_R _0923_ (.A(_0080_),
    .Y(net224));
 INVx1_ASAP7_75t_R _0924_ (.A(_0081_),
    .Y(net223));
 INVx1_ASAP7_75t_R _0925_ (.A(_0082_),
    .Y(net222));
 INVx1_ASAP7_75t_R _0926_ (.A(_0083_),
    .Y(net221));
 INVx1_ASAP7_75t_R _0927_ (.A(_0084_),
    .Y(net220));
 INVx1_ASAP7_75t_R _0928_ (.A(_0085_),
    .Y(net219));
 INVx1_ASAP7_75t_R _0929_ (.A(_0086_),
    .Y(net218));
 INVx1_ASAP7_75t_R _0930_ (.A(_0087_),
    .Y(net217));
 INVx1_ASAP7_75t_R _0931_ (.A(_0088_),
    .Y(net216));
 INVx1_ASAP7_75t_R _0932_ (.A(_0089_),
    .Y(net215));
 INVx1_ASAP7_75t_R _0933_ (.A(_0090_),
    .Y(net214));
 INVx1_ASAP7_75t_R _0934_ (.A(_0091_),
    .Y(net213));
 INVx1_ASAP7_75t_R _0935_ (.A(_0092_),
    .Y(net212));
 INVx1_ASAP7_75t_R _0936_ (.A(_0093_),
    .Y(net211));
 INVx1_ASAP7_75t_R _0937_ (.A(_0094_),
    .Y(net210));
 INVx1_ASAP7_75t_R _0938_ (.A(_0095_),
    .Y(net209));
 INVx1_ASAP7_75t_R _0939_ (.A(_0096_),
    .Y(net208));
 INVx1_ASAP7_75t_R _0940_ (.A(_0097_),
    .Y(net207));
 INVx1_ASAP7_75t_R _0941_ (.A(_0098_),
    .Y(net206));
 INVx1_ASAP7_75t_R _0942_ (.A(_0099_),
    .Y(net205));
 INVx1_ASAP7_75t_R _0943_ (.A(_0100_),
    .Y(net204));
 INVx1_ASAP7_75t_R _0944_ (.A(_0101_),
    .Y(net203));
 INVx1_ASAP7_75t_R _0945_ (.A(_0102_),
    .Y(net202));
 INVx1_ASAP7_75t_R _0946_ (.A(_0103_),
    .Y(net201));
 INVx1_ASAP7_75t_R _0947_ (.A(_0104_),
    .Y(net200));
 INVx1_ASAP7_75t_R _0948_ (.A(_0105_),
    .Y(net199));
 INVx1_ASAP7_75t_R _0949_ (.A(_0106_),
    .Y(net198));
 INVx1_ASAP7_75t_R _0950_ (.A(_0107_),
    .Y(net197));
 INVx1_ASAP7_75t_R _0951_ (.A(_0108_),
    .Y(net196));
 INVx1_ASAP7_75t_R _0952_ (.A(_0109_),
    .Y(net195));
 INVx1_ASAP7_75t_R _0953_ (.A(_0110_),
    .Y(net194));
 INVx1_ASAP7_75t_R _0954_ (.A(_0111_),
    .Y(net193));
 INVx1_ASAP7_75t_R _0955_ (.A(_0112_),
    .Y(net192));
 INVx1_ASAP7_75t_R _0956_ (.A(_0113_),
    .Y(net191));
 INVx1_ASAP7_75t_R _0957_ (.A(_0114_),
    .Y(net190));
 INVx1_ASAP7_75t_R _0958_ (.A(_0116_),
    .Y(net187));
 INVx1_ASAP7_75t_R _0959_ (.A(_0117_),
    .Y(net186));
 INVx1_ASAP7_75t_R _0960_ (.A(_0118_),
    .Y(net185));
 INVx1_ASAP7_75t_R _0961_ (.A(_0119_),
    .Y(net184));
 INVx1_ASAP7_75t_R _0962_ (.A(_0120_),
    .Y(net183));
 INVx1_ASAP7_75t_R _0963_ (.A(_0121_),
    .Y(net182));
 INVx1_ASAP7_75t_R _0964_ (.A(_0122_),
    .Y(net181));
 INVx1_ASAP7_75t_R _0965_ (.A(_0123_),
    .Y(net180));
 INVx1_ASAP7_75t_R _0966_ (.A(_0124_),
    .Y(net179));
 INVx1_ASAP7_75t_R _0967_ (.A(_0125_),
    .Y(net178));
 INVx1_ASAP7_75t_R _0968_ (.A(_0126_),
    .Y(net177));
 INVx1_ASAP7_75t_R _0969_ (.A(_0127_),
    .Y(net176));
 INVx1_ASAP7_75t_R _0970_ (.A(_0128_),
    .Y(net175));
 INVx1_ASAP7_75t_R _0971_ (.A(_0129_),
    .Y(net174));
 INVx1_ASAP7_75t_R _0972_ (.A(_0130_),
    .Y(net173));
 INVx1_ASAP7_75t_R _0973_ (.A(_0131_),
    .Y(net172));
 INVx1_ASAP7_75t_R _0974_ (.A(_0132_),
    .Y(net171));
 INVx1_ASAP7_75t_R _0975_ (.A(_0133_),
    .Y(net170));
 INVx1_ASAP7_75t_R _0976_ (.A(_0134_),
    .Y(net169));
 INVx1_ASAP7_75t_R _0977_ (.A(_0135_),
    .Y(net168));
 INVx1_ASAP7_75t_R _0978_ (.A(_0136_),
    .Y(net167));
 INVx1_ASAP7_75t_R _0979_ (.A(_0137_),
    .Y(net166));
 INVx1_ASAP7_75t_R _0980_ (.A(_0138_),
    .Y(net165));
 INVx1_ASAP7_75t_R _0981_ (.A(_0139_),
    .Y(net164));
 INVx1_ASAP7_75t_R _0982_ (.A(_0140_),
    .Y(net163));
 INVx1_ASAP7_75t_R _0983_ (.A(_0141_),
    .Y(net162));
 INVx1_ASAP7_75t_R _0984_ (.A(_0142_),
    .Y(net161));
 INVx1_ASAP7_75t_R _0985_ (.A(_0143_),
    .Y(net160));
 INVx1_ASAP7_75t_R _0986_ (.A(_0144_),
    .Y(net159));
 INVx1_ASAP7_75t_R _0987_ (.A(_0145_),
    .Y(net158));
 INVx1_ASAP7_75t_R _0988_ (.A(_0146_),
    .Y(net157));
 INVx1_ASAP7_75t_R _0989_ (.A(_0147_),
    .Y(net156));
 INVx1_ASAP7_75t_R _0990_ (.A(_0148_),
    .Y(net155));
 INVx1_ASAP7_75t_R _0991_ (.A(_0149_),
    .Y(net154));
 INVx1_ASAP7_75t_R _0992_ (.A(_0150_),
    .Y(net153));
 INVx1_ASAP7_75t_R _0993_ (.A(_0151_),
    .Y(net152));
 INVx1_ASAP7_75t_R _0994_ (.A(_0152_),
    .Y(net188));
 NAND2x1_ASAP7_75t_R _0995_ (.A(_0569_),
    .B(_0570_),
    .Y(_0636_));
 AOI22x1_ASAP7_75t_R _0996_ (.A1(_0636_),
    .A2(_0604_),
    .B1(_0593_),
    .B2(_0595_),
    .Y(_0637_));
 OR2x2_ASAP7_75t_R _0997_ (.A(_0572_),
    .B(_0605_),
    .Y(_0638_));
 BUFx6f_ASAP7_75t_R _0998_ (.A(_0638_),
    .Y(_0639_));
 OR3x1_ASAP7_75t_R _0999_ (.A(_0568_),
    .B(_0573_),
    .C(_0604_),
    .Y(_0640_));
 OA21x2_ASAP7_75t_R _1000_ (.A1(_0637_),
    .A2(_0639_),
    .B(_0640_),
    .Y(_0641_));
 AOI211x1_ASAP7_75t_R _1001_ (.A1(_0610_),
    .A2(_0611_),
    .B(_0572_),
    .C(_0636_),
    .Y(_0642_));
 AO21x1_ASAP7_75t_R _1002_ (.A1(_0565_),
    .A2(_0155_),
    .B(_0604_),
    .Y(_0643_));
 AND3x1_ASAP7_75t_R _1003_ (.A(_0595_),
    .B(_0593_),
    .C(_0610_),
    .Y(_0644_));
 AO21x1_ASAP7_75t_R _1004_ (.A1(_0636_),
    .A2(_0643_),
    .B(_0644_),
    .Y(_0645_));
 AND2x2_ASAP7_75t_R _1005_ (.A(net149),
    .B(_0567_),
    .Y(_0646_));
 AO221x1_ASAP7_75t_R _1006_ (.A1(_0641_),
    .A2(_0642_),
    .B1(_0645_),
    .B2(_0646_),
    .C(_0572_),
    .Y(_0647_));
 BUFx6f_ASAP7_75t_R _1007_ (.A(_0647_),
    .Y(_0648_));
 BUFx6f_ASAP7_75t_R _1008_ (.A(_0648_),
    .Y(_0649_));
 BUFx12f_ASAP7_75t_R _1009_ (.A(_0572_),
    .Y(_0650_));
 BUFx6f_ASAP7_75t_R _1010_ (.A(_0650_),
    .Y(_0651_));
 OA211x2_ASAP7_75t_R _1011_ (.A1(_0637_),
    .A2(_0639_),
    .B(_0640_),
    .C(_0642_),
    .Y(_0652_));
 BUFx6f_ASAP7_75t_R _1012_ (.A(_0652_),
    .Y(_0653_));
 BUFx6f_ASAP7_75t_R _1013_ (.A(_0653_),
    .Y(_0654_));
 INVx1_ASAP7_75t_R _1014_ (.A(net76),
    .Y(_0655_));
 AOI221x1_ASAP7_75t_R _1015_ (.A1(_0651_),
    .A2(_0151_),
    .B1(_0654_),
    .B2(_0655_),
    .C(_0631_),
    .Y(_0656_));
 BUFx6f_ASAP7_75t_R _1016_ (.A(_0639_),
    .Y(_0657_));
 AOI21x1_ASAP7_75t_R _1017_ (.A1(_0636_),
    .A2(_0643_),
    .B(_0644_),
    .Y(_0658_));
 BUFx6f_ASAP7_75t_R _1018_ (.A(_0658_),
    .Y(_0659_));
 OR3x1_ASAP7_75t_R _1019_ (.A(net113),
    .B(_0657_),
    .C(_0659_),
    .Y(_0660_));
 OA211x2_ASAP7_75t_R _1020_ (.A1(net38),
    .A2(_0649_),
    .B(_0656_),
    .C(_0660_),
    .Y(_0156_));
 INVx1_ASAP7_75t_R _1021_ (.A(net77),
    .Y(_0661_));
 AOI221x1_ASAP7_75t_R _1022_ (.A1(_0651_),
    .A2(_0150_),
    .B1(_0654_),
    .B2(_0661_),
    .C(_0631_),
    .Y(_0662_));
 OR3x1_ASAP7_75t_R _1023_ (.A(net114),
    .B(_0657_),
    .C(_0659_),
    .Y(_0663_));
 OA211x2_ASAP7_75t_R _1024_ (.A1(net39),
    .A2(_0649_),
    .B(_0662_),
    .C(_0663_),
    .Y(_0157_));
 INVx1_ASAP7_75t_R _1025_ (.A(net78),
    .Y(_0664_));
 AOI221x1_ASAP7_75t_R _1026_ (.A1(_0651_),
    .A2(_0149_),
    .B1(_0654_),
    .B2(_0664_),
    .C(_0631_),
    .Y(_0665_));
 OR3x1_ASAP7_75t_R _1027_ (.A(net115),
    .B(_0657_),
    .C(_0659_),
    .Y(_0666_));
 OA211x2_ASAP7_75t_R _1028_ (.A1(net40),
    .A2(_0649_),
    .B(_0665_),
    .C(_0666_),
    .Y(_0158_));
 INVx1_ASAP7_75t_R _1029_ (.A(net79),
    .Y(_0667_));
 AOI221x1_ASAP7_75t_R _1030_ (.A1(_0651_),
    .A2(_0148_),
    .B1(_0654_),
    .B2(_0667_),
    .C(_0631_),
    .Y(_0668_));
 OR3x1_ASAP7_75t_R _1031_ (.A(net116),
    .B(_0657_),
    .C(_0659_),
    .Y(_0669_));
 OA211x2_ASAP7_75t_R _1032_ (.A1(net41),
    .A2(_0649_),
    .B(_0668_),
    .C(_0669_),
    .Y(_0159_));
 INVx1_ASAP7_75t_R _1033_ (.A(net80),
    .Y(_0670_));
 AOI221x1_ASAP7_75t_R _1034_ (.A1(_0651_),
    .A2(_0147_),
    .B1(_0654_),
    .B2(_0670_),
    .C(_0631_),
    .Y(_0671_));
 OR3x1_ASAP7_75t_R _1035_ (.A(net117),
    .B(_0657_),
    .C(_0659_),
    .Y(_0672_));
 OA211x2_ASAP7_75t_R _1036_ (.A1(net42),
    .A2(_0649_),
    .B(_0671_),
    .C(_0672_),
    .Y(_0160_));
 INVx1_ASAP7_75t_R _1037_ (.A(net81),
    .Y(_0673_));
 BUFx6f_ASAP7_75t_R _1038_ (.A(_0621_),
    .Y(_0674_));
 AOI221x1_ASAP7_75t_R _1039_ (.A1(_0651_),
    .A2(_0146_),
    .B1(_0654_),
    .B2(_0673_),
    .C(_0674_),
    .Y(_0675_));
 OR3x1_ASAP7_75t_R _1040_ (.A(net118),
    .B(_0657_),
    .C(_0659_),
    .Y(_0676_));
 OA211x2_ASAP7_75t_R _1041_ (.A1(net43),
    .A2(_0649_),
    .B(_0675_),
    .C(_0676_),
    .Y(_0161_));
 INVx1_ASAP7_75t_R _1042_ (.A(net82),
    .Y(_0677_));
 AOI221x1_ASAP7_75t_R _1043_ (.A1(_0651_),
    .A2(_0145_),
    .B1(_0654_),
    .B2(_0677_),
    .C(_0674_),
    .Y(_0678_));
 OR3x1_ASAP7_75t_R _1044_ (.A(net119),
    .B(_0657_),
    .C(_0659_),
    .Y(_0679_));
 OA211x2_ASAP7_75t_R _1045_ (.A1(net44),
    .A2(_0649_),
    .B(_0678_),
    .C(_0679_),
    .Y(_0162_));
 INVx1_ASAP7_75t_R _1046_ (.A(net83),
    .Y(_0680_));
 AOI221x1_ASAP7_75t_R _1047_ (.A1(_0651_),
    .A2(_0144_),
    .B1(_0654_),
    .B2(_0680_),
    .C(_0674_),
    .Y(_0681_));
 OR3x1_ASAP7_75t_R _1048_ (.A(net120),
    .B(_0657_),
    .C(_0659_),
    .Y(_0682_));
 OA211x2_ASAP7_75t_R _1049_ (.A1(net45),
    .A2(_0649_),
    .B(_0681_),
    .C(_0682_),
    .Y(_0163_));
 BUFx6f_ASAP7_75t_R _1050_ (.A(_0650_),
    .Y(_0683_));
 INVx1_ASAP7_75t_R _1051_ (.A(net84),
    .Y(_0684_));
 AOI221x1_ASAP7_75t_R _1052_ (.A1(_0683_),
    .A2(_0143_),
    .B1(_0654_),
    .B2(_0684_),
    .C(_0674_),
    .Y(_0685_));
 OR3x1_ASAP7_75t_R _1053_ (.A(net121),
    .B(_0657_),
    .C(_0659_),
    .Y(_0686_));
 OA211x2_ASAP7_75t_R _1054_ (.A1(net46),
    .A2(_0649_),
    .B(_0685_),
    .C(_0686_),
    .Y(_0164_));
 BUFx6f_ASAP7_75t_R _1055_ (.A(_0648_),
    .Y(_0687_));
 INVx1_ASAP7_75t_R _1056_ (.A(net85),
    .Y(_0688_));
 AOI221x1_ASAP7_75t_R _1057_ (.A1(_0683_),
    .A2(_0142_),
    .B1(_0654_),
    .B2(_0688_),
    .C(_0674_),
    .Y(_0689_));
 OR3x1_ASAP7_75t_R _1058_ (.A(net122),
    .B(_0657_),
    .C(_0659_),
    .Y(_0690_));
 OA211x2_ASAP7_75t_R _1059_ (.A1(net47),
    .A2(_0687_),
    .B(_0689_),
    .C(_0690_),
    .Y(_0165_));
 BUFx6f_ASAP7_75t_R _1060_ (.A(_0653_),
    .Y(_0691_));
 INVx1_ASAP7_75t_R _1061_ (.A(net86),
    .Y(_0692_));
 AOI221x1_ASAP7_75t_R _1062_ (.A1(_0683_),
    .A2(_0141_),
    .B1(_0691_),
    .B2(_0692_),
    .C(_0674_),
    .Y(_0693_));
 BUFx6f_ASAP7_75t_R _1063_ (.A(_0639_),
    .Y(_0694_));
 BUFx6f_ASAP7_75t_R _1064_ (.A(_0658_),
    .Y(_0695_));
 OR3x1_ASAP7_75t_R _1065_ (.A(net123),
    .B(_0694_),
    .C(_0695_),
    .Y(_0696_));
 OA211x2_ASAP7_75t_R _1066_ (.A1(net48),
    .A2(_0687_),
    .B(_0693_),
    .C(_0696_),
    .Y(_0166_));
 INVx1_ASAP7_75t_R _1067_ (.A(net87),
    .Y(_0697_));
 AOI221x1_ASAP7_75t_R _1068_ (.A1(_0683_),
    .A2(_0140_),
    .B1(_0691_),
    .B2(_0697_),
    .C(_0674_),
    .Y(_0698_));
 OR3x1_ASAP7_75t_R _1069_ (.A(net124),
    .B(_0694_),
    .C(_0695_),
    .Y(_0699_));
 OA211x2_ASAP7_75t_R _1070_ (.A1(net49),
    .A2(_0687_),
    .B(_0698_),
    .C(_0699_),
    .Y(_0167_));
 INVx1_ASAP7_75t_R _1071_ (.A(net88),
    .Y(_0700_));
 AOI221x1_ASAP7_75t_R _1072_ (.A1(_0683_),
    .A2(_0139_),
    .B1(_0691_),
    .B2(_0700_),
    .C(_0674_),
    .Y(_0701_));
 OR3x1_ASAP7_75t_R _1073_ (.A(net125),
    .B(_0694_),
    .C(_0695_),
    .Y(_0702_));
 OA211x2_ASAP7_75t_R _1074_ (.A1(net50),
    .A2(_0687_),
    .B(_0701_),
    .C(_0702_),
    .Y(_0168_));
 INVx1_ASAP7_75t_R _1075_ (.A(net89),
    .Y(_0703_));
 AOI221x1_ASAP7_75t_R _1076_ (.A1(_0683_),
    .A2(_0138_),
    .B1(_0691_),
    .B2(_0703_),
    .C(_0674_),
    .Y(_0704_));
 OR3x1_ASAP7_75t_R _1077_ (.A(net126),
    .B(_0694_),
    .C(_0695_),
    .Y(_0705_));
 OA211x2_ASAP7_75t_R _1078_ (.A1(net51),
    .A2(_0687_),
    .B(_0704_),
    .C(_0705_),
    .Y(_0169_));
 INVx1_ASAP7_75t_R _1079_ (.A(net90),
    .Y(_0706_));
 AOI221x1_ASAP7_75t_R _1080_ (.A1(_0683_),
    .A2(_0137_),
    .B1(_0691_),
    .B2(_0706_),
    .C(_0674_),
    .Y(_0707_));
 OR3x1_ASAP7_75t_R _1081_ (.A(net127),
    .B(_0694_),
    .C(_0695_),
    .Y(_0708_));
 OA211x2_ASAP7_75t_R _1082_ (.A1(net52),
    .A2(_0687_),
    .B(_0707_),
    .C(_0708_),
    .Y(_0170_));
 INVx1_ASAP7_75t_R _1083_ (.A(net91),
    .Y(_0709_));
 BUFx6f_ASAP7_75t_R _1084_ (.A(_0621_),
    .Y(_0710_));
 AOI221x1_ASAP7_75t_R _1085_ (.A1(_0683_),
    .A2(_0136_),
    .B1(_0691_),
    .B2(_0709_),
    .C(_0710_),
    .Y(_0711_));
 OR3x1_ASAP7_75t_R _1086_ (.A(net128),
    .B(_0694_),
    .C(_0695_),
    .Y(_0712_));
 OA211x2_ASAP7_75t_R _1087_ (.A1(net53),
    .A2(_0687_),
    .B(_0711_),
    .C(_0712_),
    .Y(_0171_));
 INVx1_ASAP7_75t_R _1088_ (.A(net92),
    .Y(_0713_));
 AOI221x1_ASAP7_75t_R _1089_ (.A1(_0683_),
    .A2(_0135_),
    .B1(_0691_),
    .B2(_0713_),
    .C(_0710_),
    .Y(_0714_));
 OR3x1_ASAP7_75t_R _1090_ (.A(net129),
    .B(_0694_),
    .C(_0695_),
    .Y(_0715_));
 OA211x2_ASAP7_75t_R _1091_ (.A1(net54),
    .A2(_0687_),
    .B(_0714_),
    .C(_0715_),
    .Y(_0172_));
 INVx1_ASAP7_75t_R _1092_ (.A(net93),
    .Y(_0716_));
 AOI221x1_ASAP7_75t_R _1093_ (.A1(_0683_),
    .A2(_0134_),
    .B1(_0691_),
    .B2(_0716_),
    .C(_0710_),
    .Y(_0717_));
 OR3x1_ASAP7_75t_R _1094_ (.A(net130),
    .B(_0694_),
    .C(_0695_),
    .Y(_0718_));
 OA211x2_ASAP7_75t_R _1095_ (.A1(net55),
    .A2(_0687_),
    .B(_0717_),
    .C(_0718_),
    .Y(_0173_));
 BUFx6f_ASAP7_75t_R _1096_ (.A(_0650_),
    .Y(_0719_));
 INVx1_ASAP7_75t_R _1097_ (.A(net94),
    .Y(_0720_));
 AOI221x1_ASAP7_75t_R _1098_ (.A1(_0719_),
    .A2(_0133_),
    .B1(_0691_),
    .B2(_0720_),
    .C(_0710_),
    .Y(_0721_));
 OR3x1_ASAP7_75t_R _1099_ (.A(net131),
    .B(_0694_),
    .C(_0695_),
    .Y(_0722_));
 OA211x2_ASAP7_75t_R _1100_ (.A1(net56),
    .A2(_0687_),
    .B(_0721_),
    .C(_0722_),
    .Y(_0174_));
 BUFx6f_ASAP7_75t_R _1101_ (.A(_0648_),
    .Y(_0723_));
 INVx1_ASAP7_75t_R _1102_ (.A(net95),
    .Y(_0724_));
 AOI221x1_ASAP7_75t_R _1103_ (.A1(_0719_),
    .A2(_0132_),
    .B1(_0691_),
    .B2(_0724_),
    .C(_0710_),
    .Y(_0725_));
 OR3x1_ASAP7_75t_R _1104_ (.A(net132),
    .B(_0694_),
    .C(_0695_),
    .Y(_0726_));
 OA211x2_ASAP7_75t_R _1105_ (.A1(net57),
    .A2(_0723_),
    .B(_0725_),
    .C(_0726_),
    .Y(_0175_));
 BUFx6f_ASAP7_75t_R _1106_ (.A(_0653_),
    .Y(_0727_));
 INVx1_ASAP7_75t_R _1107_ (.A(net96),
    .Y(_0728_));
 AOI221x1_ASAP7_75t_R _1108_ (.A1(_0719_),
    .A2(_0131_),
    .B1(_0727_),
    .B2(_0728_),
    .C(_0710_),
    .Y(_0729_));
 BUFx6f_ASAP7_75t_R _1109_ (.A(_0639_),
    .Y(_0730_));
 BUFx6f_ASAP7_75t_R _1110_ (.A(_0658_),
    .Y(_0731_));
 OR3x1_ASAP7_75t_R _1111_ (.A(net133),
    .B(_0730_),
    .C(_0731_),
    .Y(_0732_));
 OA211x2_ASAP7_75t_R _1112_ (.A1(net58),
    .A2(_0723_),
    .B(_0729_),
    .C(_0732_),
    .Y(_0176_));
 INVx1_ASAP7_75t_R _1113_ (.A(net97),
    .Y(_0733_));
 AOI221x1_ASAP7_75t_R _1114_ (.A1(_0719_),
    .A2(_0130_),
    .B1(_0727_),
    .B2(_0733_),
    .C(_0710_),
    .Y(_0734_));
 OR3x1_ASAP7_75t_R _1115_ (.A(net134),
    .B(_0730_),
    .C(_0731_),
    .Y(_0735_));
 OA211x2_ASAP7_75t_R _1116_ (.A1(net59),
    .A2(_0723_),
    .B(_0734_),
    .C(_0735_),
    .Y(_0177_));
 INVx1_ASAP7_75t_R _1117_ (.A(net98),
    .Y(_0736_));
 AOI221x1_ASAP7_75t_R _1118_ (.A1(_0719_),
    .A2(_0129_),
    .B1(_0727_),
    .B2(_0736_),
    .C(_0710_),
    .Y(_0737_));
 OR3x1_ASAP7_75t_R _1119_ (.A(net135),
    .B(_0730_),
    .C(_0731_),
    .Y(_0738_));
 OA211x2_ASAP7_75t_R _1120_ (.A1(net60),
    .A2(_0723_),
    .B(_0737_),
    .C(_0738_),
    .Y(_0178_));
 INVx1_ASAP7_75t_R _1121_ (.A(net99),
    .Y(_0739_));
 AOI221x1_ASAP7_75t_R _1122_ (.A1(_0719_),
    .A2(_0128_),
    .B1(_0727_),
    .B2(_0739_),
    .C(_0710_),
    .Y(_0740_));
 OR3x1_ASAP7_75t_R _1123_ (.A(net136),
    .B(_0730_),
    .C(_0731_),
    .Y(_0741_));
 OA211x2_ASAP7_75t_R _1124_ (.A1(net61),
    .A2(_0723_),
    .B(_0740_),
    .C(_0741_),
    .Y(_0179_));
 INVx1_ASAP7_75t_R _1125_ (.A(net100),
    .Y(_0742_));
 AOI221x1_ASAP7_75t_R _1126_ (.A1(_0719_),
    .A2(_0127_),
    .B1(_0727_),
    .B2(_0742_),
    .C(_0710_),
    .Y(_0743_));
 OR3x1_ASAP7_75t_R _1127_ (.A(net137),
    .B(_0730_),
    .C(_0731_),
    .Y(_0744_));
 OA211x2_ASAP7_75t_R _1128_ (.A1(net62),
    .A2(_0723_),
    .B(_0743_),
    .C(_0744_),
    .Y(_0180_));
 NAND2x1_ASAP7_75t_R _1129_ (.A(net63),
    .B(_0626_),
    .Y(_0745_));
 NAND2x1_ASAP7_75t_R _1130_ (.A(_0651_),
    .B(_0624_),
    .Y(_0746_));
 OAI22x1_ASAP7_75t_R _1131_ (.A1(_0649_),
    .A2(_0745_),
    .B1(_0746_),
    .B2(_0126_),
    .Y(_0181_));
 INVx1_ASAP7_75t_R _1132_ (.A(net102),
    .Y(_0747_));
 BUFx6f_ASAP7_75t_R _1133_ (.A(_0621_),
    .Y(_0748_));
 AOI221x1_ASAP7_75t_R _1134_ (.A1(_0719_),
    .A2(_0125_),
    .B1(_0727_),
    .B2(_0747_),
    .C(_0748_),
    .Y(_0749_));
 OR3x1_ASAP7_75t_R _1135_ (.A(net139),
    .B(_0730_),
    .C(_0731_),
    .Y(_0750_));
 OA211x2_ASAP7_75t_R _1136_ (.A1(net64),
    .A2(_0723_),
    .B(_0749_),
    .C(_0750_),
    .Y(_0182_));
 INVx1_ASAP7_75t_R _1137_ (.A(net103),
    .Y(_0751_));
 AOI221x1_ASAP7_75t_R _1138_ (.A1(_0719_),
    .A2(_0124_),
    .B1(_0727_),
    .B2(_0751_),
    .C(_0748_),
    .Y(_0752_));
 OR3x1_ASAP7_75t_R _1139_ (.A(net140),
    .B(_0730_),
    .C(_0731_),
    .Y(_0753_));
 OA211x2_ASAP7_75t_R _1140_ (.A1(net65),
    .A2(_0723_),
    .B(_0752_),
    .C(_0753_),
    .Y(_0183_));
 INVx1_ASAP7_75t_R _1141_ (.A(net104),
    .Y(_0754_));
 AOI221x1_ASAP7_75t_R _1142_ (.A1(_0719_),
    .A2(_0123_),
    .B1(_0727_),
    .B2(_0754_),
    .C(_0748_),
    .Y(_0755_));
 OR3x1_ASAP7_75t_R _1143_ (.A(net141),
    .B(_0730_),
    .C(_0731_),
    .Y(_0756_));
 OA211x2_ASAP7_75t_R _1144_ (.A1(net66),
    .A2(_0723_),
    .B(_0755_),
    .C(_0756_),
    .Y(_0184_));
 INVx1_ASAP7_75t_R _1145_ (.A(net105),
    .Y(_0757_));
 AOI221x1_ASAP7_75t_R _1146_ (.A1(_0650_),
    .A2(_0122_),
    .B1(_0727_),
    .B2(_0757_),
    .C(_0748_),
    .Y(_0758_));
 OR3x1_ASAP7_75t_R _1147_ (.A(net142),
    .B(_0730_),
    .C(_0731_),
    .Y(_0759_));
 OA211x2_ASAP7_75t_R _1148_ (.A1(net67),
    .A2(_0723_),
    .B(_0758_),
    .C(_0759_),
    .Y(_0185_));
 INVx1_ASAP7_75t_R _1149_ (.A(net106),
    .Y(_0760_));
 AOI221x1_ASAP7_75t_R _1150_ (.A1(_0650_),
    .A2(_0121_),
    .B1(_0727_),
    .B2(_0760_),
    .C(_0748_),
    .Y(_0761_));
 OR3x1_ASAP7_75t_R _1151_ (.A(net143),
    .B(_0730_),
    .C(_0731_),
    .Y(_0762_));
 OA211x2_ASAP7_75t_R _1152_ (.A1(net68),
    .A2(_0648_),
    .B(_0761_),
    .C(_0762_),
    .Y(_0186_));
 INVx1_ASAP7_75t_R _1153_ (.A(net107),
    .Y(_0763_));
 AOI221x1_ASAP7_75t_R _1154_ (.A1(_0650_),
    .A2(_0120_),
    .B1(_0653_),
    .B2(_0763_),
    .C(_0748_),
    .Y(_0764_));
 OR3x1_ASAP7_75t_R _1155_ (.A(net144),
    .B(_0639_),
    .C(_0658_),
    .Y(_0765_));
 OA211x2_ASAP7_75t_R _1156_ (.A1(net69),
    .A2(_0648_),
    .B(_0764_),
    .C(_0765_),
    .Y(_0187_));
 INVx1_ASAP7_75t_R _1157_ (.A(net108),
    .Y(_0304_));
 AOI221x1_ASAP7_75t_R _1158_ (.A1(_0650_),
    .A2(_0119_),
    .B1(_0653_),
    .B2(_0304_),
    .C(_0748_),
    .Y(_0305_));
 OR3x1_ASAP7_75t_R _1159_ (.A(net145),
    .B(_0639_),
    .C(_0658_),
    .Y(_0306_));
 OA211x2_ASAP7_75t_R _1160_ (.A1(net70),
    .A2(_0648_),
    .B(_0305_),
    .C(_0306_),
    .Y(_0188_));
 INVx1_ASAP7_75t_R _1161_ (.A(net109),
    .Y(_0307_));
 AOI221x1_ASAP7_75t_R _1162_ (.A1(_0650_),
    .A2(_0118_),
    .B1(_0653_),
    .B2(_0307_),
    .C(_0748_),
    .Y(_0308_));
 OR3x1_ASAP7_75t_R _1163_ (.A(net146),
    .B(_0639_),
    .C(_0658_),
    .Y(_0309_));
 OA211x2_ASAP7_75t_R _1164_ (.A1(net71),
    .A2(_0648_),
    .B(_0308_),
    .C(_0309_),
    .Y(_0189_));
 INVx1_ASAP7_75t_R _1165_ (.A(net110),
    .Y(_0310_));
 AOI221x1_ASAP7_75t_R _1166_ (.A1(_0650_),
    .A2(_0117_),
    .B1(_0653_),
    .B2(_0310_),
    .C(_0748_),
    .Y(_0311_));
 OR3x1_ASAP7_75t_R _1167_ (.A(net147),
    .B(_0639_),
    .C(_0658_),
    .Y(_0312_));
 OA211x2_ASAP7_75t_R _1168_ (.A1(net72),
    .A2(_0648_),
    .B(_0311_),
    .C(_0312_),
    .Y(_0190_));
 INVx1_ASAP7_75t_R _1169_ (.A(net111),
    .Y(_0313_));
 AOI221x1_ASAP7_75t_R _1170_ (.A1(_0650_),
    .A2(_0116_),
    .B1(_0653_),
    .B2(_0313_),
    .C(_0748_),
    .Y(_0314_));
 OR3x1_ASAP7_75t_R _1171_ (.A(net148),
    .B(_0639_),
    .C(_0658_),
    .Y(_0315_));
 OA211x2_ASAP7_75t_R _1172_ (.A1(net73),
    .A2(_0648_),
    .B(_0314_),
    .C(_0315_),
    .Y(_0191_));
 AOI21x1_ASAP7_75t_R _1173_ (.A1(_0651_),
    .A2(net188),
    .B(_0642_),
    .Y(_0316_));
 AOI21x1_ASAP7_75t_R _1174_ (.A1(_0641_),
    .A2(_0316_),
    .B(_0631_),
    .Y(_0192_));
 BUFx6f_ASAP7_75t_R _1175_ (.A(_0594_),
    .Y(_0317_));
 OA21x2_ASAP7_75t_R _1176_ (.A1(_0317_),
    .A2(net190),
    .B(_0622_),
    .Y(_0318_));
 AO21x1_ASAP7_75t_R _1177_ (.A1(_0595_),
    .A2(_0593_),
    .B(_0599_),
    .Y(_0319_));
 AO31x2_ASAP7_75t_R _1178_ (.A1(_0595_),
    .A2(_0593_),
    .A3(_0610_),
    .B(_0597_),
    .Y(_0320_));
 OR3x1_ASAP7_75t_R _1179_ (.A(_0580_),
    .B(_0583_),
    .C(_0599_),
    .Y(_0321_));
 AND4x1_ASAP7_75t_R _1180_ (.A(_0582_),
    .B(_0319_),
    .C(_0320_),
    .D(_0321_),
    .Y(_0322_));
 BUFx6f_ASAP7_75t_R _1181_ (.A(_0322_),
    .Y(_0323_));
 OA21x2_ASAP7_75t_R _1182_ (.A1(_0609_),
    .A2(_0600_),
    .B(_0599_),
    .Y(_0324_));
 OA211x2_ASAP7_75t_R _1183_ (.A1(_0153_),
    .A2(_0599_),
    .B(_0579_),
    .C(_0594_),
    .Y(_0325_));
 AND4x1_ASAP7_75t_R _1184_ (.A(net74),
    .B(_0574_),
    .C(_0616_),
    .D(_0575_),
    .Y(_0326_));
 OR3x1_ASAP7_75t_R _1185_ (.A(_0571_),
    .B(_0600_),
    .C(_0326_),
    .Y(_0327_));
 OA211x2_ASAP7_75t_R _1186_ (.A1(_0578_),
    .A2(_0324_),
    .B(_0325_),
    .C(_0327_),
    .Y(_0328_));
 BUFx6f_ASAP7_75t_R _1187_ (.A(_0328_),
    .Y(_0329_));
 BUFx6f_ASAP7_75t_R _1188_ (.A(_0329_),
    .Y(_0330_));
 BUFx6f_ASAP7_75t_R _1189_ (.A(net75),
    .Y(_0331_));
 AO221x1_ASAP7_75t_R _1190_ (.A1(net113),
    .A2(_0323_),
    .B1(_0330_),
    .B2(net76),
    .C(_0331_),
    .Y(_0332_));
 NOR2x1_ASAP7_75t_R _1191_ (.A(_0584_),
    .B(_0599_),
    .Y(_0333_));
 AND3x1_ASAP7_75t_R _1192_ (.A(_0585_),
    .B(_0600_),
    .C(_0586_),
    .Y(_0334_));
 OA211x2_ASAP7_75t_R _1193_ (.A1(_0571_),
    .A2(_0326_),
    .B(_0582_),
    .C(_0579_),
    .Y(_0335_));
 OA21x2_ASAP7_75t_R _1194_ (.A1(_0334_),
    .A2(_0335_),
    .B(_0610_),
    .Y(_0336_));
 AOI21x1_ASAP7_75t_R _1195_ (.A1(_0582_),
    .A2(_0319_),
    .B(_0579_),
    .Y(_0337_));
 OR2x2_ASAP7_75t_R _1196_ (.A(_0597_),
    .B(_0610_),
    .Y(_0338_));
 OAI21x1_ASAP7_75t_R _1197_ (.A1(_0327_),
    .A2(_0338_),
    .B(_0317_),
    .Y(_0339_));
 OR4x1_ASAP7_75t_R _1198_ (.A(_0333_),
    .B(_0336_),
    .C(_0337_),
    .D(_0339_),
    .Y(_0340_));
 BUFx6f_ASAP7_75t_R _1199_ (.A(_0340_),
    .Y(_0341_));
 AND2x2_ASAP7_75t_R _1200_ (.A(net1),
    .B(_0318_),
    .Y(_0342_));
 AO22x1_ASAP7_75t_R _1201_ (.A1(_0318_),
    .A2(_0332_),
    .B1(_0341_),
    .B2(_0342_),
    .Y(_0193_));
 BUFx6f_ASAP7_75t_R _1202_ (.A(_0317_),
    .Y(_0343_));
 OA21x2_ASAP7_75t_R _1203_ (.A1(_0343_),
    .A2(net191),
    .B(_0623_),
    .Y(_0344_));
 AO221x1_ASAP7_75t_R _1204_ (.A1(net114),
    .A2(_0323_),
    .B1(_0330_),
    .B2(net77),
    .C(_0331_),
    .Y(_0345_));
 AND2x2_ASAP7_75t_R _1205_ (.A(net2),
    .B(_0344_),
    .Y(_0346_));
 AO22x1_ASAP7_75t_R _1206_ (.A1(_0344_),
    .A2(_0345_),
    .B1(_0346_),
    .B2(_0341_),
    .Y(_0194_));
 OA21x2_ASAP7_75t_R _1207_ (.A1(_0343_),
    .A2(net192),
    .B(_0623_),
    .Y(_0347_));
 AO221x1_ASAP7_75t_R _1208_ (.A1(net115),
    .A2(_0323_),
    .B1(_0330_),
    .B2(net78),
    .C(_0331_),
    .Y(_0348_));
 AND2x2_ASAP7_75t_R _1209_ (.A(net3),
    .B(_0347_),
    .Y(_0349_));
 AO22x1_ASAP7_75t_R _1210_ (.A1(_0347_),
    .A2(_0348_),
    .B1(_0349_),
    .B2(_0341_),
    .Y(_0195_));
 BUFx6f_ASAP7_75t_R _1211_ (.A(_0622_),
    .Y(_0350_));
 OA21x2_ASAP7_75t_R _1212_ (.A1(_0343_),
    .A2(net193),
    .B(_0350_),
    .Y(_0351_));
 AO221x1_ASAP7_75t_R _1213_ (.A1(net116),
    .A2(_0323_),
    .B1(_0330_),
    .B2(net79),
    .C(_0331_),
    .Y(_0352_));
 AND2x2_ASAP7_75t_R _1214_ (.A(net4),
    .B(_0351_),
    .Y(_0353_));
 AO22x1_ASAP7_75t_R _1215_ (.A1(_0351_),
    .A2(_0352_),
    .B1(_0353_),
    .B2(_0341_),
    .Y(_0196_));
 OA21x2_ASAP7_75t_R _1216_ (.A1(_0343_),
    .A2(net194),
    .B(_0350_),
    .Y(_0354_));
 AO221x1_ASAP7_75t_R _1217_ (.A1(net117),
    .A2(_0323_),
    .B1(_0330_),
    .B2(net80),
    .C(_0331_),
    .Y(_0355_));
 AND2x2_ASAP7_75t_R _1218_ (.A(net5),
    .B(_0354_),
    .Y(_0356_));
 AO22x1_ASAP7_75t_R _1219_ (.A1(_0354_),
    .A2(_0355_),
    .B1(_0356_),
    .B2(_0341_),
    .Y(_0197_));
 OA21x2_ASAP7_75t_R _1220_ (.A1(_0343_),
    .A2(net195),
    .B(_0350_),
    .Y(_0357_));
 AO221x1_ASAP7_75t_R _1221_ (.A1(net118),
    .A2(_0323_),
    .B1(_0330_),
    .B2(net81),
    .C(_0331_),
    .Y(_0358_));
 AND2x2_ASAP7_75t_R _1222_ (.A(net6),
    .B(_0357_),
    .Y(_0359_));
 AO22x1_ASAP7_75t_R _1223_ (.A1(_0357_),
    .A2(_0358_),
    .B1(_0359_),
    .B2(_0341_),
    .Y(_0198_));
 OA21x2_ASAP7_75t_R _1224_ (.A1(_0343_),
    .A2(net196),
    .B(_0350_),
    .Y(_0360_));
 AO221x1_ASAP7_75t_R _1225_ (.A1(net119),
    .A2(_0323_),
    .B1(_0330_),
    .B2(net82),
    .C(_0331_),
    .Y(_0361_));
 AND2x2_ASAP7_75t_R _1226_ (.A(net7),
    .B(_0360_),
    .Y(_0362_));
 AO22x1_ASAP7_75t_R _1227_ (.A1(_0360_),
    .A2(_0361_),
    .B1(_0362_),
    .B2(_0341_),
    .Y(_0199_));
 OA21x2_ASAP7_75t_R _1228_ (.A1(_0343_),
    .A2(net197),
    .B(_0350_),
    .Y(_0363_));
 BUFx6f_ASAP7_75t_R _1229_ (.A(net75),
    .Y(_0364_));
 BUFx6f_ASAP7_75t_R _1230_ (.A(_0364_),
    .Y(_0365_));
 AO221x1_ASAP7_75t_R _1231_ (.A1(net120),
    .A2(_0323_),
    .B1(_0330_),
    .B2(net83),
    .C(_0365_),
    .Y(_0366_));
 AND2x2_ASAP7_75t_R _1232_ (.A(net8),
    .B(_0363_),
    .Y(_0367_));
 AO22x1_ASAP7_75t_R _1233_ (.A1(_0363_),
    .A2(_0366_),
    .B1(_0367_),
    .B2(_0341_),
    .Y(_0200_));
 OA21x2_ASAP7_75t_R _1234_ (.A1(_0343_),
    .A2(net198),
    .B(_0350_),
    .Y(_0368_));
 AO221x1_ASAP7_75t_R _1235_ (.A1(net121),
    .A2(_0323_),
    .B1(_0330_),
    .B2(net84),
    .C(_0365_),
    .Y(_0369_));
 AND2x2_ASAP7_75t_R _1236_ (.A(net9),
    .B(_0368_),
    .Y(_0370_));
 AO22x1_ASAP7_75t_R _1237_ (.A1(_0368_),
    .A2(_0369_),
    .B1(_0370_),
    .B2(_0341_),
    .Y(_0201_));
 OA21x2_ASAP7_75t_R _1238_ (.A1(_0343_),
    .A2(net199),
    .B(_0350_),
    .Y(_0371_));
 AO221x1_ASAP7_75t_R _1239_ (.A1(net122),
    .A2(_0323_),
    .B1(_0330_),
    .B2(net85),
    .C(_0365_),
    .Y(_0372_));
 AND2x2_ASAP7_75t_R _1240_ (.A(net10),
    .B(_0371_),
    .Y(_0373_));
 AO22x1_ASAP7_75t_R _1241_ (.A1(_0371_),
    .A2(_0372_),
    .B1(_0373_),
    .B2(_0341_),
    .Y(_0202_));
 BUFx6f_ASAP7_75t_R _1242_ (.A(_0317_),
    .Y(_0374_));
 OA21x2_ASAP7_75t_R _1243_ (.A1(_0374_),
    .A2(net200),
    .B(_0350_),
    .Y(_0375_));
 BUFx6f_ASAP7_75t_R _1244_ (.A(_0322_),
    .Y(_0376_));
 BUFx6f_ASAP7_75t_R _1245_ (.A(_0329_),
    .Y(_0377_));
 AO221x1_ASAP7_75t_R _1246_ (.A1(net123),
    .A2(_0376_),
    .B1(_0377_),
    .B2(net86),
    .C(_0365_),
    .Y(_0378_));
 AND2x2_ASAP7_75t_R _1247_ (.A(net11),
    .B(_0375_),
    .Y(_0379_));
 BUFx6f_ASAP7_75t_R _1248_ (.A(_0340_),
    .Y(_0380_));
 AO22x1_ASAP7_75t_R _1249_ (.A1(_0375_),
    .A2(_0378_),
    .B1(_0379_),
    .B2(_0380_),
    .Y(_0203_));
 OA21x2_ASAP7_75t_R _1250_ (.A1(_0374_),
    .A2(net201),
    .B(_0350_),
    .Y(_0381_));
 AO221x1_ASAP7_75t_R _1251_ (.A1(net124),
    .A2(_0376_),
    .B1(_0377_),
    .B2(net87),
    .C(_0365_),
    .Y(_0382_));
 AND2x2_ASAP7_75t_R _1252_ (.A(net12),
    .B(_0381_),
    .Y(_0383_));
 AO22x1_ASAP7_75t_R _1253_ (.A1(_0381_),
    .A2(_0382_),
    .B1(_0383_),
    .B2(_0380_),
    .Y(_0204_));
 OA21x2_ASAP7_75t_R _1254_ (.A1(_0374_),
    .A2(net202),
    .B(_0350_),
    .Y(_0384_));
 AO221x1_ASAP7_75t_R _1255_ (.A1(net125),
    .A2(_0376_),
    .B1(_0377_),
    .B2(net88),
    .C(_0365_),
    .Y(_0385_));
 AND2x2_ASAP7_75t_R _1256_ (.A(net13),
    .B(_0384_),
    .Y(_0386_));
 AO22x1_ASAP7_75t_R _1257_ (.A1(_0384_),
    .A2(_0385_),
    .B1(_0386_),
    .B2(_0380_),
    .Y(_0205_));
 BUFx6f_ASAP7_75t_R _1258_ (.A(_0622_),
    .Y(_0387_));
 OA21x2_ASAP7_75t_R _1259_ (.A1(_0374_),
    .A2(net203),
    .B(_0387_),
    .Y(_0388_));
 AO221x1_ASAP7_75t_R _1260_ (.A1(net126),
    .A2(_0376_),
    .B1(_0377_),
    .B2(net89),
    .C(_0365_),
    .Y(_0389_));
 AND2x2_ASAP7_75t_R _1261_ (.A(net14),
    .B(_0388_),
    .Y(_0390_));
 AO22x1_ASAP7_75t_R _1262_ (.A1(_0388_),
    .A2(_0389_),
    .B1(_0390_),
    .B2(_0380_),
    .Y(_0206_));
 OA21x2_ASAP7_75t_R _1263_ (.A1(_0374_),
    .A2(net204),
    .B(_0387_),
    .Y(_0391_));
 AO221x1_ASAP7_75t_R _1264_ (.A1(net127),
    .A2(_0376_),
    .B1(_0377_),
    .B2(net90),
    .C(_0365_),
    .Y(_0392_));
 AND2x2_ASAP7_75t_R _1265_ (.A(net15),
    .B(_0391_),
    .Y(_0393_));
 AO22x1_ASAP7_75t_R _1266_ (.A1(_0391_),
    .A2(_0392_),
    .B1(_0393_),
    .B2(_0380_),
    .Y(_0207_));
 OA21x2_ASAP7_75t_R _1267_ (.A1(_0374_),
    .A2(net205),
    .B(_0387_),
    .Y(_0394_));
 AO221x1_ASAP7_75t_R _1268_ (.A1(net128),
    .A2(_0376_),
    .B1(_0377_),
    .B2(net91),
    .C(_0365_),
    .Y(_0395_));
 AND2x2_ASAP7_75t_R _1269_ (.A(net16),
    .B(_0394_),
    .Y(_0396_));
 AO22x1_ASAP7_75t_R _1270_ (.A1(_0394_),
    .A2(_0395_),
    .B1(_0396_),
    .B2(_0380_),
    .Y(_0208_));
 OA21x2_ASAP7_75t_R _1271_ (.A1(_0374_),
    .A2(net206),
    .B(_0387_),
    .Y(_0397_));
 AO221x1_ASAP7_75t_R _1272_ (.A1(net129),
    .A2(_0376_),
    .B1(_0377_),
    .B2(net92),
    .C(_0365_),
    .Y(_0398_));
 AND2x2_ASAP7_75t_R _1273_ (.A(net17),
    .B(_0397_),
    .Y(_0399_));
 AO22x1_ASAP7_75t_R _1274_ (.A1(_0397_),
    .A2(_0398_),
    .B1(_0399_),
    .B2(_0380_),
    .Y(_0209_));
 OA21x2_ASAP7_75t_R _1275_ (.A1(_0374_),
    .A2(net207),
    .B(_0387_),
    .Y(_0400_));
 BUFx6f_ASAP7_75t_R _1276_ (.A(_0364_),
    .Y(_0401_));
 AO221x1_ASAP7_75t_R _1277_ (.A1(net130),
    .A2(_0376_),
    .B1(_0377_),
    .B2(net93),
    .C(_0401_),
    .Y(_0402_));
 AND2x2_ASAP7_75t_R _1278_ (.A(net18),
    .B(_0400_),
    .Y(_0403_));
 AO22x1_ASAP7_75t_R _1279_ (.A1(_0400_),
    .A2(_0402_),
    .B1(_0403_),
    .B2(_0380_),
    .Y(_0210_));
 OA21x2_ASAP7_75t_R _1280_ (.A1(_0374_),
    .A2(net208),
    .B(_0387_),
    .Y(_0404_));
 AO221x1_ASAP7_75t_R _1281_ (.A1(net131),
    .A2(_0376_),
    .B1(_0377_),
    .B2(net94),
    .C(_0401_),
    .Y(_0405_));
 AND2x2_ASAP7_75t_R _1282_ (.A(net19),
    .B(_0404_),
    .Y(_0406_));
 AO22x1_ASAP7_75t_R _1283_ (.A1(_0404_),
    .A2(_0405_),
    .B1(_0406_),
    .B2(_0380_),
    .Y(_0211_));
 OA21x2_ASAP7_75t_R _1284_ (.A1(_0374_),
    .A2(net209),
    .B(_0387_),
    .Y(_0407_));
 AO221x1_ASAP7_75t_R _1285_ (.A1(net132),
    .A2(_0376_),
    .B1(_0377_),
    .B2(net95),
    .C(_0401_),
    .Y(_0408_));
 AND2x2_ASAP7_75t_R _1286_ (.A(net20),
    .B(_0407_),
    .Y(_0409_));
 AO22x1_ASAP7_75t_R _1287_ (.A1(_0407_),
    .A2(_0408_),
    .B1(_0409_),
    .B2(_0380_),
    .Y(_0212_));
 BUFx6f_ASAP7_75t_R _1288_ (.A(_0317_),
    .Y(_0410_));
 OA21x2_ASAP7_75t_R _1289_ (.A1(_0410_),
    .A2(net210),
    .B(_0387_),
    .Y(_0411_));
 BUFx3_ASAP7_75t_R _1290_ (.A(_0322_),
    .Y(_0412_));
 BUFx6f_ASAP7_75t_R _1291_ (.A(_0329_),
    .Y(_0413_));
 AO221x1_ASAP7_75t_R _1292_ (.A1(net133),
    .A2(_0412_),
    .B1(_0413_),
    .B2(net96),
    .C(_0401_),
    .Y(_0414_));
 AND2x2_ASAP7_75t_R _1293_ (.A(net21),
    .B(_0411_),
    .Y(_0415_));
 BUFx3_ASAP7_75t_R _1294_ (.A(_0340_),
    .Y(_0416_));
 AO22x1_ASAP7_75t_R _1295_ (.A1(_0411_),
    .A2(_0414_),
    .B1(_0415_),
    .B2(_0416_),
    .Y(_0213_));
 OA21x2_ASAP7_75t_R _1296_ (.A1(_0410_),
    .A2(net211),
    .B(_0387_),
    .Y(_0417_));
 AO221x1_ASAP7_75t_R _1297_ (.A1(net134),
    .A2(_0412_),
    .B1(_0413_),
    .B2(net97),
    .C(_0401_),
    .Y(_0418_));
 AND2x2_ASAP7_75t_R _1298_ (.A(net22),
    .B(_0417_),
    .Y(_0419_));
 AO22x1_ASAP7_75t_R _1299_ (.A1(_0417_),
    .A2(_0418_),
    .B1(_0419_),
    .B2(_0416_),
    .Y(_0214_));
 OA21x2_ASAP7_75t_R _1300_ (.A1(_0410_),
    .A2(net212),
    .B(_0387_),
    .Y(_0420_));
 AO221x1_ASAP7_75t_R _1301_ (.A1(net135),
    .A2(_0412_),
    .B1(_0413_),
    .B2(net98),
    .C(_0401_),
    .Y(_0421_));
 AND2x2_ASAP7_75t_R _1302_ (.A(net23),
    .B(_0420_),
    .Y(_0422_));
 AO22x1_ASAP7_75t_R _1303_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0422_),
    .B2(_0416_),
    .Y(_0215_));
 BUFx6f_ASAP7_75t_R _1304_ (.A(_0622_),
    .Y(_0423_));
 OA21x2_ASAP7_75t_R _1305_ (.A1(_0410_),
    .A2(net213),
    .B(_0423_),
    .Y(_0424_));
 AO221x1_ASAP7_75t_R _1306_ (.A1(net136),
    .A2(_0412_),
    .B1(_0413_),
    .B2(net99),
    .C(_0401_),
    .Y(_0425_));
 AND2x2_ASAP7_75t_R _1307_ (.A(net24),
    .B(_0424_),
    .Y(_0426_));
 AO22x1_ASAP7_75t_R _1308_ (.A1(_0424_),
    .A2(_0425_),
    .B1(_0426_),
    .B2(_0416_),
    .Y(_0216_));
 OA21x2_ASAP7_75t_R _1309_ (.A1(_0410_),
    .A2(net214),
    .B(_0423_),
    .Y(_0427_));
 AO221x1_ASAP7_75t_R _1310_ (.A1(net137),
    .A2(_0412_),
    .B1(_0413_),
    .B2(net100),
    .C(_0401_),
    .Y(_0428_));
 AND2x2_ASAP7_75t_R _1311_ (.A(net25),
    .B(_0427_),
    .Y(_0429_));
 AO22x1_ASAP7_75t_R _1312_ (.A1(_0427_),
    .A2(_0428_),
    .B1(_0429_),
    .B2(_0416_),
    .Y(_0217_));
 OR3x2_ASAP7_75t_R _1313_ (.A(_0336_),
    .B(_0337_),
    .C(_0339_),
    .Y(_0430_));
 NOR2x1_ASAP7_75t_R _1314_ (.A(net26),
    .B(_0331_),
    .Y(_0431_));
 AOI221x1_ASAP7_75t_R _1315_ (.A1(_0331_),
    .A2(_0089_),
    .B1(_0430_),
    .B2(_0431_),
    .C(_0631_),
    .Y(_0218_));
 OA21x2_ASAP7_75t_R _1316_ (.A1(_0410_),
    .A2(net216),
    .B(_0423_),
    .Y(_0432_));
 AO221x1_ASAP7_75t_R _1317_ (.A1(net139),
    .A2(_0412_),
    .B1(_0413_),
    .B2(net102),
    .C(_0401_),
    .Y(_0433_));
 AND2x2_ASAP7_75t_R _1318_ (.A(net27),
    .B(_0432_),
    .Y(_0434_));
 AO22x1_ASAP7_75t_R _1319_ (.A1(_0432_),
    .A2(_0433_),
    .B1(_0434_),
    .B2(_0430_),
    .Y(_0219_));
 OA21x2_ASAP7_75t_R _1320_ (.A1(_0410_),
    .A2(net217),
    .B(_0423_),
    .Y(_0435_));
 AO221x1_ASAP7_75t_R _1321_ (.A1(net140),
    .A2(_0412_),
    .B1(_0413_),
    .B2(net103),
    .C(_0401_),
    .Y(_0436_));
 AND2x2_ASAP7_75t_R _1322_ (.A(net28),
    .B(_0435_),
    .Y(_0437_));
 AO22x1_ASAP7_75t_R _1323_ (.A1(_0435_),
    .A2(_0436_),
    .B1(_0437_),
    .B2(_0430_),
    .Y(_0220_));
 OA21x2_ASAP7_75t_R _1324_ (.A1(_0410_),
    .A2(net218),
    .B(_0423_),
    .Y(_0438_));
 AO221x1_ASAP7_75t_R _1325_ (.A1(net141),
    .A2(_0412_),
    .B1(_0413_),
    .B2(net104),
    .C(_0364_),
    .Y(_0439_));
 AND2x2_ASAP7_75t_R _1326_ (.A(net29),
    .B(_0438_),
    .Y(_0440_));
 AO22x1_ASAP7_75t_R _1327_ (.A1(_0438_),
    .A2(_0439_),
    .B1(_0440_),
    .B2(_0416_),
    .Y(_0221_));
 OA21x2_ASAP7_75t_R _1328_ (.A1(_0410_),
    .A2(net219),
    .B(_0423_),
    .Y(_0441_));
 AO221x1_ASAP7_75t_R _1329_ (.A1(net142),
    .A2(_0412_),
    .B1(_0413_),
    .B2(net105),
    .C(_0364_),
    .Y(_0442_));
 AND2x2_ASAP7_75t_R _1330_ (.A(net30),
    .B(_0441_),
    .Y(_0443_));
 AO22x1_ASAP7_75t_R _1331_ (.A1(_0441_),
    .A2(_0442_),
    .B1(_0443_),
    .B2(_0416_),
    .Y(_0222_));
 OA21x2_ASAP7_75t_R _1332_ (.A1(_0410_),
    .A2(net220),
    .B(_0423_),
    .Y(_0444_));
 AO221x1_ASAP7_75t_R _1333_ (.A1(net143),
    .A2(_0412_),
    .B1(_0413_),
    .B2(net106),
    .C(_0364_),
    .Y(_0445_));
 AND2x2_ASAP7_75t_R _1334_ (.A(net31),
    .B(_0444_),
    .Y(_0446_));
 AO22x1_ASAP7_75t_R _1335_ (.A1(_0444_),
    .A2(_0445_),
    .B1(_0446_),
    .B2(_0416_),
    .Y(_0223_));
 OA21x2_ASAP7_75t_R _1336_ (.A1(_0317_),
    .A2(net221),
    .B(_0423_),
    .Y(_0447_));
 AO221x1_ASAP7_75t_R _1337_ (.A1(net144),
    .A2(_0322_),
    .B1(_0329_),
    .B2(net107),
    .C(_0364_),
    .Y(_0448_));
 AND2x2_ASAP7_75t_R _1338_ (.A(net32),
    .B(_0447_),
    .Y(_0449_));
 AO22x1_ASAP7_75t_R _1339_ (.A1(_0447_),
    .A2(_0448_),
    .B1(_0449_),
    .B2(_0416_),
    .Y(_0224_));
 OA21x2_ASAP7_75t_R _1340_ (.A1(_0317_),
    .A2(net222),
    .B(_0423_),
    .Y(_0450_));
 AO221x1_ASAP7_75t_R _1341_ (.A1(net145),
    .A2(_0322_),
    .B1(_0329_),
    .B2(net108),
    .C(_0364_),
    .Y(_0451_));
 AND2x2_ASAP7_75t_R _1342_ (.A(net33),
    .B(_0450_),
    .Y(_0452_));
 AO22x1_ASAP7_75t_R _1343_ (.A1(_0450_),
    .A2(_0451_),
    .B1(_0452_),
    .B2(_0416_),
    .Y(_0225_));
 OA21x2_ASAP7_75t_R _1344_ (.A1(_0317_),
    .A2(net223),
    .B(_0423_),
    .Y(_0453_));
 AO221x1_ASAP7_75t_R _1345_ (.A1(net146),
    .A2(_0322_),
    .B1(_0329_),
    .B2(net109),
    .C(_0364_),
    .Y(_0454_));
 AND2x2_ASAP7_75t_R _1346_ (.A(net34),
    .B(_0453_),
    .Y(_0455_));
 AO22x1_ASAP7_75t_R _1347_ (.A1(_0453_),
    .A2(_0454_),
    .B1(_0455_),
    .B2(_0340_),
    .Y(_0226_));
 OA21x2_ASAP7_75t_R _1348_ (.A1(_0317_),
    .A2(net224),
    .B(_0622_),
    .Y(_0456_));
 AO221x1_ASAP7_75t_R _1349_ (.A1(net147),
    .A2(_0322_),
    .B1(_0329_),
    .B2(net110),
    .C(_0364_),
    .Y(_0457_));
 AND2x2_ASAP7_75t_R _1350_ (.A(net35),
    .B(_0456_),
    .Y(_0458_));
 AO22x1_ASAP7_75t_R _1351_ (.A1(_0456_),
    .A2(_0457_),
    .B1(_0458_),
    .B2(_0340_),
    .Y(_0227_));
 OA21x2_ASAP7_75t_R _1352_ (.A1(_0317_),
    .A2(net225),
    .B(_0622_),
    .Y(_0459_));
 AO221x1_ASAP7_75t_R _1353_ (.A1(net148),
    .A2(_0322_),
    .B1(_0329_),
    .B2(net111),
    .C(_0364_),
    .Y(_0460_));
 AND2x2_ASAP7_75t_R _1354_ (.A(net36),
    .B(_0459_),
    .Y(_0461_));
 AO22x1_ASAP7_75t_R _1355_ (.A1(_0459_),
    .A2(_0460_),
    .B1(_0461_),
    .B2(_0340_),
    .Y(_0228_));
 AOI22x1_ASAP7_75t_R _1356_ (.A1(_0597_),
    .A2(_0599_),
    .B1(_0593_),
    .B2(_0595_),
    .Y(_0462_));
 AO21x1_ASAP7_75t_R _1357_ (.A1(_0610_),
    .A2(_0613_),
    .B(_0597_),
    .Y(_0463_));
 OA211x2_ASAP7_75t_R _1358_ (.A1(_0600_),
    .A2(_0462_),
    .B(_0463_),
    .C(_0343_),
    .Y(_0464_));
 AO21x1_ASAP7_75t_R _1359_ (.A1(_0331_),
    .A2(_0078_),
    .B(_0464_),
    .Y(_0465_));
 AOI21x1_ASAP7_75t_R _1360_ (.A1(_0321_),
    .A2(_0465_),
    .B(_0631_),
    .Y(_0229_));
 INVx4_ASAP7_75t_R _1361_ (.A(net112),
    .Y(_0466_));
 BUFx6f_ASAP7_75t_R _1362_ (.A(_0466_),
    .Y(_0467_));
 BUFx6f_ASAP7_75t_R _1363_ (.A(net112),
    .Y(_0468_));
 BUFx6f_ASAP7_75t_R _1364_ (.A(_0468_),
    .Y(_0469_));
 OR2x2_ASAP7_75t_R _1365_ (.A(_0469_),
    .B(net1),
    .Y(_0470_));
 OA211x2_ASAP7_75t_R _1366_ (.A1(_0467_),
    .A2(net228),
    .B(_0470_),
    .C(_0624_),
    .Y(_0230_));
 OR2x2_ASAP7_75t_R _1367_ (.A(_0469_),
    .B(net2),
    .Y(_0471_));
 OA211x2_ASAP7_75t_R _1368_ (.A1(_0467_),
    .A2(net229),
    .B(_0471_),
    .C(_0624_),
    .Y(_0231_));
 OR2x2_ASAP7_75t_R _1369_ (.A(_0469_),
    .B(net3),
    .Y(_0472_));
 OA211x2_ASAP7_75t_R _1370_ (.A1(_0467_),
    .A2(net230),
    .B(_0472_),
    .C(_0624_),
    .Y(_0232_));
 OR2x2_ASAP7_75t_R _1371_ (.A(_0469_),
    .B(net4),
    .Y(_0473_));
 OA211x2_ASAP7_75t_R _1372_ (.A1(_0467_),
    .A2(net231),
    .B(_0473_),
    .C(_0624_),
    .Y(_0233_));
 OR2x2_ASAP7_75t_R _1373_ (.A(_0469_),
    .B(net5),
    .Y(_0474_));
 BUFx3_ASAP7_75t_R _1374_ (.A(_0623_),
    .Y(_0475_));
 OA211x2_ASAP7_75t_R _1375_ (.A1(_0467_),
    .A2(net232),
    .B(_0474_),
    .C(_0475_),
    .Y(_0234_));
 OR2x2_ASAP7_75t_R _1376_ (.A(_0469_),
    .B(net6),
    .Y(_0476_));
 OA211x2_ASAP7_75t_R _1377_ (.A1(_0467_),
    .A2(net233),
    .B(_0476_),
    .C(_0475_),
    .Y(_0235_));
 BUFx6f_ASAP7_75t_R _1378_ (.A(_0468_),
    .Y(_0477_));
 OR2x2_ASAP7_75t_R _1379_ (.A(_0477_),
    .B(net7),
    .Y(_0478_));
 OA211x2_ASAP7_75t_R _1380_ (.A1(_0467_),
    .A2(net234),
    .B(_0478_),
    .C(_0475_),
    .Y(_0236_));
 OR2x2_ASAP7_75t_R _1381_ (.A(_0477_),
    .B(net8),
    .Y(_0479_));
 OA211x2_ASAP7_75t_R _1382_ (.A1(_0467_),
    .A2(net235),
    .B(_0479_),
    .C(_0475_),
    .Y(_0237_));
 OR2x2_ASAP7_75t_R _1383_ (.A(_0477_),
    .B(net9),
    .Y(_0480_));
 OA211x2_ASAP7_75t_R _1384_ (.A1(_0467_),
    .A2(net236),
    .B(_0480_),
    .C(_0475_),
    .Y(_0238_));
 OR2x2_ASAP7_75t_R _1385_ (.A(_0477_),
    .B(net10),
    .Y(_0481_));
 OA211x2_ASAP7_75t_R _1386_ (.A1(_0467_),
    .A2(net237),
    .B(_0481_),
    .C(_0475_),
    .Y(_0239_));
 BUFx6f_ASAP7_75t_R _1387_ (.A(_0466_),
    .Y(_0482_));
 OR2x2_ASAP7_75t_R _1388_ (.A(_0477_),
    .B(net11),
    .Y(_0483_));
 OA211x2_ASAP7_75t_R _1389_ (.A1(_0482_),
    .A2(net238),
    .B(_0483_),
    .C(_0475_),
    .Y(_0240_));
 OR2x2_ASAP7_75t_R _1390_ (.A(_0477_),
    .B(net12),
    .Y(_0484_));
 OA211x2_ASAP7_75t_R _1391_ (.A1(_0482_),
    .A2(net239),
    .B(_0484_),
    .C(_0475_),
    .Y(_0241_));
 OR2x2_ASAP7_75t_R _1392_ (.A(_0477_),
    .B(net13),
    .Y(_0485_));
 OA211x2_ASAP7_75t_R _1393_ (.A1(_0482_),
    .A2(net240),
    .B(_0485_),
    .C(_0475_),
    .Y(_0242_));
 OR2x2_ASAP7_75t_R _1394_ (.A(_0477_),
    .B(net14),
    .Y(_0486_));
 OA211x2_ASAP7_75t_R _1395_ (.A1(_0482_),
    .A2(net241),
    .B(_0486_),
    .C(_0475_),
    .Y(_0243_));
 OR2x2_ASAP7_75t_R _1396_ (.A(_0477_),
    .B(net15),
    .Y(_0487_));
 BUFx3_ASAP7_75t_R _1397_ (.A(_0623_),
    .Y(_0488_));
 OA211x2_ASAP7_75t_R _1398_ (.A1(_0482_),
    .A2(net242),
    .B(_0487_),
    .C(_0488_),
    .Y(_0244_));
 OR2x2_ASAP7_75t_R _1399_ (.A(_0477_),
    .B(net16),
    .Y(_0489_));
 OA211x2_ASAP7_75t_R _1400_ (.A1(_0482_),
    .A2(net243),
    .B(_0489_),
    .C(_0488_),
    .Y(_0245_));
 BUFx6f_ASAP7_75t_R _1401_ (.A(_0468_),
    .Y(_0490_));
 OR2x2_ASAP7_75t_R _1402_ (.A(_0490_),
    .B(net17),
    .Y(_0491_));
 OA211x2_ASAP7_75t_R _1403_ (.A1(_0482_),
    .A2(net244),
    .B(_0491_),
    .C(_0488_),
    .Y(_0246_));
 OR2x2_ASAP7_75t_R _1404_ (.A(_0490_),
    .B(net18),
    .Y(_0492_));
 OA211x2_ASAP7_75t_R _1405_ (.A1(_0482_),
    .A2(net245),
    .B(_0492_),
    .C(_0488_),
    .Y(_0247_));
 OR2x2_ASAP7_75t_R _1406_ (.A(_0490_),
    .B(net19),
    .Y(_0493_));
 OA211x2_ASAP7_75t_R _1407_ (.A1(_0482_),
    .A2(net246),
    .B(_0493_),
    .C(_0488_),
    .Y(_0248_));
 OR2x2_ASAP7_75t_R _1408_ (.A(_0490_),
    .B(net20),
    .Y(_0494_));
 OA211x2_ASAP7_75t_R _1409_ (.A1(_0482_),
    .A2(net247),
    .B(_0494_),
    .C(_0488_),
    .Y(_0249_));
 BUFx6f_ASAP7_75t_R _1410_ (.A(_0466_),
    .Y(_0495_));
 OR2x2_ASAP7_75t_R _1411_ (.A(_0490_),
    .B(net21),
    .Y(_0496_));
 OA211x2_ASAP7_75t_R _1412_ (.A1(_0495_),
    .A2(net248),
    .B(_0496_),
    .C(_0488_),
    .Y(_0250_));
 OR2x2_ASAP7_75t_R _1413_ (.A(_0490_),
    .B(net22),
    .Y(_0497_));
 OA211x2_ASAP7_75t_R _1414_ (.A1(_0495_),
    .A2(net249),
    .B(_0497_),
    .C(_0488_),
    .Y(_0251_));
 OR2x2_ASAP7_75t_R _1415_ (.A(_0490_),
    .B(net23),
    .Y(_0498_));
 OA211x2_ASAP7_75t_R _1416_ (.A1(_0495_),
    .A2(net250),
    .B(_0498_),
    .C(_0488_),
    .Y(_0252_));
 OR2x2_ASAP7_75t_R _1417_ (.A(_0490_),
    .B(net24),
    .Y(_0499_));
 OA211x2_ASAP7_75t_R _1418_ (.A1(_0495_),
    .A2(net251),
    .B(_0499_),
    .C(_0488_),
    .Y(_0253_));
 OR2x2_ASAP7_75t_R _1419_ (.A(_0490_),
    .B(net25),
    .Y(_0500_));
 BUFx3_ASAP7_75t_R _1420_ (.A(_0623_),
    .Y(_0501_));
 OA211x2_ASAP7_75t_R _1421_ (.A1(_0495_),
    .A2(net252),
    .B(_0500_),
    .C(_0501_),
    .Y(_0254_));
 OR2x2_ASAP7_75t_R _1422_ (.A(net26),
    .B(_0469_),
    .Y(_0502_));
 OA211x2_ASAP7_75t_R _1423_ (.A1(_0495_),
    .A2(net253),
    .B(_0502_),
    .C(_0501_),
    .Y(_0255_));
 OR2x2_ASAP7_75t_R _1424_ (.A(net27),
    .B(_0469_),
    .Y(_0503_));
 OA211x2_ASAP7_75t_R _1425_ (.A1(_0495_),
    .A2(net254),
    .B(_0503_),
    .C(_0501_),
    .Y(_0256_));
 OR2x2_ASAP7_75t_R _1426_ (.A(net28),
    .B(_0469_),
    .Y(_0504_));
 OA211x2_ASAP7_75t_R _1427_ (.A1(_0495_),
    .A2(net255),
    .B(_0504_),
    .C(_0501_),
    .Y(_0257_));
 OR2x2_ASAP7_75t_R _1428_ (.A(_0490_),
    .B(net29),
    .Y(_0505_));
 OA211x2_ASAP7_75t_R _1429_ (.A1(_0495_),
    .A2(net256),
    .B(_0505_),
    .C(_0501_),
    .Y(_0258_));
 OR2x2_ASAP7_75t_R _1430_ (.A(_0468_),
    .B(net30),
    .Y(_0506_));
 OA211x2_ASAP7_75t_R _1431_ (.A1(_0495_),
    .A2(net257),
    .B(_0506_),
    .C(_0501_),
    .Y(_0259_));
 OR2x2_ASAP7_75t_R _1432_ (.A(_0468_),
    .B(net31),
    .Y(_0507_));
 OA211x2_ASAP7_75t_R _1433_ (.A1(_0466_),
    .A2(net258),
    .B(_0507_),
    .C(_0501_),
    .Y(_0260_));
 OR2x2_ASAP7_75t_R _1434_ (.A(_0468_),
    .B(net32),
    .Y(_0508_));
 OA211x2_ASAP7_75t_R _1435_ (.A1(_0466_),
    .A2(net259),
    .B(_0508_),
    .C(_0501_),
    .Y(_0261_));
 OR2x2_ASAP7_75t_R _1436_ (.A(_0468_),
    .B(net33),
    .Y(_0509_));
 OA211x2_ASAP7_75t_R _1437_ (.A1(_0466_),
    .A2(net260),
    .B(_0509_),
    .C(_0501_),
    .Y(_0262_));
 OR2x2_ASAP7_75t_R _1438_ (.A(_0468_),
    .B(net34),
    .Y(_0510_));
 OA211x2_ASAP7_75t_R _1439_ (.A1(_0466_),
    .A2(net261),
    .B(_0510_),
    .C(_0501_),
    .Y(_0263_));
 OR2x2_ASAP7_75t_R _1440_ (.A(_0468_),
    .B(net35),
    .Y(_0511_));
 BUFx6f_ASAP7_75t_R _1441_ (.A(_0623_),
    .Y(_0512_));
 OA211x2_ASAP7_75t_R _1442_ (.A1(_0466_),
    .A2(net262),
    .B(_0511_),
    .C(_0512_),
    .Y(_0264_));
 OR2x2_ASAP7_75t_R _1443_ (.A(_0468_),
    .B(net36),
    .Y(_0513_));
 OA211x2_ASAP7_75t_R _1444_ (.A1(_0466_),
    .A2(net263),
    .B(_0513_),
    .C(_0512_),
    .Y(_0265_));
 AND3x1_ASAP7_75t_R _1445_ (.A(net37),
    .B(_0466_),
    .C(_0588_),
    .Y(_0514_));
 AO21x1_ASAP7_75t_R _1446_ (.A1(_0469_),
    .A2(net264),
    .B(_0514_),
    .Y(_0515_));
 AND2x2_ASAP7_75t_R _1447_ (.A(_0624_),
    .B(_0515_),
    .Y(_0266_));
 BUFx12f_ASAP7_75t_R _1448_ (.A(net150),
    .Y(_0516_));
 BUFx6f_ASAP7_75t_R _1449_ (.A(_0516_),
    .Y(_0517_));
 BUFx6f_ASAP7_75t_R _1450_ (.A(net150),
    .Y(_0518_));
 NAND2x1_ASAP7_75t_R _1451_ (.A(_0518_),
    .B(_0040_),
    .Y(_0519_));
 OA211x2_ASAP7_75t_R _1452_ (.A1(_0517_),
    .A2(net38),
    .B(_0519_),
    .C(_0512_),
    .Y(_0267_));
 NAND2x1_ASAP7_75t_R _1453_ (.A(_0518_),
    .B(_0039_),
    .Y(_0520_));
 OA211x2_ASAP7_75t_R _1454_ (.A1(_0517_),
    .A2(net39),
    .B(_0520_),
    .C(_0512_),
    .Y(_0268_));
 BUFx12f_ASAP7_75t_R _1455_ (.A(_0516_),
    .Y(_0521_));
 NAND2x1_ASAP7_75t_R _1456_ (.A(_0521_),
    .B(_0038_),
    .Y(_0522_));
 OA211x2_ASAP7_75t_R _1457_ (.A1(_0517_),
    .A2(net40),
    .B(_0522_),
    .C(_0512_),
    .Y(_0269_));
 NAND2x1_ASAP7_75t_R _1458_ (.A(_0521_),
    .B(_0037_),
    .Y(_0523_));
 OA211x2_ASAP7_75t_R _1459_ (.A1(_0517_),
    .A2(net41),
    .B(_0523_),
    .C(_0512_),
    .Y(_0270_));
 NAND2x1_ASAP7_75t_R _1460_ (.A(_0521_),
    .B(_0036_),
    .Y(_0524_));
 OA211x2_ASAP7_75t_R _1461_ (.A1(_0517_),
    .A2(net42),
    .B(_0524_),
    .C(_0512_),
    .Y(_0271_));
 NAND2x1_ASAP7_75t_R _1462_ (.A(_0521_),
    .B(_0035_),
    .Y(_0525_));
 OA211x2_ASAP7_75t_R _1463_ (.A1(_0517_),
    .A2(net43),
    .B(_0525_),
    .C(_0512_),
    .Y(_0272_));
 NAND2x1_ASAP7_75t_R _1464_ (.A(_0521_),
    .B(_0034_),
    .Y(_0526_));
 OA211x2_ASAP7_75t_R _1465_ (.A1(_0517_),
    .A2(net44),
    .B(_0526_),
    .C(_0512_),
    .Y(_0273_));
 NAND2x1_ASAP7_75t_R _1466_ (.A(_0521_),
    .B(_0033_),
    .Y(_0527_));
 OA211x2_ASAP7_75t_R _1467_ (.A1(_0517_),
    .A2(net45),
    .B(_0527_),
    .C(_0512_),
    .Y(_0274_));
 NAND2x1_ASAP7_75t_R _1468_ (.A(_0521_),
    .B(_0032_),
    .Y(_0528_));
 BUFx3_ASAP7_75t_R _1469_ (.A(_0623_),
    .Y(_0529_));
 OA211x2_ASAP7_75t_R _1470_ (.A1(_0517_),
    .A2(net46),
    .B(_0528_),
    .C(_0529_),
    .Y(_0275_));
 NAND2x1_ASAP7_75t_R _1471_ (.A(_0521_),
    .B(_0031_),
    .Y(_0530_));
 OA211x2_ASAP7_75t_R _1472_ (.A1(_0517_),
    .A2(net47),
    .B(_0530_),
    .C(_0529_),
    .Y(_0276_));
 BUFx6f_ASAP7_75t_R _1473_ (.A(_0516_),
    .Y(_0531_));
 NAND2x1_ASAP7_75t_R _1474_ (.A(_0521_),
    .B(_0030_),
    .Y(_0532_));
 OA211x2_ASAP7_75t_R _1475_ (.A1(_0531_),
    .A2(net48),
    .B(_0532_),
    .C(_0529_),
    .Y(_0277_));
 NAND2x1_ASAP7_75t_R _1476_ (.A(_0521_),
    .B(_0029_),
    .Y(_0533_));
 OA211x2_ASAP7_75t_R _1477_ (.A1(_0531_),
    .A2(net49),
    .B(_0533_),
    .C(_0529_),
    .Y(_0278_));
 BUFx12f_ASAP7_75t_R _1478_ (.A(_0516_),
    .Y(_0534_));
 NAND2x1_ASAP7_75t_R _1479_ (.A(_0534_),
    .B(_0028_),
    .Y(_0535_));
 OA211x2_ASAP7_75t_R _1480_ (.A1(_0531_),
    .A2(net50),
    .B(_0535_),
    .C(_0529_),
    .Y(_0279_));
 NAND2x1_ASAP7_75t_R _1481_ (.A(_0534_),
    .B(_0027_),
    .Y(_0536_));
 OA211x2_ASAP7_75t_R _1482_ (.A1(_0531_),
    .A2(net51),
    .B(_0536_),
    .C(_0529_),
    .Y(_0280_));
 NAND2x1_ASAP7_75t_R _1483_ (.A(_0534_),
    .B(_0026_),
    .Y(_0537_));
 OA211x2_ASAP7_75t_R _1484_ (.A1(_0531_),
    .A2(net52),
    .B(_0537_),
    .C(_0529_),
    .Y(_0281_));
 NAND2x1_ASAP7_75t_R _1485_ (.A(_0534_),
    .B(_0025_),
    .Y(_0538_));
 OA211x2_ASAP7_75t_R _1486_ (.A1(_0531_),
    .A2(net53),
    .B(_0538_),
    .C(_0529_),
    .Y(_0282_));
 NAND2x1_ASAP7_75t_R _1487_ (.A(_0534_),
    .B(_0024_),
    .Y(_0539_));
 OA211x2_ASAP7_75t_R _1488_ (.A1(_0531_),
    .A2(net54),
    .B(_0539_),
    .C(_0529_),
    .Y(_0283_));
 NAND2x1_ASAP7_75t_R _1489_ (.A(_0534_),
    .B(_0023_),
    .Y(_0540_));
 OA211x2_ASAP7_75t_R _1490_ (.A1(_0531_),
    .A2(net55),
    .B(_0540_),
    .C(_0529_),
    .Y(_0284_));
 NAND2x1_ASAP7_75t_R _1491_ (.A(_0534_),
    .B(_0022_),
    .Y(_0541_));
 BUFx6f_ASAP7_75t_R _1492_ (.A(_0623_),
    .Y(_0542_));
 OA211x2_ASAP7_75t_R _1493_ (.A1(_0531_),
    .A2(net56),
    .B(_0541_),
    .C(_0542_),
    .Y(_0285_));
 NAND2x1_ASAP7_75t_R _1494_ (.A(_0534_),
    .B(_0021_),
    .Y(_0543_));
 OA211x2_ASAP7_75t_R _1495_ (.A1(_0531_),
    .A2(net57),
    .B(_0543_),
    .C(_0542_),
    .Y(_0286_));
 BUFx6f_ASAP7_75t_R _1496_ (.A(_0516_),
    .Y(_0544_));
 NAND2x1_ASAP7_75t_R _1497_ (.A(_0534_),
    .B(_0020_),
    .Y(_0545_));
 OA211x2_ASAP7_75t_R _1498_ (.A1(_0544_),
    .A2(net58),
    .B(_0545_),
    .C(_0542_),
    .Y(_0287_));
 NAND2x1_ASAP7_75t_R _1499_ (.A(_0534_),
    .B(_0019_),
    .Y(_0546_));
 OA211x2_ASAP7_75t_R _1500_ (.A1(_0544_),
    .A2(net59),
    .B(_0546_),
    .C(_0542_),
    .Y(_0288_));
 BUFx6f_ASAP7_75t_R _1501_ (.A(_0516_),
    .Y(_0547_));
 NAND2x1_ASAP7_75t_R _1502_ (.A(_0547_),
    .B(_0018_),
    .Y(_0548_));
 OA211x2_ASAP7_75t_R _1503_ (.A1(_0544_),
    .A2(net60),
    .B(_0548_),
    .C(_0542_),
    .Y(_0289_));
 NAND2x1_ASAP7_75t_R _1504_ (.A(_0547_),
    .B(_0017_),
    .Y(_0549_));
 OA211x2_ASAP7_75t_R _1505_ (.A1(_0544_),
    .A2(net61),
    .B(_0549_),
    .C(_0542_),
    .Y(_0290_));
 NAND2x1_ASAP7_75t_R _1506_ (.A(_0547_),
    .B(_0016_),
    .Y(_0550_));
 OA211x2_ASAP7_75t_R _1507_ (.A1(_0544_),
    .A2(net62),
    .B(_0550_),
    .C(_0542_),
    .Y(_0291_));
 NAND2x1_ASAP7_75t_R _1508_ (.A(_0516_),
    .B(_0015_),
    .Y(_0551_));
 OA211x2_ASAP7_75t_R _1509_ (.A1(net63),
    .A2(_0518_),
    .B(_0624_),
    .C(_0551_),
    .Y(_0292_));
 NAND2x1_ASAP7_75t_R _1510_ (.A(_0516_),
    .B(_0014_),
    .Y(_0552_));
 OA211x2_ASAP7_75t_R _1511_ (.A1(net64),
    .A2(_0518_),
    .B(_0624_),
    .C(_0552_),
    .Y(_0293_));
 NAND2x1_ASAP7_75t_R _1512_ (.A(_0516_),
    .B(_0013_),
    .Y(_0553_));
 OA211x2_ASAP7_75t_R _1513_ (.A1(net65),
    .A2(_0518_),
    .B(_0624_),
    .C(_0553_),
    .Y(_0294_));
 NAND2x1_ASAP7_75t_R _1514_ (.A(_0547_),
    .B(_0012_),
    .Y(_0554_));
 OA211x2_ASAP7_75t_R _1515_ (.A1(_0544_),
    .A2(net66),
    .B(_0554_),
    .C(_0542_),
    .Y(_0295_));
 NAND2x1_ASAP7_75t_R _1516_ (.A(_0547_),
    .B(_0011_),
    .Y(_0555_));
 OA211x2_ASAP7_75t_R _1517_ (.A1(_0544_),
    .A2(net67),
    .B(_0555_),
    .C(_0542_),
    .Y(_0296_));
 NAND2x1_ASAP7_75t_R _1518_ (.A(_0547_),
    .B(_0010_),
    .Y(_0556_));
 OA211x2_ASAP7_75t_R _1519_ (.A1(_0544_),
    .A2(net68),
    .B(_0556_),
    .C(_0542_),
    .Y(_0297_));
 NAND2x1_ASAP7_75t_R _1520_ (.A(_0547_),
    .B(_0009_),
    .Y(_0557_));
 OA211x2_ASAP7_75t_R _1521_ (.A1(_0544_),
    .A2(net69),
    .B(_0557_),
    .C(_0626_),
    .Y(_0298_));
 NAND2x1_ASAP7_75t_R _1522_ (.A(_0547_),
    .B(_0008_),
    .Y(_0558_));
 OA211x2_ASAP7_75t_R _1523_ (.A1(_0544_),
    .A2(net70),
    .B(_0558_),
    .C(_0626_),
    .Y(_0299_));
 NAND2x1_ASAP7_75t_R _1524_ (.A(_0547_),
    .B(_0007_),
    .Y(_0559_));
 OA211x2_ASAP7_75t_R _1525_ (.A1(_0518_),
    .A2(net71),
    .B(_0559_),
    .C(_0626_),
    .Y(_0300_));
 NAND2x1_ASAP7_75t_R _1526_ (.A(_0547_),
    .B(_0006_),
    .Y(_0560_));
 OA211x2_ASAP7_75t_R _1527_ (.A1(_0518_),
    .A2(net72),
    .B(_0560_),
    .C(_0626_),
    .Y(_0301_));
 NAND2x1_ASAP7_75t_R _1528_ (.A(_0516_),
    .B(_0005_),
    .Y(_0561_));
 OA211x2_ASAP7_75t_R _1529_ (.A1(_0518_),
    .A2(net73),
    .B(_0561_),
    .C(_0626_),
    .Y(_0302_));
 NAND2x1_ASAP7_75t_R _1530_ (.A(_0518_),
    .B(net302),
    .Y(_0562_));
 OR3x1_ASAP7_75t_R _1531_ (.A(_0591_),
    .B(_0518_),
    .C(_0575_),
    .Y(_0563_));
 AOI21x1_ASAP7_75t_R _1532_ (.A1(_0562_),
    .A2(_0563_),
    .B(_0631_),
    .Y(_0303_));
 BUFx4_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx2_ASAP7_75t_R _1534_ (.A(net303),
    .Y(done));
 DFFHQNx1_ASAP7_75t_R \l_o_r[0]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0156_),
    .QN(_0151_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[10]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0157_),
    .QN(_0150_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[11]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0158_),
    .QN(_0149_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[12]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0159_),
    .QN(_0148_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[13]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0160_),
    .QN(_0147_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[14]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0161_),
    .QN(_0146_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[15]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0162_),
    .QN(_0145_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[16]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0163_),
    .QN(_0144_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[17]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0164_),
    .QN(_0143_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[18]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0165_),
    .QN(_0142_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[19]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0166_),
    .QN(_0141_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[1]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0167_),
    .QN(_0140_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[20]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0168_),
    .QN(_0139_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[21]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0169_),
    .QN(_0138_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[22]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0170_),
    .QN(_0137_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[23]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0171_),
    .QN(_0136_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[24]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0172_),
    .QN(_0135_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[25]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0173_),
    .QN(_0134_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[26]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0174_),
    .QN(_0133_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[27]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0175_),
    .QN(_0132_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[28]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0176_),
    .QN(_0131_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[29]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0177_),
    .QN(_0130_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[2]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0178_),
    .QN(_0129_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[30]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0179_),
    .QN(_0128_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[31]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0180_),
    .QN(_0127_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[32]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0181_),
    .QN(_0126_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[33]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0182_),
    .QN(_0125_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[34]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0183_),
    .QN(_0124_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[35]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0184_),
    .QN(_0123_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[3]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0185_),
    .QN(_0122_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[4]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0186_),
    .QN(_0121_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[5]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0187_),
    .QN(_0120_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[6]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0188_),
    .QN(_0119_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[7]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0189_),
    .QN(_0118_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[8]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0190_),
    .QN(_0117_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[9]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0191_),
    .QN(_0116_));
 DFFHQNx1_ASAP7_75t_R \l_o_v_r$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0192_),
    .QN(_0152_));
 DFFHQNx3_ASAP7_75t_R \r.rr[0]$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .D(_0000_),
    .QN(_0153_));
 DFFHQNx1_ASAP7_75t_R \r.rr[1]$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .D(_0001_),
    .QN(_0154_));
 DFFHQNx3_ASAP7_75t_R \r.rr[2]$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .D(_0002_),
    .QN(_0155_));
 DFFHQNx3_ASAP7_75t_R \r.rr[3]$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .D(_0003_),
    .QN(_0115_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[0]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0193_),
    .QN(_0114_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[10]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0194_),
    .QN(_0113_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[11]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0195_),
    .QN(_0112_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[12]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0196_),
    .QN(_0111_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[13]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0197_),
    .QN(_0110_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[14]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0198_),
    .QN(_0109_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[15]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0199_),
    .QN(_0108_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[16]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0200_),
    .QN(_0107_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[17]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0201_),
    .QN(_0106_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[18]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0202_),
    .QN(_0105_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[19]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0203_),
    .QN(_0104_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[1]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0204_),
    .QN(_0103_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[20]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0205_),
    .QN(_0102_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[21]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0206_),
    .QN(_0101_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[22]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0207_),
    .QN(_0100_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[23]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0208_),
    .QN(_0099_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[24]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0209_),
    .QN(_0098_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[25]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0210_),
    .QN(_0097_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[26]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0211_),
    .QN(_0096_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[27]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0212_),
    .QN(_0095_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[28]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0213_),
    .QN(_0094_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[29]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0214_),
    .QN(_0093_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[2]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0215_),
    .QN(_0092_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[30]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0216_),
    .QN(_0091_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[31]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0217_),
    .QN(_0090_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[32]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0218_),
    .QN(_0089_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[33]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0219_),
    .QN(_0088_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[34]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0220_),
    .QN(_0087_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[35]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0221_),
    .QN(_0086_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[3]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0222_),
    .QN(_0085_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[4]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0223_),
    .QN(_0084_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[5]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0224_),
    .QN(_0083_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[6]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0225_),
    .QN(_0082_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[7]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0226_),
    .QN(_0081_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[8]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0227_),
    .QN(_0080_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[9]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0228_),
    .QN(_0079_));
 DFFHQNx1_ASAP7_75t_R \r_o_v_r$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0229_),
    .QN(_0078_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[0]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0230_),
    .QN(_0077_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[10]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0231_),
    .QN(_0076_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[11]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0232_),
    .QN(_0075_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[12]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0233_),
    .QN(_0074_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[13]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0234_),
    .QN(_0073_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[14]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0235_),
    .QN(_0072_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[15]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0236_),
    .QN(_0071_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[16]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0237_),
    .QN(_0070_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[17]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0238_),
    .QN(_0069_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[18]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0239_),
    .QN(_0068_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[19]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0240_),
    .QN(_0067_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[1]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0241_),
    .QN(_0066_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[20]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0242_),
    .QN(_0065_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[21]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0243_),
    .QN(_0064_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[22]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0244_),
    .QN(_0063_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[23]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0245_),
    .QN(_0062_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[24]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0246_),
    .QN(_0061_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[25]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0247_),
    .QN(_0060_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[26]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0248_),
    .QN(_0059_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[27]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0249_),
    .QN(_0058_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[28]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0250_),
    .QN(_0057_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[29]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0251_),
    .QN(_0056_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[2]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0252_),
    .QN(_0055_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[30]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0253_),
    .QN(_0054_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[31]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0254_),
    .QN(_0053_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[32]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0255_),
    .QN(_0052_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[33]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0256_),
    .QN(_0051_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[34]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0257_),
    .QN(_0050_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[35]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0258_),
    .QN(_0049_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[3]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0259_),
    .QN(_0048_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[4]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0260_),
    .QN(_0047_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[5]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0261_),
    .QN(_0046_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[6]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0262_),
    .QN(_0045_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[7]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0263_),
    .QN(_0044_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[8]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0264_),
    .QN(_0043_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[9]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0265_),
    .QN(_0042_));
 DFFHQNx1_ASAP7_75t_R \u0_o_v_r$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0266_),
    .QN(_0041_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[0]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0267_),
    .QN(_0040_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[10]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0268_),
    .QN(_0039_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[11]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0269_),
    .QN(_0038_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[12]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0270_),
    .QN(_0037_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[13]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0271_),
    .QN(_0036_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[14]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0272_),
    .QN(_0035_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[15]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0273_),
    .QN(_0034_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[16]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0274_),
    .QN(_0033_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[17]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0275_),
    .QN(_0032_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[18]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0276_),
    .QN(_0031_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[19]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0277_),
    .QN(_0030_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[1]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0278_),
    .QN(_0029_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[20]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0279_),
    .QN(_0028_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[21]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0280_),
    .QN(_0027_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[22]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0281_),
    .QN(_0026_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[23]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0282_),
    .QN(_0025_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[24]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0283_),
    .QN(_0024_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[25]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0284_),
    .QN(_0023_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[26]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0285_),
    .QN(_0022_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[27]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0286_),
    .QN(_0021_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[28]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0287_),
    .QN(_0020_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[29]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0288_),
    .QN(_0019_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[2]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0289_),
    .QN(_0018_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[30]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0290_),
    .QN(_0017_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[31]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0291_),
    .QN(_0016_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[32]$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0292_),
    .QN(_0015_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[33]$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0293_),
    .QN(_0014_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[34]$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0294_),
    .QN(_0013_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[35]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0295_),
    .QN(_0012_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[3]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0296_),
    .QN(_0011_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[4]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0297_),
    .QN(_0010_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[5]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0298_),
    .QN(_0009_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[6]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0299_),
    .QN(_0008_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[7]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0300_),
    .QN(_0007_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[8]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0301_),
    .QN(_0006_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[9]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0302_),
    .QN(_0005_));
 DFFHQNx1_ASAP7_75t_R \u1_o_v_r$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0303_),
    .QN(_0004_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Left_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Left_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Left_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Left_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Left_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Left_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Left_123 ();
 BUFx3_ASAP7_75t_R input1 (.A(l_i[0]),
    .Y(net1));
 BUFx3_ASAP7_75t_R input2 (.A(l_i[10]),
    .Y(net2));
 BUFx3_ASAP7_75t_R input3 (.A(l_i[11]),
    .Y(net3));
 BUFx3_ASAP7_75t_R input4 (.A(l_i[12]),
    .Y(net4));
 BUFx3_ASAP7_75t_R input5 (.A(l_i[13]),
    .Y(net5));
 BUFx3_ASAP7_75t_R input6 (.A(l_i[14]),
    .Y(net6));
 BUFx3_ASAP7_75t_R input7 (.A(l_i[15]),
    .Y(net7));
 BUFx3_ASAP7_75t_R input8 (.A(l_i[16]),
    .Y(net8));
 BUFx3_ASAP7_75t_R input9 (.A(l_i[17]),
    .Y(net9));
 BUFx3_ASAP7_75t_R input10 (.A(l_i[18]),
    .Y(net10));
 BUFx3_ASAP7_75t_R input11 (.A(l_i[19]),
    .Y(net11));
 BUFx3_ASAP7_75t_R input12 (.A(l_i[1]),
    .Y(net12));
 BUFx3_ASAP7_75t_R input13 (.A(l_i[20]),
    .Y(net13));
 BUFx3_ASAP7_75t_R input14 (.A(l_i[21]),
    .Y(net14));
 BUFx3_ASAP7_75t_R input15 (.A(l_i[22]),
    .Y(net15));
 BUFx3_ASAP7_75t_R input16 (.A(l_i[23]),
    .Y(net16));
 BUFx3_ASAP7_75t_R input17 (.A(l_i[24]),
    .Y(net17));
 BUFx3_ASAP7_75t_R input18 (.A(l_i[25]),
    .Y(net18));
 BUFx3_ASAP7_75t_R input19 (.A(l_i[26]),
    .Y(net19));
 BUFx3_ASAP7_75t_R input20 (.A(l_i[27]),
    .Y(net20));
 BUFx3_ASAP7_75t_R input21 (.A(l_i[28]),
    .Y(net21));
 BUFx3_ASAP7_75t_R input22 (.A(l_i[29]),
    .Y(net22));
 BUFx3_ASAP7_75t_R input23 (.A(l_i[2]),
    .Y(net23));
 BUFx3_ASAP7_75t_R input24 (.A(l_i[30]),
    .Y(net24));
 BUFx3_ASAP7_75t_R input25 (.A(l_i[31]),
    .Y(net25));
 BUFx3_ASAP7_75t_R input26 (.A(l_i[32]),
    .Y(net26));
 BUFx3_ASAP7_75t_R input27 (.A(l_i[33]),
    .Y(net27));
 BUFx3_ASAP7_75t_R input28 (.A(l_i[34]),
    .Y(net28));
 BUFx3_ASAP7_75t_R input29 (.A(l_i[35]),
    .Y(net29));
 BUFx3_ASAP7_75t_R input30 (.A(l_i[3]),
    .Y(net30));
 BUFx3_ASAP7_75t_R input31 (.A(l_i[4]),
    .Y(net31));
 BUFx3_ASAP7_75t_R input32 (.A(l_i[5]),
    .Y(net32));
 BUFx3_ASAP7_75t_R input33 (.A(l_i[6]),
    .Y(net33));
 BUFx3_ASAP7_75t_R input34 (.A(l_i[7]),
    .Y(net34));
 BUFx3_ASAP7_75t_R input35 (.A(l_i[8]),
    .Y(net35));
 BUFx3_ASAP7_75t_R input36 (.A(l_i[9]),
    .Y(net36));
 BUFx3_ASAP7_75t_R input37 (.A(l_i_v),
    .Y(net37));
 BUFx3_ASAP7_75t_R input38 (.A(r_i[0]),
    .Y(net38));
 BUFx3_ASAP7_75t_R input39 (.A(r_i[10]),
    .Y(net39));
 BUFx3_ASAP7_75t_R input40 (.A(r_i[11]),
    .Y(net40));
 BUFx3_ASAP7_75t_R input41 (.A(r_i[12]),
    .Y(net41));
 BUFx3_ASAP7_75t_R input42 (.A(r_i[13]),
    .Y(net42));
 BUFx3_ASAP7_75t_R input43 (.A(r_i[14]),
    .Y(net43));
 BUFx3_ASAP7_75t_R input44 (.A(r_i[15]),
    .Y(net44));
 BUFx3_ASAP7_75t_R input45 (.A(r_i[16]),
    .Y(net45));
 BUFx3_ASAP7_75t_R input46 (.A(r_i[17]),
    .Y(net46));
 BUFx3_ASAP7_75t_R input47 (.A(r_i[18]),
    .Y(net47));
 BUFx3_ASAP7_75t_R input48 (.A(r_i[19]),
    .Y(net48));
 BUFx3_ASAP7_75t_R input49 (.A(r_i[1]),
    .Y(net49));
 BUFx3_ASAP7_75t_R input50 (.A(r_i[20]),
    .Y(net50));
 BUFx3_ASAP7_75t_R input51 (.A(r_i[21]),
    .Y(net51));
 BUFx3_ASAP7_75t_R input52 (.A(r_i[22]),
    .Y(net52));
 BUFx3_ASAP7_75t_R input53 (.A(r_i[23]),
    .Y(net53));
 BUFx3_ASAP7_75t_R input54 (.A(r_i[24]),
    .Y(net54));
 BUFx3_ASAP7_75t_R input55 (.A(r_i[25]),
    .Y(net55));
 BUFx3_ASAP7_75t_R input56 (.A(r_i[26]),
    .Y(net56));
 BUFx3_ASAP7_75t_R input57 (.A(r_i[27]),
    .Y(net57));
 BUFx3_ASAP7_75t_R input58 (.A(r_i[28]),
    .Y(net58));
 BUFx3_ASAP7_75t_R input59 (.A(r_i[29]),
    .Y(net59));
 BUFx3_ASAP7_75t_R input60 (.A(r_i[2]),
    .Y(net60));
 BUFx3_ASAP7_75t_R input61 (.A(r_i[30]),
    .Y(net61));
 BUFx3_ASAP7_75t_R input62 (.A(r_i[31]),
    .Y(net62));
 BUFx3_ASAP7_75t_R input63 (.A(r_i[32]),
    .Y(net63));
 BUFx3_ASAP7_75t_R input64 (.A(r_i[33]),
    .Y(net64));
 BUFx3_ASAP7_75t_R input65 (.A(r_i[34]),
    .Y(net65));
 BUFx3_ASAP7_75t_R input66 (.A(r_i[35]),
    .Y(net66));
 BUFx3_ASAP7_75t_R input67 (.A(r_i[3]),
    .Y(net67));
 BUFx3_ASAP7_75t_R input68 (.A(r_i[4]),
    .Y(net68));
 BUFx3_ASAP7_75t_R input69 (.A(r_i[5]),
    .Y(net69));
 BUFx3_ASAP7_75t_R input70 (.A(r_i[6]),
    .Y(net70));
 BUFx3_ASAP7_75t_R input71 (.A(r_i[7]),
    .Y(net71));
 BUFx3_ASAP7_75t_R input72 (.A(r_i[8]),
    .Y(net72));
 BUFx3_ASAP7_75t_R input73 (.A(r_i[9]),
    .Y(net73));
 BUFx3_ASAP7_75t_R input74 (.A(r_i_v),
    .Y(net74));
 BUFx3_ASAP7_75t_R input75 (.A(r_o_bp),
    .Y(net75));
 BUFx3_ASAP7_75t_R input76 (.A(u0_i[0]),
    .Y(net76));
 BUFx3_ASAP7_75t_R input77 (.A(u0_i[10]),
    .Y(net77));
 BUFx3_ASAP7_75t_R input78 (.A(u0_i[11]),
    .Y(net78));
 BUFx3_ASAP7_75t_R input79 (.A(u0_i[12]),
    .Y(net79));
 BUFx3_ASAP7_75t_R input80 (.A(u0_i[13]),
    .Y(net80));
 BUFx3_ASAP7_75t_R input81 (.A(u0_i[14]),
    .Y(net81));
 BUFx3_ASAP7_75t_R input82 (.A(u0_i[15]),
    .Y(net82));
 BUFx3_ASAP7_75t_R input83 (.A(u0_i[16]),
    .Y(net83));
 BUFx3_ASAP7_75t_R input84 (.A(u0_i[17]),
    .Y(net84));
 BUFx3_ASAP7_75t_R input85 (.A(u0_i[18]),
    .Y(net85));
 BUFx3_ASAP7_75t_R input86 (.A(u0_i[19]),
    .Y(net86));
 BUFx3_ASAP7_75t_R input87 (.A(u0_i[1]),
    .Y(net87));
 BUFx3_ASAP7_75t_R input88 (.A(u0_i[20]),
    .Y(net88));
 BUFx3_ASAP7_75t_R input89 (.A(u0_i[21]),
    .Y(net89));
 BUFx3_ASAP7_75t_R input90 (.A(u0_i[22]),
    .Y(net90));
 BUFx3_ASAP7_75t_R input91 (.A(u0_i[23]),
    .Y(net91));
 BUFx3_ASAP7_75t_R input92 (.A(u0_i[24]),
    .Y(net92));
 BUFx3_ASAP7_75t_R input93 (.A(u0_i[25]),
    .Y(net93));
 BUFx3_ASAP7_75t_R input94 (.A(u0_i[26]),
    .Y(net94));
 BUFx3_ASAP7_75t_R input95 (.A(u0_i[27]),
    .Y(net95));
 BUFx3_ASAP7_75t_R input96 (.A(u0_i[28]),
    .Y(net96));
 BUFx3_ASAP7_75t_R input97 (.A(u0_i[29]),
    .Y(net97));
 BUFx3_ASAP7_75t_R input98 (.A(u0_i[2]),
    .Y(net98));
 BUFx3_ASAP7_75t_R input99 (.A(u0_i[30]),
    .Y(net99));
 BUFx3_ASAP7_75t_R input100 (.A(u0_i[31]),
    .Y(net100));
 BUFx3_ASAP7_75t_R input101 (.A(u0_i[32]),
    .Y(net101));
 BUFx3_ASAP7_75t_R input102 (.A(u0_i[33]),
    .Y(net102));
 BUFx3_ASAP7_75t_R input103 (.A(u0_i[34]),
    .Y(net103));
 BUFx3_ASAP7_75t_R input104 (.A(u0_i[35]),
    .Y(net104));
 BUFx3_ASAP7_75t_R input105 (.A(u0_i[3]),
    .Y(net105));
 BUFx3_ASAP7_75t_R input106 (.A(u0_i[4]),
    .Y(net106));
 BUFx3_ASAP7_75t_R input107 (.A(u0_i[5]),
    .Y(net107));
 BUFx3_ASAP7_75t_R input108 (.A(u0_i[6]),
    .Y(net108));
 BUFx3_ASAP7_75t_R input109 (.A(u0_i[7]),
    .Y(net109));
 BUFx3_ASAP7_75t_R input110 (.A(u0_i[8]),
    .Y(net110));
 BUFx3_ASAP7_75t_R input111 (.A(u0_i[9]),
    .Y(net111));
 BUFx3_ASAP7_75t_R input112 (.A(u0_o_bp),
    .Y(net112));
 BUFx3_ASAP7_75t_R input113 (.A(u1_i[0]),
    .Y(net113));
 BUFx3_ASAP7_75t_R input114 (.A(u1_i[10]),
    .Y(net114));
 BUFx3_ASAP7_75t_R input115 (.A(u1_i[11]),
    .Y(net115));
 BUFx3_ASAP7_75t_R input116 (.A(u1_i[12]),
    .Y(net116));
 BUFx3_ASAP7_75t_R input117 (.A(u1_i[13]),
    .Y(net117));
 BUFx3_ASAP7_75t_R input118 (.A(u1_i[14]),
    .Y(net118));
 BUFx3_ASAP7_75t_R input119 (.A(u1_i[15]),
    .Y(net119));
 BUFx3_ASAP7_75t_R input120 (.A(u1_i[16]),
    .Y(net120));
 BUFx3_ASAP7_75t_R input121 (.A(u1_i[17]),
    .Y(net121));
 BUFx3_ASAP7_75t_R input122 (.A(u1_i[18]),
    .Y(net122));
 BUFx3_ASAP7_75t_R input123 (.A(u1_i[19]),
    .Y(net123));
 BUFx3_ASAP7_75t_R input124 (.A(u1_i[1]),
    .Y(net124));
 BUFx3_ASAP7_75t_R input125 (.A(u1_i[20]),
    .Y(net125));
 BUFx3_ASAP7_75t_R input126 (.A(u1_i[21]),
    .Y(net126));
 BUFx3_ASAP7_75t_R input127 (.A(u1_i[22]),
    .Y(net127));
 BUFx3_ASAP7_75t_R input128 (.A(u1_i[23]),
    .Y(net128));
 BUFx3_ASAP7_75t_R input129 (.A(u1_i[24]),
    .Y(net129));
 BUFx3_ASAP7_75t_R input130 (.A(u1_i[25]),
    .Y(net130));
 BUFx3_ASAP7_75t_R input131 (.A(u1_i[26]),
    .Y(net131));
 BUFx3_ASAP7_75t_R input132 (.A(u1_i[27]),
    .Y(net132));
 BUFx3_ASAP7_75t_R input133 (.A(u1_i[28]),
    .Y(net133));
 BUFx3_ASAP7_75t_R input134 (.A(u1_i[29]),
    .Y(net134));
 BUFx3_ASAP7_75t_R input135 (.A(u1_i[2]),
    .Y(net135));
 BUFx3_ASAP7_75t_R input136 (.A(u1_i[30]),
    .Y(net136));
 BUFx3_ASAP7_75t_R input137 (.A(u1_i[31]),
    .Y(net137));
 BUFx3_ASAP7_75t_R input138 (.A(u1_i[32]),
    .Y(net138));
 BUFx3_ASAP7_75t_R input139 (.A(u1_i[33]),
    .Y(net139));
 BUFx3_ASAP7_75t_R input140 (.A(u1_i[34]),
    .Y(net140));
 BUFx3_ASAP7_75t_R input141 (.A(u1_i[35]),
    .Y(net141));
 BUFx3_ASAP7_75t_R input142 (.A(u1_i[3]),
    .Y(net142));
 BUFx3_ASAP7_75t_R input143 (.A(u1_i[4]),
    .Y(net143));
 BUFx3_ASAP7_75t_R input144 (.A(u1_i[5]),
    .Y(net144));
 BUFx3_ASAP7_75t_R input145 (.A(u1_i[6]),
    .Y(net145));
 BUFx3_ASAP7_75t_R input146 (.A(u1_i[7]),
    .Y(net146));
 BUFx3_ASAP7_75t_R input147 (.A(u1_i[8]),
    .Y(net147));
 BUFx3_ASAP7_75t_R input148 (.A(u1_i[9]),
    .Y(net148));
 BUFx3_ASAP7_75t_R input149 (.A(u1_i_v),
    .Y(net149));
 BUFx3_ASAP7_75t_R input150 (.A(u1_o_bp),
    .Y(net150));
 BUFx3_ASAP7_75t_R output151 (.A(net151),
    .Y(l_i_bp));
 BUFx3_ASAP7_75t_R output152 (.A(net152),
    .Y(l_o[0]));
 BUFx3_ASAP7_75t_R output153 (.A(net153),
    .Y(l_o[10]));
 BUFx3_ASAP7_75t_R output154 (.A(net154),
    .Y(l_o[11]));
 BUFx3_ASAP7_75t_R output155 (.A(net155),
    .Y(l_o[12]));
 BUFx3_ASAP7_75t_R output156 (.A(net156),
    .Y(l_o[13]));
 BUFx3_ASAP7_75t_R output157 (.A(net157),
    .Y(l_o[14]));
 BUFx3_ASAP7_75t_R output158 (.A(net158),
    .Y(l_o[15]));
 BUFx3_ASAP7_75t_R output159 (.A(net159),
    .Y(l_o[16]));
 BUFx3_ASAP7_75t_R output160 (.A(net160),
    .Y(l_o[17]));
 BUFx3_ASAP7_75t_R output161 (.A(net161),
    .Y(l_o[18]));
 BUFx3_ASAP7_75t_R output162 (.A(net162),
    .Y(l_o[19]));
 BUFx3_ASAP7_75t_R output163 (.A(net163),
    .Y(l_o[1]));
 BUFx3_ASAP7_75t_R output164 (.A(net164),
    .Y(l_o[20]));
 BUFx3_ASAP7_75t_R output165 (.A(net165),
    .Y(l_o[21]));
 BUFx3_ASAP7_75t_R output166 (.A(net166),
    .Y(l_o[22]));
 BUFx3_ASAP7_75t_R output167 (.A(net167),
    .Y(l_o[23]));
 BUFx3_ASAP7_75t_R output168 (.A(net168),
    .Y(l_o[24]));
 BUFx3_ASAP7_75t_R output169 (.A(net169),
    .Y(l_o[25]));
 BUFx3_ASAP7_75t_R output170 (.A(net170),
    .Y(l_o[26]));
 BUFx3_ASAP7_75t_R output171 (.A(net171),
    .Y(l_o[27]));
 BUFx3_ASAP7_75t_R output172 (.A(net172),
    .Y(l_o[28]));
 BUFx3_ASAP7_75t_R output173 (.A(net173),
    .Y(l_o[29]));
 BUFx3_ASAP7_75t_R output174 (.A(net174),
    .Y(l_o[2]));
 BUFx3_ASAP7_75t_R output175 (.A(net175),
    .Y(l_o[30]));
 BUFx3_ASAP7_75t_R output176 (.A(net176),
    .Y(l_o[31]));
 BUFx3_ASAP7_75t_R output177 (.A(net177),
    .Y(l_o[32]));
 BUFx3_ASAP7_75t_R output178 (.A(net178),
    .Y(l_o[33]));
 BUFx3_ASAP7_75t_R output179 (.A(net179),
    .Y(l_o[34]));
 BUFx3_ASAP7_75t_R output180 (.A(net180),
    .Y(l_o[35]));
 BUFx3_ASAP7_75t_R output181 (.A(net181),
    .Y(l_o[3]));
 BUFx3_ASAP7_75t_R output182 (.A(net182),
    .Y(l_o[4]));
 BUFx3_ASAP7_75t_R output183 (.A(net183),
    .Y(l_o[5]));
 BUFx3_ASAP7_75t_R output184 (.A(net184),
    .Y(l_o[6]));
 BUFx3_ASAP7_75t_R output185 (.A(net185),
    .Y(l_o[7]));
 BUFx3_ASAP7_75t_R output186 (.A(net186),
    .Y(l_o[8]));
 BUFx3_ASAP7_75t_R output187 (.A(net187),
    .Y(l_o[9]));
 BUFx3_ASAP7_75t_R output188 (.A(net188),
    .Y(l_o_v));
 BUFx3_ASAP7_75t_R output189 (.A(net189),
    .Y(r_i_bp));
 BUFx3_ASAP7_75t_R output190 (.A(net190),
    .Y(r_o[0]));
 BUFx3_ASAP7_75t_R output191 (.A(net191),
    .Y(r_o[10]));
 BUFx3_ASAP7_75t_R output192 (.A(net192),
    .Y(r_o[11]));
 BUFx3_ASAP7_75t_R output193 (.A(net193),
    .Y(r_o[12]));
 BUFx3_ASAP7_75t_R output194 (.A(net194),
    .Y(r_o[13]));
 BUFx3_ASAP7_75t_R output195 (.A(net195),
    .Y(r_o[14]));
 BUFx3_ASAP7_75t_R output196 (.A(net196),
    .Y(r_o[15]));
 BUFx3_ASAP7_75t_R output197 (.A(net197),
    .Y(r_o[16]));
 BUFx3_ASAP7_75t_R output198 (.A(net198),
    .Y(r_o[17]));
 BUFx3_ASAP7_75t_R output199 (.A(net199),
    .Y(r_o[18]));
 BUFx3_ASAP7_75t_R output200 (.A(net200),
    .Y(r_o[19]));
 BUFx3_ASAP7_75t_R output201 (.A(net201),
    .Y(r_o[1]));
 BUFx3_ASAP7_75t_R output202 (.A(net202),
    .Y(r_o[20]));
 BUFx3_ASAP7_75t_R output203 (.A(net203),
    .Y(r_o[21]));
 BUFx3_ASAP7_75t_R output204 (.A(net204),
    .Y(r_o[22]));
 BUFx3_ASAP7_75t_R output205 (.A(net205),
    .Y(r_o[23]));
 BUFx3_ASAP7_75t_R output206 (.A(net206),
    .Y(r_o[24]));
 BUFx3_ASAP7_75t_R output207 (.A(net207),
    .Y(r_o[25]));
 BUFx3_ASAP7_75t_R output208 (.A(net208),
    .Y(r_o[26]));
 BUFx3_ASAP7_75t_R output209 (.A(net209),
    .Y(r_o[27]));
 BUFx3_ASAP7_75t_R output210 (.A(net210),
    .Y(r_o[28]));
 BUFx3_ASAP7_75t_R output211 (.A(net211),
    .Y(r_o[29]));
 BUFx3_ASAP7_75t_R output212 (.A(net212),
    .Y(r_o[2]));
 BUFx3_ASAP7_75t_R output213 (.A(net213),
    .Y(r_o[30]));
 BUFx3_ASAP7_75t_R output214 (.A(net214),
    .Y(r_o[31]));
 BUFx3_ASAP7_75t_R output215 (.A(net215),
    .Y(r_o[32]));
 BUFx3_ASAP7_75t_R output216 (.A(net216),
    .Y(r_o[33]));
 BUFx3_ASAP7_75t_R output217 (.A(net217),
    .Y(r_o[34]));
 BUFx3_ASAP7_75t_R output218 (.A(net218),
    .Y(r_o[35]));
 BUFx3_ASAP7_75t_R output219 (.A(net219),
    .Y(r_o[3]));
 BUFx3_ASAP7_75t_R output220 (.A(net220),
    .Y(r_o[4]));
 BUFx3_ASAP7_75t_R output221 (.A(net221),
    .Y(r_o[5]));
 BUFx3_ASAP7_75t_R output222 (.A(net222),
    .Y(r_o[6]));
 BUFx3_ASAP7_75t_R output223 (.A(net223),
    .Y(r_o[7]));
 BUFx3_ASAP7_75t_R output224 (.A(net224),
    .Y(r_o[8]));
 BUFx3_ASAP7_75t_R output225 (.A(net225),
    .Y(r_o[9]));
 BUFx3_ASAP7_75t_R output226 (.A(net226),
    .Y(r_o_v));
 BUFx3_ASAP7_75t_R output227 (.A(net227),
    .Y(u0_i_bp));
 BUFx3_ASAP7_75t_R output228 (.A(net228),
    .Y(u0_o[0]));
 BUFx3_ASAP7_75t_R output229 (.A(net229),
    .Y(u0_o[10]));
 BUFx3_ASAP7_75t_R output230 (.A(net230),
    .Y(u0_o[11]));
 BUFx3_ASAP7_75t_R output231 (.A(net231),
    .Y(u0_o[12]));
 BUFx3_ASAP7_75t_R output232 (.A(net232),
    .Y(u0_o[13]));
 BUFx3_ASAP7_75t_R output233 (.A(net233),
    .Y(u0_o[14]));
 BUFx3_ASAP7_75t_R output234 (.A(net234),
    .Y(u0_o[15]));
 BUFx3_ASAP7_75t_R output235 (.A(net235),
    .Y(u0_o[16]));
 BUFx3_ASAP7_75t_R output236 (.A(net236),
    .Y(u0_o[17]));
 BUFx3_ASAP7_75t_R output237 (.A(net237),
    .Y(u0_o[18]));
 BUFx3_ASAP7_75t_R output238 (.A(net238),
    .Y(u0_o[19]));
 BUFx3_ASAP7_75t_R output239 (.A(net239),
    .Y(u0_o[1]));
 BUFx3_ASAP7_75t_R output240 (.A(net240),
    .Y(u0_o[20]));
 BUFx3_ASAP7_75t_R output241 (.A(net241),
    .Y(u0_o[21]));
 BUFx3_ASAP7_75t_R output242 (.A(net242),
    .Y(u0_o[22]));
 BUFx3_ASAP7_75t_R output243 (.A(net243),
    .Y(u0_o[23]));
 BUFx3_ASAP7_75t_R output244 (.A(net244),
    .Y(u0_o[24]));
 BUFx3_ASAP7_75t_R output245 (.A(net245),
    .Y(u0_o[25]));
 BUFx3_ASAP7_75t_R output246 (.A(net246),
    .Y(u0_o[26]));
 BUFx3_ASAP7_75t_R output247 (.A(net247),
    .Y(u0_o[27]));
 BUFx3_ASAP7_75t_R output248 (.A(net248),
    .Y(u0_o[28]));
 BUFx3_ASAP7_75t_R output249 (.A(net249),
    .Y(u0_o[29]));
 BUFx3_ASAP7_75t_R output250 (.A(net250),
    .Y(u0_o[2]));
 BUFx3_ASAP7_75t_R output251 (.A(net251),
    .Y(u0_o[30]));
 BUFx3_ASAP7_75t_R output252 (.A(net252),
    .Y(u0_o[31]));
 BUFx3_ASAP7_75t_R output253 (.A(net253),
    .Y(u0_o[32]));
 BUFx3_ASAP7_75t_R output254 (.A(net254),
    .Y(u0_o[33]));
 BUFx3_ASAP7_75t_R output255 (.A(net255),
    .Y(u0_o[34]));
 BUFx3_ASAP7_75t_R output256 (.A(net256),
    .Y(u0_o[35]));
 BUFx3_ASAP7_75t_R output257 (.A(net257),
    .Y(u0_o[3]));
 BUFx3_ASAP7_75t_R output258 (.A(net258),
    .Y(u0_o[4]));
 BUFx3_ASAP7_75t_R output259 (.A(net259),
    .Y(u0_o[5]));
 BUFx3_ASAP7_75t_R output260 (.A(net260),
    .Y(u0_o[6]));
 BUFx3_ASAP7_75t_R output261 (.A(net261),
    .Y(u0_o[7]));
 BUFx3_ASAP7_75t_R output262 (.A(net262),
    .Y(u0_o[8]));
 BUFx3_ASAP7_75t_R output263 (.A(net263),
    .Y(u0_o[9]));
 BUFx3_ASAP7_75t_R output264 (.A(net264),
    .Y(u0_o_v));
 BUFx3_ASAP7_75t_R output265 (.A(net265),
    .Y(u1_i_bp));
 BUFx3_ASAP7_75t_R output266 (.A(net266),
    .Y(u1_o[0]));
 BUFx3_ASAP7_75t_R output267 (.A(net267),
    .Y(u1_o[10]));
 BUFx3_ASAP7_75t_R output268 (.A(net268),
    .Y(u1_o[11]));
 BUFx3_ASAP7_75t_R output269 (.A(net269),
    .Y(u1_o[12]));
 BUFx3_ASAP7_75t_R output270 (.A(net270),
    .Y(u1_o[13]));
 BUFx3_ASAP7_75t_R output271 (.A(net271),
    .Y(u1_o[14]));
 BUFx3_ASAP7_75t_R output272 (.A(net272),
    .Y(u1_o[15]));
 BUFx3_ASAP7_75t_R output273 (.A(net273),
    .Y(u1_o[16]));
 BUFx3_ASAP7_75t_R output274 (.A(net274),
    .Y(u1_o[17]));
 BUFx3_ASAP7_75t_R output275 (.A(net275),
    .Y(u1_o[18]));
 BUFx3_ASAP7_75t_R output276 (.A(net276),
    .Y(u1_o[19]));
 BUFx3_ASAP7_75t_R output277 (.A(net277),
    .Y(u1_o[1]));
 BUFx3_ASAP7_75t_R output278 (.A(net278),
    .Y(u1_o[20]));
 BUFx3_ASAP7_75t_R output279 (.A(net279),
    .Y(u1_o[21]));
 BUFx3_ASAP7_75t_R output280 (.A(net280),
    .Y(u1_o[22]));
 BUFx3_ASAP7_75t_R output281 (.A(net281),
    .Y(u1_o[23]));
 BUFx3_ASAP7_75t_R output282 (.A(net282),
    .Y(u1_o[24]));
 BUFx3_ASAP7_75t_R output283 (.A(net283),
    .Y(u1_o[25]));
 BUFx3_ASAP7_75t_R output284 (.A(net284),
    .Y(u1_o[26]));
 BUFx3_ASAP7_75t_R output285 (.A(net285),
    .Y(u1_o[27]));
 BUFx3_ASAP7_75t_R output286 (.A(net286),
    .Y(u1_o[28]));
 BUFx3_ASAP7_75t_R output287 (.A(net287),
    .Y(u1_o[29]));
 BUFx3_ASAP7_75t_R output288 (.A(net288),
    .Y(u1_o[2]));
 BUFx3_ASAP7_75t_R output289 (.A(net289),
    .Y(u1_o[30]));
 BUFx3_ASAP7_75t_R output290 (.A(net290),
    .Y(u1_o[31]));
 BUFx3_ASAP7_75t_R output291 (.A(net291),
    .Y(u1_o[32]));
 BUFx3_ASAP7_75t_R output292 (.A(net292),
    .Y(u1_o[33]));
 BUFx3_ASAP7_75t_R output293 (.A(net293),
    .Y(u1_o[34]));
 BUFx3_ASAP7_75t_R output294 (.A(net294),
    .Y(u1_o[35]));
 BUFx3_ASAP7_75t_R output295 (.A(net295),
    .Y(u1_o[3]));
 BUFx3_ASAP7_75t_R output296 (.A(net296),
    .Y(u1_o[4]));
 BUFx3_ASAP7_75t_R output297 (.A(net297),
    .Y(u1_o[5]));
 BUFx3_ASAP7_75t_R output298 (.A(net298),
    .Y(u1_o[6]));
 BUFx3_ASAP7_75t_R output299 (.A(net299),
    .Y(u1_o[7]));
 BUFx3_ASAP7_75t_R output300 (.A(net300),
    .Y(u1_o[8]));
 BUFx3_ASAP7_75t_R output301 (.A(net301),
    .Y(u1_o[9]));
 BUFx3_ASAP7_75t_R output302 (.A(net302),
    .Y(u1_o_v));
 TIELOx1_ASAP7_75t_R _1534__303 (.L(net303));
 BUFx10_ASAP7_75t_R clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_0_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_1_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_2_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_3_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_4_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_5_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_6_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_7_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_8_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_9_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_10_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_11_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_12_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_13_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_14_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_15_0_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload0 (.A(clknet_4_0_0_clk));
 INVx8_ASAP7_75t_R clkload1 (.A(clknet_4_1_0_clk));
 INVx6_ASAP7_75t_R clkload2 (.A(clknet_4_2_0_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload3 (.A(clknet_4_3_0_clk));
 BUFx24_ASAP7_75t_R clkload4 (.A(clknet_4_4_0_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload5 (.A(clknet_4_6_0_clk));
 INVx5_ASAP7_75t_R clkload6 (.A(clknet_4_7_0_clk));
 INVx5_ASAP7_75t_R clkload7 (.A(clknet_4_8_0_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload8 (.A(clknet_4_9_0_clk));
 INVx6_ASAP7_75t_R clkload9 (.A(clknet_4_11_0_clk));
 INVx8_ASAP7_75t_R clkload10 (.A(clknet_4_12_0_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload11 (.A(clknet_4_13_0_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload12 (.A(clknet_4_14_0_clk));
 INVx3_ASAP7_75t_R clkload13 (.A(clknet_4_15_0_clk));
 FILLERxp5_ASAP7_75t_R FILLER_0_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57 ();
 FILLER_ASAP7_75t_R FILLER_0_69 ();
 FILLER_ASAP7_75t_R FILLER_0_77 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91 ();
 FILLER_ASAP7_75t_R FILLER_0_101 ();
 DECAPx6_ASAP7_75t_R FILLER_0_109 ();
 FILLER_ASAP7_75t_R FILLER_0_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161 ();
 FILLER_ASAP7_75t_R FILLER_0_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_289 ();
 DECAPx2_ASAP7_75t_R FILLER_0_302 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx4_ASAP7_75t_R FILLER_1_46 ();
 FILLER_ASAP7_75t_R FILLER_1_56 ();
 DECAPx1_ASAP7_75t_R FILLER_1_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_85 ();
 DECAPx4_ASAP7_75t_R FILLER_1_92 ();
 FILLER_ASAP7_75t_R FILLER_1_102 ();
 DECAPx2_ASAP7_75t_R FILLER_1_114 ();
 FILLER_ASAP7_75t_R FILLER_1_120 ();
 DECAPx2_ASAP7_75t_R FILLER_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_1_258 ();
 DECAPx10_ASAP7_75t_R FILLER_1_280 ();
 DECAPx1_ASAP7_75t_R FILLER_1_302 ();
 FILLER_ASAP7_75t_R FILLER_1_312 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx6_ASAP7_75t_R FILLER_2_24 ();
 DECAPx1_ASAP7_75t_R FILLER_2_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_42 ();
 DECAPx2_ASAP7_75t_R FILLER_2_63 ();
 FILLER_ASAP7_75t_R FILLER_2_69 ();
 DECAPx10_ASAP7_75t_R FILLER_2_77 ();
 DECAPx10_ASAP7_75t_R FILLER_2_99 ();
 DECAPx6_ASAP7_75t_R FILLER_2_121 ();
 DECAPx1_ASAP7_75t_R FILLER_2_141 ();
 DECAPx10_ASAP7_75t_R FILLER_2_252 ();
 DECAPx10_ASAP7_75t_R FILLER_2_274 ();
 DECAPx6_ASAP7_75t_R FILLER_2_296 ();
 DECAPx1_ASAP7_75t_R FILLER_2_310 ();
 DECAPx6_ASAP7_75t_R FILLER_3_2 ();
 DECAPx1_ASAP7_75t_R FILLER_3_16 ();
 DECAPx6_ASAP7_75t_R FILLER_3_29 ();
 DECAPx1_ASAP7_75t_R FILLER_3_43 ();
 FILLER_ASAP7_75t_R FILLER_3_64 ();
 DECAPx10_ASAP7_75t_R FILLER_3_74 ();
 DECAPx10_ASAP7_75t_R FILLER_3_96 ();
 DECAPx6_ASAP7_75t_R FILLER_3_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_132 ();
 DECAPx2_ASAP7_75t_R FILLER_3_139 ();
 DECAPx1_ASAP7_75t_R FILLER_3_183 ();
 FILLER_ASAP7_75t_R FILLER_3_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_195 ();
 DECAPx1_ASAP7_75t_R FILLER_3_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_216 ();
 FILLER_ASAP7_75t_R FILLER_3_223 ();
 DECAPx1_ASAP7_75t_R FILLER_3_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_247 ();
 DECAPx10_ASAP7_75t_R FILLER_3_254 ();
 DECAPx10_ASAP7_75t_R FILLER_3_276 ();
 DECAPx6_ASAP7_75t_R FILLER_3_298 ();
 FILLER_ASAP7_75t_R FILLER_3_312 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_44 ();
 DECAPx6_ASAP7_75t_R FILLER_4_66 ();
 DECAPx1_ASAP7_75t_R FILLER_4_80 ();
 DECAPx1_ASAP7_75t_R FILLER_4_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_122 ();
 FILLER_ASAP7_75t_R FILLER_4_146 ();
 DECAPx1_ASAP7_75t_R FILLER_4_158 ();
 DECAPx4_ASAP7_75t_R FILLER_4_180 ();
 FILLER_ASAP7_75t_R FILLER_4_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_192 ();
 DECAPx2_ASAP7_75t_R FILLER_4_216 ();
 FILLER_ASAP7_75t_R FILLER_4_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_244 ();
 DECAPx10_ASAP7_75t_R FILLER_4_268 ();
 DECAPx10_ASAP7_75t_R FILLER_4_290 ();
 FILLER_ASAP7_75t_R FILLER_4_312 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 FILLER_ASAP7_75t_R FILLER_5_24 ();
 FILLER_ASAP7_75t_R FILLER_5_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_31 ();
 DECAPx6_ASAP7_75t_R FILLER_5_46 ();
 DECAPx1_ASAP7_75t_R FILLER_5_60 ();
 DECAPx2_ASAP7_75t_R FILLER_5_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_76 ();
 DECAPx10_ASAP7_75t_R FILLER_5_95 ();
 DECAPx2_ASAP7_75t_R FILLER_5_117 ();
 FILLER_ASAP7_75t_R FILLER_5_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_125 ();
 DECAPx2_ASAP7_75t_R FILLER_5_134 ();
 FILLER_ASAP7_75t_R FILLER_5_140 ();
 FILLER_ASAP7_75t_R FILLER_5_165 ();
 DECAPx2_ASAP7_75t_R FILLER_5_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_193 ();
 DECAPx1_ASAP7_75t_R FILLER_5_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_212 ();
 DECAPx10_ASAP7_75t_R FILLER_5_262 ();
 DECAPx10_ASAP7_75t_R FILLER_5_284 ();
 DECAPx2_ASAP7_75t_R FILLER_5_306 ();
 FILLER_ASAP7_75t_R FILLER_5_312 ();
 DECAPx6_ASAP7_75t_R FILLER_6_2 ();
 DECAPx4_ASAP7_75t_R FILLER_6_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_62 ();
 FILLER_ASAP7_75t_R FILLER_6_69 ();
 DECAPx1_ASAP7_75t_R FILLER_6_77 ();
 FILLER_ASAP7_75t_R FILLER_6_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_93 ();
 DECAPx1_ASAP7_75t_R FILLER_6_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_108 ();
 FILLER_ASAP7_75t_R FILLER_6_117 ();
 DECAPx1_ASAP7_75t_R FILLER_6_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_131 ();
 DECAPx2_ASAP7_75t_R FILLER_6_140 ();
 FILLER_ASAP7_75t_R FILLER_6_146 ();
 DECAPx6_ASAP7_75t_R FILLER_6_154 ();
 DECAPx1_ASAP7_75t_R FILLER_6_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_172 ();
 DECAPx1_ASAP7_75t_R FILLER_6_195 ();
 DECAPx6_ASAP7_75t_R FILLER_6_213 ();
 DECAPx2_ASAP7_75t_R FILLER_6_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_239 ();
 DECAPx1_ASAP7_75t_R FILLER_6_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_264 ();
 DECAPx6_ASAP7_75t_R FILLER_6_296 ();
 DECAPx1_ASAP7_75t_R FILLER_6_310 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx4_ASAP7_75t_R FILLER_7_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_34 ();
 DECAPx2_ASAP7_75t_R FILLER_7_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_61 ();
 DECAPx1_ASAP7_75t_R FILLER_7_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_74 ();
 FILLER_ASAP7_75t_R FILLER_7_101 ();
 FILLER_ASAP7_75t_R FILLER_7_115 ();
 DECAPx10_ASAP7_75t_R FILLER_7_124 ();
 DECAPx6_ASAP7_75t_R FILLER_7_146 ();
 DECAPx2_ASAP7_75t_R FILLER_7_160 ();
 DECAPx1_ASAP7_75t_R FILLER_7_183 ();
 DECAPx6_ASAP7_75t_R FILLER_7_190 ();
 DECAPx4_ASAP7_75t_R FILLER_7_207 ();
 FILLER_ASAP7_75t_R FILLER_7_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_219 ();
 DECAPx4_ASAP7_75t_R FILLER_7_228 ();
 FILLER_ASAP7_75t_R FILLER_7_238 ();
 FILLER_ASAP7_75t_R FILLER_7_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_248 ();
 DECAPx1_ASAP7_75t_R FILLER_7_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_265 ();
 DECAPx10_ASAP7_75t_R FILLER_7_272 ();
 DECAPx6_ASAP7_75t_R FILLER_7_294 ();
 DECAPx2_ASAP7_75t_R FILLER_7_308 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx6_ASAP7_75t_R FILLER_8_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_38 ();
 FILLER_ASAP7_75t_R FILLER_8_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_95 ();
 FILLER_ASAP7_75t_R FILLER_8_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_110 ();
 DECAPx2_ASAP7_75t_R FILLER_8_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_133 ();
 DECAPx4_ASAP7_75t_R FILLER_8_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_186 ();
 DECAPx4_ASAP7_75t_R FILLER_8_193 ();
 DECAPx1_ASAP7_75t_R FILLER_8_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_213 ();
 FILLER_ASAP7_75t_R FILLER_8_243 ();
 DECAPx6_ASAP7_75t_R FILLER_8_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_268 ();
 DECAPx6_ASAP7_75t_R FILLER_8_298 ();
 FILLER_ASAP7_75t_R FILLER_8_312 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx2_ASAP7_75t_R FILLER_9_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_30 ();
 DECAPx4_ASAP7_75t_R FILLER_9_41 ();
 FILLER_ASAP7_75t_R FILLER_9_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_65 ();
 FILLER_ASAP7_75t_R FILLER_9_74 ();
 DECAPx6_ASAP7_75t_R FILLER_9_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_94 ();
 DECAPx4_ASAP7_75t_R FILLER_9_101 ();
 DECAPx2_ASAP7_75t_R FILLER_9_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_123 ();
 DECAPx10_ASAP7_75t_R FILLER_9_134 ();
 DECAPx10_ASAP7_75t_R FILLER_9_156 ();
 DECAPx2_ASAP7_75t_R FILLER_9_178 ();
 FILLER_ASAP7_75t_R FILLER_9_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_213 ();
 DECAPx6_ASAP7_75t_R FILLER_9_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_245 ();
 FILLER_ASAP7_75t_R FILLER_9_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_268 ();
 DECAPx10_ASAP7_75t_R FILLER_9_278 ();
 DECAPx6_ASAP7_75t_R FILLER_9_300 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx2_ASAP7_75t_R FILLER_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_10_48 ();
 DECAPx2_ASAP7_75t_R FILLER_10_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_76 ();
 DECAPx10_ASAP7_75t_R FILLER_10_105 ();
 DECAPx2_ASAP7_75t_R FILLER_10_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_143 ();
 FILLER_ASAP7_75t_R FILLER_10_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_169 ();
 DECAPx4_ASAP7_75t_R FILLER_10_173 ();
 FILLER_ASAP7_75t_R FILLER_10_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_185 ();
 FILLER_ASAP7_75t_R FILLER_10_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_198 ();
 DECAPx2_ASAP7_75t_R FILLER_10_209 ();
 FILLER_ASAP7_75t_R FILLER_10_215 ();
 DECAPx2_ASAP7_75t_R FILLER_10_227 ();
 FILLER_ASAP7_75t_R FILLER_10_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_235 ();
 DECAPx4_ASAP7_75t_R FILLER_10_242 ();
 FILLER_ASAP7_75t_R FILLER_10_252 ();
 FILLER_ASAP7_75t_R FILLER_10_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_263 ();
 DECAPx6_ASAP7_75t_R FILLER_10_281 ();
 FILLER_ASAP7_75t_R FILLER_10_295 ();
 DECAPx6_ASAP7_75t_R FILLER_10_300 ();
 DECAPx6_ASAP7_75t_R FILLER_11_2 ();
 DECAPx1_ASAP7_75t_R FILLER_11_16 ();
 DECAPx10_ASAP7_75t_R FILLER_11_26 ();
 DECAPx1_ASAP7_75t_R FILLER_11_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_52 ();
 DECAPx1_ASAP7_75t_R FILLER_11_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_77 ();
 FILLER_ASAP7_75t_R FILLER_11_88 ();
 DECAPx1_ASAP7_75t_R FILLER_11_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_108 ();
 DECAPx4_ASAP7_75t_R FILLER_11_125 ();
 DECAPx2_ASAP7_75t_R FILLER_11_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_169 ();
 FILLER_ASAP7_75t_R FILLER_11_194 ();
 FILLER_ASAP7_75t_R FILLER_11_216 ();
 DECAPx1_ASAP7_75t_R FILLER_11_226 ();
 DECAPx10_ASAP7_75t_R FILLER_11_242 ();
 DECAPx1_ASAP7_75t_R FILLER_11_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_268 ();
 DECAPx6_ASAP7_75t_R FILLER_11_298 ();
 FILLER_ASAP7_75t_R FILLER_11_312 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx6_ASAP7_75t_R FILLER_12_24 ();
 FILLER_ASAP7_75t_R FILLER_12_38 ();
 DECAPx1_ASAP7_75t_R FILLER_12_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_52 ();
 DECAPx1_ASAP7_75t_R FILLER_12_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_83 ();
 DECAPx1_ASAP7_75t_R FILLER_12_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_104 ();
 FILLER_ASAP7_75t_R FILLER_12_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_113 ();
 FILLER_ASAP7_75t_R FILLER_12_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_126 ();
 FILLER_ASAP7_75t_R FILLER_12_135 ();
 DECAPx6_ASAP7_75t_R FILLER_12_143 ();
 DECAPx1_ASAP7_75t_R FILLER_12_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_184 ();
 DECAPx10_ASAP7_75t_R FILLER_12_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_213 ();
 FILLER_ASAP7_75t_R FILLER_12_231 ();
 DECAPx6_ASAP7_75t_R FILLER_12_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_270 ();
 DECAPx10_ASAP7_75t_R FILLER_12_283 ();
 DECAPx2_ASAP7_75t_R FILLER_12_305 ();
 FILLER_ASAP7_75t_R FILLER_12_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_313 ();
 DECAPx6_ASAP7_75t_R FILLER_13_2 ();
 FILLER_ASAP7_75t_R FILLER_13_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_18 ();
 DECAPx1_ASAP7_75t_R FILLER_13_51 ();
 DECAPx10_ASAP7_75t_R FILLER_13_63 ();
 FILLER_ASAP7_75t_R FILLER_13_85 ();
 DECAPx1_ASAP7_75t_R FILLER_13_93 ();
 DECAPx1_ASAP7_75t_R FILLER_13_111 ();
 FILLER_ASAP7_75t_R FILLER_13_128 ();
 DECAPx4_ASAP7_75t_R FILLER_13_148 ();
 FILLER_ASAP7_75t_R FILLER_13_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_160 ();
 DECAPx10_ASAP7_75t_R FILLER_13_169 ();
 DECAPx6_ASAP7_75t_R FILLER_13_191 ();
 DECAPx2_ASAP7_75t_R FILLER_13_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_211 ();
 DECAPx2_ASAP7_75t_R FILLER_13_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_234 ();
 FILLER_ASAP7_75t_R FILLER_13_242 ();
 DECAPx2_ASAP7_75t_R FILLER_13_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_273 ();
 FILLER_ASAP7_75t_R FILLER_13_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_307 ();
 DECAPx10_ASAP7_75t_R FILLER_14_2 ();
 DECAPx4_ASAP7_75t_R FILLER_14_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_34 ();
 DECAPx10_ASAP7_75t_R FILLER_14_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_69 ();
 DECAPx1_ASAP7_75t_R FILLER_14_94 ();
 DECAPx1_ASAP7_75t_R FILLER_14_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_119 ();
 DECAPx6_ASAP7_75t_R FILLER_14_132 ();
 DECAPx2_ASAP7_75t_R FILLER_14_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_152 ();
 DECAPx6_ASAP7_75t_R FILLER_14_176 ();
 FILLER_ASAP7_75t_R FILLER_14_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_192 ();
 DECAPx1_ASAP7_75t_R FILLER_14_196 ();
 DECAPx10_ASAP7_75t_R FILLER_14_220 ();
 FILLER_ASAP7_75t_R FILLER_14_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_244 ();
 FILLER_ASAP7_75t_R FILLER_14_248 ();
 DECAPx10_ASAP7_75t_R FILLER_14_259 ();
 DECAPx10_ASAP7_75t_R FILLER_14_281 ();
 DECAPx4_ASAP7_75t_R FILLER_14_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_313 ();
 DECAPx10_ASAP7_75t_R FILLER_15_2 ();
 DECAPx4_ASAP7_75t_R FILLER_15_24 ();
 FILLER_ASAP7_75t_R FILLER_15_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_53 ();
 DECAPx1_ASAP7_75t_R FILLER_15_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_70 ();
 FILLER_ASAP7_75t_R FILLER_15_81 ();
 FILLER_ASAP7_75t_R FILLER_15_97 ();
 FILLER_ASAP7_75t_R FILLER_15_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_114 ();
 DECAPx1_ASAP7_75t_R FILLER_15_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_135 ();
 DECAPx10_ASAP7_75t_R FILLER_15_139 ();
 FILLER_ASAP7_75t_R FILLER_15_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_163 ();
 DECAPx4_ASAP7_75t_R FILLER_15_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_180 ();
 DECAPx1_ASAP7_75t_R FILLER_15_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_211 ();
 FILLER_ASAP7_75t_R FILLER_15_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_224 ();
 DECAPx4_ASAP7_75t_R FILLER_15_239 ();
 FILLER_ASAP7_75t_R FILLER_15_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_258 ();
 DECAPx2_ASAP7_75t_R FILLER_15_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_272 ();
 FILLER_ASAP7_75t_R FILLER_15_279 ();
 DECAPx2_ASAP7_75t_R FILLER_15_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_307 ();
 DECAPx6_ASAP7_75t_R FILLER_16_2 ();
 DECAPx2_ASAP7_75t_R FILLER_16_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_58 ();
 DECAPx4_ASAP7_75t_R FILLER_16_66 ();
 FILLER_ASAP7_75t_R FILLER_16_76 ();
 DECAPx1_ASAP7_75t_R FILLER_16_82 ();
 DECAPx4_ASAP7_75t_R FILLER_16_94 ();
 FILLER_ASAP7_75t_R FILLER_16_104 ();
 FILLER_ASAP7_75t_R FILLER_16_118 ();
 DECAPx2_ASAP7_75t_R FILLER_16_162 ();
 FILLER_ASAP7_75t_R FILLER_16_168 ();
 DECAPx1_ASAP7_75t_R FILLER_16_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_252 ();
 DECAPx2_ASAP7_75t_R FILLER_16_262 ();
 FILLER_ASAP7_75t_R FILLER_16_268 ();
 FILLER_ASAP7_75t_R FILLER_16_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_313 ();
 DECAPx1_ASAP7_75t_R FILLER_17_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_59 ();
 DECAPx4_ASAP7_75t_R FILLER_17_76 ();
 FILLER_ASAP7_75t_R FILLER_17_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_136 ();
 DECAPx10_ASAP7_75t_R FILLER_17_151 ();
 DECAPx2_ASAP7_75t_R FILLER_17_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_179 ();
 DECAPx2_ASAP7_75t_R FILLER_17_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_197 ();
 DECAPx6_ASAP7_75t_R FILLER_17_234 ();
 DECAPx1_ASAP7_75t_R FILLER_17_248 ();
 DECAPx1_ASAP7_75t_R FILLER_17_275 ();
 DECAPx1_ASAP7_75t_R FILLER_17_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_301 ();
 DECAPx10_ASAP7_75t_R FILLER_18_2 ();
 DECAPx1_ASAP7_75t_R FILLER_18_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_28 ();
 DECAPx2_ASAP7_75t_R FILLER_18_44 ();
 FILLER_ASAP7_75t_R FILLER_18_50 ();
 DECAPx2_ASAP7_75t_R FILLER_18_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_82 ();
 FILLER_ASAP7_75t_R FILLER_18_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_101 ();
 FILLER_ASAP7_75t_R FILLER_18_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_141 ();
 DECAPx6_ASAP7_75t_R FILLER_18_148 ();
 DECAPx2_ASAP7_75t_R FILLER_18_162 ();
 DECAPx6_ASAP7_75t_R FILLER_18_178 ();
 FILLER_ASAP7_75t_R FILLER_18_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_194 ();
 DECAPx10_ASAP7_75t_R FILLER_18_232 ();
 DECAPx4_ASAP7_75t_R FILLER_18_254 ();
 FILLER_ASAP7_75t_R FILLER_18_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_266 ();
 DECAPx2_ASAP7_75t_R FILLER_18_274 ();
 DECAPx6_ASAP7_75t_R FILLER_18_300 ();
 DECAPx2_ASAP7_75t_R FILLER_19_2 ();
 FILLER_ASAP7_75t_R FILLER_19_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_16 ();
 DECAPx10_ASAP7_75t_R FILLER_19_23 ();
 DECAPx6_ASAP7_75t_R FILLER_19_45 ();
 DECAPx2_ASAP7_75t_R FILLER_19_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_65 ();
 DECAPx6_ASAP7_75t_R FILLER_19_88 ();
 DECAPx6_ASAP7_75t_R FILLER_19_166 ();
 FILLER_ASAP7_75t_R FILLER_19_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_182 ();
 FILLER_ASAP7_75t_R FILLER_19_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_205 ();
 DECAPx1_ASAP7_75t_R FILLER_19_209 ();
 DECAPx2_ASAP7_75t_R FILLER_19_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_229 ();
 FILLER_ASAP7_75t_R FILLER_19_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_242 ();
 FILLER_ASAP7_75t_R FILLER_19_249 ();
 FILLER_ASAP7_75t_R FILLER_19_262 ();
 DECAPx4_ASAP7_75t_R FILLER_19_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_289 ();
 DECAPx10_ASAP7_75t_R FILLER_20_2 ();
 DECAPx2_ASAP7_75t_R FILLER_20_24 ();
 DECAPx10_ASAP7_75t_R FILLER_20_38 ();
 DECAPx10_ASAP7_75t_R FILLER_20_60 ();
 DECAPx4_ASAP7_75t_R FILLER_20_82 ();
 DECAPx1_ASAP7_75t_R FILLER_20_108 ();
 DECAPx2_ASAP7_75t_R FILLER_20_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_152 ();
 DECAPx6_ASAP7_75t_R FILLER_20_163 ();
 DECAPx2_ASAP7_75t_R FILLER_20_177 ();
 DECAPx2_ASAP7_75t_R FILLER_20_206 ();
 FILLER_ASAP7_75t_R FILLER_20_212 ();
 DECAPx1_ASAP7_75t_R FILLER_20_237 ();
 DECAPx6_ASAP7_75t_R FILLER_20_296 ();
 DECAPx1_ASAP7_75t_R FILLER_20_310 ();
 DECAPx6_ASAP7_75t_R FILLER_21_2 ();
 FILLER_ASAP7_75t_R FILLER_21_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_66 ();
 DECAPx6_ASAP7_75t_R FILLER_21_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_87 ();
 FILLER_ASAP7_75t_R FILLER_21_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_106 ();
 FILLER_ASAP7_75t_R FILLER_21_127 ();
 DECAPx1_ASAP7_75t_R FILLER_21_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_145 ();
 DECAPx4_ASAP7_75t_R FILLER_21_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_176 ();
 DECAPx10_ASAP7_75t_R FILLER_21_187 ();
 DECAPx2_ASAP7_75t_R FILLER_21_209 ();
 FILLER_ASAP7_75t_R FILLER_21_215 ();
 DECAPx10_ASAP7_75t_R FILLER_21_240 ();
 DECAPx2_ASAP7_75t_R FILLER_21_262 ();
 FILLER_ASAP7_75t_R FILLER_21_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_2 ();
 DECAPx6_ASAP7_75t_R FILLER_22_9 ();
 DECAPx2_ASAP7_75t_R FILLER_22_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_29 ();
 DECAPx6_ASAP7_75t_R FILLER_22_39 ();
 FILLER_ASAP7_75t_R FILLER_22_53 ();
 DECAPx2_ASAP7_75t_R FILLER_22_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_88 ();
 FILLER_ASAP7_75t_R FILLER_22_111 ();
 DECAPx2_ASAP7_75t_R FILLER_22_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_180 ();
 FILLER_ASAP7_75t_R FILLER_22_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_218 ();
 DECAPx1_ASAP7_75t_R FILLER_22_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_259 ();
 DECAPx6_ASAP7_75t_R FILLER_22_263 ();
 DECAPx2_ASAP7_75t_R FILLER_22_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_283 ();
 DECAPx1_ASAP7_75t_R FILLER_22_304 ();
 FILLER_ASAP7_75t_R FILLER_23_2 ();
 DECAPx2_ASAP7_75t_R FILLER_23_16 ();
 DECAPx1_ASAP7_75t_R FILLER_23_25 ();
 DECAPx4_ASAP7_75t_R FILLER_23_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_51 ();
 DECAPx1_ASAP7_75t_R FILLER_23_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_103 ();
 DECAPx2_ASAP7_75t_R FILLER_23_113 ();
 FILLER_ASAP7_75t_R FILLER_23_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_121 ();
 FILLER_ASAP7_75t_R FILLER_23_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_138 ();
 DECAPx6_ASAP7_75t_R FILLER_23_159 ();
 DECAPx2_ASAP7_75t_R FILLER_23_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_179 ();
 FILLER_ASAP7_75t_R FILLER_23_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_202 ();
 DECAPx2_ASAP7_75t_R FILLER_23_214 ();
 DECAPx1_ASAP7_75t_R FILLER_23_242 ();
 DECAPx2_ASAP7_75t_R FILLER_23_269 ();
 FILLER_ASAP7_75t_R FILLER_23_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_277 ();
 FILLER_ASAP7_75t_R FILLER_23_304 ();
 FILLER_ASAP7_75t_R FILLER_23_312 ();
 DECAPx1_ASAP7_75t_R FILLER_24_2 ();
 DECAPx10_ASAP7_75t_R FILLER_24_68 ();
 DECAPx1_ASAP7_75t_R FILLER_24_90 ();
 FILLER_ASAP7_75t_R FILLER_24_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_106 ();
 DECAPx2_ASAP7_75t_R FILLER_24_117 ();
 FILLER_ASAP7_75t_R FILLER_24_123 ();
 DECAPx1_ASAP7_75t_R FILLER_24_131 ();
 DECAPx10_ASAP7_75t_R FILLER_24_155 ();
 DECAPx6_ASAP7_75t_R FILLER_24_177 ();
 DECAPx2_ASAP7_75t_R FILLER_24_191 ();
 DECAPx1_ASAP7_75t_R FILLER_24_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_245 ();
 DECAPx1_ASAP7_75t_R FILLER_24_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_263 ();
 DECAPx1_ASAP7_75t_R FILLER_24_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_8 ();
 FILLER_ASAP7_75t_R FILLER_25_21 ();
 DECAPx10_ASAP7_75t_R FILLER_25_41 ();
 DECAPx10_ASAP7_75t_R FILLER_25_69 ();
 DECAPx10_ASAP7_75t_R FILLER_25_91 ();
 DECAPx6_ASAP7_75t_R FILLER_25_113 ();
 DECAPx4_ASAP7_75t_R FILLER_25_141 ();
 FILLER_ASAP7_75t_R FILLER_25_151 ();
 DECAPx10_ASAP7_75t_R FILLER_25_156 ();
 DECAPx10_ASAP7_75t_R FILLER_25_196 ();
 FILLER_ASAP7_75t_R FILLER_25_218 ();
 DECAPx1_ASAP7_75t_R FILLER_25_237 ();
 DECAPx1_ASAP7_75t_R FILLER_25_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_295 ();
 FILLER_ASAP7_75t_R FILLER_26_2 ();
 DECAPx2_ASAP7_75t_R FILLER_26_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_22 ();
 DECAPx6_ASAP7_75t_R FILLER_26_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_55 ();
 FILLER_ASAP7_75t_R FILLER_26_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_72 ();
 FILLER_ASAP7_75t_R FILLER_26_92 ();
 FILLER_ASAP7_75t_R FILLER_26_100 ();
 DECAPx2_ASAP7_75t_R FILLER_26_117 ();
 FILLER_ASAP7_75t_R FILLER_26_123 ();
 FILLER_ASAP7_75t_R FILLER_26_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_133 ();
 DECAPx10_ASAP7_75t_R FILLER_26_172 ();
 DECAPx4_ASAP7_75t_R FILLER_26_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_204 ();
 DECAPx1_ASAP7_75t_R FILLER_26_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_217 ();
 DECAPx2_ASAP7_75t_R FILLER_26_234 ();
 DECAPx1_ASAP7_75t_R FILLER_26_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_280 ();
 FILLER_ASAP7_75t_R FILLER_26_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_301 ();
 DECAPx2_ASAP7_75t_R FILLER_26_308 ();
 DECAPx2_ASAP7_75t_R FILLER_27_2 ();
 DECAPx1_ASAP7_75t_R FILLER_27_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_38 ();
 FILLER_ASAP7_75t_R FILLER_27_76 ();
 DECAPx2_ASAP7_75t_R FILLER_27_121 ();
 FILLER_ASAP7_75t_R FILLER_27_127 ();
 DECAPx4_ASAP7_75t_R FILLER_27_137 ();
 DECAPx1_ASAP7_75t_R FILLER_27_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_161 ();
 DECAPx10_ASAP7_75t_R FILLER_27_172 ();
 DECAPx2_ASAP7_75t_R FILLER_27_194 ();
 FILLER_ASAP7_75t_R FILLER_27_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_202 ();
 FILLER_ASAP7_75t_R FILLER_27_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_225 ();
 DECAPx10_ASAP7_75t_R FILLER_27_252 ();
 DECAPx2_ASAP7_75t_R FILLER_27_274 ();
 FILLER_ASAP7_75t_R FILLER_27_280 ();
 DECAPx2_ASAP7_75t_R FILLER_27_308 ();
 DECAPx2_ASAP7_75t_R FILLER_28_2 ();
 DECAPx6_ASAP7_75t_R FILLER_28_29 ();
 DECAPx2_ASAP7_75t_R FILLER_28_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_72 ();
 DECAPx4_ASAP7_75t_R FILLER_28_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_109 ();
 DECAPx6_ASAP7_75t_R FILLER_28_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_127 ();
 DECAPx1_ASAP7_75t_R FILLER_28_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_155 ();
 DECAPx10_ASAP7_75t_R FILLER_28_174 ();
 DECAPx6_ASAP7_75t_R FILLER_28_196 ();
 DECAPx10_ASAP7_75t_R FILLER_28_216 ();
 DECAPx10_ASAP7_75t_R FILLER_28_238 ();
 DECAPx1_ASAP7_75t_R FILLER_28_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_264 ();
 DECAPx1_ASAP7_75t_R FILLER_28_268 ();
 DECAPx2_ASAP7_75t_R FILLER_28_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_284 ();
 DECAPx2_ASAP7_75t_R FILLER_28_291 ();
 FILLER_ASAP7_75t_R FILLER_28_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_305 ();
 FILLER_ASAP7_75t_R FILLER_28_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_2 ();
 FILLER_ASAP7_75t_R FILLER_29_35 ();
 DECAPx6_ASAP7_75t_R FILLER_29_40 ();
 DECAPx1_ASAP7_75t_R FILLER_29_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_66 ();
 DECAPx10_ASAP7_75t_R FILLER_29_73 ();
 DECAPx10_ASAP7_75t_R FILLER_29_105 ();
 DECAPx10_ASAP7_75t_R FILLER_29_127 ();
 FILLER_ASAP7_75t_R FILLER_29_149 ();
 DECAPx10_ASAP7_75t_R FILLER_29_154 ();
 DECAPx10_ASAP7_75t_R FILLER_29_176 ();
 DECAPx6_ASAP7_75t_R FILLER_29_198 ();
 DECAPx6_ASAP7_75t_R FILLER_29_218 ();
 FILLER_ASAP7_75t_R FILLER_29_232 ();
 DECAPx1_ASAP7_75t_R FILLER_29_240 ();
 DECAPx2_ASAP7_75t_R FILLER_29_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_253 ();
 DECAPx1_ASAP7_75t_R FILLER_29_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_273 ();
 DECAPx1_ASAP7_75t_R FILLER_29_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_298 ();
 DECAPx2_ASAP7_75t_R FILLER_30_23 ();
 DECAPx2_ASAP7_75t_R FILLER_30_43 ();
 FILLER_ASAP7_75t_R FILLER_30_49 ();
 DECAPx1_ASAP7_75t_R FILLER_30_68 ();
 DECAPx2_ASAP7_75t_R FILLER_30_82 ();
 FILLER_ASAP7_75t_R FILLER_30_88 ();
 FILLER_ASAP7_75t_R FILLER_30_112 ();
 DECAPx6_ASAP7_75t_R FILLER_30_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_131 ();
 FILLER_ASAP7_75t_R FILLER_30_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_148 ();
 DECAPx10_ASAP7_75t_R FILLER_30_156 ();
 DECAPx6_ASAP7_75t_R FILLER_30_178 ();
 FILLER_ASAP7_75t_R FILLER_30_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_204 ();
 DECAPx1_ASAP7_75t_R FILLER_30_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_229 ();
 FILLER_ASAP7_75t_R FILLER_30_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_252 ();
 DECAPx1_ASAP7_75t_R FILLER_30_276 ();
 DECAPx2_ASAP7_75t_R FILLER_30_300 ();
 FILLER_ASAP7_75t_R FILLER_30_312 ();
 DECAPx2_ASAP7_75t_R FILLER_31_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_26 ();
 DECAPx2_ASAP7_75t_R FILLER_31_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_49 ();
 DECAPx6_ASAP7_75t_R FILLER_31_70 ();
 FILLER_ASAP7_75t_R FILLER_31_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_86 ();
 DECAPx4_ASAP7_75t_R FILLER_31_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_139 ();
 DECAPx10_ASAP7_75t_R FILLER_31_160 ();
 DECAPx10_ASAP7_75t_R FILLER_31_182 ();
 DECAPx1_ASAP7_75t_R FILLER_31_204 ();
 DECAPx6_ASAP7_75t_R FILLER_31_216 ();
 FILLER_ASAP7_75t_R FILLER_31_230 ();
 DECAPx6_ASAP7_75t_R FILLER_31_240 ();
 DECAPx1_ASAP7_75t_R FILLER_31_254 ();
 DECAPx4_ASAP7_75t_R FILLER_31_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_293 ();
 DECAPx2_ASAP7_75t_R FILLER_31_300 ();
 FILLER_ASAP7_75t_R FILLER_31_306 ();
 FILLER_ASAP7_75t_R FILLER_32_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_10 ();
 FILLER_ASAP7_75t_R FILLER_32_34 ();
 DECAPx4_ASAP7_75t_R FILLER_32_59 ();
 DECAPx2_ASAP7_75t_R FILLER_32_79 ();
 FILLER_ASAP7_75t_R FILLER_32_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_110 ();
 DECAPx4_ASAP7_75t_R FILLER_32_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_127 ();
 DECAPx10_ASAP7_75t_R FILLER_32_148 ();
 DECAPx10_ASAP7_75t_R FILLER_32_170 ();
 DECAPx10_ASAP7_75t_R FILLER_32_202 ();
 DECAPx1_ASAP7_75t_R FILLER_32_224 ();
 DECAPx1_ASAP7_75t_R FILLER_32_256 ();
 DECAPx2_ASAP7_75t_R FILLER_32_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_272 ();
 FILLER_ASAP7_75t_R FILLER_33_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_22 ();
 DECAPx10_ASAP7_75t_R FILLER_33_32 ();
 FILLER_ASAP7_75t_R FILLER_33_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_56 ();
 DECAPx2_ASAP7_75t_R FILLER_33_67 ();
 FILLER_ASAP7_75t_R FILLER_33_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_75 ();
 DECAPx6_ASAP7_75t_R FILLER_33_102 ();
 FILLER_ASAP7_75t_R FILLER_33_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_121 ();
 FILLER_ASAP7_75t_R FILLER_33_128 ();
 DECAPx2_ASAP7_75t_R FILLER_33_138 ();
 FILLER_ASAP7_75t_R FILLER_33_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_146 ();
 DECAPx6_ASAP7_75t_R FILLER_33_150 ();
 DECAPx1_ASAP7_75t_R FILLER_33_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_179 ();
 DECAPx4_ASAP7_75t_R FILLER_33_190 ();
 FILLER_ASAP7_75t_R FILLER_33_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_202 ();
 DECAPx4_ASAP7_75t_R FILLER_33_217 ();
 DECAPx1_ASAP7_75t_R FILLER_33_230 ();
 DECAPx2_ASAP7_75t_R FILLER_33_244 ();
 FILLER_ASAP7_75t_R FILLER_33_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_252 ();
 DECAPx4_ASAP7_75t_R FILLER_33_278 ();
 FILLER_ASAP7_75t_R FILLER_33_288 ();
 DECAPx2_ASAP7_75t_R FILLER_33_308 ();
 DECAPx2_ASAP7_75t_R FILLER_34_14 ();
 FILLER_ASAP7_75t_R FILLER_34_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_22 ();
 DECAPx10_ASAP7_75t_R FILLER_34_39 ();
 FILLER_ASAP7_75t_R FILLER_34_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_63 ();
 DECAPx6_ASAP7_75t_R FILLER_34_74 ();
 DECAPx2_ASAP7_75t_R FILLER_34_88 ();
 DECAPx1_ASAP7_75t_R FILLER_34_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_124 ();
 DECAPx10_ASAP7_75t_R FILLER_34_145 ();
 FILLER_ASAP7_75t_R FILLER_34_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_209 ();
 DECAPx1_ASAP7_75t_R FILLER_34_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_236 ();
 FILLER_ASAP7_75t_R FILLER_34_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_249 ();
 DECAPx4_ASAP7_75t_R FILLER_34_270 ();
 FILLER_ASAP7_75t_R FILLER_34_280 ();
 DECAPx2_ASAP7_75t_R FILLER_35_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_20 ();
 FILLER_ASAP7_75t_R FILLER_35_55 ();
 DECAPx10_ASAP7_75t_R FILLER_35_81 ();
 DECAPx6_ASAP7_75t_R FILLER_35_103 ();
 FILLER_ASAP7_75t_R FILLER_35_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_126 ();
 DECAPx2_ASAP7_75t_R FILLER_35_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_141 ();
 DECAPx4_ASAP7_75t_R FILLER_35_145 ();
 FILLER_ASAP7_75t_R FILLER_35_155 ();
 DECAPx6_ASAP7_75t_R FILLER_35_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_181 ();
 DECAPx6_ASAP7_75t_R FILLER_35_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_206 ();
 DECAPx2_ASAP7_75t_R FILLER_35_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_234 ();
 DECAPx6_ASAP7_75t_R FILLER_35_245 ();
 FILLER_ASAP7_75t_R FILLER_35_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_269 ();
 DECAPx1_ASAP7_75t_R FILLER_35_273 ();
 FILLER_ASAP7_75t_R FILLER_35_306 ();
 DECAPx4_ASAP7_75t_R FILLER_36_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_28 ();
 FILLER_ASAP7_75t_R FILLER_36_72 ();
 FILLER_ASAP7_75t_R FILLER_36_84 ();
 DECAPx4_ASAP7_75t_R FILLER_36_92 ();
 DECAPx2_ASAP7_75t_R FILLER_36_120 ();
 FILLER_ASAP7_75t_R FILLER_36_126 ();
 DECAPx6_ASAP7_75t_R FILLER_36_138 ();
 DECAPx1_ASAP7_75t_R FILLER_36_152 ();
 DECAPx6_ASAP7_75t_R FILLER_36_166 ();
 FILLER_ASAP7_75t_R FILLER_36_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_182 ();
 DECAPx10_ASAP7_75t_R FILLER_36_193 ();
 DECAPx4_ASAP7_75t_R FILLER_36_215 ();
 DECAPx2_ASAP7_75t_R FILLER_36_252 ();
 FILLER_ASAP7_75t_R FILLER_36_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_260 ();
 DECAPx2_ASAP7_75t_R FILLER_36_276 ();
 FILLER_ASAP7_75t_R FILLER_36_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_284 ();
 DECAPx1_ASAP7_75t_R FILLER_36_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_2 ();
 DECAPx6_ASAP7_75t_R FILLER_37_9 ();
 FILLER_ASAP7_75t_R FILLER_37_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_25 ();
 DECAPx2_ASAP7_75t_R FILLER_37_32 ();
 FILLER_ASAP7_75t_R FILLER_37_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_40 ();
 DECAPx2_ASAP7_75t_R FILLER_37_44 ();
 FILLER_ASAP7_75t_R FILLER_37_50 ();
 DECAPx1_ASAP7_75t_R FILLER_37_69 ();
 DECAPx6_ASAP7_75t_R FILLER_37_83 ();
 DECAPx1_ASAP7_75t_R FILLER_37_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_101 ();
 DECAPx4_ASAP7_75t_R FILLER_37_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_118 ();
 DECAPx10_ASAP7_75t_R FILLER_37_155 ();
 DECAPx2_ASAP7_75t_R FILLER_37_177 ();
 FILLER_ASAP7_75t_R FILLER_37_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_185 ();
 DECAPx1_ASAP7_75t_R FILLER_37_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_200 ();
 FILLER_ASAP7_75t_R FILLER_37_224 ();
 FILLER_ASAP7_75t_R FILLER_37_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_262 ();
 DECAPx4_ASAP7_75t_R FILLER_37_286 ();
 FILLER_ASAP7_75t_R FILLER_37_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_304 ();
 DECAPx4_ASAP7_75t_R FILLER_38_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_25 ();
 DECAPx4_ASAP7_75t_R FILLER_38_34 ();
 FILLER_ASAP7_75t_R FILLER_38_44 ();
 DECAPx6_ASAP7_75t_R FILLER_38_68 ();
 FILLER_ASAP7_75t_R FILLER_38_82 ();
 DECAPx2_ASAP7_75t_R FILLER_38_91 ();
 FILLER_ASAP7_75t_R FILLER_38_97 ();
 DECAPx4_ASAP7_75t_R FILLER_38_130 ();
 FILLER_ASAP7_75t_R FILLER_38_140 ();
 DECAPx10_ASAP7_75t_R FILLER_38_145 ();
 DECAPx10_ASAP7_75t_R FILLER_38_167 ();
 DECAPx2_ASAP7_75t_R FILLER_38_189 ();
 DECAPx2_ASAP7_75t_R FILLER_38_203 ();
 FILLER_ASAP7_75t_R FILLER_38_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_211 ();
 DECAPx10_ASAP7_75t_R FILLER_38_232 ();
 DECAPx6_ASAP7_75t_R FILLER_38_254 ();
 DECAPx2_ASAP7_75t_R FILLER_38_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_274 ();
 DECAPx2_ASAP7_75t_R FILLER_38_306 ();
 FILLER_ASAP7_75t_R FILLER_38_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_2 ();
 DECAPx1_ASAP7_75t_R FILLER_39_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_33 ();
 FILLER_ASAP7_75t_R FILLER_39_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_59 ();
 FILLER_ASAP7_75t_R FILLER_39_63 ();
 FILLER_ASAP7_75t_R FILLER_39_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_83 ();
 FILLER_ASAP7_75t_R FILLER_39_107 ();
 DECAPx10_ASAP7_75t_R FILLER_39_149 ();
 DECAPx6_ASAP7_75t_R FILLER_39_171 ();
 FILLER_ASAP7_75t_R FILLER_39_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_202 ();
 DECAPx2_ASAP7_75t_R FILLER_39_212 ();
 DECAPx1_ASAP7_75t_R FILLER_39_242 ();
 DECAPx4_ASAP7_75t_R FILLER_39_252 ();
 FILLER_ASAP7_75t_R FILLER_39_262 ();
 DECAPx6_ASAP7_75t_R FILLER_39_279 ();
 FILLER_ASAP7_75t_R FILLER_39_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_295 ();
 DECAPx2_ASAP7_75t_R FILLER_40_2 ();
 FILLER_ASAP7_75t_R FILLER_40_23 ();
 DECAPx10_ASAP7_75t_R FILLER_40_37 ();
 FILLER_ASAP7_75t_R FILLER_40_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_61 ();
 DECAPx10_ASAP7_75t_R FILLER_40_65 ();
 DECAPx1_ASAP7_75t_R FILLER_40_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_123 ();
 DECAPx10_ASAP7_75t_R FILLER_40_132 ();
 DECAPx4_ASAP7_75t_R FILLER_40_154 ();
 DECAPx1_ASAP7_75t_R FILLER_40_174 ();
 DECAPx1_ASAP7_75t_R FILLER_40_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_192 ();
 DECAPx1_ASAP7_75t_R FILLER_40_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_238 ();
 FILLER_ASAP7_75t_R FILLER_40_259 ();
 FILLER_ASAP7_75t_R FILLER_40_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_276 ();
 DECAPx1_ASAP7_75t_R FILLER_40_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_284 ();
 DECAPx2_ASAP7_75t_R FILLER_40_288 ();
 FILLER_ASAP7_75t_R FILLER_40_294 ();
 DECAPx2_ASAP7_75t_R FILLER_40_302 ();
 FILLER_ASAP7_75t_R FILLER_41_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_4 ();
 DECAPx6_ASAP7_75t_R FILLER_41_11 ();
 FILLER_ASAP7_75t_R FILLER_41_25 ();
 DECAPx2_ASAP7_75t_R FILLER_41_35 ();
 FILLER_ASAP7_75t_R FILLER_41_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_43 ();
 DECAPx1_ASAP7_75t_R FILLER_41_52 ();
 FILLER_ASAP7_75t_R FILLER_41_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_72 ();
 DECAPx2_ASAP7_75t_R FILLER_41_79 ();
 FILLER_ASAP7_75t_R FILLER_41_85 ();
 DECAPx2_ASAP7_75t_R FILLER_41_109 ();
 DECAPx6_ASAP7_75t_R FILLER_41_144 ();
 DECAPx1_ASAP7_75t_R FILLER_41_158 ();
 DECAPx2_ASAP7_75t_R FILLER_41_182 ();
 DECAPx1_ASAP7_75t_R FILLER_41_206 ();
 DECAPx6_ASAP7_75t_R FILLER_41_248 ();
 DECAPx1_ASAP7_75t_R FILLER_41_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_266 ();
 FILLER_ASAP7_75t_R FILLER_41_287 ();
 DECAPx6_ASAP7_75t_R FILLER_41_295 ();
 DECAPx1_ASAP7_75t_R FILLER_41_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_2 ();
 FILLER_ASAP7_75t_R FILLER_42_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_38 ();
 DECAPx2_ASAP7_75t_R FILLER_42_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_68 ();
 DECAPx10_ASAP7_75t_R FILLER_42_112 ();
 DECAPx10_ASAP7_75t_R FILLER_42_134 ();
 DECAPx4_ASAP7_75t_R FILLER_42_156 ();
 FILLER_ASAP7_75t_R FILLER_42_166 ();
 FILLER_ASAP7_75t_R FILLER_42_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_184 ();
 DECAPx1_ASAP7_75t_R FILLER_42_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_203 ();
 DECAPx1_ASAP7_75t_R FILLER_42_224 ();
 DECAPx10_ASAP7_75t_R FILLER_42_234 ();
 DECAPx2_ASAP7_75t_R FILLER_42_256 ();
 FILLER_ASAP7_75t_R FILLER_42_262 ();
 DECAPx6_ASAP7_75t_R FILLER_42_271 ();
 DECAPx1_ASAP7_75t_R FILLER_42_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_289 ();
 DECAPx2_ASAP7_75t_R FILLER_42_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_299 ();
 DECAPx2_ASAP7_75t_R FILLER_42_306 ();
 FILLER_ASAP7_75t_R FILLER_42_312 ();
 DECAPx4_ASAP7_75t_R FILLER_43_8 ();
 FILLER_ASAP7_75t_R FILLER_43_18 ();
 FILLER_ASAP7_75t_R FILLER_43_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_28 ();
 DECAPx10_ASAP7_75t_R FILLER_43_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_57 ();
 DECAPx4_ASAP7_75t_R FILLER_43_72 ();
 FILLER_ASAP7_75t_R FILLER_43_82 ();
 DECAPx10_ASAP7_75t_R FILLER_43_137 ();
 DECAPx10_ASAP7_75t_R FILLER_43_159 ();
 DECAPx4_ASAP7_75t_R FILLER_43_181 ();
 FILLER_ASAP7_75t_R FILLER_43_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_193 ();
 DECAPx10_ASAP7_75t_R FILLER_43_213 ();
 DECAPx2_ASAP7_75t_R FILLER_43_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_241 ();
 DECAPx4_ASAP7_75t_R FILLER_43_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_262 ();
 FILLER_ASAP7_75t_R FILLER_43_292 ();
 DECAPx6_ASAP7_75t_R FILLER_43_300 ();
 FILLER_ASAP7_75t_R FILLER_44_8 ();
 FILLER_ASAP7_75t_R FILLER_44_38 ();
 DECAPx1_ASAP7_75t_R FILLER_44_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_81 ();
 DECAPx2_ASAP7_75t_R FILLER_44_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_121 ();
 DECAPx2_ASAP7_75t_R FILLER_44_130 ();
 FILLER_ASAP7_75t_R FILLER_44_136 ();
 DECAPx6_ASAP7_75t_R FILLER_44_144 ();
 DECAPx2_ASAP7_75t_R FILLER_44_158 ();
 DECAPx1_ASAP7_75t_R FILLER_44_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_178 ();
 DECAPx2_ASAP7_75t_R FILLER_44_193 ();
 FILLER_ASAP7_75t_R FILLER_44_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_238 ();
 FILLER_ASAP7_75t_R FILLER_44_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_249 ();
 DECAPx4_ASAP7_75t_R FILLER_44_256 ();
 FILLER_ASAP7_75t_R FILLER_44_266 ();
 DECAPx10_ASAP7_75t_R FILLER_44_280 ();
 DECAPx2_ASAP7_75t_R FILLER_44_302 ();
 FILLER_ASAP7_75t_R FILLER_45_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_16 ();
 DECAPx10_ASAP7_75t_R FILLER_45_32 ();
 DECAPx10_ASAP7_75t_R FILLER_45_54 ();
 DECAPx2_ASAP7_75t_R FILLER_45_76 ();
 DECAPx1_ASAP7_75t_R FILLER_45_92 ();
 DECAPx1_ASAP7_75t_R FILLER_45_102 ();
 FILLER_ASAP7_75t_R FILLER_45_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_122 ();
 DECAPx10_ASAP7_75t_R FILLER_45_129 ();
 DECAPx10_ASAP7_75t_R FILLER_45_151 ();
 DECAPx2_ASAP7_75t_R FILLER_45_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_241 ();
 FILLER_ASAP7_75t_R FILLER_45_268 ();
 DECAPx1_ASAP7_75t_R FILLER_45_273 ();
 FILLER_ASAP7_75t_R FILLER_45_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_287 ();
 FILLER_ASAP7_75t_R FILLER_45_294 ();
 FILLER_ASAP7_75t_R FILLER_45_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_301 ();
 DECAPx2_ASAP7_75t_R FILLER_45_308 ();
 DECAPx2_ASAP7_75t_R FILLER_46_2 ();
 FILLER_ASAP7_75t_R FILLER_46_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_10 ();
 DECAPx2_ASAP7_75t_R FILLER_46_17 ();
 FILLER_ASAP7_75t_R FILLER_46_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_25 ();
 DECAPx4_ASAP7_75t_R FILLER_46_35 ();
 FILLER_ASAP7_75t_R FILLER_46_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_47 ();
 DECAPx1_ASAP7_75t_R FILLER_46_51 ();
 DECAPx10_ASAP7_75t_R FILLER_46_72 ();
 DECAPx4_ASAP7_75t_R FILLER_46_94 ();
 FILLER_ASAP7_75t_R FILLER_46_104 ();
 DECAPx2_ASAP7_75t_R FILLER_46_114 ();
 FILLER_ASAP7_75t_R FILLER_46_120 ();
 DECAPx4_ASAP7_75t_R FILLER_46_130 ();
 FILLER_ASAP7_75t_R FILLER_46_140 ();
 DECAPx10_ASAP7_75t_R FILLER_46_145 ();
 DECAPx10_ASAP7_75t_R FILLER_46_167 ();
 FILLER_ASAP7_75t_R FILLER_46_189 ();
 DECAPx2_ASAP7_75t_R FILLER_46_211 ();
 FILLER_ASAP7_75t_R FILLER_46_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_222 ();
 FILLER_ASAP7_75t_R FILLER_46_226 ();
 DECAPx2_ASAP7_75t_R FILLER_46_238 ();
 FILLER_ASAP7_75t_R FILLER_46_244 ();
 DECAPx10_ASAP7_75t_R FILLER_46_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_277 ();
 DECAPx1_ASAP7_75t_R FILLER_46_310 ();
 FILLER_ASAP7_75t_R FILLER_47_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_4 ();
 FILLER_ASAP7_75t_R FILLER_47_39 ();
 FILLER_ASAP7_75t_R FILLER_47_94 ();
 DECAPx1_ASAP7_75t_R FILLER_47_103 ();
 DECAPx4_ASAP7_75t_R FILLER_47_114 ();
 DECAPx10_ASAP7_75t_R FILLER_47_144 ();
 DECAPx4_ASAP7_75t_R FILLER_47_166 ();
 FILLER_ASAP7_75t_R FILLER_47_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_178 ();
 DECAPx10_ASAP7_75t_R FILLER_47_207 ();
 DECAPx4_ASAP7_75t_R FILLER_47_229 ();
 FILLER_ASAP7_75t_R FILLER_47_239 ();
 DECAPx2_ASAP7_75t_R FILLER_47_271 ();
 DECAPx6_ASAP7_75t_R FILLER_47_283 ();
 DECAPx1_ASAP7_75t_R FILLER_47_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_2 ();
 DECAPx4_ASAP7_75t_R FILLER_48_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_26 ();
 DECAPx2_ASAP7_75t_R FILLER_48_33 ();
 FILLER_ASAP7_75t_R FILLER_48_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_62 ();
 FILLER_ASAP7_75t_R FILLER_48_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_68 ();
 DECAPx2_ASAP7_75t_R FILLER_48_75 ();
 FILLER_ASAP7_75t_R FILLER_48_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_118 ();
 DECAPx4_ASAP7_75t_R FILLER_48_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_155 ();
 DECAPx6_ASAP7_75t_R FILLER_48_179 ();
 FILLER_ASAP7_75t_R FILLER_48_193 ();
 DECAPx4_ASAP7_75t_R FILLER_48_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_219 ();
 DECAPx6_ASAP7_75t_R FILLER_48_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_248 ();
 DECAPx10_ASAP7_75t_R FILLER_48_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_277 ();
 DECAPx4_ASAP7_75t_R FILLER_48_286 ();
 FILLER_ASAP7_75t_R FILLER_48_296 ();
 DECAPx2_ASAP7_75t_R FILLER_48_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_2 ();
 DECAPx6_ASAP7_75t_R FILLER_49_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_51 ();
 FILLER_ASAP7_75t_R FILLER_49_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_79 ();
 FILLER_ASAP7_75t_R FILLER_49_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_101 ();
 FILLER_ASAP7_75t_R FILLER_49_125 ();
 DECAPx2_ASAP7_75t_R FILLER_49_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_141 ();
 DECAPx2_ASAP7_75t_R FILLER_49_145 ();
 FILLER_ASAP7_75t_R FILLER_49_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_153 ();
 DECAPx4_ASAP7_75t_R FILLER_49_182 ();
 FILLER_ASAP7_75t_R FILLER_49_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_226 ();
 DECAPx2_ASAP7_75t_R FILLER_49_237 ();
 DECAPx4_ASAP7_75t_R FILLER_49_246 ();
 FILLER_ASAP7_75t_R FILLER_49_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_261 ();
 DECAPx1_ASAP7_75t_R FILLER_49_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_279 ();
 DECAPx6_ASAP7_75t_R FILLER_49_300 ();
 DECAPx6_ASAP7_75t_R FILLER_50_2 ();
 DECAPx10_ASAP7_75t_R FILLER_50_22 ();
 DECAPx10_ASAP7_75t_R FILLER_50_44 ();
 DECAPx10_ASAP7_75t_R FILLER_50_66 ();
 DECAPx10_ASAP7_75t_R FILLER_50_88 ();
 DECAPx4_ASAP7_75t_R FILLER_50_110 ();
 FILLER_ASAP7_75t_R FILLER_50_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_122 ();
 DECAPx6_ASAP7_75t_R FILLER_50_129 ();
 FILLER_ASAP7_75t_R FILLER_50_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_165 ();
 DECAPx1_ASAP7_75t_R FILLER_50_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_173 ();
 FILLER_ASAP7_75t_R FILLER_50_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_179 ();
 DECAPx2_ASAP7_75t_R FILLER_50_192 ();
 FILLER_ASAP7_75t_R FILLER_50_198 ();
 DECAPx4_ASAP7_75t_R FILLER_50_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_236 ();
 DECAPx4_ASAP7_75t_R FILLER_50_251 ();
 FILLER_ASAP7_75t_R FILLER_50_261 ();
 DECAPx6_ASAP7_75t_R FILLER_50_272 ();
 DECAPx10_ASAP7_75t_R FILLER_50_289 ();
 FILLER_ASAP7_75t_R FILLER_50_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_313 ();
 DECAPx1_ASAP7_75t_R FILLER_51_2 ();
 DECAPx1_ASAP7_75t_R FILLER_51_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_19 ();
 DECAPx1_ASAP7_75t_R FILLER_51_23 ();
 DECAPx4_ASAP7_75t_R FILLER_51_33 ();
 FILLER_ASAP7_75t_R FILLER_51_63 ();
 DECAPx4_ASAP7_75t_R FILLER_51_68 ();
 FILLER_ASAP7_75t_R FILLER_51_78 ();
 FILLER_ASAP7_75t_R FILLER_51_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_92 ();
 DECAPx4_ASAP7_75t_R FILLER_51_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_119 ();
 DECAPx4_ASAP7_75t_R FILLER_51_143 ();
 DECAPx10_ASAP7_75t_R FILLER_51_161 ();
 FILLER_ASAP7_75t_R FILLER_51_183 ();
 FILLER_ASAP7_75t_R FILLER_51_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_197 ();
 DECAPx10_ASAP7_75t_R FILLER_51_208 ();
 FILLER_ASAP7_75t_R FILLER_51_230 ();
 DECAPx4_ASAP7_75t_R FILLER_51_258 ();
 DECAPx10_ASAP7_75t_R FILLER_51_288 ();
 DECAPx1_ASAP7_75t_R FILLER_51_310 ();
 FILLER_ASAP7_75t_R FILLER_52_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_4 ();
 DECAPx1_ASAP7_75t_R FILLER_52_39 ();
 DECAPx2_ASAP7_75t_R FILLER_52_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_72 ();
 DECAPx1_ASAP7_75t_R FILLER_52_89 ();
 DECAPx2_ASAP7_75t_R FILLER_52_116 ();
 DECAPx10_ASAP7_75t_R FILLER_52_130 ();
 DECAPx2_ASAP7_75t_R FILLER_52_152 ();
 FILLER_ASAP7_75t_R FILLER_52_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_186 ();
 FILLER_ASAP7_75t_R FILLER_52_197 ();
 DECAPx2_ASAP7_75t_R FILLER_52_229 ();
 FILLER_ASAP7_75t_R FILLER_52_235 ();
 DECAPx10_ASAP7_75t_R FILLER_52_265 ();
 DECAPx10_ASAP7_75t_R FILLER_52_287 ();
 DECAPx1_ASAP7_75t_R FILLER_52_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_313 ();
 DECAPx10_ASAP7_75t_R FILLER_53_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_24 ();
 DECAPx10_ASAP7_75t_R FILLER_53_31 ();
 DECAPx4_ASAP7_75t_R FILLER_53_53 ();
 DECAPx2_ASAP7_75t_R FILLER_53_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_94 ();
 DECAPx6_ASAP7_75t_R FILLER_53_101 ();
 DECAPx1_ASAP7_75t_R FILLER_53_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_119 ();
 DECAPx6_ASAP7_75t_R FILLER_53_126 ();
 DECAPx2_ASAP7_75t_R FILLER_53_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_146 ();
 DECAPx2_ASAP7_75t_R FILLER_53_167 ();
 DECAPx10_ASAP7_75t_R FILLER_53_176 ();
 FILLER_ASAP7_75t_R FILLER_53_198 ();
 DECAPx6_ASAP7_75t_R FILLER_53_216 ();
 FILLER_ASAP7_75t_R FILLER_53_230 ();
 DECAPx2_ASAP7_75t_R FILLER_53_248 ();
 DECAPx10_ASAP7_75t_R FILLER_53_257 ();
 DECAPx10_ASAP7_75t_R FILLER_53_279 ();
 DECAPx4_ASAP7_75t_R FILLER_53_301 ();
 FILLER_ASAP7_75t_R FILLER_53_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_313 ();
 DECAPx10_ASAP7_75t_R FILLER_54_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_24 ();
 DECAPx6_ASAP7_75t_R FILLER_54_41 ();
 FILLER_ASAP7_75t_R FILLER_54_55 ();
 DECAPx2_ASAP7_75t_R FILLER_54_65 ();
 DECAPx6_ASAP7_75t_R FILLER_54_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_99 ();
 DECAPx2_ASAP7_75t_R FILLER_54_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_120 ();
 DECAPx10_ASAP7_75t_R FILLER_54_124 ();
 DECAPx2_ASAP7_75t_R FILLER_54_146 ();
 DECAPx6_ASAP7_75t_R FILLER_54_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_194 ();
 DECAPx2_ASAP7_75t_R FILLER_54_204 ();
 DECAPx4_ASAP7_75t_R FILLER_54_222 ();
 DECAPx10_ASAP7_75t_R FILLER_54_255 ();
 DECAPx10_ASAP7_75t_R FILLER_54_277 ();
 DECAPx6_ASAP7_75t_R FILLER_54_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_313 ();
 DECAPx2_ASAP7_75t_R FILLER_55_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_8 ();
 DECAPx2_ASAP7_75t_R FILLER_55_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_35 ();
 DECAPx4_ASAP7_75t_R FILLER_55_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_69 ();
 FILLER_ASAP7_75t_R FILLER_55_84 ();
 DECAPx2_ASAP7_75t_R FILLER_55_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_101 ();
 FILLER_ASAP7_75t_R FILLER_55_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_134 ();
 DECAPx6_ASAP7_75t_R FILLER_55_143 ();
 DECAPx4_ASAP7_75t_R FILLER_55_163 ();
 FILLER_ASAP7_75t_R FILLER_55_173 ();
 DECAPx2_ASAP7_75t_R FILLER_55_226 ();
 FILLER_ASAP7_75t_R FILLER_55_238 ();
 FILLER_ASAP7_75t_R FILLER_55_246 ();
 DECAPx1_ASAP7_75t_R FILLER_55_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_260 ();
 DECAPx10_ASAP7_75t_R FILLER_55_264 ();
 DECAPx10_ASAP7_75t_R FILLER_55_286 ();
 DECAPx2_ASAP7_75t_R FILLER_55_308 ();
 DECAPx6_ASAP7_75t_R FILLER_56_2 ();
 DECAPx2_ASAP7_75t_R FILLER_56_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_22 ();
 DECAPx6_ASAP7_75t_R FILLER_56_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_123 ();
 DECAPx6_ASAP7_75t_R FILLER_56_147 ();
 DECAPx1_ASAP7_75t_R FILLER_56_161 ();
 DECAPx10_ASAP7_75t_R FILLER_56_168 ();
 DECAPx1_ASAP7_75t_R FILLER_56_190 ();
 FILLER_ASAP7_75t_R FILLER_56_214 ();
 DECAPx4_ASAP7_75t_R FILLER_56_239 ();
 DECAPx10_ASAP7_75t_R FILLER_56_269 ();
 DECAPx10_ASAP7_75t_R FILLER_56_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_313 ();
 DECAPx10_ASAP7_75t_R FILLER_57_2 ();
 DECAPx6_ASAP7_75t_R FILLER_57_24 ();
 DECAPx10_ASAP7_75t_R FILLER_57_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_63 ();
 DECAPx4_ASAP7_75t_R FILLER_57_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_80 ();
 DECAPx2_ASAP7_75t_R FILLER_57_104 ();
 DECAPx1_ASAP7_75t_R FILLER_57_116 ();
 DECAPx2_ASAP7_75t_R FILLER_57_126 ();
 DECAPx10_ASAP7_75t_R FILLER_57_161 ();
 DECAPx10_ASAP7_75t_R FILLER_57_183 ();
 DECAPx2_ASAP7_75t_R FILLER_57_205 ();
 DECAPx10_ASAP7_75t_R FILLER_57_214 ();
 DECAPx10_ASAP7_75t_R FILLER_57_236 ();
 DECAPx10_ASAP7_75t_R FILLER_57_258 ();
 DECAPx10_ASAP7_75t_R FILLER_57_280 ();
 DECAPx4_ASAP7_75t_R FILLER_57_302 ();
 FILLER_ASAP7_75t_R FILLER_57_312 ();
 DECAPx10_ASAP7_75t_R FILLER_58_2 ();
 DECAPx10_ASAP7_75t_R FILLER_58_24 ();
 DECAPx10_ASAP7_75t_R FILLER_58_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_68 ();
 FILLER_ASAP7_75t_R FILLER_58_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_77 ();
 FILLER_ASAP7_75t_R FILLER_58_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_92 ();
 DECAPx6_ASAP7_75t_R FILLER_58_99 ();
 FILLER_ASAP7_75t_R FILLER_58_119 ();
 DECAPx1_ASAP7_75t_R FILLER_58_127 ();
 DECAPx2_ASAP7_75t_R FILLER_58_137 ();
 FILLER_ASAP7_75t_R FILLER_58_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_145 ();
 FILLER_ASAP7_75t_R FILLER_58_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_154 ();
 DECAPx6_ASAP7_75t_R FILLER_58_161 ();
 DECAPx2_ASAP7_75t_R FILLER_58_175 ();
 DECAPx6_ASAP7_75t_R FILLER_58_187 ();
 DECAPx2_ASAP7_75t_R FILLER_58_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_207 ();
 DECAPx4_ASAP7_75t_R FILLER_58_214 ();
 FILLER_ASAP7_75t_R FILLER_58_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_226 ();
 DECAPx10_ASAP7_75t_R FILLER_58_233 ();
 DECAPx10_ASAP7_75t_R FILLER_58_255 ();
 DECAPx10_ASAP7_75t_R FILLER_58_277 ();
 DECAPx6_ASAP7_75t_R FILLER_58_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_313 ();
 DECAPx10_ASAP7_75t_R FILLER_59_2 ();
 FILLER_ASAP7_75t_R FILLER_59_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_26 ();
 DECAPx10_ASAP7_75t_R FILLER_59_33 ();
 DECAPx10_ASAP7_75t_R FILLER_59_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_84 ();
 DECAPx10_ASAP7_75t_R FILLER_59_91 ();
 FILLER_ASAP7_75t_R FILLER_59_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_127 ();
 FILLER_ASAP7_75t_R FILLER_59_134 ();
 DECAPx1_ASAP7_75t_R FILLER_59_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_158 ();
 FILLER_ASAP7_75t_R FILLER_59_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_167 ();
 FILLER_ASAP7_75t_R FILLER_59_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_182 ();
 DECAPx2_ASAP7_75t_R FILLER_59_189 ();
 FILLER_ASAP7_75t_R FILLER_59_195 ();
 DECAPx1_ASAP7_75t_R FILLER_59_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_207 ();
 DECAPx4_ASAP7_75t_R FILLER_59_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_224 ();
 DECAPx10_ASAP7_75t_R FILLER_59_237 ();
 DECAPx10_ASAP7_75t_R FILLER_59_259 ();
 DECAPx10_ASAP7_75t_R FILLER_59_281 ();
 DECAPx4_ASAP7_75t_R FILLER_59_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_313 ();
 DECAPx6_ASAP7_75t_R FILLER_60_2 ();
 FILLER_ASAP7_75t_R FILLER_60_16 ();
 DECAPx10_ASAP7_75t_R FILLER_60_24 ();
 DECAPx6_ASAP7_75t_R FILLER_60_46 ();
 DECAPx2_ASAP7_75t_R FILLER_60_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_91 ();
 DECAPx1_ASAP7_75t_R FILLER_60_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_133 ();
 DECAPx1_ASAP7_75t_R FILLER_60_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_180 ();
 DECAPx2_ASAP7_75t_R FILLER_60_217 ();
 DECAPx2_ASAP7_75t_R FILLER_60_229 ();
 DECAPx10_ASAP7_75t_R FILLER_60_253 ();
 DECAPx10_ASAP7_75t_R FILLER_60_275 ();
 DECAPx6_ASAP7_75t_R FILLER_60_297 ();
 FILLER_ASAP7_75t_R FILLER_60_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_313 ();
 DECAPx4_ASAP7_75t_R FILLER_61_2 ();
 FILLER_ASAP7_75t_R FILLER_61_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_14 ();
 DECAPx4_ASAP7_75t_R FILLER_61_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_37 ();
 DECAPx10_ASAP7_75t_R FILLER_61_44 ();
 FILLER_ASAP7_75t_R FILLER_61_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_153 ();
 FILLER_ASAP7_75t_R FILLER_61_160 ();
 FILLER_ASAP7_75t_R FILLER_61_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_213 ();
 FILLER_ASAP7_75t_R FILLER_61_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_228 ();
 FILLER_ASAP7_75t_R FILLER_61_235 ();
 DECAPx2_ASAP7_75t_R FILLER_61_249 ();
 DECAPx10_ASAP7_75t_R FILLER_61_261 ();
 DECAPx4_ASAP7_75t_R FILLER_61_289 ();
 DECAPx2_ASAP7_75t_R FILLER_61_305 ();
 FILLER_ASAP7_75t_R FILLER_61_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_313 ();
endmodule
