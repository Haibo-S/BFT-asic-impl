module credit_t_switch (clk,
    rst,
    l_i,
    l_i_bp,
    l_i_v,
    l_o,
    l_o_credit_gnt,
    l_o_v,
    r_i,
    r_i_bp,
    r_i_v,
    r_o,
    r_o_credit_gnt,
    r_o_v,
    u0_i,
    u0_i_bp,
    u0_i_v,
    u0_o,
    u0_o_credit_gnt,
    u0_o_v);
 input clk;
 input rst;
 input [73:0] l_i;
 output [1:0] l_i_bp;
 input [1:0] l_i_v;
 output [36:0] l_o;
 input [1:0] l_o_credit_gnt;
 output [1:0] l_o_v;
 input [73:0] r_i;
 output [1:0] r_i_bp;
 input [1:0] r_i_v;
 output [36:0] r_o;
 input [1:0] r_o_credit_gnt;
 output [1:0] r_o_v;
 input [73:0] u0_i;
 output [1:0] u0_i_bp;
 input [1:0] u0_i_v;
 output [36:0] u0_o;
 input [1:0] u0_o_credit_gnt;
 output [1:0] u0_o_v;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire \credit_t_route_inst.l_counters_inst.o_credits[1] ;
 wire \credit_t_route_inst.l_counters_inst.o_credits[2] ;
 wire \credit_t_route_inst.l_counters_inst.o_credits[3] ;
 wire \credit_t_route_inst.l_counters_inst.o_credits[6] ;
 wire \credit_t_route_inst.l_counters_inst.o_credits[7] ;
 wire \credit_t_route_inst.l_counters_inst.o_credits[8] ;
 wire \credit_t_route_inst.r_counters_inst.o_credits[1] ;
 wire \credit_t_route_inst.r_counters_inst.o_credits[2] ;
 wire \credit_t_route_inst.r_counters_inst.o_credits[3] ;
 wire \credit_t_route_inst.r_counters_inst.o_credits[6] ;
 wire \credit_t_route_inst.r_counters_inst.o_credits[7] ;
 wire \credit_t_route_inst.r_counters_inst.o_credits[8] ;
 wire \credit_t_route_inst.u0_counters_inst.o_credits[1] ;
 wire \credit_t_route_inst.u0_counters_inst.o_credits[2] ;
 wire \credit_t_route_inst.u0_counters_inst.o_credits[3] ;
 wire \credit_t_route_inst.u0_counters_inst.o_credits[6] ;
 wire \credit_t_route_inst.u0_counters_inst.o_credits[7] ;
 wire \credit_t_route_inst.u0_counters_inst.o_credits[8] ;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 OA21x2_ASAP7_75t_R _0709_ (.A1(_0358_),
    .A2(_0359_),
    .B(_0360_),
    .Y(_0361_));
 INVx1_ASAP7_75t_R _0710_ (.A(net153),
    .Y(_0362_));
 NOR3x1_ASAP7_75t_R _0711_ (.A(net106),
    .B(net105),
    .C(net107),
    .Y(_0363_));
 NOR3x1_ASAP7_75t_R _0712_ (.A(_0362_),
    .B(_0363_),
    .C(_0353_),
    .Y(_0364_));
 OR5x2_ASAP7_75t_R _0713_ (.A(_0356_),
    .B(_0345_),
    .C(_0357_),
    .D(_0361_),
    .E(_0364_),
    .Y(_0365_));
 OAI21x1_ASAP7_75t_R _0714_ (.A1(_0350_),
    .A2(_0355_),
    .B(_0365_),
    .Y(_0366_));
 BUFx6f_ASAP7_75t_R _0715_ (.A(_0366_),
    .Y(_0367_));
 BUFx6f_ASAP7_75t_R _0716_ (.A(_0367_),
    .Y(net358));
 INVx1_ASAP7_75t_R _0717_ (.A(net358),
    .Y(_0702_));
 AND2x2_ASAP7_75t_R _0718_ (.A(_0021_),
    .B(net154),
    .Y(_0368_));
 AOI22x1_ASAP7_75t_R _0719_ (.A1(_0346_),
    .A2(_0368_),
    .B1(_0347_),
    .B2(_0348_),
    .Y(_0369_));
 OAI21x1_ASAP7_75t_R _0720_ (.A1(_0358_),
    .A2(_0359_),
    .B(_0360_),
    .Y(_0370_));
 AO22x2_ASAP7_75t_R _0721_ (.A1(_0369_),
    .A2(_0355_),
    .B1(_0370_),
    .B2(_0364_),
    .Y(net357));
 INVx2_ASAP7_75t_R _0722_ (.A(net357),
    .Y(_0708_));
 INVx1_ASAP7_75t_R _0723_ (.A(_0699_),
    .Y(\credit_t_route_inst.l_counters_inst.o_credits[1] ));
 INVx1_ASAP7_75t_R _0724_ (.A(_0069_),
    .Y(\credit_t_route_inst.l_counters_inst.o_credits[3] ));
 INVx1_ASAP7_75t_R _0725_ (.A(_0070_),
    .Y(\credit_t_route_inst.l_counters_inst.o_credits[2] ));
 INVx1_ASAP7_75t_R _0726_ (.A(_0697_),
    .Y(\credit_t_route_inst.l_counters_inst.o_credits[6] ));
 INVx1_ASAP7_75t_R _0727_ (.A(_0066_),
    .Y(\credit_t_route_inst.l_counters_inst.o_credits[8] ));
 INVx1_ASAP7_75t_R _0728_ (.A(_0067_),
    .Y(\credit_t_route_inst.l_counters_inst.o_credits[7] ));
 OR3x1_ASAP7_75t_R _0729_ (.A(_0345_),
    .B(_0361_),
    .C(_0364_),
    .Y(_0371_));
 INVx1_ASAP7_75t_R _0730_ (.A(net144),
    .Y(_0372_));
 AND3x4_ASAP7_75t_R _0731_ (.A(net154),
    .B(_0372_),
    .C(_0357_),
    .Y(_0373_));
 AND5x2_ASAP7_75t_R _0732_ (.A(_0068_),
    .B(_0069_),
    .C(_0070_),
    .D(_0699_),
    .E(_0042_),
    .Y(_0374_));
 INVx2_ASAP7_75t_R _0733_ (.A(_0374_),
    .Y(_0375_));
 INVx1_ASAP7_75t_R _0734_ (.A(net104),
    .Y(_0376_));
 AND3x1_ASAP7_75t_R _0735_ (.A(net153),
    .B(_0376_),
    .C(_0363_),
    .Y(_0377_));
 INVx2_ASAP7_75t_R _0736_ (.A(net183),
    .Y(_0378_));
 INVx1_ASAP7_75t_R _0737_ (.A(net223),
    .Y(_0379_));
 AO22x2_ASAP7_75t_R _0738_ (.A1(net232),
    .A2(_0378_),
    .B1(net233),
    .B2(_0379_),
    .Y(_0380_));
 AND5x2_ASAP7_75t_R _0739_ (.A(_0065_),
    .B(_0066_),
    .C(_0067_),
    .D(_0697_),
    .E(_0044_),
    .Y(_0381_));
 AO221x1_ASAP7_75t_R _0740_ (.A1(_0375_),
    .A2(_0377_),
    .B1(_0380_),
    .B2(_0360_),
    .C(_0381_),
    .Y(_0382_));
 AO32x1_ASAP7_75t_R _0741_ (.A1(net154),
    .A2(_0346_),
    .A3(_0371_),
    .B1(_0373_),
    .B2(_0382_),
    .Y(_0383_));
 BUFx3_ASAP7_75t_R _0742_ (.A(_0383_),
    .Y(net278));
 AO21x1_ASAP7_75t_R _0743_ (.A1(_0360_),
    .A2(_0380_),
    .B(_0374_),
    .Y(_0384_));
 OA211x2_ASAP7_75t_R _0744_ (.A1(_0353_),
    .A2(_0361_),
    .B(net153),
    .C(_0347_),
    .Y(_0385_));
 AO21x2_ASAP7_75t_R _0745_ (.A1(_0377_),
    .A2(_0384_),
    .B(_0385_),
    .Y(net277));
 OR3x1_ASAP7_75t_R _0746_ (.A(_0345_),
    .B(_0349_),
    .C(_0355_),
    .Y(_0386_));
 AND2x4_ASAP7_75t_R _0747_ (.A(_0021_),
    .B(_0323_),
    .Y(_0387_));
 NOR3x1_ASAP7_75t_R _0748_ (.A(_0331_),
    .B(_0320_),
    .C(_0321_),
    .Y(_0388_));
 OR3x1_ASAP7_75t_R _0749_ (.A(_0387_),
    .B(_0334_),
    .C(_0388_),
    .Y(_0389_));
 AO32x2_ASAP7_75t_R _0750_ (.A1(net76),
    .A2(_0327_),
    .A3(_0386_),
    .B1(_0389_),
    .B2(_0333_),
    .Y(net237));
 OR2x2_ASAP7_75t_R _0751_ (.A(_0349_),
    .B(_0353_),
    .Y(_0390_));
 OA21x2_ASAP7_75t_R _0752_ (.A1(_0331_),
    .A2(_0387_),
    .B(_0322_),
    .Y(_0391_));
 AO21x1_ASAP7_75t_R _0753_ (.A1(_0359_),
    .A2(_0390_),
    .B(_0391_),
    .Y(net236));
 INVx1_ASAP7_75t_R _0754_ (.A(net233),
    .Y(_0392_));
 OA21x2_ASAP7_75t_R _0755_ (.A1(_0326_),
    .A2(_0329_),
    .B(_0341_),
    .Y(_0393_));
 AND2x2_ASAP7_75t_R _0756_ (.A(net232),
    .B(_0378_),
    .Y(_0394_));
 AO33x2_ASAP7_75t_R _0757_ (.A1(net154),
    .A2(_0372_),
    .A3(_0357_),
    .B1(_0363_),
    .B2(_0376_),
    .B3(net153),
    .Y(_0395_));
 OR2x2_ASAP7_75t_R _0758_ (.A(net223),
    .B(_0381_),
    .Y(_0396_));
 AOI221x1_ASAP7_75t_R _0759_ (.A1(_0375_),
    .A2(_0394_),
    .B1(_0395_),
    .B2(_0022_),
    .C(_0396_),
    .Y(_0397_));
 NOR3x1_ASAP7_75t_R _0760_ (.A(_0392_),
    .B(_0393_),
    .C(_0397_),
    .Y(net319));
 OR2x2_ASAP7_75t_R _0761_ (.A(net183),
    .B(_0374_),
    .Y(_0398_));
 AO21x1_ASAP7_75t_R _0762_ (.A1(_0022_),
    .A2(_0395_),
    .B(_0398_),
    .Y(_0399_));
 NOR2x1_ASAP7_75t_R _0763_ (.A(_0378_),
    .B(_0331_),
    .Y(_0400_));
 OAI21x1_ASAP7_75t_R _0764_ (.A1(_0326_),
    .A2(_0329_),
    .B(_0400_),
    .Y(_0401_));
 AND3x4_ASAP7_75t_R _0765_ (.A(net232),
    .B(_0399_),
    .C(_0401_),
    .Y(net318));
 INVx1_ASAP7_75t_R _0766_ (.A(_0021_),
    .Y(_0402_));
 INVx2_ASAP7_75t_R _0767_ (.A(net157),
    .Y(_0403_));
 BUFx12f_ASAP7_75t_R _0768_ (.A(_0403_),
    .Y(_0404_));
 OR2x2_ASAP7_75t_R _0769_ (.A(net278),
    .B(net277),
    .Y(_0405_));
 OR2x6_ASAP7_75t_R _0770_ (.A(net319),
    .B(net318),
    .Y(_0406_));
 NOR2x1_ASAP7_75t_R _0771_ (.A(net278),
    .B(net277),
    .Y(_0407_));
 OAI22x1_ASAP7_75t_R _0772_ (.A1(_0360_),
    .A2(_0406_),
    .B1(_0407_),
    .B2(_0022_),
    .Y(_0408_));
 OR2x6_ASAP7_75t_R _0773_ (.A(net237),
    .B(net236),
    .Y(_0409_));
 NOR2x1_ASAP7_75t_R _0774_ (.A(net157),
    .B(_0409_),
    .Y(_0410_));
 AO32x1_ASAP7_75t_R _0775_ (.A1(_0402_),
    .A2(_0404_),
    .A3(_0405_),
    .B1(_0408_),
    .B2(_0410_),
    .Y(_0002_));
 INVx1_ASAP7_75t_R _0776_ (.A(_0360_),
    .Y(_0411_));
 AO21x1_ASAP7_75t_R _0777_ (.A1(_0402_),
    .A2(_0407_),
    .B(_0411_),
    .Y(_0412_));
 AO33x2_ASAP7_75t_R _0778_ (.A1(_0326_),
    .A2(_0410_),
    .A3(_0407_),
    .B1(_0412_),
    .B2(_0406_),
    .B3(_0403_),
    .Y(_0001_));
 OR3x1_ASAP7_75t_R _0779_ (.A(_0362_),
    .B(net104),
    .C(_0347_),
    .Y(_0413_));
 AO21x2_ASAP7_75t_R _0780_ (.A1(_0360_),
    .A2(_0380_),
    .B(_0413_),
    .Y(_0414_));
 NAND2x1_ASAP7_75t_R _0781_ (.A(net232),
    .B(_0378_),
    .Y(_0415_));
 AO21x1_ASAP7_75t_R _0782_ (.A1(_0022_),
    .A2(_0395_),
    .B(_0415_),
    .Y(_0416_));
 AO21x1_ASAP7_75t_R _0783_ (.A1(_0414_),
    .A2(_0416_),
    .B(_0374_),
    .Y(_0417_));
 BUFx3_ASAP7_75t_R _0784_ (.A(_0417_),
    .Y(_0700_));
 AOI221x1_ASAP7_75t_R _0785_ (.A1(_0375_),
    .A2(_0377_),
    .B1(_0380_),
    .B2(_0360_),
    .C(_0381_),
    .Y(_0418_));
 AO22x1_ASAP7_75t_R _0786_ (.A1(_0373_),
    .A2(_0418_),
    .B1(_0397_),
    .B2(net233),
    .Y(_0419_));
 BUFx6f_ASAP7_75t_R _0787_ (.A(_0419_),
    .Y(net276));
 INVx3_ASAP7_75t_R _0788_ (.A(net276),
    .Y(_0698_));
 INVx1_ASAP7_75t_R _0789_ (.A(_0406_),
    .Y(_0420_));
 AO22x1_ASAP7_75t_R _0790_ (.A1(_0411_),
    .A2(_0409_),
    .B1(_0407_),
    .B2(_0402_),
    .Y(_0421_));
 BUFx6f_ASAP7_75t_R _0791_ (.A(net157),
    .Y(_0422_));
 AO221x1_ASAP7_75t_R _0792_ (.A1(_0326_),
    .A2(_0409_),
    .B1(_0420_),
    .B2(_0421_),
    .C(_0422_),
    .Y(_0000_));
 INVx2_ASAP7_75t_R _0793_ (.A(_0700_),
    .Y(net275));
 INVx2_ASAP7_75t_R _0794_ (.A(_0706_),
    .Y(net316));
 INVx1_ASAP7_75t_R _0795_ (.A(net77),
    .Y(_0423_));
 XNOR2x1_ASAP7_75t_R _0796_ (.B(_0700_),
    .Y(_0424_),
    .A(_0423_));
 XNOR2x2_ASAP7_75t_R _0797_ (.A(_0042_),
    .B(_0424_),
    .Y(_0425_));
 NAND2x1_ASAP7_75t_R _0798_ (.A(_0404_),
    .B(_0425_),
    .Y(_0078_));
 NAND2x1_ASAP7_75t_R _0799_ (.A(_0699_),
    .B(_0424_),
    .Y(_0426_));
 OR2x2_ASAP7_75t_R _0800_ (.A(_0043_),
    .B(_0424_),
    .Y(_0427_));
 AO21x1_ASAP7_75t_R _0801_ (.A1(_0426_),
    .A2(_0427_),
    .B(_0422_),
    .Y(_0079_));
 BUFx6f_ASAP7_75t_R _0802_ (.A(net157),
    .Y(_0428_));
 AND2x2_ASAP7_75t_R _0803_ (.A(\credit_t_route_inst.l_counters_inst.o_credits[2] ),
    .B(_0424_),
    .Y(_0429_));
 XOR2x2_ASAP7_75t_R _0804_ (.A(_0033_),
    .B(_0031_),
    .Y(_0430_));
 NOR2x1_ASAP7_75t_R _0805_ (.A(_0424_),
    .B(_0430_),
    .Y(_0431_));
 OR3x1_ASAP7_75t_R _0806_ (.A(_0428_),
    .B(_0429_),
    .C(_0431_),
    .Y(_0080_));
 NAND2x1_ASAP7_75t_R _0807_ (.A(_0069_),
    .B(_0424_),
    .Y(_0432_));
 OA21x2_ASAP7_75t_R _0808_ (.A1(_0030_),
    .A2(_0042_),
    .B(_0032_),
    .Y(_0433_));
 OA21x2_ASAP7_75t_R _0809_ (.A1(_0031_),
    .A2(_0433_),
    .B(_0035_),
    .Y(_0434_));
 XOR2x2_ASAP7_75t_R _0810_ (.A(_0034_),
    .B(_0434_),
    .Y(_0435_));
 OR2x2_ASAP7_75t_R _0811_ (.A(_0424_),
    .B(_0435_),
    .Y(_0436_));
 AO21x1_ASAP7_75t_R _0812_ (.A1(_0432_),
    .A2(_0436_),
    .B(_0422_),
    .Y(_0081_));
 INVx1_ASAP7_75t_R _0813_ (.A(_0033_),
    .Y(_0437_));
 OA21x2_ASAP7_75t_R _0814_ (.A1(_0437_),
    .A2(_0031_),
    .B(_0035_),
    .Y(_0438_));
 OAI21x1_ASAP7_75t_R _0815_ (.A1(_0034_),
    .A2(_0438_),
    .B(_0073_),
    .Y(_0439_));
 AOI211x1_ASAP7_75t_R _0816_ (.A1(_0414_),
    .A2(_0416_),
    .B(_0439_),
    .C(_0374_),
    .Y(_0440_));
 AND2x2_ASAP7_75t_R _0817_ (.A(net77),
    .B(_0439_),
    .Y(_0441_));
 AO22x1_ASAP7_75t_R _0818_ (.A1(_0423_),
    .A2(_0440_),
    .B1(_0441_),
    .B2(_0700_),
    .Y(_0442_));
 XOR2x2_ASAP7_75t_R _0819_ (.A(_0068_),
    .B(_0442_),
    .Y(_0443_));
 NAND2x1_ASAP7_75t_R _0820_ (.A(_0404_),
    .B(_0443_),
    .Y(_0082_));
 XNOR2x1_ASAP7_75t_R _0821_ (.B(_0698_),
    .Y(_0444_),
    .A(net78));
 XOR2x2_ASAP7_75t_R _0822_ (.A(_0044_),
    .B(_0444_),
    .Y(_0445_));
 NAND2x1_ASAP7_75t_R _0823_ (.A(_0404_),
    .B(_0445_),
    .Y(_0083_));
 NOR2x1_ASAP7_75t_R _0824_ (.A(_0697_),
    .B(_0444_),
    .Y(_0446_));
 AND2x2_ASAP7_75t_R _0825_ (.A(_0045_),
    .B(_0444_),
    .Y(_0447_));
 OR3x1_ASAP7_75t_R _0826_ (.A(_0428_),
    .B(_0446_),
    .C(_0447_),
    .Y(_0084_));
 NOR2x1_ASAP7_75t_R _0827_ (.A(_0067_),
    .B(_0444_),
    .Y(_0448_));
 XNOR2x2_ASAP7_75t_R _0828_ (.A(_0027_),
    .B(_0025_),
    .Y(_0449_));
 AND2x2_ASAP7_75t_R _0829_ (.A(_0444_),
    .B(_0449_),
    .Y(_0450_));
 OR3x1_ASAP7_75t_R _0830_ (.A(_0428_),
    .B(_0448_),
    .C(_0450_),
    .Y(_0085_));
 OR2x2_ASAP7_75t_R _0831_ (.A(\credit_t_route_inst.l_counters_inst.o_credits[8] ),
    .B(_0444_),
    .Y(_0451_));
 OA21x2_ASAP7_75t_R _0832_ (.A1(_0024_),
    .A2(_0044_),
    .B(_0026_),
    .Y(_0452_));
 OA21x2_ASAP7_75t_R _0833_ (.A1(_0025_),
    .A2(_0452_),
    .B(_0029_),
    .Y(_0453_));
 XNOR2x2_ASAP7_75t_R _0834_ (.A(_0028_),
    .B(_0453_),
    .Y(_0454_));
 NAND2x1_ASAP7_75t_R _0835_ (.A(_0444_),
    .B(_0454_),
    .Y(_0455_));
 AO21x1_ASAP7_75t_R _0836_ (.A1(_0451_),
    .A2(_0455_),
    .B(_0422_),
    .Y(_0086_));
 INVx1_ASAP7_75t_R _0837_ (.A(_0027_),
    .Y(_0456_));
 OA21x2_ASAP7_75t_R _0838_ (.A1(_0456_),
    .A2(_0025_),
    .B(_0029_),
    .Y(_0457_));
 OAI21x1_ASAP7_75t_R _0839_ (.A1(_0028_),
    .A2(_0457_),
    .B(_0072_),
    .Y(_0458_));
 NOR2x1_ASAP7_75t_R _0840_ (.A(net78),
    .B(_0458_),
    .Y(_0459_));
 INVx1_ASAP7_75t_R _0841_ (.A(net78),
    .Y(_0460_));
 AOI221x1_ASAP7_75t_R _0842_ (.A1(_0373_),
    .A2(_0418_),
    .B1(_0397_),
    .B2(net233),
    .C(_0460_),
    .Y(_0461_));
 AO22x1_ASAP7_75t_R _0843_ (.A1(net276),
    .A2(_0459_),
    .B1(_0461_),
    .B2(_0458_),
    .Y(_0462_));
 XOR2x2_ASAP7_75t_R _0844_ (.A(_0065_),
    .B(_0462_),
    .Y(_0463_));
 NAND2x1_ASAP7_75t_R _0845_ (.A(_0404_),
    .B(_0463_),
    .Y(_0087_));
 INVx2_ASAP7_75t_R _0846_ (.A(net155),
    .Y(_0464_));
 XNOR2x1_ASAP7_75t_R _0847_ (.B(_0706_),
    .Y(_0465_),
    .A(_0464_));
 XNOR2x2_ASAP7_75t_R _0848_ (.A(_0046_),
    .B(_0465_),
    .Y(_0466_));
 NAND2x1_ASAP7_75t_R _0849_ (.A(_0404_),
    .B(_0466_),
    .Y(_0088_));
 NAND2x1_ASAP7_75t_R _0850_ (.A(_0705_),
    .B(_0465_),
    .Y(_0467_));
 OR2x2_ASAP7_75t_R _0851_ (.A(_0047_),
    .B(_0465_),
    .Y(_0468_));
 AO21x1_ASAP7_75t_R _0852_ (.A1(_0467_),
    .A2(_0468_),
    .B(_0422_),
    .Y(_0089_));
 AND2x2_ASAP7_75t_R _0853_ (.A(\credit_t_route_inst.r_counters_inst.o_credits[2] ),
    .B(_0465_),
    .Y(_0469_));
 XOR2x2_ASAP7_75t_R _0854_ (.A(_0012_),
    .B(_0010_),
    .Y(_0470_));
 NOR2x1_ASAP7_75t_R _0855_ (.A(_0465_),
    .B(_0470_),
    .Y(_0471_));
 OR3x1_ASAP7_75t_R _0856_ (.A(_0428_),
    .B(_0469_),
    .C(_0471_),
    .Y(_0090_));
 NAND2x1_ASAP7_75t_R _0857_ (.A(_0063_),
    .B(_0465_),
    .Y(_0472_));
 OA21x2_ASAP7_75t_R _0858_ (.A1(_0009_),
    .A2(_0046_),
    .B(_0011_),
    .Y(_0473_));
 OA21x2_ASAP7_75t_R _0859_ (.A1(_0010_),
    .A2(_0473_),
    .B(_0014_),
    .Y(_0474_));
 XOR2x2_ASAP7_75t_R _0860_ (.A(_0013_),
    .B(_0474_),
    .Y(_0475_));
 OR2x2_ASAP7_75t_R _0861_ (.A(_0465_),
    .B(_0475_),
    .Y(_0476_));
 AO21x1_ASAP7_75t_R _0862_ (.A1(_0472_),
    .A2(_0476_),
    .B(_0422_),
    .Y(_0091_));
 INVx1_ASAP7_75t_R _0863_ (.A(_0012_),
    .Y(_0477_));
 OA21x2_ASAP7_75t_R _0864_ (.A1(_0477_),
    .A2(_0010_),
    .B(_0014_),
    .Y(_0478_));
 OA21x2_ASAP7_75t_R _0865_ (.A1(_0013_),
    .A2(_0478_),
    .B(_0076_),
    .Y(_0479_));
 NOR2x1_ASAP7_75t_R _0866_ (.A(_0464_),
    .B(_0479_),
    .Y(_0480_));
 OA211x2_ASAP7_75t_R _0867_ (.A1(_0325_),
    .A2(_0330_),
    .B(_0479_),
    .C(_0332_),
    .Y(_0481_));
 AO22x1_ASAP7_75t_R _0868_ (.A1(_0706_),
    .A2(_0480_),
    .B1(_0481_),
    .B2(_0464_),
    .Y(_0482_));
 XNOR2x2_ASAP7_75t_R _0869_ (.A(_0062_),
    .B(_0482_),
    .Y(_0483_));
 OR2x2_ASAP7_75t_R _0870_ (.A(_0422_),
    .B(_0483_),
    .Y(_0092_));
 XNOR2x1_ASAP7_75t_R _0871_ (.B(_0704_),
    .Y(_0484_),
    .A(net156));
 XOR2x2_ASAP7_75t_R _0872_ (.A(_0048_),
    .B(_0484_),
    .Y(_0485_));
 NAND2x1_ASAP7_75t_R _0873_ (.A(_0404_),
    .B(_0485_),
    .Y(_0093_));
 NOR2x1_ASAP7_75t_R _0874_ (.A(_0703_),
    .B(_0484_),
    .Y(_0486_));
 AND2x2_ASAP7_75t_R _0875_ (.A(_0049_),
    .B(_0484_),
    .Y(_0487_));
 OR3x1_ASAP7_75t_R _0876_ (.A(_0428_),
    .B(_0486_),
    .C(_0487_),
    .Y(_0094_));
 NOR2x1_ASAP7_75t_R _0877_ (.A(_0061_),
    .B(_0484_),
    .Y(_0488_));
 XNOR2x2_ASAP7_75t_R _0878_ (.A(_0006_),
    .B(_0004_),
    .Y(_0489_));
 AND2x2_ASAP7_75t_R _0879_ (.A(_0484_),
    .B(_0489_),
    .Y(_0490_));
 OR3x1_ASAP7_75t_R _0880_ (.A(_0428_),
    .B(_0488_),
    .C(_0490_),
    .Y(_0095_));
 OR2x2_ASAP7_75t_R _0881_ (.A(\credit_t_route_inst.r_counters_inst.o_credits[8] ),
    .B(_0484_),
    .Y(_0491_));
 OA21x2_ASAP7_75t_R _0882_ (.A1(_0003_),
    .A2(_0048_),
    .B(_0005_),
    .Y(_0492_));
 OA21x2_ASAP7_75t_R _0883_ (.A1(_0004_),
    .A2(_0492_),
    .B(_0008_),
    .Y(_0493_));
 XNOR2x2_ASAP7_75t_R _0884_ (.A(_0007_),
    .B(_0493_),
    .Y(_0494_));
 NAND2x1_ASAP7_75t_R _0885_ (.A(_0484_),
    .B(_0494_),
    .Y(_0495_));
 AO21x1_ASAP7_75t_R _0886_ (.A1(_0491_),
    .A2(_0495_),
    .B(_0422_),
    .Y(_0096_));
 INVx1_ASAP7_75t_R _0887_ (.A(_0006_),
    .Y(_0496_));
 OA21x2_ASAP7_75t_R _0888_ (.A1(_0496_),
    .A2(_0004_),
    .B(_0008_),
    .Y(_0497_));
 OAI21x1_ASAP7_75t_R _0889_ (.A1(_0007_),
    .A2(_0497_),
    .B(_0075_),
    .Y(_0498_));
 INVx1_ASAP7_75t_R _0890_ (.A(net156),
    .Y(_0499_));
 OAI21x1_ASAP7_75t_R _0891_ (.A1(_0337_),
    .A2(_0342_),
    .B(_0499_),
    .Y(_0500_));
 NAND2x1_ASAP7_75t_R _0892_ (.A(net156),
    .B(_0498_),
    .Y(_0501_));
 OAI22x1_ASAP7_75t_R _0893_ (.A1(_0498_),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net317),
    .Y(_0502_));
 XNOR2x2_ASAP7_75t_R _0894_ (.A(_0071_),
    .B(_0502_),
    .Y(_0503_));
 OR2x2_ASAP7_75t_R _0895_ (.A(_0428_),
    .B(_0503_),
    .Y(_0097_));
 XNOR2x1_ASAP7_75t_R _0896_ (.B(_0708_),
    .Y(_0504_),
    .A(net234));
 XOR2x2_ASAP7_75t_R _0897_ (.A(_0050_),
    .B(_0504_),
    .Y(_0505_));
 NAND2x1_ASAP7_75t_R _0898_ (.A(_0404_),
    .B(_0505_),
    .Y(_0098_));
 NOR2x1_ASAP7_75t_R _0899_ (.A(_0707_),
    .B(_0504_),
    .Y(_0506_));
 AND2x2_ASAP7_75t_R _0900_ (.A(_0051_),
    .B(_0504_),
    .Y(_0507_));
 OR3x1_ASAP7_75t_R _0901_ (.A(_0428_),
    .B(_0506_),
    .C(_0507_),
    .Y(_0099_));
 NOR2x1_ASAP7_75t_R _0902_ (.A(_0059_),
    .B(_0504_),
    .Y(_0508_));
 XNOR2x2_ASAP7_75t_R _0903_ (.A(_0018_),
    .B(_0016_),
    .Y(_0509_));
 AND2x2_ASAP7_75t_R _0904_ (.A(_0504_),
    .B(_0509_),
    .Y(_0510_));
 OR3x1_ASAP7_75t_R _0905_ (.A(_0428_),
    .B(_0508_),
    .C(_0510_),
    .Y(_0100_));
 OR2x2_ASAP7_75t_R _0906_ (.A(\credit_t_route_inst.u0_counters_inst.o_credits[3] ),
    .B(_0504_),
    .Y(_0511_));
 OA21x2_ASAP7_75t_R _0907_ (.A1(_0015_),
    .A2(_0050_),
    .B(_0017_),
    .Y(_0512_));
 OA21x2_ASAP7_75t_R _0908_ (.A1(_0016_),
    .A2(_0512_),
    .B(_0020_),
    .Y(_0513_));
 XNOR2x2_ASAP7_75t_R _0909_ (.A(_0019_),
    .B(_0513_),
    .Y(_0514_));
 NAND2x1_ASAP7_75t_R _0910_ (.A(_0504_),
    .B(_0514_),
    .Y(_0515_));
 AO21x1_ASAP7_75t_R _0911_ (.A1(_0511_),
    .A2(_0515_),
    .B(_0422_),
    .Y(_0101_));
 INVx1_ASAP7_75t_R _0912_ (.A(net234),
    .Y(_0516_));
 INVx1_ASAP7_75t_R _0913_ (.A(_0018_),
    .Y(_0517_));
 OA21x2_ASAP7_75t_R _0914_ (.A1(_0517_),
    .A2(_0016_),
    .B(_0020_),
    .Y(_0518_));
 OA21x2_ASAP7_75t_R _0915_ (.A1(_0019_),
    .A2(_0518_),
    .B(_0077_),
    .Y(_0519_));
 NOR2x1_ASAP7_75t_R _0916_ (.A(_0516_),
    .B(_0519_),
    .Y(_0520_));
 AND3x1_ASAP7_75t_R _0917_ (.A(_0516_),
    .B(net357),
    .C(_0519_),
    .Y(_0521_));
 AO21x1_ASAP7_75t_R _0918_ (.A1(_0708_),
    .A2(_0520_),
    .B(_0521_),
    .Y(_0522_));
 XNOR2x2_ASAP7_75t_R _0919_ (.A(_0057_),
    .B(_0522_),
    .Y(_0523_));
 OR2x2_ASAP7_75t_R _0920_ (.A(_0428_),
    .B(_0523_),
    .Y(_0102_));
 XOR2x1_ASAP7_75t_R _0921_ (.A(net235),
    .Y(_0524_),
    .B(_0366_));
 XOR2x2_ASAP7_75t_R _0922_ (.A(_0052_),
    .B(_0524_),
    .Y(_0525_));
 NAND2x1_ASAP7_75t_R _0923_ (.A(_0404_),
    .B(_0525_),
    .Y(_0103_));
 NOR2x1_ASAP7_75t_R _0924_ (.A(_0701_),
    .B(_0524_),
    .Y(_0526_));
 AND2x2_ASAP7_75t_R _0925_ (.A(_0053_),
    .B(_0524_),
    .Y(_0527_));
 OR3x1_ASAP7_75t_R _0926_ (.A(net157),
    .B(_0526_),
    .C(_0527_),
    .Y(_0104_));
 NOR2x1_ASAP7_75t_R _0927_ (.A(_0056_),
    .B(_0524_),
    .Y(_0528_));
 XNOR2x2_ASAP7_75t_R _0928_ (.A(_0039_),
    .B(_0037_),
    .Y(_0529_));
 AND2x2_ASAP7_75t_R _0929_ (.A(_0524_),
    .B(_0529_),
    .Y(_0530_));
 OR3x1_ASAP7_75t_R _0930_ (.A(net157),
    .B(_0528_),
    .C(_0530_),
    .Y(_0105_));
 OR2x2_ASAP7_75t_R _0931_ (.A(\credit_t_route_inst.u0_counters_inst.o_credits[8] ),
    .B(_0524_),
    .Y(_0531_));
 OA21x2_ASAP7_75t_R _0932_ (.A1(_0036_),
    .A2(_0052_),
    .B(_0038_),
    .Y(_0532_));
 OA21x2_ASAP7_75t_R _0933_ (.A1(_0037_),
    .A2(_0532_),
    .B(_0041_),
    .Y(_0533_));
 XNOR2x2_ASAP7_75t_R _0934_ (.A(_0040_),
    .B(_0533_),
    .Y(_0534_));
 NAND2x1_ASAP7_75t_R _0935_ (.A(_0524_),
    .B(_0534_),
    .Y(_0535_));
 AO21x1_ASAP7_75t_R _0936_ (.A1(_0531_),
    .A2(_0535_),
    .B(_0422_),
    .Y(_0106_));
 INVx1_ASAP7_75t_R _0937_ (.A(_0039_),
    .Y(_0536_));
 OA21x2_ASAP7_75t_R _0938_ (.A1(_0536_),
    .A2(_0037_),
    .B(_0041_),
    .Y(_0537_));
 OAI21x1_ASAP7_75t_R _0939_ (.A1(_0040_),
    .A2(_0537_),
    .B(_0074_),
    .Y(_0538_));
 OA211x2_ASAP7_75t_R _0940_ (.A1(_0350_),
    .A2(_0355_),
    .B(_0365_),
    .C(_0538_),
    .Y(_0539_));
 NOR2x1_ASAP7_75t_R _0941_ (.A(net235),
    .B(_0538_),
    .Y(_0540_));
 AO22x1_ASAP7_75t_R _0942_ (.A1(net235),
    .A2(_0539_),
    .B1(_0540_),
    .B2(_0366_),
    .Y(_0541_));
 XOR2x2_ASAP7_75t_R _0943_ (.A(_0054_),
    .B(_0541_),
    .Y(_0542_));
 NAND2x1_ASAP7_75t_R _0944_ (.A(_0404_),
    .B(_0542_),
    .Y(_0107_));
 NAND2x2_ASAP7_75t_R _0945_ (.A(_0373_),
    .B(_0418_),
    .Y(_0543_));
 BUFx6f_ASAP7_75t_R _0946_ (.A(_0543_),
    .Y(_0544_));
 OA21x2_ASAP7_75t_R _0947_ (.A1(_0374_),
    .A2(_0414_),
    .B(net276),
    .Y(_0545_));
 BUFx6f_ASAP7_75t_R _0948_ (.A(_0545_),
    .Y(_0546_));
 BUFx6f_ASAP7_75t_R _0949_ (.A(_0546_),
    .Y(_0547_));
 OR4x1_ASAP7_75t_R _0950_ (.A(_0356_),
    .B(net144),
    .C(_0346_),
    .D(_0381_),
    .Y(_0548_));
 OA21x2_ASAP7_75t_R _0951_ (.A1(_0374_),
    .A2(_0413_),
    .B(_0548_),
    .Y(_0549_));
 AO21x2_ASAP7_75t_R _0952_ (.A1(_0360_),
    .A2(_0380_),
    .B(_0549_),
    .Y(_0550_));
 BUFx6f_ASAP7_75t_R _0953_ (.A(_0550_),
    .Y(_0551_));
 BUFx6f_ASAP7_75t_R _0954_ (.A(_0551_),
    .Y(_0552_));
 AOI21x1_ASAP7_75t_R _0955_ (.A1(_0360_),
    .A2(_0380_),
    .B(_0549_),
    .Y(_0553_));
 BUFx6f_ASAP7_75t_R _0956_ (.A(_0553_),
    .Y(_0554_));
 AND2x2_ASAP7_75t_R _0957_ (.A(net79),
    .B(_0554_),
    .Y(_0555_));
 AO21x1_ASAP7_75t_R _0958_ (.A1(net158),
    .A2(_0552_),
    .B(_0555_),
    .Y(_0556_));
 NAND2x2_ASAP7_75t_R _0959_ (.A(net276),
    .B(_0550_),
    .Y(_0557_));
 BUFx6f_ASAP7_75t_R _0960_ (.A(_0557_),
    .Y(_0558_));
 OA222x2_ASAP7_75t_R _0961_ (.A1(net109),
    .A2(_0544_),
    .B1(_0547_),
    .B2(_0556_),
    .C1(_0558_),
    .C2(net188),
    .Y(net238));
 AND2x2_ASAP7_75t_R _0962_ (.A(net80),
    .B(_0554_),
    .Y(_0559_));
 AO21x1_ASAP7_75t_R _0963_ (.A1(net159),
    .A2(_0552_),
    .B(_0559_),
    .Y(_0560_));
 OA222x2_ASAP7_75t_R _0964_ (.A1(net120),
    .A2(_0544_),
    .B1(_0547_),
    .B2(_0560_),
    .C1(_0558_),
    .C2(net199),
    .Y(net239));
 AND2x2_ASAP7_75t_R _0965_ (.A(net81),
    .B(_0554_),
    .Y(_0561_));
 AO21x1_ASAP7_75t_R _0966_ (.A1(net160),
    .A2(_0552_),
    .B(_0561_),
    .Y(_0562_));
 OA222x2_ASAP7_75t_R _0967_ (.A1(net121),
    .A2(_0544_),
    .B1(_0547_),
    .B2(_0562_),
    .C1(_0558_),
    .C2(net200),
    .Y(net240));
 AND2x2_ASAP7_75t_R _0968_ (.A(net82),
    .B(_0554_),
    .Y(_0563_));
 AO21x1_ASAP7_75t_R _0969_ (.A1(net161),
    .A2(_0552_),
    .B(_0563_),
    .Y(_0564_));
 OA222x2_ASAP7_75t_R _0970_ (.A1(net122),
    .A2(_0544_),
    .B1(_0547_),
    .B2(_0564_),
    .C1(_0558_),
    .C2(net201),
    .Y(net241));
 AND2x2_ASAP7_75t_R _0971_ (.A(net83),
    .B(_0554_),
    .Y(_0565_));
 AO21x1_ASAP7_75t_R _0972_ (.A1(net162),
    .A2(_0552_),
    .B(_0565_),
    .Y(_0566_));
 OA222x2_ASAP7_75t_R _0973_ (.A1(net124),
    .A2(_0544_),
    .B1(_0547_),
    .B2(_0566_),
    .C1(_0558_),
    .C2(net203),
    .Y(net242));
 AND2x2_ASAP7_75t_R _0974_ (.A(net84),
    .B(_0554_),
    .Y(_0567_));
 AO21x1_ASAP7_75t_R _0975_ (.A1(net163),
    .A2(_0552_),
    .B(_0567_),
    .Y(_0568_));
 OA222x2_ASAP7_75t_R _0976_ (.A1(net125),
    .A2(_0544_),
    .B1(_0547_),
    .B2(_0568_),
    .C1(_0558_),
    .C2(net204),
    .Y(net243));
 BUFx6f_ASAP7_75t_R _0977_ (.A(_0546_),
    .Y(_0569_));
 BUFx6f_ASAP7_75t_R _0978_ (.A(_0551_),
    .Y(_0570_));
 AND2x2_ASAP7_75t_R _0979_ (.A(net85),
    .B(_0554_),
    .Y(_0571_));
 AO21x1_ASAP7_75t_R _0980_ (.A1(net164),
    .A2(_0570_),
    .B(_0571_),
    .Y(_0572_));
 OA222x2_ASAP7_75t_R _0981_ (.A1(net126),
    .A2(_0544_),
    .B1(_0569_),
    .B2(_0572_),
    .C1(_0558_),
    .C2(net205),
    .Y(net244));
 AND2x2_ASAP7_75t_R _0982_ (.A(net86),
    .B(_0554_),
    .Y(_0573_));
 AO21x1_ASAP7_75t_R _0983_ (.A1(net165),
    .A2(_0570_),
    .B(_0573_),
    .Y(_0574_));
 OA222x2_ASAP7_75t_R _0984_ (.A1(net127),
    .A2(_0544_),
    .B1(_0569_),
    .B2(_0574_),
    .C1(_0558_),
    .C2(net206),
    .Y(net245));
 AND2x2_ASAP7_75t_R _0985_ (.A(net87),
    .B(_0554_),
    .Y(_0575_));
 AO21x1_ASAP7_75t_R _0986_ (.A1(net166),
    .A2(_0570_),
    .B(_0575_),
    .Y(_0576_));
 OA222x2_ASAP7_75t_R _0987_ (.A1(net128),
    .A2(_0544_),
    .B1(_0569_),
    .B2(_0576_),
    .C1(_0558_),
    .C2(net207),
    .Y(net246));
 AND2x2_ASAP7_75t_R _0988_ (.A(net88),
    .B(_0554_),
    .Y(_0577_));
 AO21x1_ASAP7_75t_R _0989_ (.A1(net167),
    .A2(_0570_),
    .B(_0577_),
    .Y(_0578_));
 OA222x2_ASAP7_75t_R _0990_ (.A1(net129),
    .A2(_0544_),
    .B1(_0569_),
    .B2(_0578_),
    .C1(_0558_),
    .C2(net208),
    .Y(net247));
 BUFx6f_ASAP7_75t_R _0991_ (.A(_0543_),
    .Y(_0579_));
 BUFx6f_ASAP7_75t_R _0992_ (.A(_0553_),
    .Y(_0580_));
 AND2x2_ASAP7_75t_R _0993_ (.A(net89),
    .B(_0580_),
    .Y(_0581_));
 AO21x1_ASAP7_75t_R _0994_ (.A1(net168),
    .A2(_0570_),
    .B(_0581_),
    .Y(_0582_));
 BUFx6f_ASAP7_75t_R _0995_ (.A(_0557_),
    .Y(_0583_));
 OA222x2_ASAP7_75t_R _0996_ (.A1(net130),
    .A2(_0579_),
    .B1(_0569_),
    .B2(_0582_),
    .C1(_0583_),
    .C2(net209),
    .Y(net248));
 AND2x2_ASAP7_75t_R _0997_ (.A(net90),
    .B(_0580_),
    .Y(_0584_));
 AO21x1_ASAP7_75t_R _0998_ (.A1(net169),
    .A2(_0570_),
    .B(_0584_),
    .Y(_0585_));
 OA222x2_ASAP7_75t_R _0999_ (.A1(net110),
    .A2(_0579_),
    .B1(_0569_),
    .B2(_0585_),
    .C1(_0583_),
    .C2(net189),
    .Y(net249));
 AND2x2_ASAP7_75t_R _1000_ (.A(net91),
    .B(_0580_),
    .Y(_0586_));
 AO21x1_ASAP7_75t_R _1001_ (.A1(net170),
    .A2(_0570_),
    .B(_0586_),
    .Y(_0587_));
 OA222x2_ASAP7_75t_R _1002_ (.A1(net131),
    .A2(_0579_),
    .B1(_0569_),
    .B2(_0587_),
    .C1(_0583_),
    .C2(net210),
    .Y(net250));
 AND2x2_ASAP7_75t_R _1003_ (.A(net92),
    .B(_0580_),
    .Y(_0588_));
 AO21x1_ASAP7_75t_R _1004_ (.A1(net171),
    .A2(_0570_),
    .B(_0588_),
    .Y(_0589_));
 OA222x2_ASAP7_75t_R _1005_ (.A1(net132),
    .A2(_0579_),
    .B1(_0569_),
    .B2(_0589_),
    .C1(_0583_),
    .C2(net211),
    .Y(net251));
 AND2x2_ASAP7_75t_R _1006_ (.A(net93),
    .B(_0580_),
    .Y(_0590_));
 AO21x1_ASAP7_75t_R _1007_ (.A1(net172),
    .A2(_0570_),
    .B(_0590_),
    .Y(_0591_));
 OA222x2_ASAP7_75t_R _1008_ (.A1(net133),
    .A2(_0579_),
    .B1(_0569_),
    .B2(_0591_),
    .C1(_0583_),
    .C2(net212),
    .Y(net252));
 AND2x2_ASAP7_75t_R _1009_ (.A(net94),
    .B(_0580_),
    .Y(_0592_));
 AO21x1_ASAP7_75t_R _1010_ (.A1(net173),
    .A2(_0570_),
    .B(_0592_),
    .Y(_0593_));
 OA222x2_ASAP7_75t_R _1011_ (.A1(net135),
    .A2(_0579_),
    .B1(_0569_),
    .B2(_0593_),
    .C1(_0583_),
    .C2(net214),
    .Y(net253));
 BUFx6f_ASAP7_75t_R _1012_ (.A(_0546_),
    .Y(_0594_));
 BUFx6f_ASAP7_75t_R _1013_ (.A(_0551_),
    .Y(_0595_));
 AND2x2_ASAP7_75t_R _1014_ (.A(net95),
    .B(_0580_),
    .Y(_0596_));
 AO21x1_ASAP7_75t_R _1015_ (.A1(net174),
    .A2(_0595_),
    .B(_0596_),
    .Y(_0597_));
 OA222x2_ASAP7_75t_R _1016_ (.A1(net136),
    .A2(_0579_),
    .B1(_0594_),
    .B2(_0597_),
    .C1(_0583_),
    .C2(net215),
    .Y(net254));
 AND2x2_ASAP7_75t_R _1017_ (.A(net96),
    .B(_0580_),
    .Y(_0598_));
 AO21x1_ASAP7_75t_R _1018_ (.A1(net175),
    .A2(_0595_),
    .B(_0598_),
    .Y(_0599_));
 OA222x2_ASAP7_75t_R _1019_ (.A1(net137),
    .A2(_0579_),
    .B1(_0594_),
    .B2(_0599_),
    .C1(_0583_),
    .C2(net216),
    .Y(net255));
 AND2x2_ASAP7_75t_R _1020_ (.A(net97),
    .B(_0580_),
    .Y(_0600_));
 AO21x1_ASAP7_75t_R _1021_ (.A1(net176),
    .A2(_0595_),
    .B(_0600_),
    .Y(_0601_));
 OA222x2_ASAP7_75t_R _1022_ (.A1(net138),
    .A2(_0579_),
    .B1(_0594_),
    .B2(_0601_),
    .C1(_0583_),
    .C2(net217),
    .Y(net256));
 AND2x2_ASAP7_75t_R _1023_ (.A(net98),
    .B(_0580_),
    .Y(_0602_));
 AO21x1_ASAP7_75t_R _1024_ (.A1(net177),
    .A2(_0595_),
    .B(_0602_),
    .Y(_0603_));
 OA222x2_ASAP7_75t_R _1025_ (.A1(net139),
    .A2(_0579_),
    .B1(_0594_),
    .B2(_0603_),
    .C1(_0583_),
    .C2(net218),
    .Y(net257));
 BUFx6f_ASAP7_75t_R _1026_ (.A(_0543_),
    .Y(_0604_));
 BUFx6f_ASAP7_75t_R _1027_ (.A(_0553_),
    .Y(_0605_));
 AND2x2_ASAP7_75t_R _1028_ (.A(net99),
    .B(_0605_),
    .Y(_0606_));
 AO21x1_ASAP7_75t_R _1029_ (.A1(net178),
    .A2(_0595_),
    .B(_0606_),
    .Y(_0607_));
 BUFx6f_ASAP7_75t_R _1030_ (.A(_0557_),
    .Y(_0608_));
 OA222x2_ASAP7_75t_R _1031_ (.A1(net140),
    .A2(_0604_),
    .B1(_0594_),
    .B2(_0607_),
    .C1(_0608_),
    .C2(net219),
    .Y(net258));
 AND2x2_ASAP7_75t_R _1032_ (.A(net100),
    .B(_0605_),
    .Y(_0609_));
 AO21x1_ASAP7_75t_R _1033_ (.A1(net179),
    .A2(_0595_),
    .B(_0609_),
    .Y(_0610_));
 OA222x2_ASAP7_75t_R _1034_ (.A1(net141),
    .A2(_0604_),
    .B1(_0594_),
    .B2(_0610_),
    .C1(_0608_),
    .C2(net220),
    .Y(net259));
 AND2x2_ASAP7_75t_R _1035_ (.A(net101),
    .B(_0605_),
    .Y(_0611_));
 AO21x1_ASAP7_75t_R _1036_ (.A1(net180),
    .A2(_0595_),
    .B(_0611_),
    .Y(_0612_));
 OA222x2_ASAP7_75t_R _1037_ (.A1(net111),
    .A2(_0604_),
    .B1(_0594_),
    .B2(_0612_),
    .C1(_0608_),
    .C2(net190),
    .Y(net260));
 AND2x2_ASAP7_75t_R _1038_ (.A(net102),
    .B(_0605_),
    .Y(_0613_));
 AO21x1_ASAP7_75t_R _1039_ (.A1(net181),
    .A2(_0595_),
    .B(_0613_),
    .Y(_0614_));
 OA222x2_ASAP7_75t_R _1040_ (.A1(net142),
    .A2(_0604_),
    .B1(_0594_),
    .B2(_0614_),
    .C1(_0608_),
    .C2(net221),
    .Y(net261));
 AND2x2_ASAP7_75t_R _1041_ (.A(net103),
    .B(_0605_),
    .Y(_0615_));
 AO21x1_ASAP7_75t_R _1042_ (.A1(net182),
    .A2(_0595_),
    .B(_0615_),
    .Y(_0616_));
 OA222x2_ASAP7_75t_R _1043_ (.A1(net143),
    .A2(_0604_),
    .B1(_0594_),
    .B2(_0616_),
    .C1(_0608_),
    .C2(net222),
    .Y(net262));
 OA21x2_ASAP7_75t_R _1044_ (.A1(net223),
    .A2(_0698_),
    .B(_0552_),
    .Y(_0617_));
 OA21x2_ASAP7_75t_R _1045_ (.A1(net183),
    .A2(_0547_),
    .B(_0617_),
    .Y(net263));
 OA21x2_ASAP7_75t_R _1046_ (.A1(net225),
    .A2(_0698_),
    .B(_0552_),
    .Y(_0618_));
 OA21x2_ASAP7_75t_R _1047_ (.A1(net184),
    .A2(_0547_),
    .B(_0618_),
    .Y(net264));
 OA21x2_ASAP7_75t_R _1048_ (.A1(net226),
    .A2(_0698_),
    .B(_0552_),
    .Y(_0619_));
 OA21x2_ASAP7_75t_R _1049_ (.A1(net185),
    .A2(_0547_),
    .B(_0619_),
    .Y(net265));
 OA21x2_ASAP7_75t_R _1050_ (.A1(net227),
    .A2(_0698_),
    .B(_0552_),
    .Y(_0620_));
 OA21x2_ASAP7_75t_R _1051_ (.A1(net186),
    .A2(_0547_),
    .B(_0620_),
    .Y(net266));
 AND2x2_ASAP7_75t_R _1052_ (.A(net108),
    .B(_0605_),
    .Y(_0621_));
 AO21x1_ASAP7_75t_R _1053_ (.A1(net187),
    .A2(_0595_),
    .B(_0621_),
    .Y(_0622_));
 OA222x2_ASAP7_75t_R _1054_ (.A1(net149),
    .A2(_0604_),
    .B1(_0594_),
    .B2(_0622_),
    .C1(_0608_),
    .C2(net228),
    .Y(net267));
 AND2x2_ASAP7_75t_R _1055_ (.A(net112),
    .B(_0605_),
    .Y(_0623_));
 AO21x1_ASAP7_75t_R _1056_ (.A1(net191),
    .A2(_0551_),
    .B(_0623_),
    .Y(_0624_));
 OA222x2_ASAP7_75t_R _1057_ (.A1(net113),
    .A2(_0604_),
    .B1(_0546_),
    .B2(_0624_),
    .C1(_0608_),
    .C2(net192),
    .Y(net268));
 AND2x2_ASAP7_75t_R _1058_ (.A(net123),
    .B(_0605_),
    .Y(_0625_));
 AO21x1_ASAP7_75t_R _1059_ (.A1(net202),
    .A2(_0551_),
    .B(_0625_),
    .Y(_0626_));
 OA222x2_ASAP7_75t_R _1060_ (.A1(net114),
    .A2(_0604_),
    .B1(_0546_),
    .B2(_0626_),
    .C1(_0608_),
    .C2(net193),
    .Y(net269));
 AND2x2_ASAP7_75t_R _1061_ (.A(net134),
    .B(_0605_),
    .Y(_0627_));
 AO21x1_ASAP7_75t_R _1062_ (.A1(net213),
    .A2(_0551_),
    .B(_0627_),
    .Y(_0628_));
 OA222x2_ASAP7_75t_R _1063_ (.A1(net115),
    .A2(_0604_),
    .B1(_0546_),
    .B2(_0628_),
    .C1(_0608_),
    .C2(net194),
    .Y(net270));
 AND2x2_ASAP7_75t_R _1064_ (.A(net145),
    .B(_0605_),
    .Y(_0629_));
 AO21x1_ASAP7_75t_R _1065_ (.A1(net224),
    .A2(_0551_),
    .B(_0629_),
    .Y(_0630_));
 OA222x2_ASAP7_75t_R _1066_ (.A1(net116),
    .A2(_0604_),
    .B1(_0546_),
    .B2(_0630_),
    .C1(_0608_),
    .C2(net195),
    .Y(net271));
 AND2x2_ASAP7_75t_R _1067_ (.A(net150),
    .B(_0553_),
    .Y(_0631_));
 AO21x1_ASAP7_75t_R _1068_ (.A1(net229),
    .A2(_0551_),
    .B(_0631_),
    .Y(_0632_));
 OA222x2_ASAP7_75t_R _1069_ (.A1(net117),
    .A2(_0543_),
    .B1(_0546_),
    .B2(_0632_),
    .C1(_0557_),
    .C2(net196),
    .Y(net272));
 AND2x2_ASAP7_75t_R _1070_ (.A(net151),
    .B(_0553_),
    .Y(_0633_));
 AO21x1_ASAP7_75t_R _1071_ (.A1(net230),
    .A2(_0551_),
    .B(_0633_),
    .Y(_0634_));
 OA222x2_ASAP7_75t_R _1072_ (.A1(net118),
    .A2(_0543_),
    .B1(_0546_),
    .B2(_0634_),
    .C1(_0557_),
    .C2(net197),
    .Y(net273));
 AND2x2_ASAP7_75t_R _1073_ (.A(net152),
    .B(_0553_),
    .Y(_0635_));
 AO21x1_ASAP7_75t_R _1074_ (.A1(net231),
    .A2(_0551_),
    .B(_0635_),
    .Y(_0636_));
 OA222x2_ASAP7_75t_R _1075_ (.A1(net119),
    .A2(_0543_),
    .B1(_0546_),
    .B2(_0636_),
    .C1(_0557_),
    .C2(net198),
    .Y(net274));
 OR3x2_ASAP7_75t_R _1076_ (.A(_0327_),
    .B(_0328_),
    .C(_0334_),
    .Y(_0637_));
 OR3x2_ASAP7_75t_R _1077_ (.A(_0387_),
    .B(_0637_),
    .C(_0388_),
    .Y(_0638_));
 BUFx6f_ASAP7_75t_R _1078_ (.A(_0638_),
    .Y(_0639_));
 AOI21x1_ASAP7_75t_R _1079_ (.A1(_0332_),
    .A2(_0325_),
    .B(_0704_),
    .Y(_0640_));
 BUFx6f_ASAP7_75t_R _1080_ (.A(_0640_),
    .Y(_0641_));
 AO21x2_ASAP7_75t_R _1081_ (.A1(_0637_),
    .A2(_0336_),
    .B(_0387_),
    .Y(_0642_));
 BUFx6f_ASAP7_75t_R _1082_ (.A(_0642_),
    .Y(_0643_));
 BUFx6f_ASAP7_75t_R _1083_ (.A(_0643_),
    .Y(_0644_));
 AOI21x1_ASAP7_75t_R _1084_ (.A1(_0637_),
    .A2(_0336_),
    .B(_0387_),
    .Y(_0645_));
 BUFx6f_ASAP7_75t_R _1085_ (.A(_0645_),
    .Y(_0646_));
 AND2x2_ASAP7_75t_R _1086_ (.A(net1),
    .B(_0646_),
    .Y(_0647_));
 AO21x1_ASAP7_75t_R _1087_ (.A1(net158),
    .A2(_0644_),
    .B(_0647_),
    .Y(_0648_));
 NAND2x2_ASAP7_75t_R _1088_ (.A(net317),
    .B(_0642_),
    .Y(_0649_));
 BUFx6f_ASAP7_75t_R _1089_ (.A(_0649_),
    .Y(_0650_));
 OA222x2_ASAP7_75t_R _1090_ (.A1(net31),
    .A2(_0639_),
    .B1(_0641_),
    .B2(_0648_),
    .C1(_0650_),
    .C2(net188),
    .Y(net279));
 AND2x2_ASAP7_75t_R _1091_ (.A(net2),
    .B(_0646_),
    .Y(_0651_));
 AO21x1_ASAP7_75t_R _1092_ (.A1(net159),
    .A2(_0644_),
    .B(_0651_),
    .Y(_0652_));
 OA222x2_ASAP7_75t_R _1093_ (.A1(net42),
    .A2(_0639_),
    .B1(_0641_),
    .B2(_0652_),
    .C1(_0650_),
    .C2(net199),
    .Y(net280));
 AND2x2_ASAP7_75t_R _1094_ (.A(net3),
    .B(_0646_),
    .Y(_0653_));
 AO21x1_ASAP7_75t_R _1095_ (.A1(net160),
    .A2(_0644_),
    .B(_0653_),
    .Y(_0654_));
 OA222x2_ASAP7_75t_R _1096_ (.A1(net43),
    .A2(_0639_),
    .B1(_0641_),
    .B2(_0654_),
    .C1(_0650_),
    .C2(net200),
    .Y(net281));
 AND2x2_ASAP7_75t_R _1097_ (.A(net4),
    .B(_0646_),
    .Y(_0655_));
 AO21x1_ASAP7_75t_R _1098_ (.A1(net161),
    .A2(_0644_),
    .B(_0655_),
    .Y(_0656_));
 OA222x2_ASAP7_75t_R _1099_ (.A1(net44),
    .A2(_0639_),
    .B1(_0641_),
    .B2(_0656_),
    .C1(_0650_),
    .C2(net201),
    .Y(net282));
 AND2x2_ASAP7_75t_R _1100_ (.A(net5),
    .B(_0646_),
    .Y(_0657_));
 AO21x1_ASAP7_75t_R _1101_ (.A1(net162),
    .A2(_0644_),
    .B(_0657_),
    .Y(_0658_));
 OA222x2_ASAP7_75t_R _1102_ (.A1(net46),
    .A2(_0639_),
    .B1(_0641_),
    .B2(_0658_),
    .C1(_0650_),
    .C2(net203),
    .Y(net283));
 AND2x2_ASAP7_75t_R _1103_ (.A(net6),
    .B(_0646_),
    .Y(_0659_));
 AO21x1_ASAP7_75t_R _1104_ (.A1(net163),
    .A2(_0644_),
    .B(_0659_),
    .Y(_0660_));
 OA222x2_ASAP7_75t_R _1105_ (.A1(net47),
    .A2(_0639_),
    .B1(_0641_),
    .B2(_0660_),
    .C1(_0650_),
    .C2(net204),
    .Y(net284));
 BUFx6f_ASAP7_75t_R _1106_ (.A(_0643_),
    .Y(_0661_));
 AND2x2_ASAP7_75t_R _1107_ (.A(net7),
    .B(_0646_),
    .Y(_0662_));
 AO21x1_ASAP7_75t_R _1108_ (.A1(net164),
    .A2(_0661_),
    .B(_0662_),
    .Y(_0663_));
 OA222x2_ASAP7_75t_R _1109_ (.A1(net48),
    .A2(_0639_),
    .B1(_0641_),
    .B2(_0663_),
    .C1(_0650_),
    .C2(net205),
    .Y(net285));
 BUFx6f_ASAP7_75t_R _1110_ (.A(_0640_),
    .Y(_0664_));
 AND2x2_ASAP7_75t_R _1111_ (.A(net8),
    .B(_0646_),
    .Y(_0665_));
 AO21x1_ASAP7_75t_R _1112_ (.A1(net165),
    .A2(_0661_),
    .B(_0665_),
    .Y(_0666_));
 OA222x2_ASAP7_75t_R _1113_ (.A1(net49),
    .A2(_0639_),
    .B1(_0664_),
    .B2(_0666_),
    .C1(_0650_),
    .C2(net206),
    .Y(net286));
 AND2x2_ASAP7_75t_R _1114_ (.A(net9),
    .B(_0646_),
    .Y(_0667_));
 AO21x1_ASAP7_75t_R _1115_ (.A1(net166),
    .A2(_0661_),
    .B(_0667_),
    .Y(_0668_));
 OA222x2_ASAP7_75t_R _1116_ (.A1(net50),
    .A2(_0639_),
    .B1(_0664_),
    .B2(_0668_),
    .C1(_0650_),
    .C2(net207),
    .Y(net287));
 AND2x2_ASAP7_75t_R _1117_ (.A(net10),
    .B(_0646_),
    .Y(_0669_));
 AO21x1_ASAP7_75t_R _1118_ (.A1(net167),
    .A2(_0661_),
    .B(_0669_),
    .Y(_0670_));
 OA222x2_ASAP7_75t_R _1119_ (.A1(net51),
    .A2(_0639_),
    .B1(_0664_),
    .B2(_0670_),
    .C1(_0650_),
    .C2(net208),
    .Y(net288));
 BUFx6f_ASAP7_75t_R _1120_ (.A(_0638_),
    .Y(_0671_));
 BUFx6f_ASAP7_75t_R _1121_ (.A(_0645_),
    .Y(_0672_));
 AND2x2_ASAP7_75t_R _1122_ (.A(net11),
    .B(_0672_),
    .Y(_0673_));
 AO21x1_ASAP7_75t_R _1123_ (.A1(net168),
    .A2(_0661_),
    .B(_0673_),
    .Y(_0674_));
 BUFx6f_ASAP7_75t_R _1124_ (.A(_0649_),
    .Y(_0675_));
 OA222x2_ASAP7_75t_R _1125_ (.A1(net52),
    .A2(_0671_),
    .B1(_0664_),
    .B2(_0674_),
    .C1(_0675_),
    .C2(net209),
    .Y(net289));
 AND2x2_ASAP7_75t_R _1126_ (.A(net12),
    .B(_0672_),
    .Y(_0676_));
 AO21x1_ASAP7_75t_R _1127_ (.A1(net169),
    .A2(_0661_),
    .B(_0676_),
    .Y(_0677_));
 OA222x2_ASAP7_75t_R _1128_ (.A1(net32),
    .A2(_0671_),
    .B1(_0664_),
    .B2(_0677_),
    .C1(_0675_),
    .C2(net189),
    .Y(net290));
 AND2x2_ASAP7_75t_R _1129_ (.A(net13),
    .B(_0672_),
    .Y(_0678_));
 AO21x1_ASAP7_75t_R _1130_ (.A1(net170),
    .A2(_0661_),
    .B(_0678_),
    .Y(_0679_));
 OA222x2_ASAP7_75t_R _1131_ (.A1(net53),
    .A2(_0671_),
    .B1(_0664_),
    .B2(_0679_),
    .C1(_0675_),
    .C2(net210),
    .Y(net291));
 AND2x2_ASAP7_75t_R _1132_ (.A(net14),
    .B(_0672_),
    .Y(_0680_));
 AO21x1_ASAP7_75t_R _1133_ (.A1(net171),
    .A2(_0661_),
    .B(_0680_),
    .Y(_0681_));
 OA222x2_ASAP7_75t_R _1134_ (.A1(net54),
    .A2(_0671_),
    .B1(_0664_),
    .B2(_0681_),
    .C1(_0675_),
    .C2(net211),
    .Y(net292));
 AND2x2_ASAP7_75t_R _1135_ (.A(net15),
    .B(_0672_),
    .Y(_0682_));
 AO21x1_ASAP7_75t_R _1136_ (.A1(net172),
    .A2(_0661_),
    .B(_0682_),
    .Y(_0683_));
 OA222x2_ASAP7_75t_R _1137_ (.A1(net55),
    .A2(_0671_),
    .B1(_0664_),
    .B2(_0683_),
    .C1(_0675_),
    .C2(net212),
    .Y(net293));
 AND2x2_ASAP7_75t_R _1138_ (.A(net16),
    .B(_0672_),
    .Y(_0684_));
 AO21x1_ASAP7_75t_R _1139_ (.A1(net173),
    .A2(_0661_),
    .B(_0684_),
    .Y(_0685_));
 OA222x2_ASAP7_75t_R _1140_ (.A1(net57),
    .A2(_0671_),
    .B1(_0664_),
    .B2(_0685_),
    .C1(_0675_),
    .C2(net214),
    .Y(net294));
 BUFx6f_ASAP7_75t_R _1141_ (.A(_0643_),
    .Y(_0686_));
 AND2x2_ASAP7_75t_R _1142_ (.A(net17),
    .B(_0672_),
    .Y(_0687_));
 AO21x1_ASAP7_75t_R _1143_ (.A1(net174),
    .A2(_0686_),
    .B(_0687_),
    .Y(_0688_));
 OA222x2_ASAP7_75t_R _1144_ (.A1(net58),
    .A2(_0671_),
    .B1(_0664_),
    .B2(_0688_),
    .C1(_0675_),
    .C2(net215),
    .Y(net295));
 BUFx6f_ASAP7_75t_R _1145_ (.A(_0640_),
    .Y(_0689_));
 AND2x2_ASAP7_75t_R _1146_ (.A(net18),
    .B(_0672_),
    .Y(_0690_));
 AO21x1_ASAP7_75t_R _1147_ (.A1(net175),
    .A2(_0686_),
    .B(_0690_),
    .Y(_0691_));
 OA222x2_ASAP7_75t_R _1148_ (.A1(net59),
    .A2(_0671_),
    .B1(_0689_),
    .B2(_0691_),
    .C1(_0675_),
    .C2(net216),
    .Y(net296));
 AND2x2_ASAP7_75t_R _1149_ (.A(net19),
    .B(_0672_),
    .Y(_0692_));
 AO21x1_ASAP7_75t_R _1150_ (.A1(net176),
    .A2(_0686_),
    .B(_0692_),
    .Y(_0693_));
 OA222x2_ASAP7_75t_R _1151_ (.A1(net60),
    .A2(_0671_),
    .B1(_0689_),
    .B2(_0693_),
    .C1(_0675_),
    .C2(net217),
    .Y(net297));
 AND2x2_ASAP7_75t_R _1152_ (.A(net20),
    .B(_0672_),
    .Y(_0694_));
 AO21x1_ASAP7_75t_R _1153_ (.A1(net177),
    .A2(_0686_),
    .B(_0694_),
    .Y(_0695_));
 OA222x2_ASAP7_75t_R _1154_ (.A1(net61),
    .A2(_0671_),
    .B1(_0689_),
    .B2(_0695_),
    .C1(_0675_),
    .C2(net218),
    .Y(net298));
 BUFx6f_ASAP7_75t_R _1155_ (.A(_0638_),
    .Y(_0696_));
 BUFx6f_ASAP7_75t_R _1156_ (.A(_0645_),
    .Y(_0108_));
 AND2x2_ASAP7_75t_R _1157_ (.A(net21),
    .B(_0108_),
    .Y(_0109_));
 AO21x1_ASAP7_75t_R _1158_ (.A1(net178),
    .A2(_0686_),
    .B(_0109_),
    .Y(_0110_));
 BUFx6f_ASAP7_75t_R _1159_ (.A(_0649_),
    .Y(_0111_));
 OA222x2_ASAP7_75t_R _1160_ (.A1(net62),
    .A2(_0696_),
    .B1(_0689_),
    .B2(_0110_),
    .C1(_0111_),
    .C2(net219),
    .Y(net299));
 AND2x2_ASAP7_75t_R _1161_ (.A(net22),
    .B(_0108_),
    .Y(_0112_));
 AO21x1_ASAP7_75t_R _1162_ (.A1(net179),
    .A2(_0686_),
    .B(_0112_),
    .Y(_0113_));
 OA222x2_ASAP7_75t_R _1163_ (.A1(net63),
    .A2(_0696_),
    .B1(_0689_),
    .B2(_0113_),
    .C1(_0111_),
    .C2(net220),
    .Y(net300));
 AND2x2_ASAP7_75t_R _1164_ (.A(net23),
    .B(_0108_),
    .Y(_0114_));
 AO21x1_ASAP7_75t_R _1165_ (.A1(net180),
    .A2(_0686_),
    .B(_0114_),
    .Y(_0115_));
 OA222x2_ASAP7_75t_R _1166_ (.A1(net33),
    .A2(_0696_),
    .B1(_0689_),
    .B2(_0115_),
    .C1(_0111_),
    .C2(net190),
    .Y(net301));
 AND2x2_ASAP7_75t_R _1167_ (.A(net24),
    .B(_0108_),
    .Y(_0116_));
 AO21x1_ASAP7_75t_R _1168_ (.A1(net181),
    .A2(_0686_),
    .B(_0116_),
    .Y(_0117_));
 OA222x2_ASAP7_75t_R _1169_ (.A1(net64),
    .A2(_0696_),
    .B1(_0689_),
    .B2(_0117_),
    .C1(_0111_),
    .C2(net221),
    .Y(net302));
 AND2x2_ASAP7_75t_R _1170_ (.A(net25),
    .B(_0108_),
    .Y(_0118_));
 AO21x1_ASAP7_75t_R _1171_ (.A1(net182),
    .A2(_0686_),
    .B(_0118_),
    .Y(_0119_));
 OA222x2_ASAP7_75t_R _1172_ (.A1(net65),
    .A2(_0696_),
    .B1(_0689_),
    .B2(_0119_),
    .C1(_0111_),
    .C2(net222),
    .Y(net303));
 OAI22x1_ASAP7_75t_R _1173_ (.A1(net223),
    .A2(_0638_),
    .B1(_0640_),
    .B2(net183),
    .Y(_0120_));
 NAND2x1_ASAP7_75t_R _1174_ (.A(_0644_),
    .B(_0120_),
    .Y(net304));
 OA21x2_ASAP7_75t_R _1175_ (.A1(net225),
    .A2(_0704_),
    .B(_0644_),
    .Y(_0121_));
 OA21x2_ASAP7_75t_R _1176_ (.A1(net184),
    .A2(_0641_),
    .B(_0121_),
    .Y(net305));
 OA21x2_ASAP7_75t_R _1177_ (.A1(net226),
    .A2(_0704_),
    .B(_0644_),
    .Y(_0122_));
 OA21x2_ASAP7_75t_R _1178_ (.A1(net185),
    .A2(_0641_),
    .B(_0122_),
    .Y(net306));
 OA21x2_ASAP7_75t_R _1179_ (.A1(net227),
    .A2(_0704_),
    .B(_0644_),
    .Y(_0123_));
 OA21x2_ASAP7_75t_R _1180_ (.A1(net186),
    .A2(_0641_),
    .B(_0123_),
    .Y(net307));
 AND2x2_ASAP7_75t_R _1181_ (.A(net30),
    .B(_0108_),
    .Y(_0124_));
 AO21x1_ASAP7_75t_R _1182_ (.A1(net187),
    .A2(_0686_),
    .B(_0124_),
    .Y(_0125_));
 OA222x2_ASAP7_75t_R _1183_ (.A1(net71),
    .A2(_0696_),
    .B1(_0689_),
    .B2(_0125_),
    .C1(_0111_),
    .C2(net228),
    .Y(net308));
 AND2x2_ASAP7_75t_R _1184_ (.A(net34),
    .B(_0108_),
    .Y(_0126_));
 AO21x1_ASAP7_75t_R _1185_ (.A1(net191),
    .A2(_0643_),
    .B(_0126_),
    .Y(_0127_));
 OA222x2_ASAP7_75t_R _1186_ (.A1(net35),
    .A2(_0696_),
    .B1(_0689_),
    .B2(_0127_),
    .C1(_0111_),
    .C2(net192),
    .Y(net309));
 AND2x2_ASAP7_75t_R _1187_ (.A(net45),
    .B(_0108_),
    .Y(_0128_));
 AO21x1_ASAP7_75t_R _1188_ (.A1(net202),
    .A2(_0643_),
    .B(_0128_),
    .Y(_0129_));
 OA222x2_ASAP7_75t_R _1189_ (.A1(net36),
    .A2(_0696_),
    .B1(_0640_),
    .B2(_0129_),
    .C1(_0111_),
    .C2(net193),
    .Y(net310));
 AND2x2_ASAP7_75t_R _1190_ (.A(net56),
    .B(_0108_),
    .Y(_0130_));
 AO21x1_ASAP7_75t_R _1191_ (.A1(net213),
    .A2(_0643_),
    .B(_0130_),
    .Y(_0131_));
 OA222x2_ASAP7_75t_R _1192_ (.A1(net37),
    .A2(_0696_),
    .B1(_0640_),
    .B2(_0131_),
    .C1(_0111_),
    .C2(net194),
    .Y(net311));
 AND2x2_ASAP7_75t_R _1193_ (.A(net67),
    .B(_0108_),
    .Y(_0132_));
 AO21x1_ASAP7_75t_R _1194_ (.A1(net224),
    .A2(_0643_),
    .B(_0132_),
    .Y(_0133_));
 OA222x2_ASAP7_75t_R _1195_ (.A1(net38),
    .A2(_0696_),
    .B1(_0640_),
    .B2(_0133_),
    .C1(_0111_),
    .C2(net195),
    .Y(net312));
 AND2x2_ASAP7_75t_R _1196_ (.A(net72),
    .B(_0645_),
    .Y(_0134_));
 AO21x1_ASAP7_75t_R _1197_ (.A1(net229),
    .A2(_0643_),
    .B(_0134_),
    .Y(_0135_));
 OA222x2_ASAP7_75t_R _1198_ (.A1(net39),
    .A2(_0638_),
    .B1(_0640_),
    .B2(_0135_),
    .C1(_0649_),
    .C2(net196),
    .Y(net313));
 AND2x2_ASAP7_75t_R _1199_ (.A(net73),
    .B(_0645_),
    .Y(_0136_));
 AO21x1_ASAP7_75t_R _1200_ (.A1(net230),
    .A2(_0643_),
    .B(_0136_),
    .Y(_0137_));
 OA222x2_ASAP7_75t_R _1201_ (.A1(net40),
    .A2(_0638_),
    .B1(_0640_),
    .B2(_0137_),
    .C1(_0649_),
    .C2(net197),
    .Y(net314));
 AND2x2_ASAP7_75t_R _1202_ (.A(net74),
    .B(_0645_),
    .Y(_0138_));
 AO21x1_ASAP7_75t_R _1203_ (.A1(net231),
    .A2(_0643_),
    .B(_0138_),
    .Y(_0139_));
 OA222x2_ASAP7_75t_R _1204_ (.A1(net41),
    .A2(_0638_),
    .B1(_0640_),
    .B2(_0139_),
    .C1(_0649_),
    .C2(net198),
    .Y(net315));
 NAND2x2_ASAP7_75t_R _1205_ (.A(_0369_),
    .B(_0355_),
    .Y(_0140_));
 BUFx12f_ASAP7_75t_R _1206_ (.A(_0140_),
    .Y(_0141_));
 NAND2x2_ASAP7_75t_R _1207_ (.A(_0366_),
    .B(_0141_),
    .Y(_0142_));
 BUFx6f_ASAP7_75t_R _1208_ (.A(_0142_),
    .Y(_0143_));
 AND2x6_ASAP7_75t_R _1209_ (.A(_0350_),
    .B(_0140_),
    .Y(_0144_));
 BUFx6f_ASAP7_75t_R _1210_ (.A(_0144_),
    .Y(_0145_));
 NAND2x1_ASAP7_75t_R _1211_ (.A(_0350_),
    .B(_0140_),
    .Y(_0146_));
 BUFx6f_ASAP7_75t_R _1212_ (.A(_0146_),
    .Y(_0147_));
 AND2x2_ASAP7_75t_R _1213_ (.A(net31),
    .B(_0147_),
    .Y(_0148_));
 AO21x1_ASAP7_75t_R _1214_ (.A1(net109),
    .A2(_0145_),
    .B(_0148_),
    .Y(_0149_));
 BUFx3_ASAP7_75t_R _1215_ (.A(_0141_),
    .Y(_0150_));
 BUFx12f_ASAP7_75t_R _1216_ (.A(_0146_),
    .Y(_0151_));
 BUFx6f_ASAP7_75t_R _1217_ (.A(_0151_),
    .Y(_0152_));
 BUFx6f_ASAP7_75t_R _1218_ (.A(_0350_),
    .Y(_0153_));
 BUFx6f_ASAP7_75t_R _1219_ (.A(_0153_),
    .Y(_0154_));
 BUFx6f_ASAP7_75t_R _1220_ (.A(_0140_),
    .Y(_0155_));
 AND3x1_ASAP7_75t_R _1221_ (.A(net79),
    .B(_0154_),
    .C(_0155_),
    .Y(_0156_));
 AO221x1_ASAP7_75t_R _1222_ (.A1(net358),
    .A2(_0150_),
    .B1(_0152_),
    .B2(net1),
    .C(_0156_),
    .Y(_0157_));
 OA21x2_ASAP7_75t_R _1223_ (.A1(_0143_),
    .A2(_0149_),
    .B(_0157_),
    .Y(net320));
 AND2x2_ASAP7_75t_R _1224_ (.A(net42),
    .B(_0147_),
    .Y(_0158_));
 AO21x1_ASAP7_75t_R _1225_ (.A1(net120),
    .A2(_0145_),
    .B(_0158_),
    .Y(_0159_));
 AND3x1_ASAP7_75t_R _1226_ (.A(net80),
    .B(_0154_),
    .C(_0155_),
    .Y(_0160_));
 AO221x1_ASAP7_75t_R _1227_ (.A1(net358),
    .A2(_0150_),
    .B1(_0152_),
    .B2(net2),
    .C(_0160_),
    .Y(_0161_));
 OA21x2_ASAP7_75t_R _1228_ (.A1(_0143_),
    .A2(_0159_),
    .B(_0161_),
    .Y(net321));
 AND2x2_ASAP7_75t_R _1229_ (.A(net43),
    .B(_0147_),
    .Y(_0162_));
 AO21x1_ASAP7_75t_R _1230_ (.A1(net121),
    .A2(_0145_),
    .B(_0162_),
    .Y(_0163_));
 AND3x1_ASAP7_75t_R _1231_ (.A(net81),
    .B(_0154_),
    .C(_0155_),
    .Y(_0164_));
 AO221x1_ASAP7_75t_R _1232_ (.A1(net358),
    .A2(_0150_),
    .B1(_0152_),
    .B2(net3),
    .C(_0164_),
    .Y(_0165_));
 OA21x2_ASAP7_75t_R _1233_ (.A1(_0143_),
    .A2(_0163_),
    .B(_0165_),
    .Y(net322));
 BUFx6f_ASAP7_75t_R _1234_ (.A(_0151_),
    .Y(_0166_));
 AND2x2_ASAP7_75t_R _1235_ (.A(net44),
    .B(_0166_),
    .Y(_0167_));
 AO21x1_ASAP7_75t_R _1236_ (.A1(net122),
    .A2(_0145_),
    .B(_0167_),
    .Y(_0168_));
 BUFx6f_ASAP7_75t_R _1237_ (.A(_0141_),
    .Y(_0169_));
 AND3x1_ASAP7_75t_R _1238_ (.A(net82),
    .B(_0154_),
    .C(_0169_),
    .Y(_0170_));
 AO221x1_ASAP7_75t_R _1239_ (.A1(net358),
    .A2(_0150_),
    .B1(_0152_),
    .B2(net4),
    .C(_0170_),
    .Y(_0171_));
 OA21x2_ASAP7_75t_R _1240_ (.A1(_0143_),
    .A2(_0168_),
    .B(_0171_),
    .Y(net323));
 AND2x2_ASAP7_75t_R _1241_ (.A(net46),
    .B(_0166_),
    .Y(_0172_));
 AO21x1_ASAP7_75t_R _1242_ (.A1(net124),
    .A2(_0145_),
    .B(_0172_),
    .Y(_0173_));
 AND3x1_ASAP7_75t_R _1243_ (.A(net83),
    .B(_0154_),
    .C(_0169_),
    .Y(_0174_));
 AO221x1_ASAP7_75t_R _1244_ (.A1(net358),
    .A2(_0150_),
    .B1(_0152_),
    .B2(net5),
    .C(_0174_),
    .Y(_0175_));
 OA21x2_ASAP7_75t_R _1245_ (.A1(_0143_),
    .A2(_0173_),
    .B(_0175_),
    .Y(net324));
 AND2x2_ASAP7_75t_R _1246_ (.A(net47),
    .B(_0166_),
    .Y(_0176_));
 AO21x1_ASAP7_75t_R _1247_ (.A1(net125),
    .A2(_0145_),
    .B(_0176_),
    .Y(_0177_));
 AND3x1_ASAP7_75t_R _1248_ (.A(net84),
    .B(_0154_),
    .C(_0169_),
    .Y(_0178_));
 AO221x1_ASAP7_75t_R _1249_ (.A1(net358),
    .A2(_0150_),
    .B1(_0152_),
    .B2(net6),
    .C(_0178_),
    .Y(_0179_));
 OA21x2_ASAP7_75t_R _1250_ (.A1(_0143_),
    .A2(_0177_),
    .B(_0179_),
    .Y(net325));
 AND2x2_ASAP7_75t_R _1251_ (.A(net48),
    .B(_0166_),
    .Y(_0180_));
 AO21x1_ASAP7_75t_R _1252_ (.A1(net126),
    .A2(_0145_),
    .B(_0180_),
    .Y(_0181_));
 AND3x1_ASAP7_75t_R _1253_ (.A(net85),
    .B(_0154_),
    .C(_0169_),
    .Y(_0182_));
 AO221x1_ASAP7_75t_R _1254_ (.A1(net358),
    .A2(_0150_),
    .B1(_0152_),
    .B2(net7),
    .C(_0182_),
    .Y(_0183_));
 OA21x2_ASAP7_75t_R _1255_ (.A1(_0143_),
    .A2(_0181_),
    .B(_0183_),
    .Y(net326));
 AND2x2_ASAP7_75t_R _1256_ (.A(net49),
    .B(_0166_),
    .Y(_0184_));
 AO21x1_ASAP7_75t_R _1257_ (.A1(net127),
    .A2(_0145_),
    .B(_0184_),
    .Y(_0185_));
 AND3x1_ASAP7_75t_R _1258_ (.A(net86),
    .B(_0154_),
    .C(_0169_),
    .Y(_0186_));
 AO221x1_ASAP7_75t_R _1259_ (.A1(net358),
    .A2(_0150_),
    .B1(_0152_),
    .B2(net8),
    .C(_0186_),
    .Y(_0187_));
 OA21x2_ASAP7_75t_R _1260_ (.A1(_0143_),
    .A2(_0185_),
    .B(_0187_),
    .Y(net327));
 AND2x2_ASAP7_75t_R _1261_ (.A(net50),
    .B(_0166_),
    .Y(_0188_));
 AO21x1_ASAP7_75t_R _1262_ (.A1(net128),
    .A2(_0145_),
    .B(_0188_),
    .Y(_0189_));
 BUFx6f_ASAP7_75t_R _1263_ (.A(_0366_),
    .Y(_0190_));
 AND3x1_ASAP7_75t_R _1264_ (.A(net87),
    .B(_0154_),
    .C(_0169_),
    .Y(_0191_));
 AO221x1_ASAP7_75t_R _1265_ (.A1(_0190_),
    .A2(_0150_),
    .B1(_0152_),
    .B2(net9),
    .C(_0191_),
    .Y(_0192_));
 OA21x2_ASAP7_75t_R _1266_ (.A1(_0143_),
    .A2(_0189_),
    .B(_0192_),
    .Y(net328));
 AND2x2_ASAP7_75t_R _1267_ (.A(net51),
    .B(_0166_),
    .Y(_0193_));
 AO21x1_ASAP7_75t_R _1268_ (.A1(net129),
    .A2(_0145_),
    .B(_0193_),
    .Y(_0194_));
 AND3x1_ASAP7_75t_R _1269_ (.A(net88),
    .B(_0154_),
    .C(_0169_),
    .Y(_0195_));
 AO221x1_ASAP7_75t_R _1270_ (.A1(_0190_),
    .A2(_0150_),
    .B1(_0152_),
    .B2(net10),
    .C(_0195_),
    .Y(_0196_));
 OA21x2_ASAP7_75t_R _1271_ (.A1(_0143_),
    .A2(_0194_),
    .B(_0196_),
    .Y(net329));
 BUFx6f_ASAP7_75t_R _1272_ (.A(_0142_),
    .Y(_0197_));
 BUFx6f_ASAP7_75t_R _1273_ (.A(_0144_),
    .Y(_0198_));
 AND2x2_ASAP7_75t_R _1274_ (.A(net52),
    .B(_0166_),
    .Y(_0199_));
 AO21x1_ASAP7_75t_R _1275_ (.A1(net130),
    .A2(_0198_),
    .B(_0199_),
    .Y(_0200_));
 BUFx6f_ASAP7_75t_R _1276_ (.A(_0141_),
    .Y(_0201_));
 BUFx6f_ASAP7_75t_R _1277_ (.A(_0151_),
    .Y(_0202_));
 BUFx6f_ASAP7_75t_R _1278_ (.A(_0153_),
    .Y(_0203_));
 AND3x1_ASAP7_75t_R _1279_ (.A(net89),
    .B(_0203_),
    .C(_0169_),
    .Y(_0204_));
 AO221x1_ASAP7_75t_R _1280_ (.A1(_0190_),
    .A2(_0201_),
    .B1(_0202_),
    .B2(net11),
    .C(_0204_),
    .Y(_0205_));
 OA21x2_ASAP7_75t_R _1281_ (.A1(_0197_),
    .A2(_0200_),
    .B(_0205_),
    .Y(net330));
 AND2x2_ASAP7_75t_R _1282_ (.A(net32),
    .B(_0166_),
    .Y(_0206_));
 AO21x1_ASAP7_75t_R _1283_ (.A1(net110),
    .A2(_0198_),
    .B(_0206_),
    .Y(_0207_));
 AND3x1_ASAP7_75t_R _1284_ (.A(net90),
    .B(_0203_),
    .C(_0169_),
    .Y(_0208_));
 AO221x1_ASAP7_75t_R _1285_ (.A1(_0190_),
    .A2(_0201_),
    .B1(_0202_),
    .B2(net12),
    .C(_0208_),
    .Y(_0209_));
 OA21x2_ASAP7_75t_R _1286_ (.A1(_0197_),
    .A2(_0207_),
    .B(_0209_),
    .Y(net331));
 AND2x2_ASAP7_75t_R _1287_ (.A(net53),
    .B(_0166_),
    .Y(_0210_));
 AO21x1_ASAP7_75t_R _1288_ (.A1(net131),
    .A2(_0198_),
    .B(_0210_),
    .Y(_0211_));
 AND3x1_ASAP7_75t_R _1289_ (.A(net91),
    .B(_0203_),
    .C(_0169_),
    .Y(_0212_));
 AO221x1_ASAP7_75t_R _1290_ (.A1(_0190_),
    .A2(_0201_),
    .B1(_0202_),
    .B2(net13),
    .C(_0212_),
    .Y(_0213_));
 OA21x2_ASAP7_75t_R _1291_ (.A1(_0197_),
    .A2(_0211_),
    .B(_0213_),
    .Y(net332));
 BUFx6f_ASAP7_75t_R _1292_ (.A(_0151_),
    .Y(_0214_));
 AND2x2_ASAP7_75t_R _1293_ (.A(net54),
    .B(_0214_),
    .Y(_0215_));
 AO21x1_ASAP7_75t_R _1294_ (.A1(net132),
    .A2(_0198_),
    .B(_0215_),
    .Y(_0216_));
 BUFx6f_ASAP7_75t_R _1295_ (.A(_0141_),
    .Y(_0217_));
 AND3x1_ASAP7_75t_R _1296_ (.A(net92),
    .B(_0203_),
    .C(_0217_),
    .Y(_0218_));
 AO221x1_ASAP7_75t_R _1297_ (.A1(_0190_),
    .A2(_0201_),
    .B1(_0202_),
    .B2(net14),
    .C(_0218_),
    .Y(_0219_));
 OA21x2_ASAP7_75t_R _1298_ (.A1(_0197_),
    .A2(_0216_),
    .B(_0219_),
    .Y(net333));
 AND2x2_ASAP7_75t_R _1299_ (.A(net55),
    .B(_0214_),
    .Y(_0220_));
 AO21x1_ASAP7_75t_R _1300_ (.A1(net133),
    .A2(_0198_),
    .B(_0220_),
    .Y(_0221_));
 AND3x1_ASAP7_75t_R _1301_ (.A(net93),
    .B(_0203_),
    .C(_0217_),
    .Y(_0222_));
 AO221x1_ASAP7_75t_R _1302_ (.A1(_0190_),
    .A2(_0201_),
    .B1(_0202_),
    .B2(net15),
    .C(_0222_),
    .Y(_0223_));
 OA21x2_ASAP7_75t_R _1303_ (.A1(_0197_),
    .A2(_0221_),
    .B(_0223_),
    .Y(net334));
 AND2x2_ASAP7_75t_R _1304_ (.A(net57),
    .B(_0214_),
    .Y(_0224_));
 AO21x1_ASAP7_75t_R _1305_ (.A1(net135),
    .A2(_0198_),
    .B(_0224_),
    .Y(_0225_));
 AND3x1_ASAP7_75t_R _1306_ (.A(net94),
    .B(_0203_),
    .C(_0217_),
    .Y(_0226_));
 AO221x1_ASAP7_75t_R _1307_ (.A1(_0190_),
    .A2(_0201_),
    .B1(_0202_),
    .B2(net16),
    .C(_0226_),
    .Y(_0227_));
 OA21x2_ASAP7_75t_R _1308_ (.A1(_0197_),
    .A2(_0225_),
    .B(_0227_),
    .Y(net335));
 AND2x2_ASAP7_75t_R _1309_ (.A(net58),
    .B(_0214_),
    .Y(_0228_));
 AO21x1_ASAP7_75t_R _1310_ (.A1(net136),
    .A2(_0198_),
    .B(_0228_),
    .Y(_0229_));
 AND3x1_ASAP7_75t_R _1311_ (.A(net95),
    .B(_0203_),
    .C(_0217_),
    .Y(_0230_));
 AO221x1_ASAP7_75t_R _1312_ (.A1(_0190_),
    .A2(_0201_),
    .B1(_0202_),
    .B2(net17),
    .C(_0230_),
    .Y(_0231_));
 OA21x2_ASAP7_75t_R _1313_ (.A1(_0197_),
    .A2(_0229_),
    .B(_0231_),
    .Y(net336));
 AND2x2_ASAP7_75t_R _1314_ (.A(net59),
    .B(_0214_),
    .Y(_0232_));
 AO21x1_ASAP7_75t_R _1315_ (.A1(net137),
    .A2(_0198_),
    .B(_0232_),
    .Y(_0233_));
 AND3x1_ASAP7_75t_R _1316_ (.A(net96),
    .B(_0203_),
    .C(_0217_),
    .Y(_0234_));
 AO221x1_ASAP7_75t_R _1317_ (.A1(_0190_),
    .A2(_0201_),
    .B1(_0202_),
    .B2(net18),
    .C(_0234_),
    .Y(_0235_));
 OA21x2_ASAP7_75t_R _1318_ (.A1(_0197_),
    .A2(_0233_),
    .B(_0235_),
    .Y(net337));
 AND2x2_ASAP7_75t_R _1319_ (.A(net60),
    .B(_0214_),
    .Y(_0236_));
 AO21x1_ASAP7_75t_R _1320_ (.A1(net138),
    .A2(_0198_),
    .B(_0236_),
    .Y(_0237_));
 BUFx6f_ASAP7_75t_R _1321_ (.A(_0366_),
    .Y(_0238_));
 AND3x1_ASAP7_75t_R _1322_ (.A(net97),
    .B(_0203_),
    .C(_0217_),
    .Y(_0239_));
 AO221x1_ASAP7_75t_R _1323_ (.A1(_0238_),
    .A2(_0201_),
    .B1(_0202_),
    .B2(net19),
    .C(_0239_),
    .Y(_0240_));
 OA21x2_ASAP7_75t_R _1324_ (.A1(_0197_),
    .A2(_0237_),
    .B(_0240_),
    .Y(net338));
 AND2x2_ASAP7_75t_R _1325_ (.A(net61),
    .B(_0214_),
    .Y(_0241_));
 AO21x1_ASAP7_75t_R _1326_ (.A1(net139),
    .A2(_0198_),
    .B(_0241_),
    .Y(_0242_));
 AND3x1_ASAP7_75t_R _1327_ (.A(net98),
    .B(_0203_),
    .C(_0217_),
    .Y(_0243_));
 AO221x1_ASAP7_75t_R _1328_ (.A1(_0238_),
    .A2(_0201_),
    .B1(_0202_),
    .B2(net20),
    .C(_0243_),
    .Y(_0244_));
 OA21x2_ASAP7_75t_R _1329_ (.A1(_0197_),
    .A2(_0242_),
    .B(_0244_),
    .Y(net339));
 BUFx6f_ASAP7_75t_R _1330_ (.A(_0142_),
    .Y(_0245_));
 BUFx6f_ASAP7_75t_R _1331_ (.A(_0144_),
    .Y(_0246_));
 AND2x2_ASAP7_75t_R _1332_ (.A(net62),
    .B(_0214_),
    .Y(_0247_));
 AO21x1_ASAP7_75t_R _1333_ (.A1(net140),
    .A2(_0246_),
    .B(_0247_),
    .Y(_0248_));
 BUFx6f_ASAP7_75t_R _1334_ (.A(_0141_),
    .Y(_0249_));
 BUFx6f_ASAP7_75t_R _1335_ (.A(_0151_),
    .Y(_0250_));
 BUFx6f_ASAP7_75t_R _1336_ (.A(_0153_),
    .Y(_0251_));
 AND3x1_ASAP7_75t_R _1337_ (.A(net99),
    .B(_0251_),
    .C(_0217_),
    .Y(_0252_));
 AO221x1_ASAP7_75t_R _1338_ (.A1(_0238_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net21),
    .C(_0252_),
    .Y(_0253_));
 OA21x2_ASAP7_75t_R _1339_ (.A1(_0245_),
    .A2(_0248_),
    .B(_0253_),
    .Y(net340));
 AND2x2_ASAP7_75t_R _1340_ (.A(net63),
    .B(_0214_),
    .Y(_0254_));
 AO21x1_ASAP7_75t_R _1341_ (.A1(net141),
    .A2(_0246_),
    .B(_0254_),
    .Y(_0255_));
 AND3x1_ASAP7_75t_R _1342_ (.A(net100),
    .B(_0251_),
    .C(_0217_),
    .Y(_0256_));
 AO221x1_ASAP7_75t_R _1343_ (.A1(_0238_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net22),
    .C(_0256_),
    .Y(_0257_));
 OA21x2_ASAP7_75t_R _1344_ (.A1(_0245_),
    .A2(_0255_),
    .B(_0257_),
    .Y(net341));
 AND2x2_ASAP7_75t_R _1345_ (.A(net33),
    .B(_0214_),
    .Y(_0258_));
 AO21x1_ASAP7_75t_R _1346_ (.A1(net111),
    .A2(_0246_),
    .B(_0258_),
    .Y(_0259_));
 AND3x1_ASAP7_75t_R _1347_ (.A(net101),
    .B(_0251_),
    .C(_0217_),
    .Y(_0260_));
 AO221x1_ASAP7_75t_R _1348_ (.A1(_0238_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net23),
    .C(_0260_),
    .Y(_0261_));
 OA21x2_ASAP7_75t_R _1349_ (.A1(_0245_),
    .A2(_0259_),
    .B(_0261_),
    .Y(net342));
 BUFx6f_ASAP7_75t_R _1350_ (.A(_0151_),
    .Y(_0262_));
 AND2x2_ASAP7_75t_R _1351_ (.A(net64),
    .B(_0262_),
    .Y(_0263_));
 AO21x1_ASAP7_75t_R _1352_ (.A1(net142),
    .A2(_0246_),
    .B(_0263_),
    .Y(_0264_));
 BUFx6f_ASAP7_75t_R _1353_ (.A(_0140_),
    .Y(_0265_));
 AND3x1_ASAP7_75t_R _1354_ (.A(net102),
    .B(_0251_),
    .C(_0265_),
    .Y(_0266_));
 AO221x1_ASAP7_75t_R _1355_ (.A1(_0238_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net24),
    .C(_0266_),
    .Y(_0267_));
 OA21x2_ASAP7_75t_R _1356_ (.A1(_0245_),
    .A2(_0264_),
    .B(_0267_),
    .Y(net343));
 AND2x2_ASAP7_75t_R _1357_ (.A(net65),
    .B(_0262_),
    .Y(_0268_));
 AO21x1_ASAP7_75t_R _1358_ (.A1(net143),
    .A2(_0246_),
    .B(_0268_),
    .Y(_0269_));
 AND3x1_ASAP7_75t_R _1359_ (.A(net103),
    .B(_0251_),
    .C(_0265_),
    .Y(_0270_));
 AO221x1_ASAP7_75t_R _1360_ (.A1(_0238_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net25),
    .C(_0270_),
    .Y(_0271_));
 OA21x2_ASAP7_75t_R _1361_ (.A1(_0245_),
    .A2(_0269_),
    .B(_0271_),
    .Y(net344));
 AND2x2_ASAP7_75t_R _1362_ (.A(net66),
    .B(_0262_),
    .Y(_0272_));
 AO21x1_ASAP7_75t_R _1363_ (.A1(net144),
    .A2(_0246_),
    .B(_0272_),
    .Y(_0273_));
 AND3x1_ASAP7_75t_R _1364_ (.A(net104),
    .B(_0251_),
    .C(_0265_),
    .Y(_0274_));
 AO221x1_ASAP7_75t_R _1365_ (.A1(_0238_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net26),
    .C(_0274_),
    .Y(_0275_));
 OA21x2_ASAP7_75t_R _1366_ (.A1(_0245_),
    .A2(_0273_),
    .B(_0275_),
    .Y(net345));
 AND2x2_ASAP7_75t_R _1367_ (.A(net68),
    .B(_0262_),
    .Y(_0276_));
 AO21x1_ASAP7_75t_R _1368_ (.A1(net146),
    .A2(_0246_),
    .B(_0276_),
    .Y(_0277_));
 AND3x1_ASAP7_75t_R _1369_ (.A(net105),
    .B(_0251_),
    .C(_0265_),
    .Y(_0278_));
 AO221x1_ASAP7_75t_R _1370_ (.A1(_0238_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net27),
    .C(_0278_),
    .Y(_0279_));
 OA21x2_ASAP7_75t_R _1371_ (.A1(_0245_),
    .A2(_0277_),
    .B(_0279_),
    .Y(net346));
 AND2x2_ASAP7_75t_R _1372_ (.A(net69),
    .B(_0262_),
    .Y(_0280_));
 AO21x1_ASAP7_75t_R _1373_ (.A1(net147),
    .A2(_0246_),
    .B(_0280_),
    .Y(_0281_));
 AND3x1_ASAP7_75t_R _1374_ (.A(net106),
    .B(_0251_),
    .C(_0265_),
    .Y(_0282_));
 AO221x1_ASAP7_75t_R _1375_ (.A1(_0238_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net28),
    .C(_0282_),
    .Y(_0283_));
 OA21x2_ASAP7_75t_R _1376_ (.A1(_0245_),
    .A2(_0281_),
    .B(_0283_),
    .Y(net347));
 AND2x2_ASAP7_75t_R _1377_ (.A(net70),
    .B(_0262_),
    .Y(_0284_));
 AO21x1_ASAP7_75t_R _1378_ (.A1(net148),
    .A2(_0246_),
    .B(_0284_),
    .Y(_0285_));
 AND3x1_ASAP7_75t_R _1379_ (.A(net107),
    .B(_0251_),
    .C(_0265_),
    .Y(_0286_));
 AO221x1_ASAP7_75t_R _1380_ (.A1(_0367_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net29),
    .C(_0286_),
    .Y(_0287_));
 OA21x2_ASAP7_75t_R _1381_ (.A1(_0245_),
    .A2(_0285_),
    .B(_0287_),
    .Y(net348));
 AND2x2_ASAP7_75t_R _1382_ (.A(net71),
    .B(_0262_),
    .Y(_0288_));
 AO21x1_ASAP7_75t_R _1383_ (.A1(net149),
    .A2(_0246_),
    .B(_0288_),
    .Y(_0289_));
 AND3x1_ASAP7_75t_R _1384_ (.A(net108),
    .B(_0251_),
    .C(_0265_),
    .Y(_0290_));
 AO221x1_ASAP7_75t_R _1385_ (.A1(_0367_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(net30),
    .C(_0290_),
    .Y(_0291_));
 OA21x2_ASAP7_75t_R _1386_ (.A1(_0245_),
    .A2(_0289_),
    .B(_0291_),
    .Y(net349));
 AND2x2_ASAP7_75t_R _1387_ (.A(net35),
    .B(_0262_),
    .Y(_0292_));
 AO21x1_ASAP7_75t_R _1388_ (.A1(net113),
    .A2(_0144_),
    .B(_0292_),
    .Y(_0293_));
 AND3x1_ASAP7_75t_R _1389_ (.A(net112),
    .B(_0153_),
    .C(_0265_),
    .Y(_0294_));
 AO221x1_ASAP7_75t_R _1390_ (.A1(_0367_),
    .A2(_0155_),
    .B1(_0147_),
    .B2(net34),
    .C(_0294_),
    .Y(_0295_));
 OA21x2_ASAP7_75t_R _1391_ (.A1(_0142_),
    .A2(_0293_),
    .B(_0295_),
    .Y(net350));
 AND2x2_ASAP7_75t_R _1392_ (.A(net36),
    .B(_0262_),
    .Y(_0296_));
 AO21x1_ASAP7_75t_R _1393_ (.A1(net114),
    .A2(_0144_),
    .B(_0296_),
    .Y(_0297_));
 AND3x1_ASAP7_75t_R _1394_ (.A(net123),
    .B(_0153_),
    .C(_0265_),
    .Y(_0298_));
 AO221x1_ASAP7_75t_R _1395_ (.A1(_0367_),
    .A2(_0155_),
    .B1(_0147_),
    .B2(net45),
    .C(_0298_),
    .Y(_0299_));
 OA21x2_ASAP7_75t_R _1396_ (.A1(_0142_),
    .A2(_0297_),
    .B(_0299_),
    .Y(net351));
 AND2x2_ASAP7_75t_R _1397_ (.A(net37),
    .B(_0262_),
    .Y(_0300_));
 AO21x1_ASAP7_75t_R _1398_ (.A1(net115),
    .A2(_0144_),
    .B(_0300_),
    .Y(_0301_));
 AND3x1_ASAP7_75t_R _1399_ (.A(net134),
    .B(_0153_),
    .C(_0265_),
    .Y(_0302_));
 AO221x1_ASAP7_75t_R _1400_ (.A1(_0367_),
    .A2(_0155_),
    .B1(_0147_),
    .B2(net56),
    .C(_0302_),
    .Y(_0303_));
 OA21x2_ASAP7_75t_R _1401_ (.A1(_0142_),
    .A2(_0301_),
    .B(_0303_),
    .Y(net352));
 AND2x2_ASAP7_75t_R _1402_ (.A(net38),
    .B(_0151_),
    .Y(_0304_));
 AO21x1_ASAP7_75t_R _1403_ (.A1(net116),
    .A2(_0144_),
    .B(_0304_),
    .Y(_0305_));
 AND3x1_ASAP7_75t_R _1404_ (.A(net145),
    .B(_0153_),
    .C(_0141_),
    .Y(_0306_));
 AO221x1_ASAP7_75t_R _1405_ (.A1(_0367_),
    .A2(_0155_),
    .B1(_0147_),
    .B2(net67),
    .C(_0306_),
    .Y(_0307_));
 OA21x2_ASAP7_75t_R _1406_ (.A1(_0142_),
    .A2(_0305_),
    .B(_0307_),
    .Y(net353));
 AND2x2_ASAP7_75t_R _1407_ (.A(net39),
    .B(_0151_),
    .Y(_0308_));
 AO21x1_ASAP7_75t_R _1408_ (.A1(net117),
    .A2(_0144_),
    .B(_0308_),
    .Y(_0309_));
 AND3x1_ASAP7_75t_R _1409_ (.A(net150),
    .B(_0153_),
    .C(_0141_),
    .Y(_0310_));
 AO221x1_ASAP7_75t_R _1410_ (.A1(_0367_),
    .A2(_0155_),
    .B1(_0147_),
    .B2(net72),
    .C(_0310_),
    .Y(_0311_));
 OA21x2_ASAP7_75t_R _1411_ (.A1(_0142_),
    .A2(_0309_),
    .B(_0311_),
    .Y(net354));
 AND2x2_ASAP7_75t_R _1412_ (.A(net40),
    .B(_0151_),
    .Y(_0312_));
 AO21x1_ASAP7_75t_R _1413_ (.A1(net118),
    .A2(_0144_),
    .B(_0312_),
    .Y(_0313_));
 AND3x1_ASAP7_75t_R _1414_ (.A(net151),
    .B(_0153_),
    .C(_0141_),
    .Y(_0314_));
 AO221x1_ASAP7_75t_R _1415_ (.A1(_0367_),
    .A2(_0155_),
    .B1(_0147_),
    .B2(net73),
    .C(_0314_),
    .Y(_0315_));
 OA21x2_ASAP7_75t_R _1416_ (.A1(_0142_),
    .A2(_0313_),
    .B(_0315_),
    .Y(net355));
 AND2x2_ASAP7_75t_R _1417_ (.A(net41),
    .B(_0151_),
    .Y(_0316_));
 AO21x1_ASAP7_75t_R _1418_ (.A1(net119),
    .A2(_0144_),
    .B(_0316_),
    .Y(_0317_));
 AND3x1_ASAP7_75t_R _1419_ (.A(net152),
    .B(_0153_),
    .C(_0141_),
    .Y(_0318_));
 AO221x1_ASAP7_75t_R _1420_ (.A1(_0367_),
    .A2(_0155_),
    .B1(_0147_),
    .B2(net74),
    .C(_0318_),
    .Y(_0319_));
 OA21x2_ASAP7_75t_R _1421_ (.A1(_0142_),
    .A2(_0317_),
    .B(_0319_),
    .Y(net356));
 INVx1_ASAP7_75t_R _1422_ (.A(_0705_),
    .Y(\credit_t_route_inst.r_counters_inst.o_credits[1] ));
 INVx1_ASAP7_75t_R _1423_ (.A(_0063_),
    .Y(\credit_t_route_inst.r_counters_inst.o_credits[3] ));
 INVx1_ASAP7_75t_R _1424_ (.A(_0064_),
    .Y(\credit_t_route_inst.r_counters_inst.o_credits[2] ));
 OR3x2_ASAP7_75t_R _1425_ (.A(net28),
    .B(net27),
    .C(net29),
    .Y(_0320_));
 NAND2x1_ASAP7_75t_R _1426_ (.A(net75),
    .B(net26),
    .Y(_0321_));
 NOR2x1_ASAP7_75t_R _1427_ (.A(_0320_),
    .B(_0321_),
    .Y(_0322_));
 AO22x2_ASAP7_75t_R _1428_ (.A1(net232),
    .A2(net183),
    .B1(net233),
    .B2(net223),
    .Y(_0323_));
 NAND2x1_ASAP7_75t_R _1429_ (.A(_0021_),
    .B(_0323_),
    .Y(_0324_));
 AND2x4_ASAP7_75t_R _1430_ (.A(_0322_),
    .B(_0324_),
    .Y(_0325_));
 INVx2_ASAP7_75t_R _1431_ (.A(_0022_),
    .Y(_0326_));
 OR3x2_ASAP7_75t_R _1432_ (.A(net69),
    .B(net68),
    .C(net70),
    .Y(_0327_));
 NAND2x1_ASAP7_75t_R _1433_ (.A(net76),
    .B(net66),
    .Y(_0328_));
 OA22x2_ASAP7_75t_R _1434_ (.A1(_0320_),
    .A2(_0321_),
    .B1(_0327_),
    .B2(_0328_),
    .Y(_0329_));
 OA211x2_ASAP7_75t_R _1435_ (.A1(_0326_),
    .A2(_0329_),
    .B(net232),
    .C(net183),
    .Y(_0330_));
 AND5x2_ASAP7_75t_R _1436_ (.A(_0062_),
    .B(_0063_),
    .C(_0064_),
    .D(_0705_),
    .E(_0046_),
    .Y(_0331_));
 INVx2_ASAP7_75t_R _1437_ (.A(_0331_),
    .Y(_0332_));
 OAI21x1_ASAP7_75t_R _1438_ (.A1(_0325_),
    .A2(_0330_),
    .B(_0332_),
    .Y(_0706_));
 INVx1_ASAP7_75t_R _1439_ (.A(_0703_),
    .Y(\credit_t_route_inst.r_counters_inst.o_credits[6] ));
 INVx1_ASAP7_75t_R _1440_ (.A(_0060_),
    .Y(\credit_t_route_inst.r_counters_inst.o_credits[8] ));
 INVx1_ASAP7_75t_R _1441_ (.A(_0061_),
    .Y(\credit_t_route_inst.r_counters_inst.o_credits[7] ));
 NOR2x1_ASAP7_75t_R _1442_ (.A(_0327_),
    .B(_0328_),
    .Y(_0333_));
 AND5x2_ASAP7_75t_R _1443_ (.A(_0060_),
    .B(_0061_),
    .C(_0703_),
    .D(_0048_),
    .E(_0071_),
    .Y(_0334_));
 INVx1_ASAP7_75t_R _1444_ (.A(_0334_),
    .Y(_0335_));
 OR3x1_ASAP7_75t_R _1445_ (.A(_0331_),
    .B(_0320_),
    .C(_0321_),
    .Y(_0336_));
 AND4x1_ASAP7_75t_R _1446_ (.A(_0324_),
    .B(_0333_),
    .C(_0335_),
    .D(_0336_),
    .Y(_0337_));
 NAND2x1_ASAP7_75t_R _1447_ (.A(net232),
    .B(net183),
    .Y(_0338_));
 NAND2x1_ASAP7_75t_R _1448_ (.A(_0048_),
    .B(_0071_),
    .Y(_0339_));
 NAND3x1_ASAP7_75t_R _1449_ (.A(_0060_),
    .B(_0061_),
    .C(_0703_),
    .Y(_0340_));
 OA221x2_ASAP7_75t_R _1450_ (.A1(_0331_),
    .A2(_0338_),
    .B1(_0339_),
    .B2(_0340_),
    .C(net223),
    .Y(_0341_));
 OA211x2_ASAP7_75t_R _1451_ (.A1(_0326_),
    .A2(_0329_),
    .B(_0341_),
    .C(net233),
    .Y(_0342_));
 OR2x2_ASAP7_75t_R _1452_ (.A(_0337_),
    .B(_0342_),
    .Y(_0343_));
 BUFx6f_ASAP7_75t_R _1453_ (.A(_0343_),
    .Y(net317));
 INVx3_ASAP7_75t_R _1454_ (.A(net317),
    .Y(_0704_));
 INVx1_ASAP7_75t_R _1455_ (.A(_0701_),
    .Y(\credit_t_route_inst.u0_counters_inst.o_credits[6] ));
 INVx1_ASAP7_75t_R _1456_ (.A(_0055_),
    .Y(\credit_t_route_inst.u0_counters_inst.o_credits[8] ));
 INVx1_ASAP7_75t_R _1457_ (.A(_0056_),
    .Y(\credit_t_route_inst.u0_counters_inst.o_credits[7] ));
 INVx1_ASAP7_75t_R _1458_ (.A(_0707_),
    .Y(\credit_t_route_inst.u0_counters_inst.o_credits[1] ));
 INVx1_ASAP7_75t_R _1459_ (.A(_0058_),
    .Y(\credit_t_route_inst.u0_counters_inst.o_credits[3] ));
 INVx1_ASAP7_75t_R _1460_ (.A(_0059_),
    .Y(\credit_t_route_inst.u0_counters_inst.o_credits[2] ));
 NAND2x1_ASAP7_75t_R _1461_ (.A(net76),
    .B(_0327_),
    .Y(_0344_));
 AND5x2_ASAP7_75t_R _1462_ (.A(_0054_),
    .B(_0055_),
    .C(_0056_),
    .D(_0701_),
    .E(_0052_),
    .Y(_0345_));
 OR3x2_ASAP7_75t_R _1463_ (.A(net147),
    .B(net146),
    .C(net148),
    .Y(_0346_));
 OR3x2_ASAP7_75t_R _1464_ (.A(net106),
    .B(net105),
    .C(net107),
    .Y(_0347_));
 AND2x2_ASAP7_75t_R _1465_ (.A(_0021_),
    .B(net153),
    .Y(_0348_));
 AO32x2_ASAP7_75t_R _1466_ (.A1(_0021_),
    .A2(net154),
    .A3(_0346_),
    .B1(_0347_),
    .B2(_0348_),
    .Y(_0349_));
 OR3x2_ASAP7_75t_R _1467_ (.A(_0344_),
    .B(_0345_),
    .C(_0349_),
    .Y(_0350_));
 INVx1_ASAP7_75t_R _1468_ (.A(net28),
    .Y(_0351_));
 NOR2x1_ASAP7_75t_R _1469_ (.A(net27),
    .B(net29),
    .Y(_0352_));
 AND5x2_ASAP7_75t_R _1470_ (.A(_0057_),
    .B(_0058_),
    .C(_0059_),
    .D(_0707_),
    .E(_0050_),
    .Y(_0353_));
 INVx1_ASAP7_75t_R _1471_ (.A(net75),
    .Y(_0354_));
 AOI211x1_ASAP7_75t_R _1472_ (.A1(_0351_),
    .A2(_0352_),
    .B(_0353_),
    .C(_0354_),
    .Y(_0355_));
 INVx1_ASAP7_75t_R _1473_ (.A(net154),
    .Y(_0356_));
 NOR3x1_ASAP7_75t_R _1474_ (.A(net147),
    .B(net146),
    .C(net148),
    .Y(_0357_));
 OA31x2_ASAP7_75t_R _1475_ (.A1(net69),
    .A2(net68),
    .A3(net70),
    .B1(net76),
    .Y(_0358_));
 OA31x2_ASAP7_75t_R _1476_ (.A1(net28),
    .A2(net27),
    .A3(net29),
    .B1(net75),
    .Y(_0359_));
 BUFx6f_ASAP7_75t_R _1477_ (.A(_0023_),
    .Y(_0360_));
 FAx1_ASAP7_75t_R _1478_ (.SN(_0045_),
    .A(_0044_),
    .B(_0697_),
    .CI(_0698_),
    .CON(_0027_));
 FAx1_ASAP7_75t_R _1479_ (.SN(_0043_),
    .A(_0042_),
    .B(_0699_),
    .CI(_0700_),
    .CON(_0033_));
 FAx1_ASAP7_75t_R _1480_ (.SN(_0053_),
    .A(_0052_),
    .B(_0701_),
    .CI(_0702_),
    .CON(_0039_));
 FAx1_ASAP7_75t_R _1481_ (.SN(_0049_),
    .A(_0048_),
    .B(_0703_),
    .CI(_0704_),
    .CON(_0006_));
 FAx1_ASAP7_75t_R _1482_ (.SN(_0047_),
    .A(_0046_),
    .B(_0705_),
    .CI(_0706_),
    .CON(_0012_));
 FAx1_ASAP7_75t_R _1483_ (.SN(_0051_),
    .A(_0050_),
    .B(_0707_),
    .CI(_0708_),
    .CON(_0018_));
 HAxp5_ASAP7_75t_R _1484_ (.A(\credit_t_route_inst.l_counters_inst.o_credits[6] ),
    .B(net276),
    .CON(_0026_),
    .SN(_0024_));
 HAxp5_ASAP7_75t_R _1485_ (.A(\credit_t_route_inst.l_counters_inst.o_credits[7] ),
    .B(net276),
    .CON(_0029_),
    .SN(_0025_));
 HAxp5_ASAP7_75t_R _1486_ (.A(\credit_t_route_inst.l_counters_inst.o_credits[8] ),
    .B(net276),
    .CON(_0072_),
    .SN(_0028_));
 HAxp5_ASAP7_75t_R _1487_ (.A(\credit_t_route_inst.l_counters_inst.o_credits[1] ),
    .B(net275),
    .CON(_0032_),
    .SN(_0030_));
 HAxp5_ASAP7_75t_R _1488_ (.A(\credit_t_route_inst.l_counters_inst.o_credits[2] ),
    .B(net275),
    .CON(_0035_),
    .SN(_0031_));
 HAxp5_ASAP7_75t_R _1489_ (.A(\credit_t_route_inst.l_counters_inst.o_credits[3] ),
    .B(net275),
    .CON(_0073_),
    .SN(_0034_));
 HAxp5_ASAP7_75t_R _1490_ (.A(\credit_t_route_inst.u0_counters_inst.o_credits[6] ),
    .B(net358),
    .CON(_0038_),
    .SN(_0036_));
 HAxp5_ASAP7_75t_R _1491_ (.A(\credit_t_route_inst.u0_counters_inst.o_credits[7] ),
    .B(net358),
    .CON(_0041_),
    .SN(_0037_));
 HAxp5_ASAP7_75t_R _1492_ (.A(\credit_t_route_inst.u0_counters_inst.o_credits[8] ),
    .B(net358),
    .CON(_0074_),
    .SN(_0040_));
 HAxp5_ASAP7_75t_R _1493_ (.A(\credit_t_route_inst.r_counters_inst.o_credits[6] ),
    .B(net317),
    .CON(_0005_),
    .SN(_0003_));
 HAxp5_ASAP7_75t_R _1494_ (.A(\credit_t_route_inst.r_counters_inst.o_credits[7] ),
    .B(net317),
    .CON(_0008_),
    .SN(_0004_));
 HAxp5_ASAP7_75t_R _1495_ (.A(\credit_t_route_inst.r_counters_inst.o_credits[8] ),
    .B(net317),
    .CON(_0075_),
    .SN(_0007_));
 HAxp5_ASAP7_75t_R _1496_ (.A(\credit_t_route_inst.r_counters_inst.o_credits[1] ),
    .B(net316),
    .CON(_0011_),
    .SN(_0009_));
 HAxp5_ASAP7_75t_R _1497_ (.A(\credit_t_route_inst.r_counters_inst.o_credits[2] ),
    .B(net316),
    .CON(_0014_),
    .SN(_0010_));
 HAxp5_ASAP7_75t_R _1498_ (.A(\credit_t_route_inst.r_counters_inst.o_credits[3] ),
    .B(net316),
    .CON(_0076_),
    .SN(_0013_));
 HAxp5_ASAP7_75t_R _1499_ (.A(\credit_t_route_inst.u0_counters_inst.o_credits[1] ),
    .B(net357),
    .CON(_0017_),
    .SN(_0015_));
 HAxp5_ASAP7_75t_R _1500_ (.A(\credit_t_route_inst.u0_counters_inst.o_credits[2] ),
    .B(net357),
    .CON(_0020_),
    .SN(_0016_));
 HAxp5_ASAP7_75t_R _1501_ (.A(\credit_t_route_inst.u0_counters_inst.o_credits[3] ),
    .B(net357),
    .CON(_0077_),
    .SN(_0019_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.l_counters_inst.o_credits[0]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0078_),
    .QN(_0042_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.l_counters_inst.o_credits[1]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0079_),
    .QN(_0699_));
 DFFHQNx1_ASAP7_75t_R \credit_t_route_inst.l_counters_inst.o_credits[2]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0080_),
    .QN(_0070_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.l_counters_inst.o_credits[3]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0081_),
    .QN(_0069_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.l_counters_inst.o_credits[4]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0082_),
    .QN(_0068_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.l_counters_inst.o_credits[5]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0083_),
    .QN(_0044_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.l_counters_inst.o_credits[6]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0084_),
    .QN(_0697_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.l_counters_inst.o_credits[7]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0085_),
    .QN(_0067_));
 DFFHQNx1_ASAP7_75t_R \credit_t_route_inst.l_counters_inst.o_credits[8]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0086_),
    .QN(_0066_));
 DFFHQNx1_ASAP7_75t_R \credit_t_route_inst.l_counters_inst.o_credits[9]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0087_),
    .QN(_0065_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.r_counters_inst.o_credits[0]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0088_),
    .QN(_0046_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.r_counters_inst.o_credits[1]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0089_),
    .QN(_0705_));
 DFFHQNx1_ASAP7_75t_R \credit_t_route_inst.r_counters_inst.o_credits[2]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0090_),
    .QN(_0064_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.r_counters_inst.o_credits[3]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0091_),
    .QN(_0063_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.r_counters_inst.o_credits[4]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0092_),
    .QN(_0062_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.r_counters_inst.o_credits[5]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0093_),
    .QN(_0048_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.r_counters_inst.o_credits[6]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0094_),
    .QN(_0703_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.r_counters_inst.o_credits[7]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0095_),
    .QN(_0061_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.r_counters_inst.o_credits[8]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0096_),
    .QN(_0060_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.r_counters_inst.o_credits[9]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0097_),
    .QN(_0071_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.state[0]$_DFF_P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0000_),
    .QN(_0021_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.state[1]$_DFF_P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0001_),
    .QN(_0022_));
 DFFHQNx1_ASAP7_75t_R \credit_t_route_inst.state[2]$_DFF_P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0002_),
    .QN(_0023_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.u0_counters_inst.o_credits[0]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0098_),
    .QN(_0050_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.u0_counters_inst.o_credits[1]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0099_),
    .QN(_0707_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.u0_counters_inst.o_credits[2]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0100_),
    .QN(_0059_));
 DFFHQNx1_ASAP7_75t_R \credit_t_route_inst.u0_counters_inst.o_credits[3]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0101_),
    .QN(_0058_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.u0_counters_inst.o_credits[4]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0102_),
    .QN(_0057_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.u0_counters_inst.o_credits[5]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0103_),
    .QN(_0052_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.u0_counters_inst.o_credits[6]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0104_),
    .QN(_0701_));
 DFFHQNx3_ASAP7_75t_R \credit_t_route_inst.u0_counters_inst.o_credits[7]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0105_),
    .QN(_0056_));
 DFFHQNx1_ASAP7_75t_R \credit_t_route_inst.u0_counters_inst.o_credits[8]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0106_),
    .QN(_0055_));
 DFFHQNx1_ASAP7_75t_R \credit_t_route_inst.u0_counters_inst.o_credits[9]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0107_),
    .QN(_0054_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_109 ();
 BUFx3_ASAP7_75t_R input1 (.A(l_i[0]),
    .Y(net1));
 BUFx3_ASAP7_75t_R input2 (.A(l_i[10]),
    .Y(net2));
 BUFx3_ASAP7_75t_R input3 (.A(l_i[11]),
    .Y(net3));
 BUFx3_ASAP7_75t_R input4 (.A(l_i[12]),
    .Y(net4));
 BUFx3_ASAP7_75t_R input5 (.A(l_i[13]),
    .Y(net5));
 BUFx3_ASAP7_75t_R input6 (.A(l_i[14]),
    .Y(net6));
 BUFx3_ASAP7_75t_R input7 (.A(l_i[15]),
    .Y(net7));
 BUFx3_ASAP7_75t_R input8 (.A(l_i[16]),
    .Y(net8));
 BUFx3_ASAP7_75t_R input9 (.A(l_i[17]),
    .Y(net9));
 BUFx3_ASAP7_75t_R input10 (.A(l_i[18]),
    .Y(net10));
 BUFx3_ASAP7_75t_R input11 (.A(l_i[19]),
    .Y(net11));
 BUFx3_ASAP7_75t_R input12 (.A(l_i[1]),
    .Y(net12));
 BUFx3_ASAP7_75t_R input13 (.A(l_i[20]),
    .Y(net13));
 BUFx3_ASAP7_75t_R input14 (.A(l_i[21]),
    .Y(net14));
 BUFx3_ASAP7_75t_R input15 (.A(l_i[22]),
    .Y(net15));
 BUFx3_ASAP7_75t_R input16 (.A(l_i[23]),
    .Y(net16));
 BUFx3_ASAP7_75t_R input17 (.A(l_i[24]),
    .Y(net17));
 BUFx3_ASAP7_75t_R input18 (.A(l_i[25]),
    .Y(net18));
 BUFx3_ASAP7_75t_R input19 (.A(l_i[26]),
    .Y(net19));
 BUFx3_ASAP7_75t_R input20 (.A(l_i[27]),
    .Y(net20));
 BUFx3_ASAP7_75t_R input21 (.A(l_i[28]),
    .Y(net21));
 BUFx3_ASAP7_75t_R input22 (.A(l_i[29]),
    .Y(net22));
 BUFx3_ASAP7_75t_R input23 (.A(l_i[2]),
    .Y(net23));
 BUFx3_ASAP7_75t_R input24 (.A(l_i[30]),
    .Y(net24));
 BUFx3_ASAP7_75t_R input25 (.A(l_i[31]),
    .Y(net25));
 BUFx3_ASAP7_75t_R input26 (.A(l_i[32]),
    .Y(net26));
 BUFx3_ASAP7_75t_R input27 (.A(l_i[33]),
    .Y(net27));
 BUFx3_ASAP7_75t_R input28 (.A(l_i[34]),
    .Y(net28));
 BUFx3_ASAP7_75t_R input29 (.A(l_i[35]),
    .Y(net29));
 BUFx3_ASAP7_75t_R input30 (.A(l_i[36]),
    .Y(net30));
 BUFx3_ASAP7_75t_R input31 (.A(l_i[37]),
    .Y(net31));
 BUFx3_ASAP7_75t_R input32 (.A(l_i[38]),
    .Y(net32));
 BUFx3_ASAP7_75t_R input33 (.A(l_i[39]),
    .Y(net33));
 BUFx3_ASAP7_75t_R input34 (.A(l_i[3]),
    .Y(net34));
 BUFx3_ASAP7_75t_R input35 (.A(l_i[40]),
    .Y(net35));
 BUFx3_ASAP7_75t_R input36 (.A(l_i[41]),
    .Y(net36));
 BUFx3_ASAP7_75t_R input37 (.A(l_i[42]),
    .Y(net37));
 BUFx3_ASAP7_75t_R input38 (.A(l_i[43]),
    .Y(net38));
 BUFx3_ASAP7_75t_R input39 (.A(l_i[44]),
    .Y(net39));
 BUFx3_ASAP7_75t_R input40 (.A(l_i[45]),
    .Y(net40));
 BUFx3_ASAP7_75t_R input41 (.A(l_i[46]),
    .Y(net41));
 BUFx3_ASAP7_75t_R input42 (.A(l_i[47]),
    .Y(net42));
 BUFx3_ASAP7_75t_R input43 (.A(l_i[48]),
    .Y(net43));
 BUFx3_ASAP7_75t_R input44 (.A(l_i[49]),
    .Y(net44));
 BUFx3_ASAP7_75t_R input45 (.A(l_i[4]),
    .Y(net45));
 BUFx3_ASAP7_75t_R input46 (.A(l_i[50]),
    .Y(net46));
 BUFx3_ASAP7_75t_R input47 (.A(l_i[51]),
    .Y(net47));
 BUFx3_ASAP7_75t_R input48 (.A(l_i[52]),
    .Y(net48));
 BUFx3_ASAP7_75t_R input49 (.A(l_i[53]),
    .Y(net49));
 BUFx3_ASAP7_75t_R input50 (.A(l_i[54]),
    .Y(net50));
 BUFx3_ASAP7_75t_R input51 (.A(l_i[55]),
    .Y(net51));
 BUFx3_ASAP7_75t_R input52 (.A(l_i[56]),
    .Y(net52));
 BUFx3_ASAP7_75t_R input53 (.A(l_i[57]),
    .Y(net53));
 BUFx3_ASAP7_75t_R input54 (.A(l_i[58]),
    .Y(net54));
 BUFx3_ASAP7_75t_R input55 (.A(l_i[59]),
    .Y(net55));
 BUFx3_ASAP7_75t_R input56 (.A(l_i[5]),
    .Y(net56));
 BUFx3_ASAP7_75t_R input57 (.A(l_i[60]),
    .Y(net57));
 BUFx3_ASAP7_75t_R input58 (.A(l_i[61]),
    .Y(net58));
 BUFx3_ASAP7_75t_R input59 (.A(l_i[62]),
    .Y(net59));
 BUFx3_ASAP7_75t_R input60 (.A(l_i[63]),
    .Y(net60));
 BUFx3_ASAP7_75t_R input61 (.A(l_i[64]),
    .Y(net61));
 BUFx3_ASAP7_75t_R input62 (.A(l_i[65]),
    .Y(net62));
 BUFx3_ASAP7_75t_R input63 (.A(l_i[66]),
    .Y(net63));
 BUFx3_ASAP7_75t_R input64 (.A(l_i[67]),
    .Y(net64));
 BUFx3_ASAP7_75t_R input65 (.A(l_i[68]),
    .Y(net65));
 BUFx3_ASAP7_75t_R input66 (.A(l_i[69]),
    .Y(net66));
 BUFx3_ASAP7_75t_R input67 (.A(l_i[6]),
    .Y(net67));
 BUFx3_ASAP7_75t_R input68 (.A(l_i[70]),
    .Y(net68));
 BUFx3_ASAP7_75t_R input69 (.A(l_i[71]),
    .Y(net69));
 BUFx3_ASAP7_75t_R input70 (.A(l_i[72]),
    .Y(net70));
 BUFx3_ASAP7_75t_R input71 (.A(l_i[73]),
    .Y(net71));
 BUFx3_ASAP7_75t_R input72 (.A(l_i[7]),
    .Y(net72));
 BUFx3_ASAP7_75t_R input73 (.A(l_i[8]),
    .Y(net73));
 BUFx3_ASAP7_75t_R input74 (.A(l_i[9]),
    .Y(net74));
 BUFx3_ASAP7_75t_R input75 (.A(l_i_v[0]),
    .Y(net75));
 BUFx3_ASAP7_75t_R input76 (.A(l_i_v[1]),
    .Y(net76));
 BUFx3_ASAP7_75t_R input77 (.A(l_o_credit_gnt[0]),
    .Y(net77));
 BUFx3_ASAP7_75t_R input78 (.A(l_o_credit_gnt[1]),
    .Y(net78));
 BUFx3_ASAP7_75t_R input79 (.A(r_i[0]),
    .Y(net79));
 BUFx3_ASAP7_75t_R input80 (.A(r_i[10]),
    .Y(net80));
 BUFx3_ASAP7_75t_R input81 (.A(r_i[11]),
    .Y(net81));
 BUFx3_ASAP7_75t_R input82 (.A(r_i[12]),
    .Y(net82));
 BUFx3_ASAP7_75t_R input83 (.A(r_i[13]),
    .Y(net83));
 BUFx3_ASAP7_75t_R input84 (.A(r_i[14]),
    .Y(net84));
 BUFx3_ASAP7_75t_R input85 (.A(r_i[15]),
    .Y(net85));
 BUFx3_ASAP7_75t_R input86 (.A(r_i[16]),
    .Y(net86));
 BUFx3_ASAP7_75t_R input87 (.A(r_i[17]),
    .Y(net87));
 BUFx3_ASAP7_75t_R input88 (.A(r_i[18]),
    .Y(net88));
 BUFx3_ASAP7_75t_R input89 (.A(r_i[19]),
    .Y(net89));
 BUFx3_ASAP7_75t_R input90 (.A(r_i[1]),
    .Y(net90));
 BUFx3_ASAP7_75t_R input91 (.A(r_i[20]),
    .Y(net91));
 BUFx3_ASAP7_75t_R input92 (.A(r_i[21]),
    .Y(net92));
 BUFx3_ASAP7_75t_R input93 (.A(r_i[22]),
    .Y(net93));
 BUFx3_ASAP7_75t_R input94 (.A(r_i[23]),
    .Y(net94));
 BUFx3_ASAP7_75t_R input95 (.A(r_i[24]),
    .Y(net95));
 BUFx3_ASAP7_75t_R input96 (.A(r_i[25]),
    .Y(net96));
 BUFx3_ASAP7_75t_R input97 (.A(r_i[26]),
    .Y(net97));
 BUFx3_ASAP7_75t_R input98 (.A(r_i[27]),
    .Y(net98));
 BUFx3_ASAP7_75t_R input99 (.A(r_i[28]),
    .Y(net99));
 BUFx3_ASAP7_75t_R input100 (.A(r_i[29]),
    .Y(net100));
 BUFx3_ASAP7_75t_R input101 (.A(r_i[2]),
    .Y(net101));
 BUFx3_ASAP7_75t_R input102 (.A(r_i[30]),
    .Y(net102));
 BUFx3_ASAP7_75t_R input103 (.A(r_i[31]),
    .Y(net103));
 BUFx3_ASAP7_75t_R input104 (.A(r_i[32]),
    .Y(net104));
 BUFx3_ASAP7_75t_R input105 (.A(r_i[33]),
    .Y(net105));
 BUFx3_ASAP7_75t_R input106 (.A(r_i[34]),
    .Y(net106));
 BUFx3_ASAP7_75t_R input107 (.A(r_i[35]),
    .Y(net107));
 BUFx3_ASAP7_75t_R input108 (.A(r_i[36]),
    .Y(net108));
 BUFx3_ASAP7_75t_R input109 (.A(r_i[37]),
    .Y(net109));
 BUFx3_ASAP7_75t_R input110 (.A(r_i[38]),
    .Y(net110));
 BUFx3_ASAP7_75t_R input111 (.A(r_i[39]),
    .Y(net111));
 BUFx3_ASAP7_75t_R input112 (.A(r_i[3]),
    .Y(net112));
 BUFx3_ASAP7_75t_R input113 (.A(r_i[40]),
    .Y(net113));
 BUFx3_ASAP7_75t_R input114 (.A(r_i[41]),
    .Y(net114));
 BUFx3_ASAP7_75t_R input115 (.A(r_i[42]),
    .Y(net115));
 BUFx3_ASAP7_75t_R input116 (.A(r_i[43]),
    .Y(net116));
 BUFx3_ASAP7_75t_R input117 (.A(r_i[44]),
    .Y(net117));
 BUFx3_ASAP7_75t_R input118 (.A(r_i[45]),
    .Y(net118));
 BUFx3_ASAP7_75t_R input119 (.A(r_i[46]),
    .Y(net119));
 BUFx3_ASAP7_75t_R input120 (.A(r_i[47]),
    .Y(net120));
 BUFx3_ASAP7_75t_R input121 (.A(r_i[48]),
    .Y(net121));
 BUFx3_ASAP7_75t_R input122 (.A(r_i[49]),
    .Y(net122));
 BUFx3_ASAP7_75t_R input123 (.A(r_i[4]),
    .Y(net123));
 BUFx3_ASAP7_75t_R input124 (.A(r_i[50]),
    .Y(net124));
 BUFx3_ASAP7_75t_R input125 (.A(r_i[51]),
    .Y(net125));
 BUFx3_ASAP7_75t_R input126 (.A(r_i[52]),
    .Y(net126));
 BUFx3_ASAP7_75t_R input127 (.A(r_i[53]),
    .Y(net127));
 BUFx3_ASAP7_75t_R input128 (.A(r_i[54]),
    .Y(net128));
 BUFx3_ASAP7_75t_R input129 (.A(r_i[55]),
    .Y(net129));
 BUFx3_ASAP7_75t_R input130 (.A(r_i[56]),
    .Y(net130));
 BUFx3_ASAP7_75t_R input131 (.A(r_i[57]),
    .Y(net131));
 BUFx3_ASAP7_75t_R input132 (.A(r_i[58]),
    .Y(net132));
 BUFx3_ASAP7_75t_R input133 (.A(r_i[59]),
    .Y(net133));
 BUFx3_ASAP7_75t_R input134 (.A(r_i[5]),
    .Y(net134));
 BUFx3_ASAP7_75t_R input135 (.A(r_i[60]),
    .Y(net135));
 BUFx3_ASAP7_75t_R input136 (.A(r_i[61]),
    .Y(net136));
 BUFx3_ASAP7_75t_R input137 (.A(r_i[62]),
    .Y(net137));
 BUFx3_ASAP7_75t_R input138 (.A(r_i[63]),
    .Y(net138));
 BUFx3_ASAP7_75t_R input139 (.A(r_i[64]),
    .Y(net139));
 BUFx3_ASAP7_75t_R input140 (.A(r_i[65]),
    .Y(net140));
 BUFx3_ASAP7_75t_R input141 (.A(r_i[66]),
    .Y(net141));
 BUFx3_ASAP7_75t_R input142 (.A(r_i[67]),
    .Y(net142));
 BUFx3_ASAP7_75t_R input143 (.A(r_i[68]),
    .Y(net143));
 BUFx3_ASAP7_75t_R input144 (.A(r_i[69]),
    .Y(net144));
 BUFx3_ASAP7_75t_R input145 (.A(r_i[6]),
    .Y(net145));
 BUFx3_ASAP7_75t_R input146 (.A(r_i[70]),
    .Y(net146));
 BUFx3_ASAP7_75t_R input147 (.A(r_i[71]),
    .Y(net147));
 BUFx3_ASAP7_75t_R input148 (.A(r_i[72]),
    .Y(net148));
 BUFx3_ASAP7_75t_R input149 (.A(r_i[73]),
    .Y(net149));
 BUFx3_ASAP7_75t_R input150 (.A(r_i[7]),
    .Y(net150));
 BUFx3_ASAP7_75t_R input151 (.A(r_i[8]),
    .Y(net151));
 BUFx3_ASAP7_75t_R input152 (.A(r_i[9]),
    .Y(net152));
 BUFx3_ASAP7_75t_R input153 (.A(r_i_v[0]),
    .Y(net153));
 BUFx3_ASAP7_75t_R input154 (.A(r_i_v[1]),
    .Y(net154));
 BUFx3_ASAP7_75t_R input155 (.A(r_o_credit_gnt[0]),
    .Y(net155));
 BUFx3_ASAP7_75t_R input156 (.A(r_o_credit_gnt[1]),
    .Y(net156));
 BUFx6f_ASAP7_75t_R input157 (.A(rst),
    .Y(net157));
 BUFx3_ASAP7_75t_R input158 (.A(u0_i[0]),
    .Y(net158));
 BUFx3_ASAP7_75t_R input159 (.A(u0_i[10]),
    .Y(net159));
 BUFx3_ASAP7_75t_R input160 (.A(u0_i[11]),
    .Y(net160));
 BUFx3_ASAP7_75t_R input161 (.A(u0_i[12]),
    .Y(net161));
 BUFx3_ASAP7_75t_R input162 (.A(u0_i[13]),
    .Y(net162));
 BUFx3_ASAP7_75t_R input163 (.A(u0_i[14]),
    .Y(net163));
 BUFx3_ASAP7_75t_R input164 (.A(u0_i[15]),
    .Y(net164));
 BUFx3_ASAP7_75t_R input165 (.A(u0_i[16]),
    .Y(net165));
 BUFx3_ASAP7_75t_R input166 (.A(u0_i[17]),
    .Y(net166));
 BUFx3_ASAP7_75t_R input167 (.A(u0_i[18]),
    .Y(net167));
 BUFx3_ASAP7_75t_R input168 (.A(u0_i[19]),
    .Y(net168));
 BUFx3_ASAP7_75t_R input169 (.A(u0_i[1]),
    .Y(net169));
 BUFx3_ASAP7_75t_R input170 (.A(u0_i[20]),
    .Y(net170));
 BUFx3_ASAP7_75t_R input171 (.A(u0_i[21]),
    .Y(net171));
 BUFx3_ASAP7_75t_R input172 (.A(u0_i[22]),
    .Y(net172));
 BUFx3_ASAP7_75t_R input173 (.A(u0_i[23]),
    .Y(net173));
 BUFx3_ASAP7_75t_R input174 (.A(u0_i[24]),
    .Y(net174));
 BUFx3_ASAP7_75t_R input175 (.A(u0_i[25]),
    .Y(net175));
 BUFx3_ASAP7_75t_R input176 (.A(u0_i[26]),
    .Y(net176));
 BUFx3_ASAP7_75t_R input177 (.A(u0_i[27]),
    .Y(net177));
 BUFx3_ASAP7_75t_R input178 (.A(u0_i[28]),
    .Y(net178));
 BUFx3_ASAP7_75t_R input179 (.A(u0_i[29]),
    .Y(net179));
 BUFx3_ASAP7_75t_R input180 (.A(u0_i[2]),
    .Y(net180));
 BUFx3_ASAP7_75t_R input181 (.A(u0_i[30]),
    .Y(net181));
 BUFx3_ASAP7_75t_R input182 (.A(u0_i[31]),
    .Y(net182));
 BUFx6f_ASAP7_75t_R input183 (.A(u0_i[32]),
    .Y(net183));
 BUFx3_ASAP7_75t_R input184 (.A(u0_i[33]),
    .Y(net184));
 BUFx3_ASAP7_75t_R input185 (.A(u0_i[34]),
    .Y(net185));
 BUFx3_ASAP7_75t_R input186 (.A(u0_i[35]),
    .Y(net186));
 BUFx3_ASAP7_75t_R input187 (.A(u0_i[36]),
    .Y(net187));
 BUFx3_ASAP7_75t_R input188 (.A(u0_i[37]),
    .Y(net188));
 BUFx3_ASAP7_75t_R input189 (.A(u0_i[38]),
    .Y(net189));
 BUFx3_ASAP7_75t_R input190 (.A(u0_i[39]),
    .Y(net190));
 BUFx3_ASAP7_75t_R input191 (.A(u0_i[3]),
    .Y(net191));
 BUFx3_ASAP7_75t_R input192 (.A(u0_i[40]),
    .Y(net192));
 BUFx3_ASAP7_75t_R input193 (.A(u0_i[41]),
    .Y(net193));
 BUFx3_ASAP7_75t_R input194 (.A(u0_i[42]),
    .Y(net194));
 BUFx3_ASAP7_75t_R input195 (.A(u0_i[43]),
    .Y(net195));
 BUFx3_ASAP7_75t_R input196 (.A(u0_i[44]),
    .Y(net196));
 BUFx3_ASAP7_75t_R input197 (.A(u0_i[45]),
    .Y(net197));
 BUFx3_ASAP7_75t_R input198 (.A(u0_i[46]),
    .Y(net198));
 BUFx3_ASAP7_75t_R input199 (.A(u0_i[47]),
    .Y(net199));
 BUFx3_ASAP7_75t_R input200 (.A(u0_i[48]),
    .Y(net200));
 BUFx3_ASAP7_75t_R input201 (.A(u0_i[49]),
    .Y(net201));
 BUFx3_ASAP7_75t_R input202 (.A(u0_i[4]),
    .Y(net202));
 BUFx3_ASAP7_75t_R input203 (.A(u0_i[50]),
    .Y(net203));
 BUFx3_ASAP7_75t_R input204 (.A(u0_i[51]),
    .Y(net204));
 BUFx3_ASAP7_75t_R input205 (.A(u0_i[52]),
    .Y(net205));
 BUFx3_ASAP7_75t_R input206 (.A(u0_i[53]),
    .Y(net206));
 BUFx3_ASAP7_75t_R input207 (.A(u0_i[54]),
    .Y(net207));
 BUFx3_ASAP7_75t_R input208 (.A(u0_i[55]),
    .Y(net208));
 BUFx3_ASAP7_75t_R input209 (.A(u0_i[56]),
    .Y(net209));
 BUFx3_ASAP7_75t_R input210 (.A(u0_i[57]),
    .Y(net210));
 BUFx3_ASAP7_75t_R input211 (.A(u0_i[58]),
    .Y(net211));
 BUFx3_ASAP7_75t_R input212 (.A(u0_i[59]),
    .Y(net212));
 BUFx3_ASAP7_75t_R input213 (.A(u0_i[5]),
    .Y(net213));
 BUFx3_ASAP7_75t_R input214 (.A(u0_i[60]),
    .Y(net214));
 BUFx3_ASAP7_75t_R input215 (.A(u0_i[61]),
    .Y(net215));
 BUFx3_ASAP7_75t_R input216 (.A(u0_i[62]),
    .Y(net216));
 BUFx3_ASAP7_75t_R input217 (.A(u0_i[63]),
    .Y(net217));
 BUFx3_ASAP7_75t_R input218 (.A(u0_i[64]),
    .Y(net218));
 BUFx3_ASAP7_75t_R input219 (.A(u0_i[65]),
    .Y(net219));
 BUFx3_ASAP7_75t_R input220 (.A(u0_i[66]),
    .Y(net220));
 BUFx3_ASAP7_75t_R input221 (.A(u0_i[67]),
    .Y(net221));
 BUFx3_ASAP7_75t_R input222 (.A(u0_i[68]),
    .Y(net222));
 BUFx6f_ASAP7_75t_R input223 (.A(u0_i[69]),
    .Y(net223));
 BUFx3_ASAP7_75t_R input224 (.A(u0_i[6]),
    .Y(net224));
 BUFx3_ASAP7_75t_R input225 (.A(u0_i[70]),
    .Y(net225));
 BUFx3_ASAP7_75t_R input226 (.A(u0_i[71]),
    .Y(net226));
 BUFx3_ASAP7_75t_R input227 (.A(u0_i[72]),
    .Y(net227));
 BUFx3_ASAP7_75t_R input228 (.A(u0_i[73]),
    .Y(net228));
 BUFx3_ASAP7_75t_R input229 (.A(u0_i[7]),
    .Y(net229));
 BUFx3_ASAP7_75t_R input230 (.A(u0_i[8]),
    .Y(net230));
 BUFx3_ASAP7_75t_R input231 (.A(u0_i[9]),
    .Y(net231));
 BUFx6f_ASAP7_75t_R input232 (.A(u0_i_v[0]),
    .Y(net232));
 BUFx3_ASAP7_75t_R input233 (.A(u0_i_v[1]),
    .Y(net233));
 BUFx3_ASAP7_75t_R input234 (.A(u0_o_credit_gnt[0]),
    .Y(net234));
 BUFx3_ASAP7_75t_R input235 (.A(u0_o_credit_gnt[1]),
    .Y(net235));
 BUFx3_ASAP7_75t_R output236 (.A(net236),
    .Y(l_i_bp[0]));
 BUFx3_ASAP7_75t_R output237 (.A(net237),
    .Y(l_i_bp[1]));
 BUFx3_ASAP7_75t_R output238 (.A(net238),
    .Y(l_o[0]));
 BUFx3_ASAP7_75t_R output239 (.A(net239),
    .Y(l_o[10]));
 BUFx3_ASAP7_75t_R output240 (.A(net240),
    .Y(l_o[11]));
 BUFx3_ASAP7_75t_R output241 (.A(net241),
    .Y(l_o[12]));
 BUFx3_ASAP7_75t_R output242 (.A(net242),
    .Y(l_o[13]));
 BUFx3_ASAP7_75t_R output243 (.A(net243),
    .Y(l_o[14]));
 BUFx3_ASAP7_75t_R output244 (.A(net244),
    .Y(l_o[15]));
 BUFx3_ASAP7_75t_R output245 (.A(net245),
    .Y(l_o[16]));
 BUFx3_ASAP7_75t_R output246 (.A(net246),
    .Y(l_o[17]));
 BUFx3_ASAP7_75t_R output247 (.A(net247),
    .Y(l_o[18]));
 BUFx3_ASAP7_75t_R output248 (.A(net248),
    .Y(l_o[19]));
 BUFx3_ASAP7_75t_R output249 (.A(net249),
    .Y(l_o[1]));
 BUFx3_ASAP7_75t_R output250 (.A(net250),
    .Y(l_o[20]));
 BUFx3_ASAP7_75t_R output251 (.A(net251),
    .Y(l_o[21]));
 BUFx3_ASAP7_75t_R output252 (.A(net252),
    .Y(l_o[22]));
 BUFx3_ASAP7_75t_R output253 (.A(net253),
    .Y(l_o[23]));
 BUFx3_ASAP7_75t_R output254 (.A(net254),
    .Y(l_o[24]));
 BUFx3_ASAP7_75t_R output255 (.A(net255),
    .Y(l_o[25]));
 BUFx3_ASAP7_75t_R output256 (.A(net256),
    .Y(l_o[26]));
 BUFx3_ASAP7_75t_R output257 (.A(net257),
    .Y(l_o[27]));
 BUFx3_ASAP7_75t_R output258 (.A(net258),
    .Y(l_o[28]));
 BUFx3_ASAP7_75t_R output259 (.A(net259),
    .Y(l_o[29]));
 BUFx3_ASAP7_75t_R output260 (.A(net260),
    .Y(l_o[2]));
 BUFx3_ASAP7_75t_R output261 (.A(net261),
    .Y(l_o[30]));
 BUFx3_ASAP7_75t_R output262 (.A(net262),
    .Y(l_o[31]));
 BUFx3_ASAP7_75t_R output263 (.A(net263),
    .Y(l_o[32]));
 BUFx3_ASAP7_75t_R output264 (.A(net264),
    .Y(l_o[33]));
 BUFx3_ASAP7_75t_R output265 (.A(net265),
    .Y(l_o[34]));
 BUFx3_ASAP7_75t_R output266 (.A(net266),
    .Y(l_o[35]));
 BUFx3_ASAP7_75t_R output267 (.A(net267),
    .Y(l_o[36]));
 BUFx3_ASAP7_75t_R output268 (.A(net268),
    .Y(l_o[3]));
 BUFx3_ASAP7_75t_R output269 (.A(net269),
    .Y(l_o[4]));
 BUFx3_ASAP7_75t_R output270 (.A(net270),
    .Y(l_o[5]));
 BUFx3_ASAP7_75t_R output271 (.A(net271),
    .Y(l_o[6]));
 BUFx3_ASAP7_75t_R output272 (.A(net272),
    .Y(l_o[7]));
 BUFx3_ASAP7_75t_R output273 (.A(net273),
    .Y(l_o[8]));
 BUFx3_ASAP7_75t_R output274 (.A(net274),
    .Y(l_o[9]));
 BUFx3_ASAP7_75t_R output275 (.A(net275),
    .Y(l_o_v[0]));
 BUFx3_ASAP7_75t_R output276 (.A(net276),
    .Y(l_o_v[1]));
 BUFx3_ASAP7_75t_R output277 (.A(net277),
    .Y(r_i_bp[0]));
 BUFx3_ASAP7_75t_R output278 (.A(net278),
    .Y(r_i_bp[1]));
 BUFx3_ASAP7_75t_R output279 (.A(net279),
    .Y(r_o[0]));
 BUFx3_ASAP7_75t_R output280 (.A(net280),
    .Y(r_o[10]));
 BUFx3_ASAP7_75t_R output281 (.A(net281),
    .Y(r_o[11]));
 BUFx3_ASAP7_75t_R output282 (.A(net282),
    .Y(r_o[12]));
 BUFx3_ASAP7_75t_R output283 (.A(net283),
    .Y(r_o[13]));
 BUFx3_ASAP7_75t_R output284 (.A(net284),
    .Y(r_o[14]));
 BUFx3_ASAP7_75t_R output285 (.A(net285),
    .Y(r_o[15]));
 BUFx3_ASAP7_75t_R output286 (.A(net286),
    .Y(r_o[16]));
 BUFx3_ASAP7_75t_R output287 (.A(net287),
    .Y(r_o[17]));
 BUFx3_ASAP7_75t_R output288 (.A(net288),
    .Y(r_o[18]));
 BUFx3_ASAP7_75t_R output289 (.A(net289),
    .Y(r_o[19]));
 BUFx3_ASAP7_75t_R output290 (.A(net290),
    .Y(r_o[1]));
 BUFx3_ASAP7_75t_R output291 (.A(net291),
    .Y(r_o[20]));
 BUFx3_ASAP7_75t_R output292 (.A(net292),
    .Y(r_o[21]));
 BUFx3_ASAP7_75t_R output293 (.A(net293),
    .Y(r_o[22]));
 BUFx3_ASAP7_75t_R output294 (.A(net294),
    .Y(r_o[23]));
 BUFx3_ASAP7_75t_R output295 (.A(net295),
    .Y(r_o[24]));
 BUFx3_ASAP7_75t_R output296 (.A(net296),
    .Y(r_o[25]));
 BUFx3_ASAP7_75t_R output297 (.A(net297),
    .Y(r_o[26]));
 BUFx3_ASAP7_75t_R output298 (.A(net298),
    .Y(r_o[27]));
 BUFx3_ASAP7_75t_R output299 (.A(net299),
    .Y(r_o[28]));
 BUFx3_ASAP7_75t_R output300 (.A(net300),
    .Y(r_o[29]));
 BUFx3_ASAP7_75t_R output301 (.A(net301),
    .Y(r_o[2]));
 BUFx3_ASAP7_75t_R output302 (.A(net302),
    .Y(r_o[30]));
 BUFx3_ASAP7_75t_R output303 (.A(net303),
    .Y(r_o[31]));
 BUFx3_ASAP7_75t_R output304 (.A(net304),
    .Y(r_o[32]));
 BUFx3_ASAP7_75t_R output305 (.A(net305),
    .Y(r_o[33]));
 BUFx3_ASAP7_75t_R output306 (.A(net306),
    .Y(r_o[34]));
 BUFx3_ASAP7_75t_R output307 (.A(net307),
    .Y(r_o[35]));
 BUFx3_ASAP7_75t_R output308 (.A(net308),
    .Y(r_o[36]));
 BUFx3_ASAP7_75t_R output309 (.A(net309),
    .Y(r_o[3]));
 BUFx3_ASAP7_75t_R output310 (.A(net310),
    .Y(r_o[4]));
 BUFx3_ASAP7_75t_R output311 (.A(net311),
    .Y(r_o[5]));
 BUFx3_ASAP7_75t_R output312 (.A(net312),
    .Y(r_o[6]));
 BUFx3_ASAP7_75t_R output313 (.A(net313),
    .Y(r_o[7]));
 BUFx3_ASAP7_75t_R output314 (.A(net314),
    .Y(r_o[8]));
 BUFx3_ASAP7_75t_R output315 (.A(net315),
    .Y(r_o[9]));
 BUFx3_ASAP7_75t_R output316 (.A(net316),
    .Y(r_o_v[0]));
 BUFx3_ASAP7_75t_R output317 (.A(net317),
    .Y(r_o_v[1]));
 BUFx3_ASAP7_75t_R output318 (.A(net318),
    .Y(u0_i_bp[0]));
 BUFx3_ASAP7_75t_R output319 (.A(net319),
    .Y(u0_i_bp[1]));
 BUFx3_ASAP7_75t_R output320 (.A(net320),
    .Y(u0_o[0]));
 BUFx3_ASAP7_75t_R output321 (.A(net321),
    .Y(u0_o[10]));
 BUFx3_ASAP7_75t_R output322 (.A(net322),
    .Y(u0_o[11]));
 BUFx3_ASAP7_75t_R output323 (.A(net323),
    .Y(u0_o[12]));
 BUFx3_ASAP7_75t_R output324 (.A(net324),
    .Y(u0_o[13]));
 BUFx3_ASAP7_75t_R output325 (.A(net325),
    .Y(u0_o[14]));
 BUFx3_ASAP7_75t_R output326 (.A(net326),
    .Y(u0_o[15]));
 BUFx3_ASAP7_75t_R output327 (.A(net327),
    .Y(u0_o[16]));
 BUFx3_ASAP7_75t_R output328 (.A(net328),
    .Y(u0_o[17]));
 BUFx3_ASAP7_75t_R output329 (.A(net329),
    .Y(u0_o[18]));
 BUFx3_ASAP7_75t_R output330 (.A(net330),
    .Y(u0_o[19]));
 BUFx3_ASAP7_75t_R output331 (.A(net331),
    .Y(u0_o[1]));
 BUFx3_ASAP7_75t_R output332 (.A(net332),
    .Y(u0_o[20]));
 BUFx3_ASAP7_75t_R output333 (.A(net333),
    .Y(u0_o[21]));
 BUFx3_ASAP7_75t_R output334 (.A(net334),
    .Y(u0_o[22]));
 BUFx3_ASAP7_75t_R output335 (.A(net335),
    .Y(u0_o[23]));
 BUFx3_ASAP7_75t_R output336 (.A(net336),
    .Y(u0_o[24]));
 BUFx3_ASAP7_75t_R output337 (.A(net337),
    .Y(u0_o[25]));
 BUFx3_ASAP7_75t_R output338 (.A(net338),
    .Y(u0_o[26]));
 BUFx3_ASAP7_75t_R output339 (.A(net339),
    .Y(u0_o[27]));
 BUFx3_ASAP7_75t_R output340 (.A(net340),
    .Y(u0_o[28]));
 BUFx3_ASAP7_75t_R output341 (.A(net341),
    .Y(u0_o[29]));
 BUFx3_ASAP7_75t_R output342 (.A(net342),
    .Y(u0_o[2]));
 BUFx3_ASAP7_75t_R output343 (.A(net343),
    .Y(u0_o[30]));
 BUFx3_ASAP7_75t_R output344 (.A(net344),
    .Y(u0_o[31]));
 BUFx3_ASAP7_75t_R output345 (.A(net345),
    .Y(u0_o[32]));
 BUFx3_ASAP7_75t_R output346 (.A(net346),
    .Y(u0_o[33]));
 BUFx3_ASAP7_75t_R output347 (.A(net347),
    .Y(u0_o[34]));
 BUFx3_ASAP7_75t_R output348 (.A(net348),
    .Y(u0_o[35]));
 BUFx3_ASAP7_75t_R output349 (.A(net349),
    .Y(u0_o[36]));
 BUFx3_ASAP7_75t_R output350 (.A(net350),
    .Y(u0_o[3]));
 BUFx3_ASAP7_75t_R output351 (.A(net351),
    .Y(u0_o[4]));
 BUFx3_ASAP7_75t_R output352 (.A(net352),
    .Y(u0_o[5]));
 BUFx3_ASAP7_75t_R output353 (.A(net353),
    .Y(u0_o[6]));
 BUFx3_ASAP7_75t_R output354 (.A(net354),
    .Y(u0_o[7]));
 BUFx3_ASAP7_75t_R output355 (.A(net355),
    .Y(u0_o[8]));
 BUFx3_ASAP7_75t_R output356 (.A(net356),
    .Y(u0_o[9]));
 BUFx3_ASAP7_75t_R output357 (.A(net357),
    .Y(u0_o_v[0]));
 BUFx3_ASAP7_75t_R output358 (.A(net358),
    .Y(u0_o_v[1]));
 BUFx4_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_0__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_1__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_2__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_3__leaf_clk));
 BUFx12_ASAP7_75t_R clkload0 (.A(clknet_2_1__leaf_clk));
 INVxp67_ASAP7_75t_R clkload1 (.A(clknet_2_2__leaf_clk));
 BUFx12_ASAP7_75t_R clkload2 (.A(clknet_2_3__leaf_clk));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24 ();
 DECAPx4_ASAP7_75t_R FILLER_0_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100 ();
 FILLER_ASAP7_75t_R FILLER_0_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112 ();
 FILLER_ASAP7_75t_R FILLER_0_123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153 ();
 DECAPx1_ASAP7_75t_R FILLER_0_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242 ();
 DECAPx6_ASAP7_75t_R FILLER_0_264 ();
 DECAPx4_ASAP7_75t_R FILLER_1_2 ();
 FILLER_ASAP7_75t_R FILLER_1_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_18 ();
 FILLER_ASAP7_75t_R FILLER_1_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_60 ();
 DECAPx2_ASAP7_75t_R FILLER_1_67 ();
 FILLER_ASAP7_75t_R FILLER_1_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_75 ();
 DECAPx1_ASAP7_75t_R FILLER_1_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_90 ();
 DECAPx6_ASAP7_75t_R FILLER_1_103 ();
 DECAPx10_ASAP7_75t_R FILLER_1_123 ();
 DECAPx10_ASAP7_75t_R FILLER_1_145 ();
 DECAPx4_ASAP7_75t_R FILLER_1_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_177 ();
 DECAPx10_ASAP7_75t_R FILLER_1_184 ();
 DECAPx10_ASAP7_75t_R FILLER_1_206 ();
 DECAPx10_ASAP7_75t_R FILLER_1_228 ();
 DECAPx6_ASAP7_75t_R FILLER_1_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_277 ();
 DECAPx1_ASAP7_75t_R FILLER_2_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_6 ();
 DECAPx1_ASAP7_75t_R FILLER_2_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_35 ();
 FILLER_ASAP7_75t_R FILLER_2_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_49 ();
 FILLER_ASAP7_75t_R FILLER_2_56 ();
 DECAPx2_ASAP7_75t_R FILLER_2_70 ();
 FILLER_ASAP7_75t_R FILLER_2_76 ();
 DECAPx2_ASAP7_75t_R FILLER_2_120 ();
 DECAPx2_ASAP7_75t_R FILLER_2_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_143 ();
 DECAPx4_ASAP7_75t_R FILLER_2_151 ();
 DECAPx10_ASAP7_75t_R FILLER_2_189 ();
 DECAPx10_ASAP7_75t_R FILLER_2_211 ();
 DECAPx6_ASAP7_75t_R FILLER_2_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_247 ();
 DECAPx1_ASAP7_75t_R FILLER_2_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_265 ();
 DECAPx2_ASAP7_75t_R FILLER_2_272 ();
 DECAPx2_ASAP7_75t_R FILLER_3_2 ();
 FILLER_ASAP7_75t_R FILLER_3_8 ();
 DECAPx1_ASAP7_75t_R FILLER_3_14 ();
 DECAPx2_ASAP7_75t_R FILLER_3_24 ();
 FILLER_ASAP7_75t_R FILLER_3_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_32 ();
 DECAPx1_ASAP7_75t_R FILLER_3_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_47 ();
 DECAPx4_ASAP7_75t_R FILLER_3_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_78 ();
 DECAPx2_ASAP7_75t_R FILLER_3_91 ();
 FILLER_ASAP7_75t_R FILLER_3_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_99 ();
 DECAPx6_ASAP7_75t_R FILLER_3_106 ();
 FILLER_ASAP7_75t_R FILLER_3_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_122 ();
 DECAPx2_ASAP7_75t_R FILLER_3_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_138 ();
 DECAPx1_ASAP7_75t_R FILLER_3_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_155 ();
 DECAPx10_ASAP7_75t_R FILLER_3_168 ();
 DECAPx10_ASAP7_75t_R FILLER_3_190 ();
 DECAPx10_ASAP7_75t_R FILLER_3_212 ();
 DECAPx10_ASAP7_75t_R FILLER_3_234 ();
 DECAPx1_ASAP7_75t_R FILLER_3_256 ();
 DECAPx2_ASAP7_75t_R FILLER_3_266 ();
 DECAPx6_ASAP7_75t_R FILLER_4_2 ();
 DECAPx1_ASAP7_75t_R FILLER_4_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_20 ();
 DECAPx2_ASAP7_75t_R FILLER_4_28 ();
 FILLER_ASAP7_75t_R FILLER_4_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_36 ();
 DECAPx4_ASAP7_75t_R FILLER_4_49 ();
 FILLER_ASAP7_75t_R FILLER_4_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_61 ();
 FILLER_ASAP7_75t_R FILLER_4_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_92 ();
 FILLER_ASAP7_75t_R FILLER_4_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_98 ();
 DECAPx2_ASAP7_75t_R FILLER_4_111 ();
 FILLER_ASAP7_75t_R FILLER_4_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_119 ();
 DECAPx1_ASAP7_75t_R FILLER_4_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_149 ();
 DECAPx10_ASAP7_75t_R FILLER_4_167 ();
 DECAPx10_ASAP7_75t_R FILLER_4_189 ();
 DECAPx10_ASAP7_75t_R FILLER_4_211 ();
 DECAPx6_ASAP7_75t_R FILLER_4_233 ();
 DECAPx2_ASAP7_75t_R FILLER_4_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_277 ();
 DECAPx6_ASAP7_75t_R FILLER_5_2 ();
 FILLER_ASAP7_75t_R FILLER_5_16 ();
 DECAPx6_ASAP7_75t_R FILLER_5_65 ();
 DECAPx1_ASAP7_75t_R FILLER_5_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_89 ();
 DECAPx2_ASAP7_75t_R FILLER_5_108 ();
 FILLER_ASAP7_75t_R FILLER_5_114 ();
 DECAPx1_ASAP7_75t_R FILLER_5_128 ();
 DECAPx2_ASAP7_75t_R FILLER_5_151 ();
 FILLER_ASAP7_75t_R FILLER_5_157 ();
 DECAPx10_ASAP7_75t_R FILLER_5_171 ();
 DECAPx10_ASAP7_75t_R FILLER_5_193 ();
 DECAPx10_ASAP7_75t_R FILLER_5_215 ();
 DECAPx6_ASAP7_75t_R FILLER_5_237 ();
 FILLER_ASAP7_75t_R FILLER_5_251 ();
 DECAPx2_ASAP7_75t_R FILLER_5_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_271 ();
 DECAPx2_ASAP7_75t_R FILLER_6_2 ();
 DECAPx2_ASAP7_75t_R FILLER_6_14 ();
 FILLER_ASAP7_75t_R FILLER_6_20 ();
 DECAPx2_ASAP7_75t_R FILLER_6_25 ();
 DECAPx2_ASAP7_75t_R FILLER_6_37 ();
 FILLER_ASAP7_75t_R FILLER_6_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_45 ();
 DECAPx2_ASAP7_75t_R FILLER_6_65 ();
 FILLER_ASAP7_75t_R FILLER_6_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_94 ();
 DECAPx4_ASAP7_75t_R FILLER_6_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_117 ();
 DECAPx4_ASAP7_75t_R FILLER_6_141 ();
 FILLER_ASAP7_75t_R FILLER_6_151 ();
 DECAPx10_ASAP7_75t_R FILLER_6_173 ();
 DECAPx10_ASAP7_75t_R FILLER_6_195 ();
 DECAPx10_ASAP7_75t_R FILLER_6_217 ();
 DECAPx4_ASAP7_75t_R FILLER_6_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_249 ();
 DECAPx2_ASAP7_75t_R FILLER_6_262 ();
 DECAPx1_ASAP7_75t_R FILLER_6_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_22 ();
 DECAPx2_ASAP7_75t_R FILLER_7_35 ();
 DECAPx10_ASAP7_75t_R FILLER_7_52 ();
 DECAPx2_ASAP7_75t_R FILLER_7_74 ();
 FILLER_ASAP7_75t_R FILLER_7_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_92 ();
 DECAPx10_ASAP7_75t_R FILLER_7_100 ();
 FILLER_ASAP7_75t_R FILLER_7_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_124 ();
 DECAPx1_ASAP7_75t_R FILLER_7_137 ();
 FILLER_ASAP7_75t_R FILLER_7_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_163 ();
 DECAPx10_ASAP7_75t_R FILLER_7_186 ();
 DECAPx10_ASAP7_75t_R FILLER_7_208 ();
 DECAPx6_ASAP7_75t_R FILLER_7_230 ();
 DECAPx2_ASAP7_75t_R FILLER_7_244 ();
 DECAPx4_ASAP7_75t_R FILLER_7_256 ();
 DECAPx2_ASAP7_75t_R FILLER_7_272 ();
 FILLER_ASAP7_75t_R FILLER_8_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_4 ();
 DECAPx6_ASAP7_75t_R FILLER_8_27 ();
 DECAPx1_ASAP7_75t_R FILLER_8_41 ();
 DECAPx2_ASAP7_75t_R FILLER_8_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_73 ();
 DECAPx10_ASAP7_75t_R FILLER_8_95 ();
 DECAPx4_ASAP7_75t_R FILLER_8_117 ();
 FILLER_ASAP7_75t_R FILLER_8_127 ();
 DECAPx6_ASAP7_75t_R FILLER_8_134 ();
 DECAPx2_ASAP7_75t_R FILLER_8_148 ();
 DECAPx10_ASAP7_75t_R FILLER_8_165 ();
 DECAPx10_ASAP7_75t_R FILLER_8_187 ();
 DECAPx10_ASAP7_75t_R FILLER_8_209 ();
 DECAPx6_ASAP7_75t_R FILLER_8_231 ();
 FILLER_ASAP7_75t_R FILLER_8_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_247 ();
 DECAPx2_ASAP7_75t_R FILLER_8_260 ();
 DECAPx2_ASAP7_75t_R FILLER_9_2 ();
 FILLER_ASAP7_75t_R FILLER_9_14 ();
 DECAPx4_ASAP7_75t_R FILLER_9_36 ();
 DECAPx10_ASAP7_75t_R FILLER_9_52 ();
 DECAPx6_ASAP7_75t_R FILLER_9_109 ();
 DECAPx2_ASAP7_75t_R FILLER_9_123 ();
 DECAPx10_ASAP7_75t_R FILLER_9_149 ();
 DECAPx10_ASAP7_75t_R FILLER_9_171 ();
 DECAPx10_ASAP7_75t_R FILLER_9_193 ();
 DECAPx10_ASAP7_75t_R FILLER_9_215 ();
 DECAPx2_ASAP7_75t_R FILLER_9_237 ();
 FILLER_ASAP7_75t_R FILLER_9_243 ();
 FILLER_ASAP7_75t_R FILLER_9_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_253 ();
 DECAPx6_ASAP7_75t_R FILLER_9_260 ();
 DECAPx1_ASAP7_75t_R FILLER_9_274 ();
 FILLER_ASAP7_75t_R FILLER_10_2 ();
 FILLER_ASAP7_75t_R FILLER_10_15 ();
 FILLER_ASAP7_75t_R FILLER_10_35 ();
 DECAPx6_ASAP7_75t_R FILLER_10_43 ();
 DECAPx2_ASAP7_75t_R FILLER_10_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_70 ();
 FILLER_ASAP7_75t_R FILLER_10_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_79 ();
 DECAPx4_ASAP7_75t_R FILLER_10_83 ();
 FILLER_ASAP7_75t_R FILLER_10_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_99 ();
 DECAPx4_ASAP7_75t_R FILLER_10_117 ();
 DECAPx1_ASAP7_75t_R FILLER_10_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_137 ();
 DECAPx10_ASAP7_75t_R FILLER_10_180 ();
 DECAPx10_ASAP7_75t_R FILLER_10_202 ();
 DECAPx6_ASAP7_75t_R FILLER_10_224 ();
 FILLER_ASAP7_75t_R FILLER_10_238 ();
 DECAPx4_ASAP7_75t_R FILLER_10_246 ();
 DECAPx4_ASAP7_75t_R FILLER_10_262 ();
 DECAPx1_ASAP7_75t_R FILLER_11_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_6 ();
 FILLER_ASAP7_75t_R FILLER_11_21 ();
 DECAPx10_ASAP7_75t_R FILLER_11_40 ();
 DECAPx2_ASAP7_75t_R FILLER_11_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_75 ();
 DECAPx2_ASAP7_75t_R FILLER_11_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_104 ();
 DECAPx1_ASAP7_75t_R FILLER_11_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_141 ();
 DECAPx4_ASAP7_75t_R FILLER_11_148 ();
 FILLER_ASAP7_75t_R FILLER_11_158 ();
 DECAPx10_ASAP7_75t_R FILLER_11_166 ();
 DECAPx10_ASAP7_75t_R FILLER_11_188 ();
 DECAPx10_ASAP7_75t_R FILLER_11_210 ();
 DECAPx6_ASAP7_75t_R FILLER_11_232 ();
 FILLER_ASAP7_75t_R FILLER_11_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_248 ();
 DECAPx2_ASAP7_75t_R FILLER_11_255 ();
 DECAPx1_ASAP7_75t_R FILLER_11_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_271 ();
 FILLER_ASAP7_75t_R FILLER_12_2 ();
 FILLER_ASAP7_75t_R FILLER_12_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_25 ();
 DECAPx1_ASAP7_75t_R FILLER_12_29 ();
 DECAPx1_ASAP7_75t_R FILLER_12_78 ();
 DECAPx6_ASAP7_75t_R FILLER_12_103 ();
 DECAPx1_ASAP7_75t_R FILLER_12_117 ();
 DECAPx2_ASAP7_75t_R FILLER_12_131 ();
 DECAPx10_ASAP7_75t_R FILLER_12_159 ();
 DECAPx10_ASAP7_75t_R FILLER_12_181 ();
 DECAPx10_ASAP7_75t_R FILLER_12_203 ();
 DECAPx6_ASAP7_75t_R FILLER_12_225 ();
 DECAPx1_ASAP7_75t_R FILLER_12_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_243 ();
 DECAPx2_ASAP7_75t_R FILLER_12_256 ();
 FILLER_ASAP7_75t_R FILLER_12_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_264 ();
 DECAPx2_ASAP7_75t_R FILLER_12_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_277 ();
 DECAPx6_ASAP7_75t_R FILLER_13_2 ();
 DECAPx6_ASAP7_75t_R FILLER_13_41 ();
 FILLER_ASAP7_75t_R FILLER_13_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_57 ();
 DECAPx1_ASAP7_75t_R FILLER_13_80 ();
 DECAPx2_ASAP7_75t_R FILLER_13_88 ();
 DECAPx2_ASAP7_75t_R FILLER_13_122 ();
 FILLER_ASAP7_75t_R FILLER_13_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_152 ();
 DECAPx10_ASAP7_75t_R FILLER_13_164 ();
 DECAPx10_ASAP7_75t_R FILLER_13_186 ();
 DECAPx10_ASAP7_75t_R FILLER_13_208 ();
 DECAPx4_ASAP7_75t_R FILLER_13_230 ();
 FILLER_ASAP7_75t_R FILLER_13_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_242 ();
 DECAPx6_ASAP7_75t_R FILLER_13_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_263 ();
 FILLER_ASAP7_75t_R FILLER_13_276 ();
 DECAPx4_ASAP7_75t_R FILLER_14_2 ();
 FILLER_ASAP7_75t_R FILLER_14_12 ();
 FILLER_ASAP7_75t_R FILLER_14_18 ();
 DECAPx10_ASAP7_75t_R FILLER_14_41 ();
 DECAPx1_ASAP7_75t_R FILLER_14_63 ();
 DECAPx6_ASAP7_75t_R FILLER_14_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_87 ();
 DECAPx6_ASAP7_75t_R FILLER_14_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_118 ();
 DECAPx2_ASAP7_75t_R FILLER_14_134 ();
 FILLER_ASAP7_75t_R FILLER_14_140 ();
 DECAPx4_ASAP7_75t_R FILLER_14_148 ();
 DECAPx10_ASAP7_75t_R FILLER_14_186 ();
 DECAPx10_ASAP7_75t_R FILLER_14_208 ();
 DECAPx6_ASAP7_75t_R FILLER_14_230 ();
 FILLER_ASAP7_75t_R FILLER_14_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_246 ();
 DECAPx2_ASAP7_75t_R FILLER_14_253 ();
 DECAPx2_ASAP7_75t_R FILLER_14_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_277 ();
 FILLER_ASAP7_75t_R FILLER_15_2 ();
 DECAPx1_ASAP7_75t_R FILLER_15_16 ();
 DECAPx1_ASAP7_75t_R FILLER_15_28 ();
 DECAPx2_ASAP7_75t_R FILLER_15_47 ();
 DECAPx6_ASAP7_75t_R FILLER_15_60 ();
 DECAPx1_ASAP7_75t_R FILLER_15_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_78 ();
 DECAPx6_ASAP7_75t_R FILLER_15_92 ();
 DECAPx1_ASAP7_75t_R FILLER_15_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_110 ();
 DECAPx4_ASAP7_75t_R FILLER_15_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_161 ();
 DECAPx10_ASAP7_75t_R FILLER_15_184 ();
 DECAPx10_ASAP7_75t_R FILLER_15_206 ();
 DECAPx10_ASAP7_75t_R FILLER_15_228 ();
 DECAPx4_ASAP7_75t_R FILLER_15_250 ();
 DECAPx2_ASAP7_75t_R FILLER_16_2 ();
 DECAPx4_ASAP7_75t_R FILLER_16_20 ();
 FILLER_ASAP7_75t_R FILLER_16_30 ();
 DECAPx1_ASAP7_75t_R FILLER_16_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_77 ();
 FILLER_ASAP7_75t_R FILLER_16_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_102 ();
 DECAPx2_ASAP7_75t_R FILLER_16_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_140 ();
 DECAPx6_ASAP7_75t_R FILLER_16_152 ();
 DECAPx2_ASAP7_75t_R FILLER_16_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_172 ();
 DECAPx6_ASAP7_75t_R FILLER_16_180 ();
 DECAPx2_ASAP7_75t_R FILLER_16_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_200 ();
 DECAPx10_ASAP7_75t_R FILLER_16_208 ();
 DECAPx6_ASAP7_75t_R FILLER_16_230 ();
 DECAPx1_ASAP7_75t_R FILLER_16_244 ();
 DECAPx2_ASAP7_75t_R FILLER_16_254 ();
 FILLER_ASAP7_75t_R FILLER_17_2 ();
 FILLER_ASAP7_75t_R FILLER_17_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_12 ();
 DECAPx4_ASAP7_75t_R FILLER_17_45 ();
 FILLER_ASAP7_75t_R FILLER_17_55 ();
 DECAPx6_ASAP7_75t_R FILLER_17_71 ();
 FILLER_ASAP7_75t_R FILLER_17_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_87 ();
 DECAPx4_ASAP7_75t_R FILLER_17_105 ();
 FILLER_ASAP7_75t_R FILLER_17_127 ();
 DECAPx1_ASAP7_75t_R FILLER_17_148 ();
 DECAPx6_ASAP7_75t_R FILLER_17_158 ();
 DECAPx1_ASAP7_75t_R FILLER_17_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_191 ();
 FILLER_ASAP7_75t_R FILLER_17_199 ();
 DECAPx10_ASAP7_75t_R FILLER_17_208 ();
 DECAPx4_ASAP7_75t_R FILLER_17_230 ();
 FILLER_ASAP7_75t_R FILLER_17_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_261 ();
 DECAPx1_ASAP7_75t_R FILLER_17_268 ();
 DECAPx2_ASAP7_75t_R FILLER_18_2 ();
 FILLER_ASAP7_75t_R FILLER_18_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_10 ();
 DECAPx2_ASAP7_75t_R FILLER_18_22 ();
 FILLER_ASAP7_75t_R FILLER_18_28 ();
 DECAPx4_ASAP7_75t_R FILLER_18_42 ();
 FILLER_ASAP7_75t_R FILLER_18_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_54 ();
 DECAPx4_ASAP7_75t_R FILLER_18_74 ();
 DECAPx1_ASAP7_75t_R FILLER_18_106 ();
 DECAPx1_ASAP7_75t_R FILLER_18_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_145 ();
 DECAPx6_ASAP7_75t_R FILLER_18_160 ();
 DECAPx1_ASAP7_75t_R FILLER_18_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_178 ();
 DECAPx2_ASAP7_75t_R FILLER_18_193 ();
 FILLER_ASAP7_75t_R FILLER_18_199 ();
 DECAPx2_ASAP7_75t_R FILLER_18_225 ();
 FILLER_ASAP7_75t_R FILLER_18_231 ();
 FILLER_ASAP7_75t_R FILLER_18_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_247 ();
 DECAPx4_ASAP7_75t_R FILLER_19_2 ();
 DECAPx2_ASAP7_75t_R FILLER_19_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_24 ();
 DECAPx1_ASAP7_75t_R FILLER_19_37 ();
 DECAPx1_ASAP7_75t_R FILLER_19_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_51 ();
 DECAPx1_ASAP7_75t_R FILLER_19_58 ();
 FILLER_ASAP7_75t_R FILLER_19_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_90 ();
 DECAPx4_ASAP7_75t_R FILLER_19_132 ();
 DECAPx4_ASAP7_75t_R FILLER_19_154 ();
 FILLER_ASAP7_75t_R FILLER_19_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_181 ();
 FILLER_ASAP7_75t_R FILLER_19_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_233 ();
 DECAPx2_ASAP7_75t_R FILLER_19_264 ();
 FILLER_ASAP7_75t_R FILLER_19_270 ();
 DECAPx2_ASAP7_75t_R FILLER_20_2 ();
 DECAPx1_ASAP7_75t_R FILLER_20_30 ();
 FILLER_ASAP7_75t_R FILLER_20_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_67 ();
 DECAPx6_ASAP7_75t_R FILLER_20_71 ();
 DECAPx2_ASAP7_75t_R FILLER_20_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_91 ();
 FILLER_ASAP7_75t_R FILLER_20_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_104 ();
 DECAPx4_ASAP7_75t_R FILLER_20_108 ();
 DECAPx10_ASAP7_75t_R FILLER_20_136 ();
 DECAPx6_ASAP7_75t_R FILLER_20_158 ();
 DECAPx2_ASAP7_75t_R FILLER_20_186 ();
 FILLER_ASAP7_75t_R FILLER_20_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_194 ();
 DECAPx4_ASAP7_75t_R FILLER_20_201 ();
 DECAPx2_ASAP7_75t_R FILLER_20_223 ();
 DECAPx1_ASAP7_75t_R FILLER_20_235 ();
 DECAPx1_ASAP7_75t_R FILLER_20_251 ();
 DECAPx1_ASAP7_75t_R FILLER_20_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_271 ();
 DECAPx2_ASAP7_75t_R FILLER_21_2 ();
 FILLER_ASAP7_75t_R FILLER_21_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_10 ();
 DECAPx4_ASAP7_75t_R FILLER_21_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_43 ();
 FILLER_ASAP7_75t_R FILLER_21_48 ();
 FILLER_ASAP7_75t_R FILLER_21_56 ();
 FILLER_ASAP7_75t_R FILLER_21_94 ();
 DECAPx10_ASAP7_75t_R FILLER_21_104 ();
 DECAPx10_ASAP7_75t_R FILLER_21_126 ();
 DECAPx10_ASAP7_75t_R FILLER_21_148 ();
 DECAPx1_ASAP7_75t_R FILLER_21_170 ();
 DECAPx2_ASAP7_75t_R FILLER_21_181 ();
 FILLER_ASAP7_75t_R FILLER_21_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_189 ();
 DECAPx1_ASAP7_75t_R FILLER_21_202 ();
 DECAPx4_ASAP7_75t_R FILLER_21_218 ();
 FILLER_ASAP7_75t_R FILLER_21_228 ();
 DECAPx2_ASAP7_75t_R FILLER_21_236 ();
 FILLER_ASAP7_75t_R FILLER_21_254 ();
 DECAPx1_ASAP7_75t_R FILLER_21_268 ();
 DECAPx1_ASAP7_75t_R FILLER_22_14 ();
 FILLER_ASAP7_75t_R FILLER_22_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_60 ();
 DECAPx1_ASAP7_75t_R FILLER_22_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_71 ();
 DECAPx10_ASAP7_75t_R FILLER_22_88 ();
 FILLER_ASAP7_75t_R FILLER_22_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_131 ();
 DECAPx1_ASAP7_75t_R FILLER_22_166 ();
 DECAPx4_ASAP7_75t_R FILLER_22_180 ();
 DECAPx1_ASAP7_75t_R FILLER_22_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_231 ();
 FILLER_ASAP7_75t_R FILLER_22_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_240 ();
 FILLER_ASAP7_75t_R FILLER_22_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_261 ();
 DECAPx1_ASAP7_75t_R FILLER_22_274 ();
 FILLER_ASAP7_75t_R FILLER_23_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_26 ();
 FILLER_ASAP7_75t_R FILLER_23_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_35 ();
 DECAPx2_ASAP7_75t_R FILLER_23_58 ();
 DECAPx4_ASAP7_75t_R FILLER_23_76 ();
 DECAPx2_ASAP7_75t_R FILLER_23_102 ();
 FILLER_ASAP7_75t_R FILLER_23_108 ();
 DECAPx2_ASAP7_75t_R FILLER_23_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_138 ();
 DECAPx10_ASAP7_75t_R FILLER_23_145 ();
 DECAPx6_ASAP7_75t_R FILLER_23_167 ();
 DECAPx2_ASAP7_75t_R FILLER_23_181 ();
 FILLER_ASAP7_75t_R FILLER_23_206 ();
 FILLER_ASAP7_75t_R FILLER_23_214 ();
 FILLER_ASAP7_75t_R FILLER_23_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_253 ();
 DECAPx6_ASAP7_75t_R FILLER_24_2 ();
 DECAPx1_ASAP7_75t_R FILLER_24_16 ();
 DECAPx10_ASAP7_75t_R FILLER_24_30 ();
 DECAPx10_ASAP7_75t_R FILLER_24_52 ();
 DECAPx4_ASAP7_75t_R FILLER_24_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_101 ();
 DECAPx10_ASAP7_75t_R FILLER_24_105 ();
 DECAPx2_ASAP7_75t_R FILLER_24_127 ();
 FILLER_ASAP7_75t_R FILLER_24_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_135 ();
 FILLER_ASAP7_75t_R FILLER_24_142 ();
 DECAPx10_ASAP7_75t_R FILLER_24_170 ();
 FILLER_ASAP7_75t_R FILLER_24_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_194 ();
 DECAPx1_ASAP7_75t_R FILLER_24_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_209 ();
 DECAPx2_ASAP7_75t_R FILLER_24_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_277 ();
 FILLER_ASAP7_75t_R FILLER_25_14 ();
 DECAPx1_ASAP7_75t_R FILLER_25_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_40 ();
 FILLER_ASAP7_75t_R FILLER_25_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_65 ();
 FILLER_ASAP7_75t_R FILLER_25_73 ();
 DECAPx2_ASAP7_75t_R FILLER_25_82 ();
 FILLER_ASAP7_75t_R FILLER_25_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_90 ();
 DECAPx4_ASAP7_75t_R FILLER_25_108 ();
 DECAPx2_ASAP7_75t_R FILLER_25_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_130 ();
 DECAPx4_ASAP7_75t_R FILLER_25_169 ();
 FILLER_ASAP7_75t_R FILLER_25_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_181 ();
 DECAPx10_ASAP7_75t_R FILLER_25_192 ();
 DECAPx4_ASAP7_75t_R FILLER_25_226 ();
 FILLER_ASAP7_75t_R FILLER_25_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_238 ();
 FILLER_ASAP7_75t_R FILLER_25_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_277 ();
 DECAPx4_ASAP7_75t_R FILLER_26_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_12 ();
 DECAPx2_ASAP7_75t_R FILLER_26_36 ();
 FILLER_ASAP7_75t_R FILLER_26_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_44 ();
 DECAPx4_ASAP7_75t_R FILLER_26_69 ();
 DECAPx1_ASAP7_75t_R FILLER_26_85 ();
 FILLER_ASAP7_75t_R FILLER_26_97 ();
 DECAPx2_ASAP7_75t_R FILLER_26_149 ();
 FILLER_ASAP7_75t_R FILLER_26_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_161 ();
 DECAPx6_ASAP7_75t_R FILLER_26_169 ();
 FILLER_ASAP7_75t_R FILLER_26_183 ();
 DECAPx2_ASAP7_75t_R FILLER_26_195 ();
 FILLER_ASAP7_75t_R FILLER_26_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_221 ();
 FILLER_ASAP7_75t_R FILLER_26_234 ();
 FILLER_ASAP7_75t_R FILLER_26_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_257 ();
 FILLER_ASAP7_75t_R FILLER_26_276 ();
 FILLER_ASAP7_75t_R FILLER_27_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_22 ();
 DECAPx2_ASAP7_75t_R FILLER_27_46 ();
 DECAPx1_ASAP7_75t_R FILLER_27_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_63 ();
 FILLER_ASAP7_75t_R FILLER_27_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_72 ();
 FILLER_ASAP7_75t_R FILLER_27_90 ();
 DECAPx6_ASAP7_75t_R FILLER_27_99 ();
 DECAPx6_ASAP7_75t_R FILLER_27_124 ();
 FILLER_ASAP7_75t_R FILLER_27_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_157 ();
 DECAPx6_ASAP7_75t_R FILLER_27_167 ();
 FILLER_ASAP7_75t_R FILLER_27_181 ();
 DECAPx6_ASAP7_75t_R FILLER_27_193 ();
 DECAPx1_ASAP7_75t_R FILLER_27_207 ();
 DECAPx6_ASAP7_75t_R FILLER_27_217 ();
 DECAPx1_ASAP7_75t_R FILLER_27_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_241 ();
 DECAPx2_ASAP7_75t_R FILLER_27_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_268 ();
 FILLER_ASAP7_75t_R FILLER_27_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_277 ();
 FILLER_ASAP7_75t_R FILLER_28_2 ();
 DECAPx2_ASAP7_75t_R FILLER_28_10 ();
 DECAPx2_ASAP7_75t_R FILLER_28_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_42 ();
 FILLER_ASAP7_75t_R FILLER_28_58 ();
 DECAPx2_ASAP7_75t_R FILLER_28_68 ();
 FILLER_ASAP7_75t_R FILLER_28_74 ();
 FILLER_ASAP7_75t_R FILLER_28_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_88 ();
 DECAPx6_ASAP7_75t_R FILLER_28_96 ();
 DECAPx2_ASAP7_75t_R FILLER_28_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_116 ();
 DECAPx2_ASAP7_75t_R FILLER_28_143 ();
 FILLER_ASAP7_75t_R FILLER_28_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_151 ();
 DECAPx6_ASAP7_75t_R FILLER_28_162 ();
 DECAPx1_ASAP7_75t_R FILLER_28_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_180 ();
 DECAPx4_ASAP7_75t_R FILLER_28_191 ();
 DECAPx1_ASAP7_75t_R FILLER_28_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_211 ();
 DECAPx4_ASAP7_75t_R FILLER_28_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_234 ();
 FILLER_ASAP7_75t_R FILLER_28_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_277 ();
 DECAPx2_ASAP7_75t_R FILLER_29_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_14 ();
 DECAPx2_ASAP7_75t_R FILLER_29_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_27 ();
 DECAPx1_ASAP7_75t_R FILLER_29_39 ();
 DECAPx2_ASAP7_75t_R FILLER_29_50 ();
 FILLER_ASAP7_75t_R FILLER_29_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_58 ();
 DECAPx2_ASAP7_75t_R FILLER_29_69 ();
 FILLER_ASAP7_75t_R FILLER_29_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_83 ();
 DECAPx6_ASAP7_75t_R FILLER_29_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_107 ();
 DECAPx1_ASAP7_75t_R FILLER_29_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_141 ();
 DECAPx4_ASAP7_75t_R FILLER_29_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_158 ();
 DECAPx6_ASAP7_75t_R FILLER_29_170 ();
 DECAPx10_ASAP7_75t_R FILLER_29_221 ();
 DECAPx2_ASAP7_75t_R FILLER_29_243 ();
 FILLER_ASAP7_75t_R FILLER_29_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_251 ();
 DECAPx1_ASAP7_75t_R FILLER_29_265 ();
 FILLER_ASAP7_75t_R FILLER_29_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_277 ();
 DECAPx1_ASAP7_75t_R FILLER_30_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_6 ();
 DECAPx4_ASAP7_75t_R FILLER_30_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_23 ();
 DECAPx1_ASAP7_75t_R FILLER_30_30 ();
 DECAPx2_ASAP7_75t_R FILLER_30_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_43 ();
 FILLER_ASAP7_75t_R FILLER_30_58 ();
 DECAPx4_ASAP7_75t_R FILLER_30_67 ();
 FILLER_ASAP7_75t_R FILLER_30_77 ();
 DECAPx1_ASAP7_75t_R FILLER_30_85 ();
 DECAPx6_ASAP7_75t_R FILLER_30_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_119 ();
 DECAPx10_ASAP7_75t_R FILLER_30_132 ();
 DECAPx4_ASAP7_75t_R FILLER_30_163 ();
 DECAPx10_ASAP7_75t_R FILLER_30_183 ();
 DECAPx10_ASAP7_75t_R FILLER_30_205 ();
 DECAPx4_ASAP7_75t_R FILLER_30_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_237 ();
 DECAPx1_ASAP7_75t_R FILLER_30_268 ();
 FILLER_ASAP7_75t_R FILLER_31_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_10 ();
 DECAPx2_ASAP7_75t_R FILLER_31_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_47 ();
 FILLER_ASAP7_75t_R FILLER_31_60 ();
 FILLER_ASAP7_75t_R FILLER_31_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_70 ();
 FILLER_ASAP7_75t_R FILLER_31_77 ();
 FILLER_ASAP7_75t_R FILLER_31_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_94 ();
 DECAPx10_ASAP7_75t_R FILLER_31_117 ();
 DECAPx2_ASAP7_75t_R FILLER_31_139 ();
 FILLER_ASAP7_75t_R FILLER_31_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_147 ();
 DECAPx2_ASAP7_75t_R FILLER_31_162 ();
 DECAPx10_ASAP7_75t_R FILLER_31_180 ();
 DECAPx10_ASAP7_75t_R FILLER_31_202 ();
 DECAPx4_ASAP7_75t_R FILLER_31_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_271 ();
 DECAPx2_ASAP7_75t_R FILLER_32_2 ();
 FILLER_ASAP7_75t_R FILLER_32_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_33 ();
 FILLER_ASAP7_75t_R FILLER_32_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_42 ();
 DECAPx1_ASAP7_75t_R FILLER_32_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_56 ();
 DECAPx4_ASAP7_75t_R FILLER_32_72 ();
 FILLER_ASAP7_75t_R FILLER_32_82 ();
 DECAPx10_ASAP7_75t_R FILLER_32_90 ();
 DECAPx6_ASAP7_75t_R FILLER_32_112 ();
 FILLER_ASAP7_75t_R FILLER_32_126 ();
 DECAPx4_ASAP7_75t_R FILLER_32_156 ();
 FILLER_ASAP7_75t_R FILLER_32_166 ();
 DECAPx2_ASAP7_75t_R FILLER_32_180 ();
 FILLER_ASAP7_75t_R FILLER_32_186 ();
 DECAPx10_ASAP7_75t_R FILLER_32_208 ();
 DECAPx6_ASAP7_75t_R FILLER_32_230 ();
 DECAPx2_ASAP7_75t_R FILLER_32_256 ();
 DECAPx1_ASAP7_75t_R FILLER_32_274 ();
 DECAPx2_ASAP7_75t_R FILLER_33_8 ();
 FILLER_ASAP7_75t_R FILLER_33_29 ();
 DECAPx1_ASAP7_75t_R FILLER_33_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_41 ();
 FILLER_ASAP7_75t_R FILLER_33_52 ();
 FILLER_ASAP7_75t_R FILLER_33_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_65 ();
 DECAPx1_ASAP7_75t_R FILLER_33_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_87 ();
 DECAPx2_ASAP7_75t_R FILLER_33_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_104 ();
 DECAPx2_ASAP7_75t_R FILLER_33_125 ();
 FILLER_ASAP7_75t_R FILLER_33_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_133 ();
 FILLER_ASAP7_75t_R FILLER_33_150 ();
 DECAPx1_ASAP7_75t_R FILLER_33_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_166 ();
 DECAPx4_ASAP7_75t_R FILLER_33_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_221 ();
 FILLER_ASAP7_75t_R FILLER_33_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_240 ();
 FILLER_ASAP7_75t_R FILLER_33_257 ();
 DECAPx2_ASAP7_75t_R FILLER_34_2 ();
 DECAPx4_ASAP7_75t_R FILLER_34_38 ();
 DECAPx6_ASAP7_75t_R FILLER_34_63 ();
 FILLER_ASAP7_75t_R FILLER_34_77 ();
 DECAPx2_ASAP7_75t_R FILLER_34_86 ();
 FILLER_ASAP7_75t_R FILLER_34_92 ();
 DECAPx4_ASAP7_75t_R FILLER_34_112 ();
 DECAPx10_ASAP7_75t_R FILLER_34_132 ();
 DECAPx1_ASAP7_75t_R FILLER_34_160 ();
 DECAPx4_ASAP7_75t_R FILLER_34_170 ();
 FILLER_ASAP7_75t_R FILLER_34_180 ();
 FILLER_ASAP7_75t_R FILLER_34_192 ();
 DECAPx1_ASAP7_75t_R FILLER_34_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_208 ();
 FILLER_ASAP7_75t_R FILLER_34_215 ();
 DECAPx1_ASAP7_75t_R FILLER_34_224 ();
 DECAPx1_ASAP7_75t_R FILLER_34_234 ();
 FILLER_ASAP7_75t_R FILLER_34_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_277 ();
 DECAPx2_ASAP7_75t_R FILLER_35_2 ();
 DECAPx2_ASAP7_75t_R FILLER_35_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_26 ();
 FILLER_ASAP7_75t_R FILLER_35_33 ();
 DECAPx6_ASAP7_75t_R FILLER_35_68 ();
 DECAPx6_ASAP7_75t_R FILLER_35_135 ();
 DECAPx2_ASAP7_75t_R FILLER_35_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_179 ();
 DECAPx4_ASAP7_75t_R FILLER_35_192 ();
 FILLER_ASAP7_75t_R FILLER_35_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_204 ();
 DECAPx4_ASAP7_75t_R FILLER_35_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_253 ();
 DECAPx2_ASAP7_75t_R FILLER_36_2 ();
 FILLER_ASAP7_75t_R FILLER_36_8 ();
 DECAPx1_ASAP7_75t_R FILLER_36_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_20 ();
 FILLER_ASAP7_75t_R FILLER_36_50 ();
 FILLER_ASAP7_75t_R FILLER_36_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_66 ();
 FILLER_ASAP7_75t_R FILLER_36_83 ();
 DECAPx10_ASAP7_75t_R FILLER_36_95 ();
 DECAPx10_ASAP7_75t_R FILLER_36_117 ();
 DECAPx4_ASAP7_75t_R FILLER_36_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_179 ();
 DECAPx6_ASAP7_75t_R FILLER_36_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_219 ();
 FILLER_ASAP7_75t_R FILLER_36_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_234 ();
 DECAPx1_ASAP7_75t_R FILLER_36_241 ();
 FILLER_ASAP7_75t_R FILLER_36_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_271 ();
 DECAPx4_ASAP7_75t_R FILLER_37_2 ();
 DECAPx4_ASAP7_75t_R FILLER_37_24 ();
 FILLER_ASAP7_75t_R FILLER_37_40 ();
 DECAPx10_ASAP7_75t_R FILLER_37_75 ();
 DECAPx4_ASAP7_75t_R FILLER_37_97 ();
 FILLER_ASAP7_75t_R FILLER_37_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_109 ();
 DECAPx10_ASAP7_75t_R FILLER_37_116 ();
 DECAPx10_ASAP7_75t_R FILLER_37_138 ();
 DECAPx2_ASAP7_75t_R FILLER_37_160 ();
 FILLER_ASAP7_75t_R FILLER_37_166 ();
 DECAPx1_ASAP7_75t_R FILLER_37_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_179 ();
 DECAPx2_ASAP7_75t_R FILLER_37_190 ();
 FILLER_ASAP7_75t_R FILLER_37_196 ();
 FILLER_ASAP7_75t_R FILLER_37_214 ();
 DECAPx1_ASAP7_75t_R FILLER_37_252 ();
 DECAPx1_ASAP7_75t_R FILLER_37_274 ();
 FILLER_ASAP7_75t_R FILLER_38_2 ();
 DECAPx2_ASAP7_75t_R FILLER_38_10 ();
 DECAPx6_ASAP7_75t_R FILLER_38_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_36 ();
 DECAPx10_ASAP7_75t_R FILLER_38_47 ();
 DECAPx4_ASAP7_75t_R FILLER_38_69 ();
 FILLER_ASAP7_75t_R FILLER_38_79 ();
 DECAPx4_ASAP7_75t_R FILLER_38_91 ();
 FILLER_ASAP7_75t_R FILLER_38_107 ();
 DECAPx4_ASAP7_75t_R FILLER_38_115 ();
 FILLER_ASAP7_75t_R FILLER_38_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_127 ();
 DECAPx4_ASAP7_75t_R FILLER_38_138 ();
 FILLER_ASAP7_75t_R FILLER_38_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_206 ();
 DECAPx2_ASAP7_75t_R FILLER_38_225 ();
 FILLER_ASAP7_75t_R FILLER_38_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_233 ();
 FILLER_ASAP7_75t_R FILLER_38_252 ();
 DECAPx1_ASAP7_75t_R FILLER_39_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_6 ();
 DECAPx10_ASAP7_75t_R FILLER_39_13 ();
 DECAPx4_ASAP7_75t_R FILLER_39_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_52 ();
 DECAPx4_ASAP7_75t_R FILLER_39_59 ();
 FILLER_ASAP7_75t_R FILLER_39_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_89 ();
 FILLER_ASAP7_75t_R FILLER_39_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_147 ();
 FILLER_ASAP7_75t_R FILLER_39_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_172 ();
 DECAPx6_ASAP7_75t_R FILLER_39_179 ();
 DECAPx6_ASAP7_75t_R FILLER_39_203 ();
 FILLER_ASAP7_75t_R FILLER_39_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_231 ();
 FILLER_ASAP7_75t_R FILLER_39_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_277 ();
 DECAPx10_ASAP7_75t_R FILLER_40_2 ();
 DECAPx6_ASAP7_75t_R FILLER_40_24 ();
 DECAPx1_ASAP7_75t_R FILLER_40_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_42 ();
 DECAPx10_ASAP7_75t_R FILLER_40_50 ();
 FILLER_ASAP7_75t_R FILLER_40_72 ();
 DECAPx2_ASAP7_75t_R FILLER_40_94 ();
 FILLER_ASAP7_75t_R FILLER_40_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_112 ();
 DECAPx4_ASAP7_75t_R FILLER_40_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_145 ();
 DECAPx1_ASAP7_75t_R FILLER_40_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_183 ();
 FILLER_ASAP7_75t_R FILLER_40_228 ();
 FILLER_ASAP7_75t_R FILLER_40_242 ();
 DECAPx1_ASAP7_75t_R FILLER_40_268 ();
 DECAPx10_ASAP7_75t_R FILLER_41_2 ();
 DECAPx10_ASAP7_75t_R FILLER_41_24 ();
 DECAPx2_ASAP7_75t_R FILLER_41_46 ();
 DECAPx10_ASAP7_75t_R FILLER_41_62 ();
 DECAPx4_ASAP7_75t_R FILLER_41_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_94 ();
 DECAPx2_ASAP7_75t_R FILLER_41_107 ();
 FILLER_ASAP7_75t_R FILLER_41_113 ();
 DECAPx4_ASAP7_75t_R FILLER_41_121 ();
 DECAPx10_ASAP7_75t_R FILLER_41_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_159 ();
 DECAPx4_ASAP7_75t_R FILLER_41_170 ();
 DECAPx4_ASAP7_75t_R FILLER_41_190 ();
 FILLER_ASAP7_75t_R FILLER_41_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_202 ();
 FILLER_ASAP7_75t_R FILLER_41_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_235 ();
 DECAPx10_ASAP7_75t_R FILLER_42_2 ();
 DECAPx6_ASAP7_75t_R FILLER_42_24 ();
 DECAPx2_ASAP7_75t_R FILLER_42_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_44 ();
 DECAPx4_ASAP7_75t_R FILLER_42_52 ();
 FILLER_ASAP7_75t_R FILLER_42_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_70 ();
 FILLER_ASAP7_75t_R FILLER_42_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_83 ();
 DECAPx2_ASAP7_75t_R FILLER_42_94 ();
 FILLER_ASAP7_75t_R FILLER_42_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_102 ();
 DECAPx2_ASAP7_75t_R FILLER_42_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_123 ();
 DECAPx1_ASAP7_75t_R FILLER_42_136 ();
 DECAPx2_ASAP7_75t_R FILLER_42_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_156 ();
 DECAPx4_ASAP7_75t_R FILLER_42_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_241 ();
 FILLER_ASAP7_75t_R FILLER_42_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_256 ();
 FILLER_ASAP7_75t_R FILLER_42_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_277 ();
 DECAPx10_ASAP7_75t_R FILLER_43_2 ();
 DECAPx6_ASAP7_75t_R FILLER_43_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_48 ();
 DECAPx2_ASAP7_75t_R FILLER_43_55 ();
 DECAPx6_ASAP7_75t_R FILLER_43_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_81 ();
 FILLER_ASAP7_75t_R FILLER_43_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_105 ();
 FILLER_ASAP7_75t_R FILLER_43_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_150 ();
 DECAPx6_ASAP7_75t_R FILLER_43_158 ();
 FILLER_ASAP7_75t_R FILLER_43_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_174 ();
 DECAPx1_ASAP7_75t_R FILLER_43_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_189 ();
 DECAPx1_ASAP7_75t_R FILLER_43_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_200 ();
 DECAPx2_ASAP7_75t_R FILLER_43_219 ();
 FILLER_ASAP7_75t_R FILLER_43_225 ();
 FILLER_ASAP7_75t_R FILLER_43_237 ();
 FILLER_ASAP7_75t_R FILLER_43_276 ();
 DECAPx10_ASAP7_75t_R FILLER_44_2 ();
 DECAPx2_ASAP7_75t_R FILLER_44_24 ();
 FILLER_ASAP7_75t_R FILLER_44_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_45 ();
 DECAPx1_ASAP7_75t_R FILLER_44_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_68 ();
 DECAPx4_ASAP7_75t_R FILLER_44_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_92 ();
 DECAPx2_ASAP7_75t_R FILLER_44_99 ();
 FILLER_ASAP7_75t_R FILLER_44_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_107 ();
 DECAPx6_ASAP7_75t_R FILLER_44_114 ();
 FILLER_ASAP7_75t_R FILLER_44_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_130 ();
 FILLER_ASAP7_75t_R FILLER_44_143 ();
 DECAPx10_ASAP7_75t_R FILLER_44_151 ();
 FILLER_ASAP7_75t_R FILLER_44_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_175 ();
 DECAPx4_ASAP7_75t_R FILLER_44_183 ();
 FILLER_ASAP7_75t_R FILLER_44_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_213 ();
 FILLER_ASAP7_75t_R FILLER_44_239 ();
 FILLER_ASAP7_75t_R FILLER_44_247 ();
 DECAPx1_ASAP7_75t_R FILLER_44_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_271 ();
 DECAPx10_ASAP7_75t_R FILLER_45_2 ();
 DECAPx6_ASAP7_75t_R FILLER_45_24 ();
 DECAPx1_ASAP7_75t_R FILLER_45_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_68 ();
 FILLER_ASAP7_75t_R FILLER_45_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_99 ();
 FILLER_ASAP7_75t_R FILLER_45_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_108 ();
 DECAPx10_ASAP7_75t_R FILLER_45_121 ();
 FILLER_ASAP7_75t_R FILLER_45_143 ();
 DECAPx1_ASAP7_75t_R FILLER_45_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_199 ();
 FILLER_ASAP7_75t_R FILLER_45_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_230 ();
 FILLER_ASAP7_75t_R FILLER_45_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_269 ();
 FILLER_ASAP7_75t_R FILLER_45_276 ();
 DECAPx10_ASAP7_75t_R FILLER_46_2 ();
 DECAPx2_ASAP7_75t_R FILLER_46_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_30 ();
 DECAPx2_ASAP7_75t_R FILLER_46_43 ();
 FILLER_ASAP7_75t_R FILLER_46_49 ();
 FILLER_ASAP7_75t_R FILLER_46_57 ();
 FILLER_ASAP7_75t_R FILLER_46_71 ();
 DECAPx6_ASAP7_75t_R FILLER_46_79 ();
 FILLER_ASAP7_75t_R FILLER_46_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_95 ();
 DECAPx1_ASAP7_75t_R FILLER_46_108 ();
 DECAPx1_ASAP7_75t_R FILLER_46_118 ();
 DECAPx1_ASAP7_75t_R FILLER_46_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_138 ();
 DECAPx1_ASAP7_75t_R FILLER_46_155 ();
 FILLER_ASAP7_75t_R FILLER_46_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_179 ();
 FILLER_ASAP7_75t_R FILLER_46_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_202 ();
 FILLER_ASAP7_75t_R FILLER_46_243 ();
 DECAPx2_ASAP7_75t_R FILLER_46_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_271 ();
 DECAPx10_ASAP7_75t_R FILLER_47_2 ();
 DECAPx2_ASAP7_75t_R FILLER_47_24 ();
 FILLER_ASAP7_75t_R FILLER_47_30 ();
 FILLER_ASAP7_75t_R FILLER_47_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_52 ();
 DECAPx2_ASAP7_75t_R FILLER_47_65 ();
 FILLER_ASAP7_75t_R FILLER_47_71 ();
 FILLER_ASAP7_75t_R FILLER_47_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_101 ();
 FILLER_ASAP7_75t_R FILLER_47_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_116 ();
 FILLER_ASAP7_75t_R FILLER_47_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_131 ();
 DECAPx2_ASAP7_75t_R FILLER_47_142 ();
 FILLER_ASAP7_75t_R FILLER_47_160 ();
 FILLER_ASAP7_75t_R FILLER_47_168 ();
 DECAPx4_ASAP7_75t_R FILLER_47_176 ();
 FILLER_ASAP7_75t_R FILLER_47_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_247 ();
 DECAPx6_ASAP7_75t_R FILLER_48_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_16 ();
 FILLER_ASAP7_75t_R FILLER_48_100 ();
 FILLER_ASAP7_75t_R FILLER_48_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_134 ();
 FILLER_ASAP7_75t_R FILLER_48_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_153 ();
 FILLER_ASAP7_75t_R FILLER_48_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_174 ();
 DECAPx1_ASAP7_75t_R FILLER_48_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_192 ();
 FILLER_ASAP7_75t_R FILLER_48_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_232 ();
 FILLER_ASAP7_75t_R FILLER_48_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_271 ();
 DECAPx6_ASAP7_75t_R FILLER_49_2 ();
 FILLER_ASAP7_75t_R FILLER_49_16 ();
 FILLER_ASAP7_75t_R FILLER_49_42 ();
 FILLER_ASAP7_75t_R FILLER_49_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_90 ();
 DECAPx2_ASAP7_75t_R FILLER_49_121 ();
 FILLER_ASAP7_75t_R FILLER_49_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_193 ();
 DECAPx1_ASAP7_75t_R FILLER_49_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_234 ();
 FILLER_ASAP7_75t_R FILLER_49_247 ();
 DECAPx1_ASAP7_75t_R FILLER_49_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_271 ();
 DECAPx4_ASAP7_75t_R FILLER_50_2 ();
 DECAPx2_ASAP7_75t_R FILLER_50_18 ();
 FILLER_ASAP7_75t_R FILLER_50_36 ();
 FILLER_ASAP7_75t_R FILLER_50_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_83 ();
 FILLER_ASAP7_75t_R FILLER_50_90 ();
 FILLER_ASAP7_75t_R FILLER_50_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_106 ();
 DECAPx2_ASAP7_75t_R FILLER_50_125 ();
 FILLER_ASAP7_75t_R FILLER_50_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_182 ();
 FILLER_ASAP7_75t_R FILLER_50_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_197 ();
 FILLER_ASAP7_75t_R FILLER_50_204 ();
 DECAPx1_ASAP7_75t_R FILLER_50_224 ();
 FILLER_ASAP7_75t_R FILLER_50_270 ();
 DECAPx2_ASAP7_75t_R FILLER_51_2 ();
 FILLER_ASAP7_75t_R FILLER_51_110 ();
 DECAPx1_ASAP7_75t_R FILLER_51_136 ();
 DECAPx1_ASAP7_75t_R FILLER_51_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_162 ();
 FILLER_ASAP7_75t_R FILLER_51_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_250 ();
 FILLER_ASAP7_75t_R FILLER_51_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_271 ();
 DECAPx1_ASAP7_75t_R FILLER_52_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_62 ();
 FILLER_ASAP7_75t_R FILLER_52_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_94 ();
 FILLER_ASAP7_75t_R FILLER_52_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_192 ();
 FILLER_ASAP7_75t_R FILLER_52_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_236 ();
 DECAPx2_ASAP7_75t_R FILLER_52_269 ();
 FILLER_ASAP7_75t_R FILLER_52_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_277 ();
 FILLER_ASAP7_75t_R FILLER_53_2 ();
 FILLER_ASAP7_75t_R FILLER_53_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_12 ();
 FILLER_ASAP7_75t_R FILLER_53_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_62 ();
 FILLER_ASAP7_75t_R FILLER_53_69 ();
 FILLER_ASAP7_75t_R FILLER_53_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_83 ();
 FILLER_ASAP7_75t_R FILLER_53_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_93 ();
 DECAPx2_ASAP7_75t_R FILLER_53_100 ();
 FILLER_ASAP7_75t_R FILLER_53_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_152 ();
 FILLER_ASAP7_75t_R FILLER_53_159 ();
 FILLER_ASAP7_75t_R FILLER_53_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_169 ();
 FILLER_ASAP7_75t_R FILLER_53_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_182 ();
 FILLER_ASAP7_75t_R FILLER_53_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_262 ();
 FILLER_ASAP7_75t_R FILLER_53_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_277 ();
 DECAPx2_ASAP7_75t_R FILLER_54_2 ();
endmodule
