module credit_pi_switch (clk,
    rst,
    l_i,
    l_i_bp,
    l_i_v,
    l_o,
    l_o_credit_gnt,
    l_o_v,
    r_i,
    r_i_bp,
    r_i_v,
    r_o,
    r_o_credit_gnt,
    r_o_v,
    u0_i,
    u0_i_bp,
    u0_i_v,
    u0_o,
    u0_o_credit_gnt,
    u0_o_v,
    u1_i,
    u1_i_bp,
    u1_i_v,
    u1_o,
    u1_o_credit_gnt,
    u1_o_v);
 input clk;
 input rst;
 input [73:0] l_i;
 output [1:0] l_i_bp;
 input [1:0] l_i_v;
 output [36:0] l_o;
 input [1:0] l_o_credit_gnt;
 output [1:0] l_o_v;
 input [73:0] r_i;
 output [1:0] r_i_bp;
 input [1:0] r_i_v;
 output [36:0] r_o;
 input [1:0] r_o_credit_gnt;
 output [1:0] r_o_v;
 input [73:0] u0_i;
 output [1:0] u0_i_bp;
 input [1:0] u0_i_v;
 output [36:0] u0_o;
 input [1:0] u0_o_credit_gnt;
 output [1:0] u0_o_v;
 input [73:0] u1_i;
 output [1:0] u1_i_bp;
 input [1:0] u1_i_v;
 output [36:0] u1_o;
 input [1:0] u1_o_credit_gnt;
 output [1:0] u1_o_v;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire \credit_pi_route_inst.l_counters_inst.o_credits[1] ;
 wire \credit_pi_route_inst.l_counters_inst.o_credits[2] ;
 wire \credit_pi_route_inst.l_counters_inst.o_credits[3] ;
 wire \credit_pi_route_inst.l_counters_inst.o_credits[6] ;
 wire \credit_pi_route_inst.l_counters_inst.o_credits[7] ;
 wire \credit_pi_route_inst.l_counters_inst.o_credits[8] ;
 wire \credit_pi_route_inst.r_counters_inst.o_credits[1] ;
 wire \credit_pi_route_inst.r_counters_inst.o_credits[2] ;
 wire \credit_pi_route_inst.r_counters_inst.o_credits[3] ;
 wire \credit_pi_route_inst.r_counters_inst.o_credits[6] ;
 wire \credit_pi_route_inst.r_counters_inst.o_credits[7] ;
 wire \credit_pi_route_inst.r_counters_inst.o_credits[8] ;
 wire \credit_pi_route_inst.u0_counters_inst.o_credits[1] ;
 wire \credit_pi_route_inst.u0_counters_inst.o_credits[2] ;
 wire \credit_pi_route_inst.u0_counters_inst.o_credits[3] ;
 wire \credit_pi_route_inst.u0_counters_inst.o_credits[5] ;
 wire \credit_pi_route_inst.u0_counters_inst.o_credits[6] ;
 wire \credit_pi_route_inst.u0_counters_inst.o_credits[7] ;
 wire \credit_pi_route_inst.u0_counters_inst.o_credits[8] ;
 wire \credit_pi_route_inst.u1_counters_inst.o_credits[1] ;
 wire \credit_pi_route_inst.u1_counters_inst.o_credits[2] ;
 wire \credit_pi_route_inst.u1_counters_inst.o_credits[3] ;
 wire \credit_pi_route_inst.u1_counters_inst.o_credits[5] ;
 wire \credit_pi_route_inst.u1_counters_inst.o_credits[6] ;
 wire \credit_pi_route_inst.u1_counters_inst.o_credits[7] ;
 wire \credit_pi_route_inst.u1_counters_inst.o_credits[8] ;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 INVx1_ASAP7_75t_R _1181_ (.A(_1171_),
    .Y(\credit_pi_route_inst.l_counters_inst.o_credits[6] ));
 INVx1_ASAP7_75t_R _1182_ (.A(_0092_),
    .Y(\credit_pi_route_inst.l_counters_inst.o_credits[8] ));
 INVx1_ASAP7_75t_R _1183_ (.A(_0093_),
    .Y(\credit_pi_route_inst.l_counters_inst.o_credits[7] ));
 INVx1_ASAP7_75t_R _1184_ (.A(_1173_),
    .Y(\credit_pi_route_inst.l_counters_inst.o_credits[1] ));
 INVx1_ASAP7_75t_R _1185_ (.A(_0095_),
    .Y(\credit_pi_route_inst.l_counters_inst.o_credits[3] ));
 INVx1_ASAP7_75t_R _1186_ (.A(_0096_),
    .Y(\credit_pi_route_inst.l_counters_inst.o_credits[2] ));
 INVx1_ASAP7_75t_R _1187_ (.A(net261),
    .Y(_0916_));
 INVx1_ASAP7_75t_R _1188_ (.A(net301),
    .Y(_0917_));
 AO22x2_ASAP7_75t_R _1189_ (.A1(_0916_),
    .A2(net310),
    .B1(net311),
    .B2(_0917_),
    .Y(_0918_));
 INVx1_ASAP7_75t_R _1190_ (.A(net183),
    .Y(_0919_));
 INVx1_ASAP7_75t_R _1191_ (.A(net223),
    .Y(_0920_));
 AO22x2_ASAP7_75t_R _1192_ (.A1(_0919_),
    .A2(net232),
    .B1(net233),
    .B2(_0920_),
    .Y(_0921_));
 OA21x2_ASAP7_75t_R _1193_ (.A1(_0918_),
    .A2(_0921_),
    .B(_0099_),
    .Y(_0922_));
 INVx1_ASAP7_75t_R _1194_ (.A(net154),
    .Y(_0923_));
 OR3x2_ASAP7_75t_R _1195_ (.A(net148),
    .B(net147),
    .C(net146),
    .Y(_0924_));
 OR3x2_ASAP7_75t_R _1196_ (.A(net144),
    .B(_0923_),
    .C(_0924_),
    .Y(_0925_));
 AND5x2_ASAP7_75t_R _1197_ (.A(_0091_),
    .B(_0092_),
    .C(_0093_),
    .D(_1171_),
    .E(_0062_),
    .Y(_0926_));
 AND5x2_ASAP7_75t_R _1198_ (.A(_0094_),
    .B(_0095_),
    .C(_0096_),
    .D(_1173_),
    .E(_0060_),
    .Y(_0927_));
 INVx2_ASAP7_75t_R _1199_ (.A(_0927_),
    .Y(_0928_));
 INVx1_ASAP7_75t_R _1200_ (.A(net104),
    .Y(_0929_));
 NOR3x1_ASAP7_75t_R _1201_ (.A(net107),
    .B(net106),
    .C(net105),
    .Y(_0930_));
 AND3x1_ASAP7_75t_R _1202_ (.A(net153),
    .B(_0929_),
    .C(_0930_),
    .Y(_0931_));
 AND2x4_ASAP7_75t_R _1203_ (.A(_0928_),
    .B(_0931_),
    .Y(_0932_));
 OR4x1_ASAP7_75t_R _1204_ (.A(_0922_),
    .B(_0925_),
    .C(_0926_),
    .D(_0932_),
    .Y(_0933_));
 BUFx12f_ASAP7_75t_R _1205_ (.A(_0933_),
    .Y(_0934_));
 INVx1_ASAP7_75t_R _1206_ (.A(net233),
    .Y(_0935_));
 INVx1_ASAP7_75t_R _1207_ (.A(net144),
    .Y(_0936_));
 NOR3x1_ASAP7_75t_R _1208_ (.A(net148),
    .B(net147),
    .C(net146),
    .Y(_0937_));
 AO33x2_ASAP7_75t_R _1209_ (.A1(_0936_),
    .A2(net154),
    .A3(_0937_),
    .B1(_0930_),
    .B2(net153),
    .B3(_0929_),
    .Y(_0938_));
 BUFx6f_ASAP7_75t_R _1210_ (.A(_0056_),
    .Y(_0939_));
 OA21x2_ASAP7_75t_R _1211_ (.A1(_0918_),
    .A2(_0938_),
    .B(_0939_),
    .Y(_0940_));
 AND3x4_ASAP7_75t_R _1212_ (.A(_0919_),
    .B(net232),
    .C(_0928_),
    .Y(_0941_));
 OR5x2_ASAP7_75t_R _1213_ (.A(_0935_),
    .B(net223),
    .C(_0926_),
    .D(_0940_),
    .E(_0941_),
    .Y(_0942_));
 OAI21x1_ASAP7_75t_R _1214_ (.A1(_0921_),
    .A2(_0938_),
    .B(_0057_),
    .Y(_0943_));
 NAND2x1_ASAP7_75t_R _1215_ (.A(_0916_),
    .B(net310),
    .Y(_0944_));
 INVx1_ASAP7_75t_R _1216_ (.A(_0926_),
    .Y(_0945_));
 AND2x2_ASAP7_75t_R _1217_ (.A(net311),
    .B(_0917_),
    .Y(_0946_));
 OA211x2_ASAP7_75t_R _1218_ (.A1(_0944_),
    .A2(_0927_),
    .B(_0945_),
    .C(_0946_),
    .Y(_0947_));
 NAND2x2_ASAP7_75t_R _1219_ (.A(_0943_),
    .B(_0947_),
    .Y(_0948_));
 NAND3x2_ASAP7_75t_R _1220_ (.B(_0942_),
    .C(_0948_),
    .Y(net354),
    .A(_0934_));
 INVx2_ASAP7_75t_R _1221_ (.A(net354),
    .Y(_1172_));
 NAND2x1_ASAP7_75t_R _1222_ (.A(_0928_),
    .B(_0943_),
    .Y(_0949_));
 OAI21x1_ASAP7_75t_R _1223_ (.A1(_0918_),
    .A2(_0921_),
    .B(_0099_),
    .Y(_0950_));
 OAI21x1_ASAP7_75t_R _1224_ (.A1(_0918_),
    .A2(_0938_),
    .B(_0939_),
    .Y(_0951_));
 AOI22x1_ASAP7_75t_R _1225_ (.A1(_0950_),
    .A2(_0932_),
    .B1(_0951_),
    .B2(_0941_),
    .Y(_0952_));
 OAI21x1_ASAP7_75t_R _1226_ (.A1(_0944_),
    .A2(_0949_),
    .B(_0952_),
    .Y(net353));
 INVx1_ASAP7_75t_R _1227_ (.A(net353),
    .Y(_1174_));
 INVx1_ASAP7_75t_R _1228_ (.A(_1175_),
    .Y(\credit_pi_route_inst.r_counters_inst.o_credits[6] ));
 INVx1_ASAP7_75t_R _1229_ (.A(_0086_),
    .Y(\credit_pi_route_inst.r_counters_inst.o_credits[8] ));
 INVx1_ASAP7_75t_R _1230_ (.A(_0087_),
    .Y(\credit_pi_route_inst.r_counters_inst.o_credits[7] ));
 INVx1_ASAP7_75t_R _1231_ (.A(_1177_),
    .Y(\credit_pi_route_inst.r_counters_inst.o_credits[1] ));
 INVx1_ASAP7_75t_R _1232_ (.A(_0089_),
    .Y(\credit_pi_route_inst.r_counters_inst.o_credits[3] ));
 INVx1_ASAP7_75t_R _1233_ (.A(_0090_),
    .Y(\credit_pi_route_inst.r_counters_inst.o_credits[2] ));
 AO22x1_ASAP7_75t_R _1234_ (.A1(net261),
    .A2(net310),
    .B1(net311),
    .B2(net301),
    .Y(_0953_));
 AO22x1_ASAP7_75t_R _1235_ (.A1(net183),
    .A2(net232),
    .B1(net233),
    .B2(net223),
    .Y(_0954_));
 OA21x2_ASAP7_75t_R _1236_ (.A1(_0953_),
    .A2(_0954_),
    .B(_0098_),
    .Y(_0955_));
 OR3x1_ASAP7_75t_R _1237_ (.A(net70),
    .B(net69),
    .C(net68),
    .Y(_0956_));
 NAND2x1_ASAP7_75t_R _1238_ (.A(net76),
    .B(net66),
    .Y(_0957_));
 AND5x2_ASAP7_75t_R _1239_ (.A(_0086_),
    .B(_0087_),
    .C(_1175_),
    .D(_0066_),
    .E(_0097_),
    .Y(_0958_));
 OR3x1_ASAP7_75t_R _1240_ (.A(_0956_),
    .B(_0957_),
    .C(_0958_),
    .Y(_0959_));
 AND5x2_ASAP7_75t_R _1241_ (.A(_0088_),
    .B(_0089_),
    .C(_0090_),
    .D(_1177_),
    .E(_0064_),
    .Y(_0960_));
 OR3x2_ASAP7_75t_R _1242_ (.A(net29),
    .B(net28),
    .C(net27),
    .Y(_0961_));
 NAND2x1_ASAP7_75t_R _1243_ (.A(net75),
    .B(net26),
    .Y(_0962_));
 NOR3x1_ASAP7_75t_R _1244_ (.A(_0960_),
    .B(_0961_),
    .C(_0962_),
    .Y(_0963_));
 OR3x2_ASAP7_75t_R _1245_ (.A(_0955_),
    .B(_0959_),
    .C(_0963_),
    .Y(_0964_));
 BUFx12f_ASAP7_75t_R _1246_ (.A(_0964_),
    .Y(_0965_));
 AND4x1_ASAP7_75t_R _1247_ (.A(_0089_),
    .B(_0090_),
    .C(_1177_),
    .D(_0064_),
    .Y(_0966_));
 NAND2x1_ASAP7_75t_R _1248_ (.A(_0088_),
    .B(_0966_),
    .Y(_0967_));
 AND3x4_ASAP7_75t_R _1249_ (.A(net183),
    .B(net232),
    .C(_0967_),
    .Y(_0968_));
 NOR3x1_ASAP7_75t_R _1250_ (.A(net70),
    .B(net69),
    .C(net68),
    .Y(_0969_));
 AND2x2_ASAP7_75t_R _1251_ (.A(net76),
    .B(net66),
    .Y(_0970_));
 NOR3x1_ASAP7_75t_R _1252_ (.A(net29),
    .B(net28),
    .C(net27),
    .Y(_0971_));
 AND2x2_ASAP7_75t_R _1253_ (.A(net75),
    .B(net26),
    .Y(_0972_));
 AO221x1_ASAP7_75t_R _1254_ (.A1(_0969_),
    .A2(_0970_),
    .B1(_0971_),
    .B2(_0972_),
    .C(_0953_),
    .Y(_0973_));
 OR3x1_ASAP7_75t_R _1255_ (.A(_0935_),
    .B(_0920_),
    .C(_0958_),
    .Y(_0974_));
 AO21x1_ASAP7_75t_R _1256_ (.A1(_0939_),
    .A2(_0973_),
    .B(_0974_),
    .Y(_0975_));
 BUFx6f_ASAP7_75t_R _1257_ (.A(_0975_),
    .Y(_0976_));
 AND2x4_ASAP7_75t_R _1258_ (.A(net261),
    .B(net310),
    .Y(_0977_));
 AO221x1_ASAP7_75t_R _1259_ (.A1(_0969_),
    .A2(_0970_),
    .B1(_0971_),
    .B2(_0972_),
    .C(_0954_),
    .Y(_0978_));
 INVx1_ASAP7_75t_R _1260_ (.A(net311),
    .Y(_0979_));
 OR3x1_ASAP7_75t_R _1261_ (.A(_0979_),
    .B(_0917_),
    .C(_0958_),
    .Y(_0980_));
 AO221x1_ASAP7_75t_R _1262_ (.A1(_0977_),
    .A2(_0967_),
    .B1(_0978_),
    .B2(_0057_),
    .C(_0980_),
    .Y(_0981_));
 OA21x2_ASAP7_75t_R _1263_ (.A1(_0968_),
    .A2(_0976_),
    .B(_0981_),
    .Y(_0982_));
 NAND2x2_ASAP7_75t_R _1264_ (.A(_0965_),
    .B(_0982_),
    .Y(net395));
 INVx2_ASAP7_75t_R _1265_ (.A(net395),
    .Y(_1176_));
 INVx1_ASAP7_75t_R _1266_ (.A(_0955_),
    .Y(_0983_));
 NAND2x2_ASAP7_75t_R _1267_ (.A(_0939_),
    .B(_0973_),
    .Y(_0984_));
 AOI21x1_ASAP7_75t_R _1268_ (.A1(_0057_),
    .A2(_0978_),
    .B(_0960_),
    .Y(_0985_));
 AO222x2_ASAP7_75t_R _1269_ (.A1(_0983_),
    .A2(_0963_),
    .B1(_0984_),
    .B2(_0968_),
    .C1(_0985_),
    .C2(_0977_),
    .Y(_0986_));
 BUFx6f_ASAP7_75t_R _1270_ (.A(_0986_),
    .Y(net394));
 INVx1_ASAP7_75t_R _1271_ (.A(net394),
    .Y(_1178_));
 INVx2_ASAP7_75t_R _1272_ (.A(_0083_),
    .Y(\credit_pi_route_inst.u0_counters_inst.o_credits[6] ));
 INVx1_ASAP7_75t_R _1273_ (.A(_0070_),
    .Y(\credit_pi_route_inst.u0_counters_inst.o_credits[5] ));
 INVx1_ASAP7_75t_R _1274_ (.A(_0081_),
    .Y(\credit_pi_route_inst.u0_counters_inst.o_credits[8] ));
 INVx1_ASAP7_75t_R _1275_ (.A(_0082_),
    .Y(\credit_pi_route_inst.u0_counters_inst.o_credits[7] ));
 INVx1_ASAP7_75t_R _1276_ (.A(_1180_),
    .Y(\credit_pi_route_inst.u0_counters_inst.o_credits[1] ));
 INVx1_ASAP7_75t_R _1277_ (.A(_0084_),
    .Y(\credit_pi_route_inst.u0_counters_inst.o_credits[3] ));
 INVx1_ASAP7_75t_R _1278_ (.A(_0085_),
    .Y(\credit_pi_route_inst.u0_counters_inst.o_credits[2] ));
 INVx1_ASAP7_75t_R _1279_ (.A(net75),
    .Y(_0987_));
 AND5x2_ASAP7_75t_R _1280_ (.A(_0058_),
    .B(_0084_),
    .C(_0085_),
    .D(_1180_),
    .E(_0068_),
    .Y(_0988_));
 OR3x2_ASAP7_75t_R _1281_ (.A(_0987_),
    .B(_0971_),
    .C(_0988_),
    .Y(_0989_));
 INVx4_ASAP7_75t_R _1282_ (.A(_0989_),
    .Y(_0990_));
 BUFx12f_ASAP7_75t_R _1283_ (.A(_0990_),
    .Y(net435));
 INVx2_ASAP7_75t_R _1284_ (.A(_0077_),
    .Y(\credit_pi_route_inst.u1_counters_inst.o_credits[6] ));
 INVx1_ASAP7_75t_R _1285_ (.A(_0073_),
    .Y(\credit_pi_route_inst.u1_counters_inst.o_credits[5] ));
 INVx1_ASAP7_75t_R _1286_ (.A(_0075_),
    .Y(\credit_pi_route_inst.u1_counters_inst.o_credits[8] ));
 INVx1_ASAP7_75t_R _1287_ (.A(_0076_),
    .Y(\credit_pi_route_inst.u1_counters_inst.o_credits[7] ));
 INVx1_ASAP7_75t_R _1288_ (.A(_1170_),
    .Y(\credit_pi_route_inst.u1_counters_inst.o_credits[1] ));
 INVx1_ASAP7_75t_R _1289_ (.A(_0078_),
    .Y(\credit_pi_route_inst.u1_counters_inst.o_credits[3] ));
 INVx1_ASAP7_75t_R _1290_ (.A(_0079_),
    .Y(\credit_pi_route_inst.u1_counters_inst.o_credits[2] ));
 INVx1_ASAP7_75t_R _1291_ (.A(net153),
    .Y(_0991_));
 AND5x1_ASAP7_75t_R _1292_ (.A(_0059_),
    .B(_0078_),
    .C(_0079_),
    .D(_1170_),
    .E(_0071_),
    .Y(_0992_));
 OR3x2_ASAP7_75t_R _1293_ (.A(_0991_),
    .B(_0930_),
    .C(_0992_),
    .Y(_1169_));
 INVx3_ASAP7_75t_R _1294_ (.A(_1169_),
    .Y(net476));
 AND2x2_ASAP7_75t_R _1295_ (.A(_0969_),
    .B(_0970_),
    .Y(_0993_));
 BUFx6f_ASAP7_75t_R _1296_ (.A(_0965_),
    .Y(_0994_));
 BUFx6f_ASAP7_75t_R _1297_ (.A(_0994_),
    .Y(_0995_));
 AND5x2_ASAP7_75t_R _1298_ (.A(_0080_),
    .B(_0081_),
    .C(_0082_),
    .D(_0083_),
    .E(_0070_),
    .Y(_0996_));
 OA211x2_ASAP7_75t_R _1299_ (.A1(_0990_),
    .A2(_0996_),
    .B(net76),
    .C(_0956_),
    .Y(_0997_));
 AO21x1_ASAP7_75t_R _1300_ (.A1(_0993_),
    .A2(_0995_),
    .B(_0997_),
    .Y(net315));
 AND2x2_ASAP7_75t_R _1301_ (.A(_0971_),
    .B(_0972_),
    .Y(_0998_));
 AO32x1_ASAP7_75t_R _1302_ (.A1(net75),
    .A2(_0961_),
    .A3(_0988_),
    .B1(_0998_),
    .B2(_0960_),
    .Y(_0999_));
 AO21x1_ASAP7_75t_R _1303_ (.A1(_0955_),
    .A2(_0998_),
    .B(_0999_),
    .Y(net314));
 BUFx6f_ASAP7_75t_R _1304_ (.A(_0934_),
    .Y(_1000_));
 AND2x2_ASAP7_75t_R _1305_ (.A(_0936_),
    .B(_0937_),
    .Y(_1001_));
 AND4x1_ASAP7_75t_R _1306_ (.A(_0075_),
    .B(_0076_),
    .C(_0077_),
    .D(_0073_),
    .Y(_1002_));
 AO21x2_ASAP7_75t_R _1307_ (.A1(_0074_),
    .A2(_1002_),
    .B(net476),
    .Y(_1003_));
 AO22x1_ASAP7_75t_R _1308_ (.A1(_1000_),
    .A2(_1001_),
    .B1(_1003_),
    .B2(_0924_),
    .Y(_1004_));
 AND2x2_ASAP7_75t_R _1309_ (.A(net154),
    .B(_1004_),
    .Y(net356));
 OR3x1_ASAP7_75t_R _1310_ (.A(net107),
    .B(net106),
    .C(net105),
    .Y(_1005_));
 AO32x1_ASAP7_75t_R _1311_ (.A1(net153),
    .A2(_1005_),
    .A3(_0992_),
    .B1(_0931_),
    .B2(_0927_),
    .Y(_1006_));
 AO21x1_ASAP7_75t_R _1312_ (.A1(_0922_),
    .A2(_0931_),
    .B(_1006_),
    .Y(net355));
 OA211x2_ASAP7_75t_R _1313_ (.A1(_0968_),
    .A2(_0976_),
    .B(net233),
    .C(_0942_),
    .Y(_1007_));
 BUFx3_ASAP7_75t_R _1314_ (.A(_1007_),
    .Y(net397));
 INVx1_ASAP7_75t_R _1315_ (.A(net232),
    .Y(_1008_));
 AO32x1_ASAP7_75t_R _1316_ (.A1(net183),
    .A2(_0967_),
    .A3(_0984_),
    .B1(_0951_),
    .B2(_0941_),
    .Y(_1009_));
 NOR2x1_ASAP7_75t_R _1317_ (.A(_1008_),
    .B(_1009_),
    .Y(net396));
 AND3x4_ASAP7_75t_R _1318_ (.A(net311),
    .B(_0948_),
    .C(_0981_),
    .Y(net438));
 INVx1_ASAP7_75t_R _1319_ (.A(_0977_),
    .Y(_1010_));
 AO21x1_ASAP7_75t_R _1320_ (.A1(_0928_),
    .A2(_0943_),
    .B(_0944_),
    .Y(_1011_));
 OAI21x1_ASAP7_75t_R _1321_ (.A1(_1010_),
    .A2(_0985_),
    .B(_1011_),
    .Y(net437));
 BUFx6f_ASAP7_75t_R _1322_ (.A(net157),
    .Y(_1012_));
 NOR2x1_ASAP7_75t_R _1323_ (.A(net438),
    .B(net437),
    .Y(_1013_));
 OR2x2_ASAP7_75t_R _1324_ (.A(_1012_),
    .B(_1013_),
    .Y(_1014_));
 OR2x6_ASAP7_75t_R _1325_ (.A(net397),
    .B(net396),
    .Y(_1015_));
 INVx1_ASAP7_75t_R _1326_ (.A(_0925_),
    .Y(_1016_));
 AND2x2_ASAP7_75t_R _1327_ (.A(net154),
    .B(_0924_),
    .Y(_1017_));
 AO221x1_ASAP7_75t_R _1328_ (.A1(_1016_),
    .A2(_0934_),
    .B1(_1003_),
    .B2(_1017_),
    .C(net355),
    .Y(_1018_));
 OA211x2_ASAP7_75t_R _1329_ (.A1(_0098_),
    .A2(_1018_),
    .B(_0099_),
    .C(_0939_),
    .Y(_1019_));
 AO21x1_ASAP7_75t_R _1330_ (.A1(_0939_),
    .A2(_1015_),
    .B(_1019_),
    .Y(_1020_));
 AO21x1_ASAP7_75t_R _1331_ (.A1(_0955_),
    .A2(_0998_),
    .B(_0993_),
    .Y(_1021_));
 AO211x2_ASAP7_75t_R _1332_ (.A1(_0965_),
    .A2(_1021_),
    .B(_0999_),
    .C(_0997_),
    .Y(_1022_));
 OR5x1_ASAP7_75t_R _1333_ (.A(_0057_),
    .B(_1012_),
    .C(_1018_),
    .D(_1022_),
    .E(_1015_),
    .Y(_1023_));
 OAI21x1_ASAP7_75t_R _1334_ (.A1(_1014_),
    .A2(_1020_),
    .B(_1023_),
    .Y(_0003_));
 OR4x1_ASAP7_75t_R _1335_ (.A(net157),
    .B(net438),
    .C(net437),
    .D(_1022_),
    .Y(_1024_));
 OR3x1_ASAP7_75t_R _1336_ (.A(_0099_),
    .B(net397),
    .C(net396),
    .Y(_1025_));
 OA21x2_ASAP7_75t_R _1337_ (.A1(_0057_),
    .A2(_1022_),
    .B(_0098_),
    .Y(_1026_));
 OA22x2_ASAP7_75t_R _1338_ (.A1(_0939_),
    .A2(_1024_),
    .B1(_1026_),
    .B2(_1012_),
    .Y(_1027_));
 INVx1_ASAP7_75t_R _1339_ (.A(_1018_),
    .Y(_1028_));
 OAI22x1_ASAP7_75t_R _1340_ (.A1(_1024_),
    .A2(_1025_),
    .B1(_1027_),
    .B2(_1028_),
    .Y(_0002_));
 INVx4_ASAP7_75t_R _1341_ (.A(net157),
    .Y(_1029_));
 OAI21x1_ASAP7_75t_R _1342_ (.A1(_1018_),
    .A2(_1026_),
    .B(_0099_),
    .Y(_1030_));
 NOR2x1_ASAP7_75t_R _1343_ (.A(_0939_),
    .B(_1024_),
    .Y(_1031_));
 AO32x1_ASAP7_75t_R _1344_ (.A1(_1029_),
    .A2(_1015_),
    .A3(_1030_),
    .B1(_1031_),
    .B2(_1028_),
    .Y(_0001_));
 INVx1_ASAP7_75t_R _1345_ (.A(_0057_),
    .Y(_1032_));
 INVx1_ASAP7_75t_R _1346_ (.A(_1022_),
    .Y(_1033_));
 OA22x2_ASAP7_75t_R _1347_ (.A1(_0098_),
    .A2(_1018_),
    .B1(_1033_),
    .B2(_0099_),
    .Y(_1034_));
 OAI22x1_ASAP7_75t_R _1348_ (.A1(_0939_),
    .A2(_1033_),
    .B1(_1015_),
    .B2(_1034_),
    .Y(_1035_));
 BUFx6f_ASAP7_75t_R _1349_ (.A(net157),
    .Y(_1036_));
 AO221x1_ASAP7_75t_R _1350_ (.A1(_1032_),
    .A2(_1022_),
    .B1(_1013_),
    .B2(_1035_),
    .C(_1036_),
    .Y(_0000_));
 BUFx6f_ASAP7_75t_R _1351_ (.A(_0989_),
    .Y(_1179_));
 NAND2x1_ASAP7_75t_R _1352_ (.A(net154),
    .B(_0924_),
    .Y(_1037_));
 OR2x6_ASAP7_75t_R _1353_ (.A(_1003_),
    .B(_1037_),
    .Y(_1038_));
 INVx3_ASAP7_75t_R _1354_ (.A(_1038_),
    .Y(_1039_));
 BUFx12f_ASAP7_75t_R _1355_ (.A(_1039_),
    .Y(net477));
 NAND2x1_ASAP7_75t_R _1356_ (.A(net76),
    .B(_0956_),
    .Y(_1040_));
 NOR2x1_ASAP7_75t_R _1357_ (.A(_1040_),
    .B(_0996_),
    .Y(_1041_));
 AND2x6_ASAP7_75t_R _1358_ (.A(_0989_),
    .B(_1041_),
    .Y(net436));
 BUFx12f_ASAP7_75t_R _1359_ (.A(_1029_),
    .Y(_1042_));
 XOR2x1_ASAP7_75t_R _1360_ (.A(net77),
    .Y(_1043_),
    .B(net353));
 XOR2x2_ASAP7_75t_R _1361_ (.A(_0060_),
    .B(_1043_),
    .Y(_1044_));
 NAND2x1_ASAP7_75t_R _1362_ (.A(_1042_),
    .B(_1044_),
    .Y(_0106_));
 NOR2x1_ASAP7_75t_R _1363_ (.A(_1173_),
    .B(_1043_),
    .Y(_1045_));
 AND2x2_ASAP7_75t_R _1364_ (.A(_0061_),
    .B(_1043_),
    .Y(_1046_));
 OR3x1_ASAP7_75t_R _1365_ (.A(_1036_),
    .B(_1045_),
    .C(_1046_),
    .Y(_0107_));
 NOR2x1_ASAP7_75t_R _1366_ (.A(_0096_),
    .B(_1043_),
    .Y(_1047_));
 XNOR2x2_ASAP7_75t_R _1367_ (.A(_0026_),
    .B(_0024_),
    .Y(_1048_));
 AND2x2_ASAP7_75t_R _1368_ (.A(_1043_),
    .B(_1048_),
    .Y(_1049_));
 OR3x1_ASAP7_75t_R _1369_ (.A(_1036_),
    .B(_1047_),
    .C(_1049_),
    .Y(_0108_));
 OR2x2_ASAP7_75t_R _1370_ (.A(\credit_pi_route_inst.l_counters_inst.o_credits[3] ),
    .B(_1043_),
    .Y(_1050_));
 OA21x2_ASAP7_75t_R _1371_ (.A1(_0023_),
    .A2(_0060_),
    .B(_0025_),
    .Y(_1051_));
 OA21x2_ASAP7_75t_R _1372_ (.A1(_0024_),
    .A2(_1051_),
    .B(_0028_),
    .Y(_1052_));
 XNOR2x2_ASAP7_75t_R _1373_ (.A(_0027_),
    .B(_1052_),
    .Y(_1053_));
 NAND2x1_ASAP7_75t_R _1374_ (.A(_1043_),
    .B(_1053_),
    .Y(_1054_));
 BUFx6f_ASAP7_75t_R _1375_ (.A(_1012_),
    .Y(_1055_));
 AO21x1_ASAP7_75t_R _1376_ (.A1(_1050_),
    .A2(_1054_),
    .B(_1055_),
    .Y(_0109_));
 INVx1_ASAP7_75t_R _1377_ (.A(_0026_),
    .Y(_1056_));
 OA21x2_ASAP7_75t_R _1378_ (.A1(_1056_),
    .A2(_0024_),
    .B(_0028_),
    .Y(_1057_));
 OAI21x1_ASAP7_75t_R _1379_ (.A1(_0027_),
    .A2(_1057_),
    .B(_0029_),
    .Y(_1058_));
 OA211x2_ASAP7_75t_R _1380_ (.A1(_0944_),
    .A2(_0949_),
    .B(_1058_),
    .C(_0952_),
    .Y(_1059_));
 NOR2x1_ASAP7_75t_R _1381_ (.A(net77),
    .B(_1058_),
    .Y(_1060_));
 AO22x1_ASAP7_75t_R _1382_ (.A1(net77),
    .A2(_1059_),
    .B1(_1060_),
    .B2(net353),
    .Y(_1061_));
 XNOR2x2_ASAP7_75t_R _1383_ (.A(_0094_),
    .B(_1061_),
    .Y(_1062_));
 OR2x2_ASAP7_75t_R _1384_ (.A(_1036_),
    .B(_1062_),
    .Y(_0110_));
 XNOR2x1_ASAP7_75t_R _1385_ (.B(_1172_),
    .Y(_1063_),
    .A(net78));
 XOR2x2_ASAP7_75t_R _1386_ (.A(_0062_),
    .B(_1063_),
    .Y(_1064_));
 NAND2x1_ASAP7_75t_R _1387_ (.A(_1042_),
    .B(_1064_),
    .Y(_0111_));
 NOR2x1_ASAP7_75t_R _1388_ (.A(_1171_),
    .B(_1063_),
    .Y(_1065_));
 AND2x2_ASAP7_75t_R _1389_ (.A(_0063_),
    .B(_1063_),
    .Y(_1066_));
 OR3x1_ASAP7_75t_R _1390_ (.A(_1036_),
    .B(_1065_),
    .C(_1066_),
    .Y(_0112_));
 NOR2x1_ASAP7_75t_R _1391_ (.A(_0093_),
    .B(_1063_),
    .Y(_1067_));
 XNOR2x2_ASAP7_75t_R _1392_ (.A(_0020_),
    .B(_0018_),
    .Y(_1068_));
 AND2x2_ASAP7_75t_R _1393_ (.A(_1063_),
    .B(_1068_),
    .Y(_1069_));
 OR3x1_ASAP7_75t_R _1394_ (.A(_1036_),
    .B(_1067_),
    .C(_1069_),
    .Y(_0113_));
 OR2x2_ASAP7_75t_R _1395_ (.A(\credit_pi_route_inst.l_counters_inst.o_credits[8] ),
    .B(_1063_),
    .Y(_1070_));
 OA21x2_ASAP7_75t_R _1396_ (.A1(_0017_),
    .A2(_0062_),
    .B(_0019_),
    .Y(_1071_));
 OA21x2_ASAP7_75t_R _1397_ (.A1(_0018_),
    .A2(_1071_),
    .B(_0022_),
    .Y(_1072_));
 XNOR2x2_ASAP7_75t_R _1398_ (.A(_0021_),
    .B(_1072_),
    .Y(_1073_));
 NAND2x1_ASAP7_75t_R _1399_ (.A(_1063_),
    .B(_1073_),
    .Y(_1074_));
 AO21x1_ASAP7_75t_R _1400_ (.A1(_1070_),
    .A2(_1074_),
    .B(_1055_),
    .Y(_0114_));
 INVx1_ASAP7_75t_R _1401_ (.A(_0020_),
    .Y(_1075_));
 OA21x2_ASAP7_75t_R _1402_ (.A1(_1075_),
    .A2(_0018_),
    .B(_0022_),
    .Y(_1076_));
 OAI21x1_ASAP7_75t_R _1403_ (.A1(_0021_),
    .A2(_1076_),
    .B(_0104_),
    .Y(_1077_));
 NOR2x1_ASAP7_75t_R _1404_ (.A(net78),
    .B(_1077_),
    .Y(_1078_));
 AND5x1_ASAP7_75t_R _1405_ (.A(net78),
    .B(_0934_),
    .C(_0942_),
    .D(_0948_),
    .E(_1077_),
    .Y(_1079_));
 AO21x1_ASAP7_75t_R _1406_ (.A1(net354),
    .A2(_1078_),
    .B(_1079_),
    .Y(_1080_));
 XOR2x2_ASAP7_75t_R _1407_ (.A(_0091_),
    .B(_1080_),
    .Y(_1081_));
 NAND2x1_ASAP7_75t_R _1408_ (.A(_1042_),
    .B(_1081_),
    .Y(_0115_));
 INVx1_ASAP7_75t_R _1409_ (.A(net155),
    .Y(_1082_));
 XNOR2x1_ASAP7_75t_R _1410_ (.B(net394),
    .Y(_1083_),
    .A(_1082_));
 XOR2x2_ASAP7_75t_R _1411_ (.A(_0064_),
    .B(_1083_),
    .Y(_1084_));
 NAND2x1_ASAP7_75t_R _1412_ (.A(_1042_),
    .B(_1084_),
    .Y(_0116_));
 NOR2x1_ASAP7_75t_R _1413_ (.A(_1177_),
    .B(_1083_),
    .Y(_1085_));
 AND2x2_ASAP7_75t_R _1414_ (.A(_0065_),
    .B(_1083_),
    .Y(_1086_));
 OR3x1_ASAP7_75t_R _1415_ (.A(_1012_),
    .B(_1085_),
    .C(_1086_),
    .Y(_0117_));
 NOR2x1_ASAP7_75t_R _1416_ (.A(_0090_),
    .B(_1083_),
    .Y(_1087_));
 XNOR2x2_ASAP7_75t_R _1417_ (.A(_0039_),
    .B(_0037_),
    .Y(_1088_));
 AND2x2_ASAP7_75t_R _1418_ (.A(_1083_),
    .B(_1088_),
    .Y(_1089_));
 OR3x1_ASAP7_75t_R _1419_ (.A(_1012_),
    .B(_1087_),
    .C(_1089_),
    .Y(_0118_));
 OR2x2_ASAP7_75t_R _1420_ (.A(\credit_pi_route_inst.r_counters_inst.o_credits[3] ),
    .B(_1083_),
    .Y(_1090_));
 OA21x2_ASAP7_75t_R _1421_ (.A1(_0036_),
    .A2(_0064_),
    .B(_0038_),
    .Y(_1091_));
 OA21x2_ASAP7_75t_R _1422_ (.A1(_0037_),
    .A2(_1091_),
    .B(_0041_),
    .Y(_1092_));
 XNOR2x2_ASAP7_75t_R _1423_ (.A(_0040_),
    .B(_1092_),
    .Y(_1093_));
 NAND2x1_ASAP7_75t_R _1424_ (.A(_1083_),
    .B(_1093_),
    .Y(_1094_));
 AO21x1_ASAP7_75t_R _1425_ (.A1(_1090_),
    .A2(_1094_),
    .B(_1055_),
    .Y(_0119_));
 INVx1_ASAP7_75t_R _1426_ (.A(_0039_),
    .Y(_1095_));
 OA21x2_ASAP7_75t_R _1427_ (.A1(_1095_),
    .A2(_0037_),
    .B(_0041_),
    .Y(_1096_));
 OA21x2_ASAP7_75t_R _1428_ (.A1(_0040_),
    .A2(_1096_),
    .B(_0042_),
    .Y(_1097_));
 NOR2x1_ASAP7_75t_R _1429_ (.A(net394),
    .B(_1097_),
    .Y(_1098_));
 AND3x1_ASAP7_75t_R _1430_ (.A(_1082_),
    .B(net394),
    .C(_1097_),
    .Y(_1099_));
 AO21x1_ASAP7_75t_R _1431_ (.A1(net155),
    .A2(_1098_),
    .B(_1099_),
    .Y(_1100_));
 XOR2x2_ASAP7_75t_R _1432_ (.A(_0088_),
    .B(_1100_),
    .Y(_1101_));
 NAND2x1_ASAP7_75t_R _1433_ (.A(_1042_),
    .B(_1101_),
    .Y(_0120_));
 XNOR2x1_ASAP7_75t_R _1434_ (.B(_1176_),
    .Y(_1102_),
    .A(net156));
 XOR2x2_ASAP7_75t_R _1435_ (.A(_0066_),
    .B(_1102_),
    .Y(_1103_));
 NAND2x1_ASAP7_75t_R _1436_ (.A(_1042_),
    .B(_1103_),
    .Y(_0121_));
 NOR2x1_ASAP7_75t_R _1437_ (.A(_1175_),
    .B(_1102_),
    .Y(_1104_));
 AND2x2_ASAP7_75t_R _1438_ (.A(_0067_),
    .B(_1102_),
    .Y(_1105_));
 OR3x1_ASAP7_75t_R _1439_ (.A(_1012_),
    .B(_1104_),
    .C(_1105_),
    .Y(_0122_));
 NOR2x1_ASAP7_75t_R _1440_ (.A(_0087_),
    .B(_1102_),
    .Y(_1106_));
 XNOR2x2_ASAP7_75t_R _1441_ (.A(_0033_),
    .B(_0031_),
    .Y(_1107_));
 AND2x2_ASAP7_75t_R _1442_ (.A(_1102_),
    .B(_1107_),
    .Y(_1108_));
 OR3x1_ASAP7_75t_R _1443_ (.A(_1012_),
    .B(_1106_),
    .C(_1108_),
    .Y(_0123_));
 OR2x2_ASAP7_75t_R _1444_ (.A(\credit_pi_route_inst.r_counters_inst.o_credits[8] ),
    .B(_1102_),
    .Y(_1109_));
 OA21x2_ASAP7_75t_R _1445_ (.A1(_0030_),
    .A2(_0066_),
    .B(_0032_),
    .Y(_1110_));
 OA21x2_ASAP7_75t_R _1446_ (.A1(_0031_),
    .A2(_1110_),
    .B(_0035_),
    .Y(_1111_));
 XNOR2x2_ASAP7_75t_R _1447_ (.A(_0034_),
    .B(_1111_),
    .Y(_1112_));
 NAND2x1_ASAP7_75t_R _1448_ (.A(_1102_),
    .B(_1112_),
    .Y(_1113_));
 AO21x1_ASAP7_75t_R _1449_ (.A1(_1109_),
    .A2(_1113_),
    .B(_1055_),
    .Y(_0124_));
 INVx1_ASAP7_75t_R _1450_ (.A(_0033_),
    .Y(_1114_));
 OA21x2_ASAP7_75t_R _1451_ (.A1(_1114_),
    .A2(_0031_),
    .B(_0035_),
    .Y(_1115_));
 OAI21x1_ASAP7_75t_R _1452_ (.A1(_0034_),
    .A2(_1115_),
    .B(_0105_),
    .Y(_1116_));
 NOR2x1_ASAP7_75t_R _1453_ (.A(net156),
    .B(_1116_),
    .Y(_1117_));
 AND3x1_ASAP7_75t_R _1454_ (.A(net156),
    .B(_1176_),
    .C(_1116_),
    .Y(_1118_));
 AO21x1_ASAP7_75t_R _1455_ (.A1(net395),
    .A2(_1117_),
    .B(_1118_),
    .Y(_1119_));
 XOR2x2_ASAP7_75t_R _1456_ (.A(_0097_),
    .B(_1119_),
    .Y(_1120_));
 NAND2x1_ASAP7_75t_R _1457_ (.A(_1042_),
    .B(_1120_),
    .Y(_0125_));
 XNOR2x1_ASAP7_75t_R _1458_ (.B(_0990_),
    .Y(_1121_),
    .A(net234));
 XNOR2x2_ASAP7_75t_R _1459_ (.A(_0068_),
    .B(_1121_),
    .Y(_1122_));
 NAND2x1_ASAP7_75t_R _1460_ (.A(_1042_),
    .B(_1122_),
    .Y(_0126_));
 NAND2x1_ASAP7_75t_R _1461_ (.A(_1180_),
    .B(_1121_),
    .Y(_1123_));
 OR2x2_ASAP7_75t_R _1462_ (.A(_0069_),
    .B(_1121_),
    .Y(_1124_));
 AO21x1_ASAP7_75t_R _1463_ (.A1(_1123_),
    .A2(_1124_),
    .B(_1055_),
    .Y(_0127_));
 AND2x2_ASAP7_75t_R _1464_ (.A(\credit_pi_route_inst.u0_counters_inst.o_credits[2] ),
    .B(_1121_),
    .Y(_1125_));
 XOR2x2_ASAP7_75t_R _1465_ (.A(_0051_),
    .B(_0103_),
    .Y(_1126_));
 NOR2x1_ASAP7_75t_R _1466_ (.A(_1121_),
    .B(_1126_),
    .Y(_1127_));
 OR3x1_ASAP7_75t_R _1467_ (.A(_1012_),
    .B(_1125_),
    .C(_1127_),
    .Y(_0128_));
 NAND2x1_ASAP7_75t_R _1468_ (.A(_0084_),
    .B(_1121_),
    .Y(_1128_));
 OA21x2_ASAP7_75t_R _1469_ (.A1(_0050_),
    .A2(_0068_),
    .B(_0052_),
    .Y(_1129_));
 OA21x2_ASAP7_75t_R _1470_ (.A1(_0051_),
    .A2(_1129_),
    .B(_0054_),
    .Y(_1130_));
 XOR2x2_ASAP7_75t_R _1471_ (.A(_0053_),
    .B(_1130_),
    .Y(_1131_));
 OR2x2_ASAP7_75t_R _1472_ (.A(_1121_),
    .B(_1131_),
    .Y(_1132_));
 AO21x1_ASAP7_75t_R _1473_ (.A1(_1128_),
    .A2(_1132_),
    .B(_1055_),
    .Y(_0129_));
 INVx1_ASAP7_75t_R _1474_ (.A(_0103_),
    .Y(_1133_));
 OA21x2_ASAP7_75t_R _1475_ (.A1(_0051_),
    .A2(_1133_),
    .B(_0054_),
    .Y(_1134_));
 OAI21x1_ASAP7_75t_R _1476_ (.A1(_0053_),
    .A2(_1134_),
    .B(_0055_),
    .Y(_1135_));
 NOR2x1_ASAP7_75t_R _1477_ (.A(net234),
    .B(_1135_),
    .Y(_1136_));
 AND3x1_ASAP7_75t_R _1478_ (.A(net234),
    .B(_0989_),
    .C(_1135_),
    .Y(_1137_));
 AO21x1_ASAP7_75t_R _1479_ (.A1(_0990_),
    .A2(_1136_),
    .B(_1137_),
    .Y(_1138_));
 XOR2x2_ASAP7_75t_R _1480_ (.A(_0058_),
    .B(_1138_),
    .Y(_1139_));
 NAND2x1_ASAP7_75t_R _1481_ (.A(_1042_),
    .B(_1139_),
    .Y(_0130_));
 XNOR2x1_ASAP7_75t_R _1482_ (.B(net436),
    .Y(_1140_),
    .A(net235));
 XNOR2x2_ASAP7_75t_R _1483_ (.A(_0070_),
    .B(_1140_),
    .Y(_1141_));
 NAND2x1_ASAP7_75t_R _1484_ (.A(_1042_),
    .B(_1141_),
    .Y(_0131_));
 NAND2x1_ASAP7_75t_R _1485_ (.A(_0083_),
    .B(_1140_),
    .Y(_1142_));
 INVx1_ASAP7_75t_R _1486_ (.A(_0102_),
    .Y(_1143_));
 OR2x2_ASAP7_75t_R _1487_ (.A(_1143_),
    .B(_1140_),
    .Y(_1144_));
 AO21x1_ASAP7_75t_R _1488_ (.A1(_1142_),
    .A2(_1144_),
    .B(_1055_),
    .Y(_0132_));
 NAND2x1_ASAP7_75t_R _1489_ (.A(_0082_),
    .B(_1140_),
    .Y(_1145_));
 XOR2x2_ASAP7_75t_R _1490_ (.A(_0046_),
    .B(_0044_),
    .Y(_1146_));
 OR2x2_ASAP7_75t_R _1491_ (.A(_1140_),
    .B(_1146_),
    .Y(_1147_));
 AO21x1_ASAP7_75t_R _1492_ (.A1(_1145_),
    .A2(_1147_),
    .B(_1055_),
    .Y(_0133_));
 NAND2x1_ASAP7_75t_R _1493_ (.A(_0081_),
    .B(_1140_),
    .Y(_1148_));
 OA21x2_ASAP7_75t_R _1494_ (.A1(_0043_),
    .A2(_0070_),
    .B(_0045_),
    .Y(_1149_));
 OA21x2_ASAP7_75t_R _1495_ (.A1(_0044_),
    .A2(_1149_),
    .B(_0048_),
    .Y(_1150_));
 XOR2x2_ASAP7_75t_R _1496_ (.A(_0047_),
    .B(_1150_),
    .Y(_1151_));
 OR2x2_ASAP7_75t_R _1497_ (.A(_1140_),
    .B(_1151_),
    .Y(_1152_));
 AO21x1_ASAP7_75t_R _1498_ (.A1(_1148_),
    .A2(_1152_),
    .B(_1055_),
    .Y(_0134_));
 OR2x2_ASAP7_75t_R _1499_ (.A(_1040_),
    .B(_0996_),
    .Y(_1153_));
 OR3x1_ASAP7_75t_R _1500_ (.A(net235),
    .B(_0990_),
    .C(_1153_),
    .Y(_1154_));
 OA21x2_ASAP7_75t_R _1501_ (.A1(_0046_),
    .A2(_0044_),
    .B(_0048_),
    .Y(_1155_));
 OAI21x1_ASAP7_75t_R _1502_ (.A1(_0047_),
    .A2(_1155_),
    .B(_0049_),
    .Y(_1156_));
 NAND2x1_ASAP7_75t_R _1503_ (.A(net235),
    .B(_1156_),
    .Y(_1157_));
 OAI22x1_ASAP7_75t_R _1504_ (.A1(_1154_),
    .A2(_1156_),
    .B1(_1157_),
    .B2(net436),
    .Y(_1158_));
 XOR2x2_ASAP7_75t_R _1505_ (.A(_0080_),
    .B(_1158_),
    .Y(_1159_));
 NAND2x1_ASAP7_75t_R _1506_ (.A(_1029_),
    .B(_1159_),
    .Y(_0135_));
 XNOR2x1_ASAP7_75t_R _1507_ (.B(net476),
    .Y(_1160_),
    .A(net312));
 XNOR2x2_ASAP7_75t_R _1508_ (.A(_0071_),
    .B(_1160_),
    .Y(_1161_));
 NAND2x1_ASAP7_75t_R _1509_ (.A(_1029_),
    .B(_1161_),
    .Y(_0136_));
 NAND2x1_ASAP7_75t_R _1510_ (.A(_1170_),
    .B(_1160_),
    .Y(_1162_));
 OR2x2_ASAP7_75t_R _1511_ (.A(_0072_),
    .B(_1160_),
    .Y(_1163_));
 AO21x1_ASAP7_75t_R _1512_ (.A1(_1162_),
    .A2(_1163_),
    .B(_1055_),
    .Y(_0137_));
 AND2x2_ASAP7_75t_R _1513_ (.A(\credit_pi_route_inst.u1_counters_inst.o_credits[2] ),
    .B(_1160_),
    .Y(_1164_));
 XOR2x2_ASAP7_75t_R _1514_ (.A(_0005_),
    .B(_0100_),
    .Y(_1165_));
 NOR2x1_ASAP7_75t_R _1515_ (.A(_1160_),
    .B(_1165_),
    .Y(_1166_));
 OR3x1_ASAP7_75t_R _1516_ (.A(_1012_),
    .B(_1164_),
    .C(_1166_),
    .Y(_0138_));
 NAND2x1_ASAP7_75t_R _1517_ (.A(_0078_),
    .B(_1160_),
    .Y(_1167_));
 OA21x2_ASAP7_75t_R _1518_ (.A1(_0004_),
    .A2(_0071_),
    .B(_0006_),
    .Y(_1168_));
 OA21x2_ASAP7_75t_R _1519_ (.A1(_0005_),
    .A2(_1168_),
    .B(_0008_),
    .Y(_0146_));
 XOR2x2_ASAP7_75t_R _1520_ (.A(_0007_),
    .B(_0146_),
    .Y(_0147_));
 OR2x2_ASAP7_75t_R _1521_ (.A(_1160_),
    .B(_0147_),
    .Y(_0148_));
 AO21x1_ASAP7_75t_R _1522_ (.A1(_1167_),
    .A2(_0148_),
    .B(_1036_),
    .Y(_0139_));
 INVx1_ASAP7_75t_R _1523_ (.A(_0100_),
    .Y(_0149_));
 OA21x2_ASAP7_75t_R _1524_ (.A1(_0005_),
    .A2(_0149_),
    .B(_0008_),
    .Y(_0150_));
 OAI21x1_ASAP7_75t_R _1525_ (.A1(_0007_),
    .A2(_0150_),
    .B(_0009_),
    .Y(_0151_));
 NOR2x1_ASAP7_75t_R _1526_ (.A(net312),
    .B(_0151_),
    .Y(_0152_));
 AND3x1_ASAP7_75t_R _1527_ (.A(net312),
    .B(_1169_),
    .C(_0151_),
    .Y(_0153_));
 AO21x1_ASAP7_75t_R _1528_ (.A1(net476),
    .A2(_0152_),
    .B(_0153_),
    .Y(_0154_));
 XOR2x2_ASAP7_75t_R _1529_ (.A(_0059_),
    .B(_0154_),
    .Y(_0155_));
 NAND2x1_ASAP7_75t_R _1530_ (.A(_1029_),
    .B(_0155_),
    .Y(_0140_));
 XNOR2x1_ASAP7_75t_R _1531_ (.B(_1039_),
    .Y(_0156_),
    .A(net313));
 XNOR2x2_ASAP7_75t_R _1532_ (.A(_0073_),
    .B(_0156_),
    .Y(_0157_));
 NAND2x1_ASAP7_75t_R _1533_ (.A(_1029_),
    .B(_0157_),
    .Y(_0141_));
 NAND2x1_ASAP7_75t_R _1534_ (.A(_0077_),
    .B(_0156_),
    .Y(_0158_));
 INVx1_ASAP7_75t_R _1535_ (.A(_0101_),
    .Y(_0159_));
 OR2x2_ASAP7_75t_R _1536_ (.A(_0159_),
    .B(_0156_),
    .Y(_0160_));
 AO21x1_ASAP7_75t_R _1537_ (.A1(_0158_),
    .A2(_0160_),
    .B(_1036_),
    .Y(_0142_));
 NAND2x1_ASAP7_75t_R _1538_ (.A(_0076_),
    .B(_0156_),
    .Y(_0161_));
 XOR2x2_ASAP7_75t_R _1539_ (.A(_0013_),
    .B(_0011_),
    .Y(_0162_));
 OR2x2_ASAP7_75t_R _1540_ (.A(_0156_),
    .B(_0162_),
    .Y(_0163_));
 AO21x1_ASAP7_75t_R _1541_ (.A1(_0161_),
    .A2(_0163_),
    .B(_1036_),
    .Y(_0143_));
 NAND2x1_ASAP7_75t_R _1542_ (.A(_0075_),
    .B(_0156_),
    .Y(_0164_));
 OA21x2_ASAP7_75t_R _1543_ (.A1(_0010_),
    .A2(_0073_),
    .B(_0012_),
    .Y(_0165_));
 OA21x2_ASAP7_75t_R _1544_ (.A1(_0011_),
    .A2(_0165_),
    .B(_0015_),
    .Y(_0166_));
 XOR2x2_ASAP7_75t_R _1545_ (.A(_0014_),
    .B(_0166_),
    .Y(_0167_));
 OR2x2_ASAP7_75t_R _1546_ (.A(_0156_),
    .B(_0167_),
    .Y(_0168_));
 AO21x1_ASAP7_75t_R _1547_ (.A1(_0164_),
    .A2(_0168_),
    .B(_1036_),
    .Y(_0144_));
 OA21x2_ASAP7_75t_R _1548_ (.A1(_0013_),
    .A2(_0011_),
    .B(_0015_),
    .Y(_0169_));
 OAI21x1_ASAP7_75t_R _1549_ (.A1(_0014_),
    .A2(_0169_),
    .B(_0016_),
    .Y(_0170_));
 NOR2x1_ASAP7_75t_R _1550_ (.A(net313),
    .B(_0170_),
    .Y(_0171_));
 AND3x1_ASAP7_75t_R _1551_ (.A(net313),
    .B(_1038_),
    .C(_0170_),
    .Y(_0172_));
 AO21x1_ASAP7_75t_R _1552_ (.A1(_1039_),
    .A2(_0171_),
    .B(_0172_),
    .Y(_0173_));
 XOR2x2_ASAP7_75t_R _1553_ (.A(_0074_),
    .B(_0173_),
    .Y(_0174_));
 NAND2x1_ASAP7_75t_R _1554_ (.A(_1029_),
    .B(_0174_),
    .Y(_0145_));
 AND3x1_ASAP7_75t_R _1555_ (.A(net233),
    .B(_0920_),
    .C(_0945_),
    .Y(_0175_));
 AO22x1_ASAP7_75t_R _1556_ (.A1(_0951_),
    .A2(_0175_),
    .B1(_0943_),
    .B2(_0947_),
    .Y(_0176_));
 BUFx6f_ASAP7_75t_R _1557_ (.A(_0176_),
    .Y(_0177_));
 OR3x1_ASAP7_75t_R _1558_ (.A(_0991_),
    .B(net104),
    .C(_1005_),
    .Y(_0178_));
 NOR2x1_ASAP7_75t_R _1559_ (.A(_0925_),
    .B(_0926_),
    .Y(_0179_));
 OA211x2_ASAP7_75t_R _1560_ (.A1(_0927_),
    .A2(_0178_),
    .B(_0950_),
    .C(_0179_),
    .Y(_0180_));
 AOI21x1_ASAP7_75t_R _1561_ (.A1(_0952_),
    .A2(_0177_),
    .B(_0180_),
    .Y(_0181_));
 BUFx6f_ASAP7_75t_R _1562_ (.A(_0181_),
    .Y(_0182_));
 AND2x2_ASAP7_75t_R _1563_ (.A(net158),
    .B(_0182_),
    .Y(_0183_));
 AO21x2_ASAP7_75t_R _1564_ (.A1(_0952_),
    .A2(_0177_),
    .B(_0180_),
    .Y(_0184_));
 BUFx6f_ASAP7_75t_R _1565_ (.A(_0184_),
    .Y(_0185_));
 AND2x2_ASAP7_75t_R _1566_ (.A(net188),
    .B(_0185_),
    .Y(_0186_));
 OAI21x1_ASAP7_75t_R _1567_ (.A1(_0179_),
    .A2(_0932_),
    .B(_0950_),
    .Y(_0187_));
 INVx2_ASAP7_75t_R _1568_ (.A(_0187_),
    .Y(_0188_));
 OAI21x1_ASAP7_75t_R _1569_ (.A1(_0941_),
    .A2(_0175_),
    .B(_0951_),
    .Y(_0189_));
 NOR2x1_ASAP7_75t_R _1570_ (.A(_0188_),
    .B(_0189_),
    .Y(_0190_));
 OA21x2_ASAP7_75t_R _1571_ (.A1(_0183_),
    .A2(_0186_),
    .B(_0190_),
    .Y(_0191_));
 AND2x2_ASAP7_75t_R _1572_ (.A(net79),
    .B(_0182_),
    .Y(_0192_));
 AND2x2_ASAP7_75t_R _1573_ (.A(net109),
    .B(_0185_),
    .Y(_0193_));
 OA21x2_ASAP7_75t_R _1574_ (.A1(_0192_),
    .A2(_0193_),
    .B(_0188_),
    .Y(_0194_));
 BUFx6f_ASAP7_75t_R _1575_ (.A(_0184_),
    .Y(_0195_));
 BUFx6f_ASAP7_75t_R _1576_ (.A(_0195_),
    .Y(_0196_));
 AND2x4_ASAP7_75t_R _1577_ (.A(_0187_),
    .B(_0189_),
    .Y(_0197_));
 AND3x1_ASAP7_75t_R _1578_ (.A(net266),
    .B(_0196_),
    .C(_0197_),
    .Y(_0198_));
 BUFx6f_ASAP7_75t_R _1579_ (.A(_0181_),
    .Y(_0199_));
 BUFx6f_ASAP7_75t_R _1580_ (.A(_0199_),
    .Y(_0200_));
 AND3x1_ASAP7_75t_R _1581_ (.A(net236),
    .B(_0200_),
    .C(_0197_),
    .Y(_0201_));
 OR4x1_ASAP7_75t_R _1582_ (.A(_0191_),
    .B(_0194_),
    .C(_0198_),
    .D(_0201_),
    .Y(net316));
 BUFx12f_ASAP7_75t_R _1583_ (.A(_0187_),
    .Y(_0202_));
 BUFx6f_ASAP7_75t_R _1584_ (.A(_0202_),
    .Y(_0203_));
 BUFx6f_ASAP7_75t_R _1585_ (.A(_0182_),
    .Y(_0204_));
 OR3x1_ASAP7_75t_R _1586_ (.A(net120),
    .B(_0203_),
    .C(_0204_),
    .Y(_0205_));
 BUFx6f_ASAP7_75t_R _1587_ (.A(_0202_),
    .Y(_0206_));
 BUFx6f_ASAP7_75t_R _1588_ (.A(_0185_),
    .Y(_0207_));
 OR3x1_ASAP7_75t_R _1589_ (.A(net80),
    .B(_0206_),
    .C(_0207_),
    .Y(_0208_));
 NAND2x2_ASAP7_75t_R _1590_ (.A(_0187_),
    .B(_0189_),
    .Y(_0209_));
 BUFx6f_ASAP7_75t_R _1591_ (.A(_0209_),
    .Y(_0210_));
 AND2x2_ASAP7_75t_R _1592_ (.A(net237),
    .B(_0182_),
    .Y(_0211_));
 AND2x2_ASAP7_75t_R _1593_ (.A(net277),
    .B(_0185_),
    .Y(_0212_));
 BUFx6f_ASAP7_75t_R _1594_ (.A(_0952_),
    .Y(_0213_));
 BUFx6f_ASAP7_75t_R _1595_ (.A(_0177_),
    .Y(_0214_));
 AND3x1_ASAP7_75t_R _1596_ (.A(net199),
    .B(_0213_),
    .C(_0214_),
    .Y(_0215_));
 NAND2x2_ASAP7_75t_R _1597_ (.A(_0952_),
    .B(_0177_),
    .Y(_0216_));
 BUFx6f_ASAP7_75t_R _1598_ (.A(_0216_),
    .Y(_0217_));
 AND3x1_ASAP7_75t_R _1599_ (.A(net159),
    .B(_1000_),
    .C(_0217_),
    .Y(_0218_));
 OR2x6_ASAP7_75t_R _1600_ (.A(_0188_),
    .B(_0189_),
    .Y(_0219_));
 BUFx6f_ASAP7_75t_R _1601_ (.A(_0219_),
    .Y(_0220_));
 OA33x2_ASAP7_75t_R _1602_ (.A1(_0210_),
    .A2(_0211_),
    .A3(_0212_),
    .B1(_0215_),
    .B2(_0218_),
    .B3(_0220_),
    .Y(_0221_));
 AND3x1_ASAP7_75t_R _1603_ (.A(_0205_),
    .B(_0208_),
    .C(_0221_),
    .Y(net317));
 OR3x1_ASAP7_75t_R _1604_ (.A(net121),
    .B(_0203_),
    .C(_0204_),
    .Y(_0222_));
 OR3x1_ASAP7_75t_R _1605_ (.A(net81),
    .B(_0206_),
    .C(_0207_),
    .Y(_0223_));
 AND2x2_ASAP7_75t_R _1606_ (.A(net238),
    .B(_0182_),
    .Y(_0224_));
 AND2x2_ASAP7_75t_R _1607_ (.A(net278),
    .B(_0185_),
    .Y(_0225_));
 AND3x1_ASAP7_75t_R _1608_ (.A(net200),
    .B(_0213_),
    .C(_0214_),
    .Y(_0226_));
 AND3x1_ASAP7_75t_R _1609_ (.A(net160),
    .B(_1000_),
    .C(_0217_),
    .Y(_0227_));
 OA33x2_ASAP7_75t_R _1610_ (.A1(_0210_),
    .A2(_0224_),
    .A3(_0225_),
    .B1(_0226_),
    .B2(_0227_),
    .B3(_0220_),
    .Y(_0228_));
 AND3x1_ASAP7_75t_R _1611_ (.A(_0222_),
    .B(_0223_),
    .C(_0228_),
    .Y(net318));
 OR3x1_ASAP7_75t_R _1612_ (.A(net122),
    .B(_0203_),
    .C(_0204_),
    .Y(_0229_));
 OR3x1_ASAP7_75t_R _1613_ (.A(net82),
    .B(_0206_),
    .C(_0207_),
    .Y(_0230_));
 AND2x2_ASAP7_75t_R _1614_ (.A(net239),
    .B(_0182_),
    .Y(_0231_));
 AND2x2_ASAP7_75t_R _1615_ (.A(net279),
    .B(_0185_),
    .Y(_0232_));
 AND3x1_ASAP7_75t_R _1616_ (.A(net201),
    .B(_0213_),
    .C(_0214_),
    .Y(_0233_));
 AND3x1_ASAP7_75t_R _1617_ (.A(net161),
    .B(_1000_),
    .C(_0217_),
    .Y(_0234_));
 OA33x2_ASAP7_75t_R _1618_ (.A1(_0210_),
    .A2(_0231_),
    .A3(_0232_),
    .B1(_0233_),
    .B2(_0234_),
    .B3(_0220_),
    .Y(_0235_));
 AND3x1_ASAP7_75t_R _1619_ (.A(_0229_),
    .B(_0230_),
    .C(_0235_),
    .Y(net319));
 OR3x1_ASAP7_75t_R _1620_ (.A(net124),
    .B(_0203_),
    .C(_0204_),
    .Y(_0236_));
 BUFx6f_ASAP7_75t_R _1621_ (.A(_0185_),
    .Y(_0237_));
 OR3x1_ASAP7_75t_R _1622_ (.A(net83),
    .B(_0206_),
    .C(_0237_),
    .Y(_0238_));
 AND2x2_ASAP7_75t_R _1623_ (.A(net240),
    .B(_0182_),
    .Y(_0239_));
 AND2x2_ASAP7_75t_R _1624_ (.A(net281),
    .B(_0185_),
    .Y(_0240_));
 AND3x1_ASAP7_75t_R _1625_ (.A(net203),
    .B(_0213_),
    .C(_0214_),
    .Y(_0241_));
 AND3x1_ASAP7_75t_R _1626_ (.A(net162),
    .B(_1000_),
    .C(_0217_),
    .Y(_0242_));
 OA33x2_ASAP7_75t_R _1627_ (.A1(_0210_),
    .A2(_0239_),
    .A3(_0240_),
    .B1(_0241_),
    .B2(_0242_),
    .B3(_0220_),
    .Y(_0243_));
 AND3x1_ASAP7_75t_R _1628_ (.A(_0236_),
    .B(_0238_),
    .C(_0243_),
    .Y(net320));
 OR3x1_ASAP7_75t_R _1629_ (.A(net125),
    .B(_0203_),
    .C(_0204_),
    .Y(_0244_));
 OR3x1_ASAP7_75t_R _1630_ (.A(net84),
    .B(_0206_),
    .C(_0237_),
    .Y(_0245_));
 AND2x2_ASAP7_75t_R _1631_ (.A(net241),
    .B(_0182_),
    .Y(_0246_));
 AND2x2_ASAP7_75t_R _1632_ (.A(net282),
    .B(_0185_),
    .Y(_0247_));
 AND3x1_ASAP7_75t_R _1633_ (.A(net204),
    .B(_0213_),
    .C(_0214_),
    .Y(_0248_));
 AND3x1_ASAP7_75t_R _1634_ (.A(net163),
    .B(_1000_),
    .C(_0217_),
    .Y(_0249_));
 OA33x2_ASAP7_75t_R _1635_ (.A1(_0210_),
    .A2(_0246_),
    .A3(_0247_),
    .B1(_0248_),
    .B2(_0249_),
    .B3(_0220_),
    .Y(_0250_));
 AND3x1_ASAP7_75t_R _1636_ (.A(_0244_),
    .B(_0245_),
    .C(_0250_),
    .Y(net321));
 OR3x1_ASAP7_75t_R _1637_ (.A(net126),
    .B(_0203_),
    .C(_0204_),
    .Y(_0251_));
 OR3x1_ASAP7_75t_R _1638_ (.A(net85),
    .B(_0206_),
    .C(_0237_),
    .Y(_0252_));
 BUFx6f_ASAP7_75t_R _1639_ (.A(_0199_),
    .Y(_0253_));
 AND2x2_ASAP7_75t_R _1640_ (.A(net242),
    .B(_0253_),
    .Y(_0254_));
 BUFx6f_ASAP7_75t_R _1641_ (.A(_0195_),
    .Y(_0255_));
 AND2x2_ASAP7_75t_R _1642_ (.A(net283),
    .B(_0255_),
    .Y(_0256_));
 AND3x1_ASAP7_75t_R _1643_ (.A(net205),
    .B(_0213_),
    .C(_0214_),
    .Y(_0257_));
 AND3x1_ASAP7_75t_R _1644_ (.A(net164),
    .B(_1000_),
    .C(_0217_),
    .Y(_0258_));
 OA33x2_ASAP7_75t_R _1645_ (.A1(_0210_),
    .A2(_0254_),
    .A3(_0256_),
    .B1(_0257_),
    .B2(_0258_),
    .B3(_0220_),
    .Y(_0259_));
 AND3x1_ASAP7_75t_R _1646_ (.A(_0251_),
    .B(_0252_),
    .C(_0259_),
    .Y(net322));
 OR3x1_ASAP7_75t_R _1647_ (.A(net127),
    .B(_0203_),
    .C(_0204_),
    .Y(_0260_));
 OR3x1_ASAP7_75t_R _1648_ (.A(net86),
    .B(_0206_),
    .C(_0237_),
    .Y(_0261_));
 AND2x2_ASAP7_75t_R _1649_ (.A(net243),
    .B(_0253_),
    .Y(_0262_));
 AND2x2_ASAP7_75t_R _1650_ (.A(net284),
    .B(_0255_),
    .Y(_0263_));
 AND3x1_ASAP7_75t_R _1651_ (.A(net206),
    .B(_0213_),
    .C(_0214_),
    .Y(_0264_));
 AND3x1_ASAP7_75t_R _1652_ (.A(net165),
    .B(_1000_),
    .C(_0217_),
    .Y(_0265_));
 OA33x2_ASAP7_75t_R _1653_ (.A1(_0210_),
    .A2(_0262_),
    .A3(_0263_),
    .B1(_0264_),
    .B2(_0265_),
    .B3(_0220_),
    .Y(_0266_));
 AND3x1_ASAP7_75t_R _1654_ (.A(_0260_),
    .B(_0261_),
    .C(_0266_),
    .Y(net323));
 OR3x1_ASAP7_75t_R _1655_ (.A(net128),
    .B(_0203_),
    .C(_0204_),
    .Y(_0267_));
 OR3x1_ASAP7_75t_R _1656_ (.A(net87),
    .B(_0206_),
    .C(_0237_),
    .Y(_0268_));
 AND2x2_ASAP7_75t_R _1657_ (.A(net244),
    .B(_0253_),
    .Y(_0269_));
 AND2x2_ASAP7_75t_R _1658_ (.A(net285),
    .B(_0255_),
    .Y(_0270_));
 AND3x1_ASAP7_75t_R _1659_ (.A(net207),
    .B(_0213_),
    .C(_0214_),
    .Y(_0271_));
 AND3x1_ASAP7_75t_R _1660_ (.A(net166),
    .B(_1000_),
    .C(_0217_),
    .Y(_0272_));
 OA33x2_ASAP7_75t_R _1661_ (.A1(_0210_),
    .A2(_0269_),
    .A3(_0270_),
    .B1(_0271_),
    .B2(_0272_),
    .B3(_0220_),
    .Y(_0273_));
 AND3x1_ASAP7_75t_R _1662_ (.A(_0267_),
    .B(_0268_),
    .C(_0273_),
    .Y(net324));
 OR3x1_ASAP7_75t_R _1663_ (.A(net129),
    .B(_0203_),
    .C(_0204_),
    .Y(_0274_));
 BUFx6f_ASAP7_75t_R _1664_ (.A(_0202_),
    .Y(_0275_));
 OR3x1_ASAP7_75t_R _1665_ (.A(net88),
    .B(_0275_),
    .C(_0237_),
    .Y(_0276_));
 AND2x2_ASAP7_75t_R _1666_ (.A(net245),
    .B(_0253_),
    .Y(_0277_));
 AND2x2_ASAP7_75t_R _1667_ (.A(net286),
    .B(_0255_),
    .Y(_0278_));
 AND3x1_ASAP7_75t_R _1668_ (.A(net208),
    .B(_0213_),
    .C(_0214_),
    .Y(_0279_));
 AND3x1_ASAP7_75t_R _1669_ (.A(net167),
    .B(_1000_),
    .C(_0217_),
    .Y(_0280_));
 OA33x2_ASAP7_75t_R _1670_ (.A1(_0210_),
    .A2(_0277_),
    .A3(_0278_),
    .B1(_0279_),
    .B2(_0280_),
    .B3(_0220_),
    .Y(_0281_));
 AND3x1_ASAP7_75t_R _1671_ (.A(_0274_),
    .B(_0276_),
    .C(_0281_),
    .Y(net325));
 OR3x1_ASAP7_75t_R _1672_ (.A(net130),
    .B(_0203_),
    .C(_0204_),
    .Y(_0282_));
 OR3x1_ASAP7_75t_R _1673_ (.A(net89),
    .B(_0275_),
    .C(_0237_),
    .Y(_0283_));
 AND2x2_ASAP7_75t_R _1674_ (.A(net246),
    .B(_0253_),
    .Y(_0284_));
 AND2x2_ASAP7_75t_R _1675_ (.A(net287),
    .B(_0255_),
    .Y(_0285_));
 AND3x1_ASAP7_75t_R _1676_ (.A(net209),
    .B(_0213_),
    .C(_0214_),
    .Y(_0286_));
 BUFx6f_ASAP7_75t_R _1677_ (.A(_0934_),
    .Y(_0287_));
 AND3x1_ASAP7_75t_R _1678_ (.A(net168),
    .B(_0287_),
    .C(_0217_),
    .Y(_0288_));
 OA33x2_ASAP7_75t_R _1679_ (.A1(_0210_),
    .A2(_0284_),
    .A3(_0285_),
    .B1(_0286_),
    .B2(_0288_),
    .B3(_0220_),
    .Y(_0289_));
 AND3x1_ASAP7_75t_R _1680_ (.A(_0282_),
    .B(_0283_),
    .C(_0289_),
    .Y(net326));
 BUFx6f_ASAP7_75t_R _1681_ (.A(_0202_),
    .Y(_0290_));
 BUFx6f_ASAP7_75t_R _1682_ (.A(_0182_),
    .Y(_0291_));
 OR3x1_ASAP7_75t_R _1683_ (.A(net110),
    .B(_0290_),
    .C(_0291_),
    .Y(_0292_));
 OR3x1_ASAP7_75t_R _1684_ (.A(net90),
    .B(_0275_),
    .C(_0237_),
    .Y(_0293_));
 BUFx6f_ASAP7_75t_R _1685_ (.A(_0209_),
    .Y(_0294_));
 AND2x2_ASAP7_75t_R _1686_ (.A(net247),
    .B(_0253_),
    .Y(_0295_));
 AND2x2_ASAP7_75t_R _1687_ (.A(net267),
    .B(_0255_),
    .Y(_0296_));
 BUFx6f_ASAP7_75t_R _1688_ (.A(_0952_),
    .Y(_0297_));
 BUFx6f_ASAP7_75t_R _1689_ (.A(_0177_),
    .Y(_0298_));
 AND3x1_ASAP7_75t_R _1690_ (.A(net189),
    .B(_0297_),
    .C(_0298_),
    .Y(_0299_));
 BUFx6f_ASAP7_75t_R _1691_ (.A(_0216_),
    .Y(_0300_));
 AND3x1_ASAP7_75t_R _1692_ (.A(net169),
    .B(_0287_),
    .C(_0300_),
    .Y(_0301_));
 BUFx6f_ASAP7_75t_R _1693_ (.A(_0219_),
    .Y(_0302_));
 OA33x2_ASAP7_75t_R _1694_ (.A1(_0294_),
    .A2(_0295_),
    .A3(_0296_),
    .B1(_0299_),
    .B2(_0301_),
    .B3(_0302_),
    .Y(_0303_));
 AND3x1_ASAP7_75t_R _1695_ (.A(_0292_),
    .B(_0293_),
    .C(_0303_),
    .Y(net327));
 OR3x1_ASAP7_75t_R _1696_ (.A(net131),
    .B(_0290_),
    .C(_0291_),
    .Y(_0304_));
 OR3x1_ASAP7_75t_R _1697_ (.A(net91),
    .B(_0275_),
    .C(_0237_),
    .Y(_0305_));
 AND2x2_ASAP7_75t_R _1698_ (.A(net248),
    .B(_0253_),
    .Y(_0306_));
 AND2x2_ASAP7_75t_R _1699_ (.A(net288),
    .B(_0255_),
    .Y(_0307_));
 AND3x1_ASAP7_75t_R _1700_ (.A(net210),
    .B(_0297_),
    .C(_0298_),
    .Y(_0308_));
 AND3x1_ASAP7_75t_R _1701_ (.A(net170),
    .B(_0287_),
    .C(_0300_),
    .Y(_0309_));
 OA33x2_ASAP7_75t_R _1702_ (.A1(_0294_),
    .A2(_0306_),
    .A3(_0307_),
    .B1(_0308_),
    .B2(_0309_),
    .B3(_0302_),
    .Y(_0310_));
 AND3x1_ASAP7_75t_R _1703_ (.A(_0304_),
    .B(_0305_),
    .C(_0310_),
    .Y(net328));
 OR3x1_ASAP7_75t_R _1704_ (.A(net132),
    .B(_0290_),
    .C(_0291_),
    .Y(_0311_));
 OR3x1_ASAP7_75t_R _1705_ (.A(net92),
    .B(_0275_),
    .C(_0237_),
    .Y(_0312_));
 AND2x2_ASAP7_75t_R _1706_ (.A(net249),
    .B(_0253_),
    .Y(_0313_));
 AND2x2_ASAP7_75t_R _1707_ (.A(net289),
    .B(_0255_),
    .Y(_0314_));
 AND3x1_ASAP7_75t_R _1708_ (.A(net211),
    .B(_0297_),
    .C(_0298_),
    .Y(_0315_));
 AND3x1_ASAP7_75t_R _1709_ (.A(net171),
    .B(_0287_),
    .C(_0300_),
    .Y(_0316_));
 OA33x2_ASAP7_75t_R _1710_ (.A1(_0294_),
    .A2(_0313_),
    .A3(_0314_),
    .B1(_0315_),
    .B2(_0316_),
    .B3(_0302_),
    .Y(_0317_));
 AND3x1_ASAP7_75t_R _1711_ (.A(_0311_),
    .B(_0312_),
    .C(_0317_),
    .Y(net329));
 OR3x1_ASAP7_75t_R _1712_ (.A(net133),
    .B(_0290_),
    .C(_0291_),
    .Y(_0318_));
 BUFx6f_ASAP7_75t_R _1713_ (.A(_0185_),
    .Y(_0319_));
 OR3x1_ASAP7_75t_R _1714_ (.A(net93),
    .B(_0275_),
    .C(_0319_),
    .Y(_0320_));
 AND2x2_ASAP7_75t_R _1715_ (.A(net250),
    .B(_0253_),
    .Y(_0321_));
 AND2x2_ASAP7_75t_R _1716_ (.A(net290),
    .B(_0255_),
    .Y(_0322_));
 AND3x1_ASAP7_75t_R _1717_ (.A(net212),
    .B(_0297_),
    .C(_0298_),
    .Y(_0323_));
 AND3x1_ASAP7_75t_R _1718_ (.A(net172),
    .B(_0287_),
    .C(_0300_),
    .Y(_0324_));
 OA33x2_ASAP7_75t_R _1719_ (.A1(_0294_),
    .A2(_0321_),
    .A3(_0322_),
    .B1(_0323_),
    .B2(_0324_),
    .B3(_0302_),
    .Y(_0325_));
 AND3x1_ASAP7_75t_R _1720_ (.A(_0318_),
    .B(_0320_),
    .C(_0325_),
    .Y(net330));
 OR3x1_ASAP7_75t_R _1721_ (.A(net135),
    .B(_0290_),
    .C(_0291_),
    .Y(_0326_));
 OR3x1_ASAP7_75t_R _1722_ (.A(net94),
    .B(_0275_),
    .C(_0319_),
    .Y(_0327_));
 AND2x2_ASAP7_75t_R _1723_ (.A(net251),
    .B(_0253_),
    .Y(_0328_));
 AND2x2_ASAP7_75t_R _1724_ (.A(net292),
    .B(_0255_),
    .Y(_0329_));
 AND3x1_ASAP7_75t_R _1725_ (.A(net214),
    .B(_0297_),
    .C(_0298_),
    .Y(_0330_));
 AND3x1_ASAP7_75t_R _1726_ (.A(net173),
    .B(_0287_),
    .C(_0300_),
    .Y(_0331_));
 OA33x2_ASAP7_75t_R _1727_ (.A1(_0294_),
    .A2(_0328_),
    .A3(_0329_),
    .B1(_0330_),
    .B2(_0331_),
    .B3(_0302_),
    .Y(_0332_));
 AND3x1_ASAP7_75t_R _1728_ (.A(_0326_),
    .B(_0327_),
    .C(_0332_),
    .Y(net331));
 OR3x1_ASAP7_75t_R _1729_ (.A(net136),
    .B(_0290_),
    .C(_0291_),
    .Y(_0333_));
 OR3x1_ASAP7_75t_R _1730_ (.A(net95),
    .B(_0275_),
    .C(_0319_),
    .Y(_0334_));
 BUFx6f_ASAP7_75t_R _1731_ (.A(_0199_),
    .Y(_0335_));
 AND2x2_ASAP7_75t_R _1732_ (.A(net252),
    .B(_0335_),
    .Y(_0336_));
 BUFx6f_ASAP7_75t_R _1733_ (.A(_0195_),
    .Y(_0337_));
 AND2x2_ASAP7_75t_R _1734_ (.A(net293),
    .B(_0337_),
    .Y(_0338_));
 AND3x1_ASAP7_75t_R _1735_ (.A(net215),
    .B(_0297_),
    .C(_0298_),
    .Y(_0339_));
 AND3x1_ASAP7_75t_R _1736_ (.A(net174),
    .B(_0287_),
    .C(_0300_),
    .Y(_0340_));
 OA33x2_ASAP7_75t_R _1737_ (.A1(_0294_),
    .A2(_0336_),
    .A3(_0338_),
    .B1(_0339_),
    .B2(_0340_),
    .B3(_0302_),
    .Y(_0341_));
 AND3x1_ASAP7_75t_R _1738_ (.A(_0333_),
    .B(_0334_),
    .C(_0341_),
    .Y(net332));
 OR3x1_ASAP7_75t_R _1739_ (.A(net137),
    .B(_0290_),
    .C(_0291_),
    .Y(_0342_));
 OR3x1_ASAP7_75t_R _1740_ (.A(net96),
    .B(_0275_),
    .C(_0319_),
    .Y(_0343_));
 AND2x2_ASAP7_75t_R _1741_ (.A(net253),
    .B(_0335_),
    .Y(_0344_));
 AND2x2_ASAP7_75t_R _1742_ (.A(net294),
    .B(_0337_),
    .Y(_0345_));
 AND3x1_ASAP7_75t_R _1743_ (.A(net216),
    .B(_0297_),
    .C(_0298_),
    .Y(_0346_));
 AND3x1_ASAP7_75t_R _1744_ (.A(net175),
    .B(_0287_),
    .C(_0300_),
    .Y(_0347_));
 OA33x2_ASAP7_75t_R _1745_ (.A1(_0294_),
    .A2(_0344_),
    .A3(_0345_),
    .B1(_0346_),
    .B2(_0347_),
    .B3(_0302_),
    .Y(_0348_));
 AND3x1_ASAP7_75t_R _1746_ (.A(_0342_),
    .B(_0343_),
    .C(_0348_),
    .Y(net333));
 OR3x1_ASAP7_75t_R _1747_ (.A(net138),
    .B(_0290_),
    .C(_0291_),
    .Y(_0349_));
 OR3x1_ASAP7_75t_R _1748_ (.A(net97),
    .B(_0275_),
    .C(_0319_),
    .Y(_0350_));
 AND2x2_ASAP7_75t_R _1749_ (.A(net254),
    .B(_0335_),
    .Y(_0351_));
 AND2x2_ASAP7_75t_R _1750_ (.A(net295),
    .B(_0337_),
    .Y(_0352_));
 AND3x1_ASAP7_75t_R _1751_ (.A(net217),
    .B(_0297_),
    .C(_0298_),
    .Y(_0353_));
 AND3x1_ASAP7_75t_R _1752_ (.A(net176),
    .B(_0287_),
    .C(_0300_),
    .Y(_0354_));
 OA33x2_ASAP7_75t_R _1753_ (.A1(_0294_),
    .A2(_0351_),
    .A3(_0352_),
    .B1(_0353_),
    .B2(_0354_),
    .B3(_0302_),
    .Y(_0355_));
 AND3x1_ASAP7_75t_R _1754_ (.A(_0349_),
    .B(_0350_),
    .C(_0355_),
    .Y(net334));
 OR3x1_ASAP7_75t_R _1755_ (.A(net139),
    .B(_0290_),
    .C(_0291_),
    .Y(_0356_));
 BUFx6f_ASAP7_75t_R _1756_ (.A(_0202_),
    .Y(_0357_));
 OR3x1_ASAP7_75t_R _1757_ (.A(net98),
    .B(_0357_),
    .C(_0319_),
    .Y(_0358_));
 AND2x2_ASAP7_75t_R _1758_ (.A(net255),
    .B(_0335_),
    .Y(_0359_));
 AND2x2_ASAP7_75t_R _1759_ (.A(net296),
    .B(_0337_),
    .Y(_0360_));
 AND3x1_ASAP7_75t_R _1760_ (.A(net218),
    .B(_0297_),
    .C(_0298_),
    .Y(_0361_));
 AND3x1_ASAP7_75t_R _1761_ (.A(net177),
    .B(_0287_),
    .C(_0300_),
    .Y(_0362_));
 OA33x2_ASAP7_75t_R _1762_ (.A1(_0294_),
    .A2(_0359_),
    .A3(_0360_),
    .B1(_0361_),
    .B2(_0362_),
    .B3(_0302_),
    .Y(_0363_));
 AND3x1_ASAP7_75t_R _1763_ (.A(_0356_),
    .B(_0358_),
    .C(_0363_),
    .Y(net335));
 OR3x1_ASAP7_75t_R _1764_ (.A(net140),
    .B(_0290_),
    .C(_0291_),
    .Y(_0364_));
 OR3x1_ASAP7_75t_R _1765_ (.A(net99),
    .B(_0357_),
    .C(_0319_),
    .Y(_0365_));
 AND2x2_ASAP7_75t_R _1766_ (.A(net256),
    .B(_0335_),
    .Y(_0366_));
 AND2x2_ASAP7_75t_R _1767_ (.A(net297),
    .B(_0337_),
    .Y(_0367_));
 AND3x1_ASAP7_75t_R _1768_ (.A(net219),
    .B(_0297_),
    .C(_0298_),
    .Y(_0368_));
 BUFx6f_ASAP7_75t_R _1769_ (.A(_0934_),
    .Y(_0369_));
 AND3x1_ASAP7_75t_R _1770_ (.A(net178),
    .B(_0369_),
    .C(_0300_),
    .Y(_0370_));
 OA33x2_ASAP7_75t_R _1771_ (.A1(_0294_),
    .A2(_0366_),
    .A3(_0367_),
    .B1(_0368_),
    .B2(_0370_),
    .B3(_0302_),
    .Y(_0371_));
 AND3x1_ASAP7_75t_R _1772_ (.A(_0364_),
    .B(_0365_),
    .C(_0371_),
    .Y(net336));
 BUFx6f_ASAP7_75t_R _1773_ (.A(_0202_),
    .Y(_0372_));
 BUFx6f_ASAP7_75t_R _1774_ (.A(_0182_),
    .Y(_0373_));
 OR3x1_ASAP7_75t_R _1775_ (.A(net141),
    .B(_0372_),
    .C(_0373_),
    .Y(_0374_));
 OR3x1_ASAP7_75t_R _1776_ (.A(net100),
    .B(_0357_),
    .C(_0319_),
    .Y(_0375_));
 BUFx6f_ASAP7_75t_R _1777_ (.A(_0209_),
    .Y(_0376_));
 AND2x2_ASAP7_75t_R _1778_ (.A(net257),
    .B(_0335_),
    .Y(_0377_));
 AND2x2_ASAP7_75t_R _1779_ (.A(net298),
    .B(_0337_),
    .Y(_0378_));
 BUFx6f_ASAP7_75t_R _1780_ (.A(_0952_),
    .Y(_0379_));
 BUFx6f_ASAP7_75t_R _1781_ (.A(_0177_),
    .Y(_0380_));
 AND3x1_ASAP7_75t_R _1782_ (.A(net220),
    .B(_0379_),
    .C(_0380_),
    .Y(_0381_));
 BUFx6f_ASAP7_75t_R _1783_ (.A(_0216_),
    .Y(_0382_));
 AND3x1_ASAP7_75t_R _1784_ (.A(net179),
    .B(_0369_),
    .C(_0382_),
    .Y(_0383_));
 BUFx6f_ASAP7_75t_R _1785_ (.A(_0219_),
    .Y(_0384_));
 OA33x2_ASAP7_75t_R _1786_ (.A1(_0376_),
    .A2(_0377_),
    .A3(_0378_),
    .B1(_0381_),
    .B2(_0383_),
    .B3(_0384_),
    .Y(_0385_));
 AND3x1_ASAP7_75t_R _1787_ (.A(_0374_),
    .B(_0375_),
    .C(_0385_),
    .Y(net337));
 OR3x1_ASAP7_75t_R _1788_ (.A(net111),
    .B(_0372_),
    .C(_0373_),
    .Y(_0386_));
 OR3x1_ASAP7_75t_R _1789_ (.A(net101),
    .B(_0357_),
    .C(_0319_),
    .Y(_0387_));
 AND2x2_ASAP7_75t_R _1790_ (.A(net258),
    .B(_0335_),
    .Y(_0388_));
 AND2x2_ASAP7_75t_R _1791_ (.A(net268),
    .B(_0337_),
    .Y(_0389_));
 AND3x1_ASAP7_75t_R _1792_ (.A(net190),
    .B(_0379_),
    .C(_0380_),
    .Y(_0390_));
 AND3x1_ASAP7_75t_R _1793_ (.A(net180),
    .B(_0369_),
    .C(_0382_),
    .Y(_0391_));
 OA33x2_ASAP7_75t_R _1794_ (.A1(_0376_),
    .A2(_0388_),
    .A3(_0389_),
    .B1(_0390_),
    .B2(_0391_),
    .B3(_0384_),
    .Y(_0392_));
 AND3x1_ASAP7_75t_R _1795_ (.A(_0386_),
    .B(_0387_),
    .C(_0392_),
    .Y(net338));
 OR3x1_ASAP7_75t_R _1796_ (.A(net142),
    .B(_0372_),
    .C(_0373_),
    .Y(_0393_));
 OR3x1_ASAP7_75t_R _1797_ (.A(net102),
    .B(_0357_),
    .C(_0319_),
    .Y(_0394_));
 AND2x2_ASAP7_75t_R _1798_ (.A(net259),
    .B(_0335_),
    .Y(_0395_));
 AND2x2_ASAP7_75t_R _1799_ (.A(net299),
    .B(_0337_),
    .Y(_0396_));
 AND3x1_ASAP7_75t_R _1800_ (.A(net221),
    .B(_0379_),
    .C(_0380_),
    .Y(_0397_));
 AND3x1_ASAP7_75t_R _1801_ (.A(net181),
    .B(_0369_),
    .C(_0382_),
    .Y(_0398_));
 OA33x2_ASAP7_75t_R _1802_ (.A1(_0376_),
    .A2(_0395_),
    .A3(_0396_),
    .B1(_0397_),
    .B2(_0398_),
    .B3(_0384_),
    .Y(_0399_));
 AND3x1_ASAP7_75t_R _1803_ (.A(_0393_),
    .B(_0394_),
    .C(_0399_),
    .Y(net339));
 OR3x1_ASAP7_75t_R _1804_ (.A(net143),
    .B(_0372_),
    .C(_0373_),
    .Y(_0400_));
 OR3x1_ASAP7_75t_R _1805_ (.A(net103),
    .B(_0357_),
    .C(_0196_),
    .Y(_0401_));
 AND2x2_ASAP7_75t_R _1806_ (.A(net260),
    .B(_0335_),
    .Y(_0402_));
 AND2x2_ASAP7_75t_R _1807_ (.A(net300),
    .B(_0337_),
    .Y(_0403_));
 AND3x1_ASAP7_75t_R _1808_ (.A(net222),
    .B(_0379_),
    .C(_0380_),
    .Y(_0404_));
 AND3x1_ASAP7_75t_R _1809_ (.A(net182),
    .B(_0369_),
    .C(_0382_),
    .Y(_0405_));
 OA33x2_ASAP7_75t_R _1810_ (.A1(_0376_),
    .A2(_0402_),
    .A3(_0403_),
    .B1(_0404_),
    .B2(_0405_),
    .B3(_0384_),
    .Y(_0406_));
 AND3x1_ASAP7_75t_R _1811_ (.A(_0400_),
    .B(_0401_),
    .C(_0406_),
    .Y(net340));
 AND2x2_ASAP7_75t_R _1812_ (.A(net261),
    .B(_0200_),
    .Y(_0407_));
 AO21x1_ASAP7_75t_R _1813_ (.A1(net301),
    .A2(_0207_),
    .B(_0407_),
    .Y(_0408_));
 AND2x2_ASAP7_75t_R _1814_ (.A(_0197_),
    .B(_0408_),
    .Y(net341));
 AND2x2_ASAP7_75t_R _1815_ (.A(net262),
    .B(_0200_),
    .Y(_0409_));
 AO21x1_ASAP7_75t_R _1816_ (.A1(net303),
    .A2(_0207_),
    .B(_0409_),
    .Y(_0410_));
 AND2x2_ASAP7_75t_R _1817_ (.A(net184),
    .B(_0200_),
    .Y(_0411_));
 AO21x1_ASAP7_75t_R _1818_ (.A1(net225),
    .A2(_0207_),
    .B(_0411_),
    .Y(_0412_));
 AO22x1_ASAP7_75t_R _1819_ (.A1(_0197_),
    .A2(_0410_),
    .B1(_0412_),
    .B2(_0190_),
    .Y(net342));
 AND2x2_ASAP7_75t_R _1820_ (.A(net263),
    .B(_0200_),
    .Y(_0413_));
 AO21x1_ASAP7_75t_R _1821_ (.A1(net304),
    .A2(_0207_),
    .B(_0413_),
    .Y(_0414_));
 AND2x2_ASAP7_75t_R _1822_ (.A(net185),
    .B(_0200_),
    .Y(_0415_));
 AO21x1_ASAP7_75t_R _1823_ (.A1(net226),
    .A2(_0207_),
    .B(_0415_),
    .Y(_0416_));
 AO22x1_ASAP7_75t_R _1824_ (.A1(_0197_),
    .A2(_0414_),
    .B1(_0416_),
    .B2(_0190_),
    .Y(net343));
 AND2x2_ASAP7_75t_R _1825_ (.A(net264),
    .B(_0200_),
    .Y(_0417_));
 AO21x1_ASAP7_75t_R _1826_ (.A1(net305),
    .A2(_0207_),
    .B(_0417_),
    .Y(_0418_));
 AND2x2_ASAP7_75t_R _1827_ (.A(net186),
    .B(_0200_),
    .Y(_0419_));
 AO21x1_ASAP7_75t_R _1828_ (.A1(net227),
    .A2(_0207_),
    .B(_0419_),
    .Y(_0420_));
 AO22x1_ASAP7_75t_R _1829_ (.A1(_0197_),
    .A2(_0418_),
    .B1(_0420_),
    .B2(_0190_),
    .Y(net344));
 OR3x1_ASAP7_75t_R _1830_ (.A(net149),
    .B(_0372_),
    .C(_0373_),
    .Y(_0421_));
 OR3x1_ASAP7_75t_R _1831_ (.A(net108),
    .B(_0357_),
    .C(_0196_),
    .Y(_0422_));
 AND2x2_ASAP7_75t_R _1832_ (.A(net265),
    .B(_0335_),
    .Y(_0423_));
 AND2x2_ASAP7_75t_R _1833_ (.A(net306),
    .B(_0337_),
    .Y(_0424_));
 AND3x1_ASAP7_75t_R _1834_ (.A(net228),
    .B(_0379_),
    .C(_0380_),
    .Y(_0425_));
 AND3x1_ASAP7_75t_R _1835_ (.A(net187),
    .B(_0369_),
    .C(_0382_),
    .Y(_0426_));
 OA33x2_ASAP7_75t_R _1836_ (.A1(_0376_),
    .A2(_0423_),
    .A3(_0424_),
    .B1(_0425_),
    .B2(_0426_),
    .B3(_0384_),
    .Y(_0427_));
 AND3x1_ASAP7_75t_R _1837_ (.A(_0421_),
    .B(_0422_),
    .C(_0427_),
    .Y(net345));
 OR3x1_ASAP7_75t_R _1838_ (.A(net113),
    .B(_0372_),
    .C(_0373_),
    .Y(_0428_));
 OR3x1_ASAP7_75t_R _1839_ (.A(net112),
    .B(_0357_),
    .C(_0196_),
    .Y(_0429_));
 AND2x2_ASAP7_75t_R _1840_ (.A(net269),
    .B(_0199_),
    .Y(_0430_));
 AND2x2_ASAP7_75t_R _1841_ (.A(net270),
    .B(_0195_),
    .Y(_0431_));
 AND3x1_ASAP7_75t_R _1842_ (.A(net192),
    .B(_0379_),
    .C(_0380_),
    .Y(_0432_));
 AND3x1_ASAP7_75t_R _1843_ (.A(net191),
    .B(_0369_),
    .C(_0382_),
    .Y(_0433_));
 OA33x2_ASAP7_75t_R _1844_ (.A1(_0376_),
    .A2(_0430_),
    .A3(_0431_),
    .B1(_0432_),
    .B2(_0433_),
    .B3(_0384_),
    .Y(_0434_));
 AND3x1_ASAP7_75t_R _1845_ (.A(_0428_),
    .B(_0429_),
    .C(_0434_),
    .Y(net346));
 OR3x1_ASAP7_75t_R _1846_ (.A(net114),
    .B(_0372_),
    .C(_0373_),
    .Y(_0435_));
 OR3x1_ASAP7_75t_R _1847_ (.A(net123),
    .B(_0357_),
    .C(_0196_),
    .Y(_0436_));
 AND2x2_ASAP7_75t_R _1848_ (.A(net280),
    .B(_0199_),
    .Y(_0437_));
 AND2x2_ASAP7_75t_R _1849_ (.A(net271),
    .B(_0195_),
    .Y(_0438_));
 AND3x1_ASAP7_75t_R _1850_ (.A(net193),
    .B(_0379_),
    .C(_0380_),
    .Y(_0439_));
 AND3x1_ASAP7_75t_R _1851_ (.A(net202),
    .B(_0369_),
    .C(_0382_),
    .Y(_0440_));
 OA33x2_ASAP7_75t_R _1852_ (.A1(_0376_),
    .A2(_0437_),
    .A3(_0438_),
    .B1(_0439_),
    .B2(_0440_),
    .B3(_0384_),
    .Y(_0441_));
 AND3x1_ASAP7_75t_R _1853_ (.A(_0435_),
    .B(_0436_),
    .C(_0441_),
    .Y(net347));
 OR3x1_ASAP7_75t_R _1854_ (.A(net115),
    .B(_0372_),
    .C(_0373_),
    .Y(_0442_));
 OR3x1_ASAP7_75t_R _1855_ (.A(net134),
    .B(_0357_),
    .C(_0196_),
    .Y(_0443_));
 AND2x2_ASAP7_75t_R _1856_ (.A(net291),
    .B(_0199_),
    .Y(_0444_));
 AND2x2_ASAP7_75t_R _1857_ (.A(net272),
    .B(_0195_),
    .Y(_0445_));
 AND3x1_ASAP7_75t_R _1858_ (.A(net194),
    .B(_0379_),
    .C(_0380_),
    .Y(_0446_));
 AND3x1_ASAP7_75t_R _1859_ (.A(net213),
    .B(_0369_),
    .C(_0382_),
    .Y(_0447_));
 OA33x2_ASAP7_75t_R _1860_ (.A1(_0376_),
    .A2(_0444_),
    .A3(_0445_),
    .B1(_0446_),
    .B2(_0447_),
    .B3(_0384_),
    .Y(_0448_));
 AND3x1_ASAP7_75t_R _1861_ (.A(_0442_),
    .B(_0443_),
    .C(_0448_),
    .Y(net348));
 OR3x1_ASAP7_75t_R _1862_ (.A(net116),
    .B(_0372_),
    .C(_0373_),
    .Y(_0449_));
 OR3x1_ASAP7_75t_R _1863_ (.A(net145),
    .B(_0202_),
    .C(_0196_),
    .Y(_0450_));
 AND2x2_ASAP7_75t_R _1864_ (.A(net302),
    .B(_0199_),
    .Y(_0451_));
 AND2x2_ASAP7_75t_R _1865_ (.A(net273),
    .B(_0195_),
    .Y(_0452_));
 AND3x1_ASAP7_75t_R _1866_ (.A(net195),
    .B(_0379_),
    .C(_0380_),
    .Y(_0453_));
 AND3x1_ASAP7_75t_R _1867_ (.A(net224),
    .B(_0369_),
    .C(_0382_),
    .Y(_0454_));
 OA33x2_ASAP7_75t_R _1868_ (.A1(_0376_),
    .A2(_0451_),
    .A3(_0452_),
    .B1(_0453_),
    .B2(_0454_),
    .B3(_0384_),
    .Y(_0455_));
 AND3x1_ASAP7_75t_R _1869_ (.A(_0449_),
    .B(_0450_),
    .C(_0455_),
    .Y(net349));
 OR3x1_ASAP7_75t_R _1870_ (.A(net117),
    .B(_0372_),
    .C(_0373_),
    .Y(_0456_));
 OR3x1_ASAP7_75t_R _1871_ (.A(net150),
    .B(_0202_),
    .C(_0196_),
    .Y(_0457_));
 AND2x2_ASAP7_75t_R _1872_ (.A(net307),
    .B(_0199_),
    .Y(_0458_));
 AND2x2_ASAP7_75t_R _1873_ (.A(net274),
    .B(_0195_),
    .Y(_0459_));
 AND3x1_ASAP7_75t_R _1874_ (.A(net196),
    .B(_0379_),
    .C(_0380_),
    .Y(_0460_));
 AND3x1_ASAP7_75t_R _1875_ (.A(net229),
    .B(_0934_),
    .C(_0382_),
    .Y(_0461_));
 OA33x2_ASAP7_75t_R _1876_ (.A1(_0376_),
    .A2(_0458_),
    .A3(_0459_),
    .B1(_0460_),
    .B2(_0461_),
    .B3(_0384_),
    .Y(_0462_));
 AND3x1_ASAP7_75t_R _1877_ (.A(_0456_),
    .B(_0457_),
    .C(_0462_),
    .Y(net350));
 OR3x1_ASAP7_75t_R _1878_ (.A(net118),
    .B(_0206_),
    .C(_0200_),
    .Y(_0463_));
 OR3x1_ASAP7_75t_R _1879_ (.A(net151),
    .B(_0202_),
    .C(_0196_),
    .Y(_0464_));
 AND2x2_ASAP7_75t_R _1880_ (.A(net308),
    .B(_0199_),
    .Y(_0465_));
 AND2x2_ASAP7_75t_R _1881_ (.A(net275),
    .B(_0195_),
    .Y(_0466_));
 AND3x1_ASAP7_75t_R _1882_ (.A(net197),
    .B(_0952_),
    .C(_0177_),
    .Y(_0467_));
 AND3x1_ASAP7_75t_R _1883_ (.A(net230),
    .B(_0934_),
    .C(_0216_),
    .Y(_0468_));
 OA33x2_ASAP7_75t_R _1884_ (.A1(_0209_),
    .A2(_0465_),
    .A3(_0466_),
    .B1(_0467_),
    .B2(_0468_),
    .B3(_0219_),
    .Y(_0469_));
 AND3x1_ASAP7_75t_R _1885_ (.A(_0463_),
    .B(_0464_),
    .C(_0469_),
    .Y(net351));
 OR3x1_ASAP7_75t_R _1886_ (.A(net119),
    .B(_0206_),
    .C(_0200_),
    .Y(_0470_));
 OR3x1_ASAP7_75t_R _1887_ (.A(net152),
    .B(_0202_),
    .C(_0196_),
    .Y(_0471_));
 AND2x2_ASAP7_75t_R _1888_ (.A(net309),
    .B(_0199_),
    .Y(_0472_));
 AND2x2_ASAP7_75t_R _1889_ (.A(net276),
    .B(_0195_),
    .Y(_0473_));
 AND3x1_ASAP7_75t_R _1890_ (.A(net198),
    .B(_0952_),
    .C(_0177_),
    .Y(_0474_));
 AND3x1_ASAP7_75t_R _1891_ (.A(net231),
    .B(_0934_),
    .C(_0216_),
    .Y(_0475_));
 OA33x2_ASAP7_75t_R _1892_ (.A1(_0209_),
    .A2(_0472_),
    .A3(_0473_),
    .B1(_0474_),
    .B2(_0475_),
    .B3(_0219_),
    .Y(_0476_));
 AND3x1_ASAP7_75t_R _1893_ (.A(_0470_),
    .B(_0471_),
    .C(_0476_),
    .Y(net352));
 AO222x2_ASAP7_75t_R _1894_ (.A1(_0983_),
    .A2(_0963_),
    .B1(_0984_),
    .B2(_0968_),
    .C1(_0976_),
    .C2(_0981_),
    .Y(_0477_));
 BUFx6f_ASAP7_75t_R _1895_ (.A(_0477_),
    .Y(_0478_));
 BUFx6f_ASAP7_75t_R _1896_ (.A(_0478_),
    .Y(_0479_));
 AND3x1_ASAP7_75t_R _1897_ (.A(net158),
    .B(_0994_),
    .C(_0479_),
    .Y(_0480_));
 NAND2x1_ASAP7_75t_R _1898_ (.A(_0965_),
    .B(_0478_),
    .Y(_0481_));
 BUFx12f_ASAP7_75t_R _1899_ (.A(_0481_),
    .Y(_0482_));
 AND2x2_ASAP7_75t_R _1900_ (.A(net188),
    .B(_0482_),
    .Y(_0483_));
 OR3x1_ASAP7_75t_R _1901_ (.A(_0960_),
    .B(_0961_),
    .C(_0962_),
    .Y(_0484_));
 AO21x2_ASAP7_75t_R _1902_ (.A1(_0959_),
    .A2(_0484_),
    .B(_0955_),
    .Y(_0485_));
 BUFx12f_ASAP7_75t_R _1903_ (.A(_0485_),
    .Y(_0486_));
 NAND2x2_ASAP7_75t_R _1904_ (.A(_0984_),
    .B(_0968_),
    .Y(_0487_));
 NAND2x1_ASAP7_75t_R _1905_ (.A(_0976_),
    .B(_0487_),
    .Y(_0488_));
 AND2x4_ASAP7_75t_R _1906_ (.A(_0486_),
    .B(_0488_),
    .Y(_0489_));
 OA21x2_ASAP7_75t_R _1907_ (.A1(_0480_),
    .A2(_0483_),
    .B(_0489_),
    .Y(_0490_));
 AND2x2_ASAP7_75t_R _1908_ (.A(_0994_),
    .B(_0479_),
    .Y(_0491_));
 NAND2x1_ASAP7_75t_R _1909_ (.A(net1),
    .B(_0491_),
    .Y(_0492_));
 NAND2x1_ASAP7_75t_R _1910_ (.A(net31),
    .B(_0482_),
    .Y(_0493_));
 AOI21x1_ASAP7_75t_R _1911_ (.A1(_0492_),
    .A2(_0493_),
    .B(_0486_),
    .Y(_0494_));
 AND3x4_ASAP7_75t_R _1912_ (.A(_0976_),
    .B(_0487_),
    .C(_0486_),
    .Y(_0495_));
 AND3x1_ASAP7_75t_R _1913_ (.A(net266),
    .B(_0482_),
    .C(_0495_),
    .Y(_0496_));
 AND3x1_ASAP7_75t_R _1914_ (.A(net236),
    .B(_0491_),
    .C(_0495_),
    .Y(_0497_));
 OR4x1_ASAP7_75t_R _1915_ (.A(_0490_),
    .B(_0494_),
    .C(_0496_),
    .D(_0497_),
    .Y(net357));
 NAND2x2_ASAP7_75t_R _1916_ (.A(_0486_),
    .B(_0488_),
    .Y(_0498_));
 BUFx6f_ASAP7_75t_R _1917_ (.A(_0498_),
    .Y(_0499_));
 OR2x2_ASAP7_75t_R _1918_ (.A(_0955_),
    .B(_0484_),
    .Y(_0500_));
 NAND2x1_ASAP7_75t_R _1919_ (.A(_0976_),
    .B(_0981_),
    .Y(_0501_));
 AND3x4_ASAP7_75t_R _1920_ (.A(_0487_),
    .B(_0500_),
    .C(_0501_),
    .Y(_0502_));
 BUFx6f_ASAP7_75t_R _1921_ (.A(_0502_),
    .Y(_0503_));
 BUFx6f_ASAP7_75t_R _1922_ (.A(_0479_),
    .Y(_0504_));
 AND3x1_ASAP7_75t_R _1923_ (.A(net159),
    .B(_0995_),
    .C(_0504_),
    .Y(_0505_));
 AO21x1_ASAP7_75t_R _1924_ (.A1(net199),
    .A2(_0503_),
    .B(_0505_),
    .Y(_0506_));
 BUFx6f_ASAP7_75t_R _1925_ (.A(_0482_),
    .Y(_0507_));
 BUFx6f_ASAP7_75t_R _1926_ (.A(_0965_),
    .Y(_0508_));
 BUFx6f_ASAP7_75t_R _1927_ (.A(_0479_),
    .Y(_0509_));
 AND3x1_ASAP7_75t_R _1928_ (.A(net237),
    .B(_0508_),
    .C(_0509_),
    .Y(_0510_));
 AO21x1_ASAP7_75t_R _1929_ (.A1(net277),
    .A2(_0507_),
    .B(_0510_),
    .Y(_0511_));
 NAND3x2_ASAP7_75t_R _1930_ (.B(_0487_),
    .C(_0486_),
    .Y(_0512_),
    .A(_0976_));
 BUFx6f_ASAP7_75t_R _1931_ (.A(_0512_),
    .Y(_0513_));
 BUFx6f_ASAP7_75t_R _1932_ (.A(_0482_),
    .Y(_0514_));
 BUFx6f_ASAP7_75t_R _1933_ (.A(_0965_),
    .Y(_0515_));
 BUFx6f_ASAP7_75t_R _1934_ (.A(_0478_),
    .Y(_0516_));
 AND3x1_ASAP7_75t_R _1935_ (.A(net2),
    .B(_0515_),
    .C(_0516_),
    .Y(_0517_));
 AO21x1_ASAP7_75t_R _1936_ (.A1(net42),
    .A2(_0514_),
    .B(_0517_),
    .Y(_0518_));
 BUFx6f_ASAP7_75t_R _1937_ (.A(_0486_),
    .Y(_0519_));
 OA222x2_ASAP7_75t_R _1938_ (.A1(_0499_),
    .A2(_0506_),
    .B1(_0511_),
    .B2(_0513_),
    .C1(_0518_),
    .C2(_0519_),
    .Y(net358));
 AND3x1_ASAP7_75t_R _1939_ (.A(net160),
    .B(_0995_),
    .C(_0504_),
    .Y(_0520_));
 AO21x1_ASAP7_75t_R _1940_ (.A1(net200),
    .A2(_0503_),
    .B(_0520_),
    .Y(_0521_));
 BUFx6f_ASAP7_75t_R _1941_ (.A(_0479_),
    .Y(_0522_));
 AND3x1_ASAP7_75t_R _1942_ (.A(net238),
    .B(_0508_),
    .C(_0522_),
    .Y(_0523_));
 AO21x1_ASAP7_75t_R _1943_ (.A1(net278),
    .A2(_0507_),
    .B(_0523_),
    .Y(_0524_));
 AND3x1_ASAP7_75t_R _1944_ (.A(net3),
    .B(_0515_),
    .C(_0516_),
    .Y(_0525_));
 AO21x1_ASAP7_75t_R _1945_ (.A1(net43),
    .A2(_0514_),
    .B(_0525_),
    .Y(_0526_));
 OA222x2_ASAP7_75t_R _1946_ (.A1(_0499_),
    .A2(_0521_),
    .B1(_0524_),
    .B2(_0513_),
    .C1(_0526_),
    .C2(_0519_),
    .Y(net359));
 BUFx6f_ASAP7_75t_R _1947_ (.A(_0994_),
    .Y(_0527_));
 AND3x1_ASAP7_75t_R _1948_ (.A(net161),
    .B(_0527_),
    .C(_0504_),
    .Y(_0528_));
 AO21x1_ASAP7_75t_R _1949_ (.A1(net201),
    .A2(_0503_),
    .B(_0528_),
    .Y(_0529_));
 AND3x1_ASAP7_75t_R _1950_ (.A(net239),
    .B(_0508_),
    .C(_0522_),
    .Y(_0530_));
 AO21x1_ASAP7_75t_R _1951_ (.A1(net279),
    .A2(_0507_),
    .B(_0530_),
    .Y(_0531_));
 BUFx6f_ASAP7_75t_R _1952_ (.A(_0482_),
    .Y(_0532_));
 AND3x1_ASAP7_75t_R _1953_ (.A(net4),
    .B(_0515_),
    .C(_0516_),
    .Y(_0533_));
 AO21x1_ASAP7_75t_R _1954_ (.A1(net44),
    .A2(_0532_),
    .B(_0533_),
    .Y(_0534_));
 OA222x2_ASAP7_75t_R _1955_ (.A1(_0499_),
    .A2(_0529_),
    .B1(_0531_),
    .B2(_0513_),
    .C1(_0534_),
    .C2(_0519_),
    .Y(net360));
 BUFx6f_ASAP7_75t_R _1956_ (.A(_0479_),
    .Y(_0535_));
 AND3x1_ASAP7_75t_R _1957_ (.A(net162),
    .B(_0527_),
    .C(_0535_),
    .Y(_0536_));
 AO21x1_ASAP7_75t_R _1958_ (.A1(net203),
    .A2(_0503_),
    .B(_0536_),
    .Y(_0537_));
 AND3x1_ASAP7_75t_R _1959_ (.A(net240),
    .B(_0508_),
    .C(_0522_),
    .Y(_0538_));
 AO21x1_ASAP7_75t_R _1960_ (.A1(net281),
    .A2(_0507_),
    .B(_0538_),
    .Y(_0539_));
 AND3x1_ASAP7_75t_R _1961_ (.A(net5),
    .B(_0515_),
    .C(_0516_),
    .Y(_0540_));
 AO21x1_ASAP7_75t_R _1962_ (.A1(net46),
    .A2(_0532_),
    .B(_0540_),
    .Y(_0541_));
 OA222x2_ASAP7_75t_R _1963_ (.A1(_0499_),
    .A2(_0537_),
    .B1(_0539_),
    .B2(_0513_),
    .C1(_0541_),
    .C2(_0519_),
    .Y(net361));
 AND3x1_ASAP7_75t_R _1964_ (.A(net163),
    .B(_0527_),
    .C(_0535_),
    .Y(_0542_));
 AO21x1_ASAP7_75t_R _1965_ (.A1(net204),
    .A2(_0503_),
    .B(_0542_),
    .Y(_0543_));
 BUFx6f_ASAP7_75t_R _1966_ (.A(_0482_),
    .Y(_0544_));
 AND3x1_ASAP7_75t_R _1967_ (.A(net241),
    .B(_0508_),
    .C(_0522_),
    .Y(_0545_));
 AO21x1_ASAP7_75t_R _1968_ (.A1(net282),
    .A2(_0544_),
    .B(_0545_),
    .Y(_0546_));
 AND3x1_ASAP7_75t_R _1969_ (.A(net6),
    .B(_0515_),
    .C(_0516_),
    .Y(_0547_));
 AO21x1_ASAP7_75t_R _1970_ (.A1(net47),
    .A2(_0532_),
    .B(_0547_),
    .Y(_0548_));
 OA222x2_ASAP7_75t_R _1971_ (.A1(_0499_),
    .A2(_0543_),
    .B1(_0546_),
    .B2(_0513_),
    .C1(_0548_),
    .C2(_0519_),
    .Y(net362));
 AND3x1_ASAP7_75t_R _1972_ (.A(net164),
    .B(_0527_),
    .C(_0535_),
    .Y(_0549_));
 AO21x1_ASAP7_75t_R _1973_ (.A1(net205),
    .A2(_0503_),
    .B(_0549_),
    .Y(_0550_));
 AND3x1_ASAP7_75t_R _1974_ (.A(net242),
    .B(_0508_),
    .C(_0522_),
    .Y(_0551_));
 AO21x1_ASAP7_75t_R _1975_ (.A1(net283),
    .A2(_0544_),
    .B(_0551_),
    .Y(_0552_));
 AND3x1_ASAP7_75t_R _1976_ (.A(net7),
    .B(_0515_),
    .C(_0516_),
    .Y(_0553_));
 AO21x1_ASAP7_75t_R _1977_ (.A1(net48),
    .A2(_0532_),
    .B(_0553_),
    .Y(_0554_));
 OA222x2_ASAP7_75t_R _1978_ (.A1(_0499_),
    .A2(_0550_),
    .B1(_0552_),
    .B2(_0513_),
    .C1(_0554_),
    .C2(_0519_),
    .Y(net363));
 AND3x1_ASAP7_75t_R _1979_ (.A(net165),
    .B(_0527_),
    .C(_0535_),
    .Y(_0555_));
 AO21x1_ASAP7_75t_R _1980_ (.A1(net206),
    .A2(_0503_),
    .B(_0555_),
    .Y(_0556_));
 AND3x1_ASAP7_75t_R _1981_ (.A(net243),
    .B(_0508_),
    .C(_0522_),
    .Y(_0557_));
 AO21x1_ASAP7_75t_R _1982_ (.A1(net284),
    .A2(_0544_),
    .B(_0557_),
    .Y(_0558_));
 AND3x1_ASAP7_75t_R _1983_ (.A(net8),
    .B(_0515_),
    .C(_0516_),
    .Y(_0559_));
 AO21x1_ASAP7_75t_R _1984_ (.A1(net49),
    .A2(_0532_),
    .B(_0559_),
    .Y(_0560_));
 OA222x2_ASAP7_75t_R _1985_ (.A1(_0499_),
    .A2(_0556_),
    .B1(_0558_),
    .B2(_0513_),
    .C1(_0560_),
    .C2(_0519_),
    .Y(net364));
 AND3x1_ASAP7_75t_R _1986_ (.A(net166),
    .B(_0527_),
    .C(_0535_),
    .Y(_0561_));
 AO21x1_ASAP7_75t_R _1987_ (.A1(net207),
    .A2(_0503_),
    .B(_0561_),
    .Y(_0562_));
 AND3x1_ASAP7_75t_R _1988_ (.A(net244),
    .B(_0508_),
    .C(_0522_),
    .Y(_0563_));
 AO21x1_ASAP7_75t_R _1989_ (.A1(net285),
    .A2(_0544_),
    .B(_0563_),
    .Y(_0564_));
 AND3x1_ASAP7_75t_R _1990_ (.A(net9),
    .B(_0515_),
    .C(_0516_),
    .Y(_0565_));
 AO21x1_ASAP7_75t_R _1991_ (.A1(net50),
    .A2(_0532_),
    .B(_0565_),
    .Y(_0566_));
 OA222x2_ASAP7_75t_R _1992_ (.A1(_0499_),
    .A2(_0562_),
    .B1(_0564_),
    .B2(_0513_),
    .C1(_0566_),
    .C2(_0519_),
    .Y(net365));
 AND3x1_ASAP7_75t_R _1993_ (.A(net167),
    .B(_0527_),
    .C(_0535_),
    .Y(_0567_));
 AO21x1_ASAP7_75t_R _1994_ (.A1(net208),
    .A2(_0503_),
    .B(_0567_),
    .Y(_0568_));
 AND3x1_ASAP7_75t_R _1995_ (.A(net245),
    .B(_0508_),
    .C(_0522_),
    .Y(_0569_));
 AO21x1_ASAP7_75t_R _1996_ (.A1(net286),
    .A2(_0544_),
    .B(_0569_),
    .Y(_0570_));
 BUFx6f_ASAP7_75t_R _1997_ (.A(_0965_),
    .Y(_0571_));
 AND3x1_ASAP7_75t_R _1998_ (.A(net10),
    .B(_0571_),
    .C(_0516_),
    .Y(_0572_));
 AO21x1_ASAP7_75t_R _1999_ (.A1(net51),
    .A2(_0532_),
    .B(_0572_),
    .Y(_0573_));
 OA222x2_ASAP7_75t_R _2000_ (.A1(_0499_),
    .A2(_0568_),
    .B1(_0570_),
    .B2(_0513_),
    .C1(_0573_),
    .C2(_0519_),
    .Y(net366));
 AND3x1_ASAP7_75t_R _2001_ (.A(net168),
    .B(_0527_),
    .C(_0535_),
    .Y(_0574_));
 AO21x1_ASAP7_75t_R _2002_ (.A1(net209),
    .A2(_0503_),
    .B(_0574_),
    .Y(_0575_));
 AND3x1_ASAP7_75t_R _2003_ (.A(net246),
    .B(_0508_),
    .C(_0522_),
    .Y(_0576_));
 AO21x1_ASAP7_75t_R _2004_ (.A1(net287),
    .A2(_0544_),
    .B(_0576_),
    .Y(_0577_));
 BUFx6f_ASAP7_75t_R _2005_ (.A(_0512_),
    .Y(_0578_));
 BUFx6f_ASAP7_75t_R _2006_ (.A(_0478_),
    .Y(_0579_));
 AND3x1_ASAP7_75t_R _2007_ (.A(net11),
    .B(_0571_),
    .C(_0579_),
    .Y(_0580_));
 AO21x1_ASAP7_75t_R _2008_ (.A1(net52),
    .A2(_0532_),
    .B(_0580_),
    .Y(_0581_));
 OA222x2_ASAP7_75t_R _2009_ (.A1(_0499_),
    .A2(_0575_),
    .B1(_0577_),
    .B2(_0578_),
    .C1(_0581_),
    .C2(_0519_),
    .Y(net367));
 BUFx6f_ASAP7_75t_R _2010_ (.A(_0498_),
    .Y(_0582_));
 BUFx6f_ASAP7_75t_R _2011_ (.A(_0502_),
    .Y(_0583_));
 AND3x1_ASAP7_75t_R _2012_ (.A(net169),
    .B(_0527_),
    .C(_0535_),
    .Y(_0584_));
 AO21x1_ASAP7_75t_R _2013_ (.A1(net189),
    .A2(_0583_),
    .B(_0584_),
    .Y(_0585_));
 BUFx6f_ASAP7_75t_R _2014_ (.A(_0965_),
    .Y(_0586_));
 AND3x1_ASAP7_75t_R _2015_ (.A(net247),
    .B(_0586_),
    .C(_0522_),
    .Y(_0587_));
 AO21x1_ASAP7_75t_R _2016_ (.A1(net267),
    .A2(_0544_),
    .B(_0587_),
    .Y(_0588_));
 AND3x1_ASAP7_75t_R _2017_ (.A(net12),
    .B(_0571_),
    .C(_0579_),
    .Y(_0589_));
 AO21x1_ASAP7_75t_R _2018_ (.A1(net32),
    .A2(_0532_),
    .B(_0589_),
    .Y(_0590_));
 BUFx6f_ASAP7_75t_R _2019_ (.A(_0486_),
    .Y(_0591_));
 OA222x2_ASAP7_75t_R _2020_ (.A1(_0582_),
    .A2(_0585_),
    .B1(_0588_),
    .B2(_0578_),
    .C1(_0590_),
    .C2(_0591_),
    .Y(net368));
 AND3x1_ASAP7_75t_R _2021_ (.A(net170),
    .B(_0527_),
    .C(_0535_),
    .Y(_0592_));
 AO21x1_ASAP7_75t_R _2022_ (.A1(net210),
    .A2(_0583_),
    .B(_0592_),
    .Y(_0593_));
 BUFx6f_ASAP7_75t_R _2023_ (.A(_0478_),
    .Y(_0594_));
 AND3x1_ASAP7_75t_R _2024_ (.A(net248),
    .B(_0586_),
    .C(_0594_),
    .Y(_0595_));
 AO21x1_ASAP7_75t_R _2025_ (.A1(net288),
    .A2(_0544_),
    .B(_0595_),
    .Y(_0596_));
 AND3x1_ASAP7_75t_R _2026_ (.A(net13),
    .B(_0571_),
    .C(_0579_),
    .Y(_0597_));
 AO21x1_ASAP7_75t_R _2027_ (.A1(net53),
    .A2(_0532_),
    .B(_0597_),
    .Y(_0598_));
 OA222x2_ASAP7_75t_R _2028_ (.A1(_0582_),
    .A2(_0593_),
    .B1(_0596_),
    .B2(_0578_),
    .C1(_0598_),
    .C2(_0591_),
    .Y(net369));
 BUFx6f_ASAP7_75t_R _2029_ (.A(_0994_),
    .Y(_0599_));
 AND3x1_ASAP7_75t_R _2030_ (.A(net171),
    .B(_0599_),
    .C(_0535_),
    .Y(_0600_));
 AO21x1_ASAP7_75t_R _2031_ (.A1(net211),
    .A2(_0583_),
    .B(_0600_),
    .Y(_0601_));
 AND3x1_ASAP7_75t_R _2032_ (.A(net249),
    .B(_0586_),
    .C(_0594_),
    .Y(_0602_));
 AO21x1_ASAP7_75t_R _2033_ (.A1(net289),
    .A2(_0544_),
    .B(_0602_),
    .Y(_0603_));
 BUFx6f_ASAP7_75t_R _2034_ (.A(_0482_),
    .Y(_0604_));
 AND3x1_ASAP7_75t_R _2035_ (.A(net14),
    .B(_0571_),
    .C(_0579_),
    .Y(_0605_));
 AO21x1_ASAP7_75t_R _2036_ (.A1(net54),
    .A2(_0604_),
    .B(_0605_),
    .Y(_0606_));
 OA222x2_ASAP7_75t_R _2037_ (.A1(_0582_),
    .A2(_0601_),
    .B1(_0603_),
    .B2(_0578_),
    .C1(_0606_),
    .C2(_0591_),
    .Y(net370));
 BUFx6f_ASAP7_75t_R _2038_ (.A(_0479_),
    .Y(_0607_));
 AND3x1_ASAP7_75t_R _2039_ (.A(net172),
    .B(_0599_),
    .C(_0607_),
    .Y(_0608_));
 AO21x1_ASAP7_75t_R _2040_ (.A1(net212),
    .A2(_0583_),
    .B(_0608_),
    .Y(_0609_));
 AND3x1_ASAP7_75t_R _2041_ (.A(net250),
    .B(_0586_),
    .C(_0594_),
    .Y(_0610_));
 AO21x1_ASAP7_75t_R _2042_ (.A1(net290),
    .A2(_0544_),
    .B(_0610_),
    .Y(_0611_));
 AND3x1_ASAP7_75t_R _2043_ (.A(net15),
    .B(_0571_),
    .C(_0579_),
    .Y(_0612_));
 AO21x1_ASAP7_75t_R _2044_ (.A1(net55),
    .A2(_0604_),
    .B(_0612_),
    .Y(_0613_));
 OA222x2_ASAP7_75t_R _2045_ (.A1(_0582_),
    .A2(_0609_),
    .B1(_0611_),
    .B2(_0578_),
    .C1(_0613_),
    .C2(_0591_),
    .Y(net371));
 AND3x1_ASAP7_75t_R _2046_ (.A(net173),
    .B(_0599_),
    .C(_0607_),
    .Y(_0614_));
 AO21x1_ASAP7_75t_R _2047_ (.A1(net214),
    .A2(_0583_),
    .B(_0614_),
    .Y(_0615_));
 BUFx6f_ASAP7_75t_R _2048_ (.A(_0482_),
    .Y(_0616_));
 AND3x1_ASAP7_75t_R _2049_ (.A(net251),
    .B(_0586_),
    .C(_0594_),
    .Y(_0617_));
 AO21x1_ASAP7_75t_R _2050_ (.A1(net292),
    .A2(_0616_),
    .B(_0617_),
    .Y(_0618_));
 AND3x1_ASAP7_75t_R _2051_ (.A(net16),
    .B(_0571_),
    .C(_0579_),
    .Y(_0619_));
 AO21x1_ASAP7_75t_R _2052_ (.A1(net57),
    .A2(_0604_),
    .B(_0619_),
    .Y(_0620_));
 OA222x2_ASAP7_75t_R _2053_ (.A1(_0582_),
    .A2(_0615_),
    .B1(_0618_),
    .B2(_0578_),
    .C1(_0620_),
    .C2(_0591_),
    .Y(net372));
 AND3x1_ASAP7_75t_R _2054_ (.A(net174),
    .B(_0599_),
    .C(_0607_),
    .Y(_0621_));
 AO21x1_ASAP7_75t_R _2055_ (.A1(net215),
    .A2(_0583_),
    .B(_0621_),
    .Y(_0622_));
 AND3x1_ASAP7_75t_R _2056_ (.A(net252),
    .B(_0586_),
    .C(_0594_),
    .Y(_0623_));
 AO21x1_ASAP7_75t_R _2057_ (.A1(net293),
    .A2(_0616_),
    .B(_0623_),
    .Y(_0624_));
 AND3x1_ASAP7_75t_R _2058_ (.A(net17),
    .B(_0571_),
    .C(_0579_),
    .Y(_0625_));
 AO21x1_ASAP7_75t_R _2059_ (.A1(net58),
    .A2(_0604_),
    .B(_0625_),
    .Y(_0626_));
 OA222x2_ASAP7_75t_R _2060_ (.A1(_0582_),
    .A2(_0622_),
    .B1(_0624_),
    .B2(_0578_),
    .C1(_0626_),
    .C2(_0591_),
    .Y(net373));
 AND3x1_ASAP7_75t_R _2061_ (.A(net175),
    .B(_0599_),
    .C(_0607_),
    .Y(_0627_));
 AO21x1_ASAP7_75t_R _2062_ (.A1(net216),
    .A2(_0583_),
    .B(_0627_),
    .Y(_0628_));
 AND3x1_ASAP7_75t_R _2063_ (.A(net253),
    .B(_0586_),
    .C(_0594_),
    .Y(_0629_));
 AO21x1_ASAP7_75t_R _2064_ (.A1(net294),
    .A2(_0616_),
    .B(_0629_),
    .Y(_0630_));
 AND3x1_ASAP7_75t_R _2065_ (.A(net18),
    .B(_0571_),
    .C(_0579_),
    .Y(_0631_));
 AO21x1_ASAP7_75t_R _2066_ (.A1(net59),
    .A2(_0604_),
    .B(_0631_),
    .Y(_0632_));
 OA222x2_ASAP7_75t_R _2067_ (.A1(_0582_),
    .A2(_0628_),
    .B1(_0630_),
    .B2(_0578_),
    .C1(_0632_),
    .C2(_0591_),
    .Y(net374));
 AND3x1_ASAP7_75t_R _2068_ (.A(net176),
    .B(_0599_),
    .C(_0607_),
    .Y(_0633_));
 AO21x1_ASAP7_75t_R _2069_ (.A1(net217),
    .A2(_0583_),
    .B(_0633_),
    .Y(_0634_));
 AND3x1_ASAP7_75t_R _2070_ (.A(net254),
    .B(_0586_),
    .C(_0594_),
    .Y(_0635_));
 AO21x1_ASAP7_75t_R _2071_ (.A1(net295),
    .A2(_0616_),
    .B(_0635_),
    .Y(_0636_));
 AND3x1_ASAP7_75t_R _2072_ (.A(net19),
    .B(_0571_),
    .C(_0579_),
    .Y(_0637_));
 AO21x1_ASAP7_75t_R _2073_ (.A1(net60),
    .A2(_0604_),
    .B(_0637_),
    .Y(_0638_));
 OA222x2_ASAP7_75t_R _2074_ (.A1(_0582_),
    .A2(_0634_),
    .B1(_0636_),
    .B2(_0578_),
    .C1(_0638_),
    .C2(_0591_),
    .Y(net375));
 AND3x1_ASAP7_75t_R _2075_ (.A(net177),
    .B(_0599_),
    .C(_0607_),
    .Y(_0639_));
 AO21x1_ASAP7_75t_R _2076_ (.A1(net218),
    .A2(_0583_),
    .B(_0639_),
    .Y(_0640_));
 AND3x1_ASAP7_75t_R _2077_ (.A(net255),
    .B(_0586_),
    .C(_0594_),
    .Y(_0641_));
 AO21x1_ASAP7_75t_R _2078_ (.A1(net296),
    .A2(_0616_),
    .B(_0641_),
    .Y(_0642_));
 BUFx6f_ASAP7_75t_R _2079_ (.A(_0965_),
    .Y(_0643_));
 AND3x1_ASAP7_75t_R _2080_ (.A(net20),
    .B(_0643_),
    .C(_0579_),
    .Y(_0644_));
 AO21x1_ASAP7_75t_R _2081_ (.A1(net61),
    .A2(_0604_),
    .B(_0644_),
    .Y(_0645_));
 OA222x2_ASAP7_75t_R _2082_ (.A1(_0582_),
    .A2(_0640_),
    .B1(_0642_),
    .B2(_0578_),
    .C1(_0645_),
    .C2(_0591_),
    .Y(net376));
 AND3x1_ASAP7_75t_R _2083_ (.A(net178),
    .B(_0599_),
    .C(_0607_),
    .Y(_0646_));
 AO21x1_ASAP7_75t_R _2084_ (.A1(net219),
    .A2(_0583_),
    .B(_0646_),
    .Y(_0647_));
 AND3x1_ASAP7_75t_R _2085_ (.A(net256),
    .B(_0586_),
    .C(_0594_),
    .Y(_0648_));
 AO21x1_ASAP7_75t_R _2086_ (.A1(net297),
    .A2(_0616_),
    .B(_0648_),
    .Y(_0649_));
 BUFx6f_ASAP7_75t_R _2087_ (.A(_0512_),
    .Y(_0650_));
 BUFx6f_ASAP7_75t_R _2088_ (.A(_0478_),
    .Y(_0651_));
 AND3x1_ASAP7_75t_R _2089_ (.A(net21),
    .B(_0643_),
    .C(_0651_),
    .Y(_0652_));
 AO21x1_ASAP7_75t_R _2090_ (.A1(net62),
    .A2(_0604_),
    .B(_0652_),
    .Y(_0653_));
 OA222x2_ASAP7_75t_R _2091_ (.A1(_0582_),
    .A2(_0647_),
    .B1(_0649_),
    .B2(_0650_),
    .C1(_0653_),
    .C2(_0591_),
    .Y(net377));
 BUFx6f_ASAP7_75t_R _2092_ (.A(_0498_),
    .Y(_0654_));
 BUFx6f_ASAP7_75t_R _2093_ (.A(_0502_),
    .Y(_0655_));
 AND3x1_ASAP7_75t_R _2094_ (.A(net179),
    .B(_0599_),
    .C(_0607_),
    .Y(_0656_));
 AO21x1_ASAP7_75t_R _2095_ (.A1(net220),
    .A2(_0655_),
    .B(_0656_),
    .Y(_0657_));
 BUFx6f_ASAP7_75t_R _2096_ (.A(_0965_),
    .Y(_0658_));
 AND3x1_ASAP7_75t_R _2097_ (.A(net257),
    .B(_0658_),
    .C(_0594_),
    .Y(_0659_));
 AO21x1_ASAP7_75t_R _2098_ (.A1(net298),
    .A2(_0616_),
    .B(_0659_),
    .Y(_0660_));
 AND3x1_ASAP7_75t_R _2099_ (.A(net22),
    .B(_0643_),
    .C(_0651_),
    .Y(_0661_));
 AO21x1_ASAP7_75t_R _2100_ (.A1(net63),
    .A2(_0604_),
    .B(_0661_),
    .Y(_0662_));
 BUFx6f_ASAP7_75t_R _2101_ (.A(_0486_),
    .Y(_0663_));
 OA222x2_ASAP7_75t_R _2102_ (.A1(_0654_),
    .A2(_0657_),
    .B1(_0660_),
    .B2(_0650_),
    .C1(_0662_),
    .C2(_0663_),
    .Y(net378));
 AND3x1_ASAP7_75t_R _2103_ (.A(net180),
    .B(_0599_),
    .C(_0607_),
    .Y(_0664_));
 AO21x1_ASAP7_75t_R _2104_ (.A1(net190),
    .A2(_0655_),
    .B(_0664_),
    .Y(_0665_));
 BUFx6f_ASAP7_75t_R _2105_ (.A(_0478_),
    .Y(_0666_));
 AND3x1_ASAP7_75t_R _2106_ (.A(net258),
    .B(_0658_),
    .C(_0666_),
    .Y(_0667_));
 AO21x1_ASAP7_75t_R _2107_ (.A1(net268),
    .A2(_0616_),
    .B(_0667_),
    .Y(_0668_));
 AND3x1_ASAP7_75t_R _2108_ (.A(net23),
    .B(_0643_),
    .C(_0651_),
    .Y(_0669_));
 AO21x1_ASAP7_75t_R _2109_ (.A1(net33),
    .A2(_0604_),
    .B(_0669_),
    .Y(_0670_));
 OA222x2_ASAP7_75t_R _2110_ (.A1(_0654_),
    .A2(_0665_),
    .B1(_0668_),
    .B2(_0650_),
    .C1(_0670_),
    .C2(_0663_),
    .Y(net379));
 BUFx6f_ASAP7_75t_R _2111_ (.A(_0994_),
    .Y(_0671_));
 AND3x1_ASAP7_75t_R _2112_ (.A(net181),
    .B(_0671_),
    .C(_0607_),
    .Y(_0672_));
 AO21x1_ASAP7_75t_R _2113_ (.A1(net221),
    .A2(_0655_),
    .B(_0672_),
    .Y(_0673_));
 AND3x1_ASAP7_75t_R _2114_ (.A(net259),
    .B(_0658_),
    .C(_0666_),
    .Y(_0674_));
 AO21x1_ASAP7_75t_R _2115_ (.A1(net299),
    .A2(_0616_),
    .B(_0674_),
    .Y(_0675_));
 BUFx6f_ASAP7_75t_R _2116_ (.A(_0481_),
    .Y(_0676_));
 AND3x1_ASAP7_75t_R _2117_ (.A(net24),
    .B(_0643_),
    .C(_0651_),
    .Y(_0677_));
 AO21x1_ASAP7_75t_R _2118_ (.A1(net64),
    .A2(_0676_),
    .B(_0677_),
    .Y(_0678_));
 OA222x2_ASAP7_75t_R _2119_ (.A1(_0654_),
    .A2(_0673_),
    .B1(_0675_),
    .B2(_0650_),
    .C1(_0678_),
    .C2(_0663_),
    .Y(net380));
 AND3x1_ASAP7_75t_R _2120_ (.A(net182),
    .B(_0671_),
    .C(_0509_),
    .Y(_0679_));
 AO21x1_ASAP7_75t_R _2121_ (.A1(net222),
    .A2(_0655_),
    .B(_0679_),
    .Y(_0680_));
 AND3x1_ASAP7_75t_R _2122_ (.A(net260),
    .B(_0658_),
    .C(_0666_),
    .Y(_0681_));
 AO21x1_ASAP7_75t_R _2123_ (.A1(net300),
    .A2(_0616_),
    .B(_0681_),
    .Y(_0682_));
 AND3x1_ASAP7_75t_R _2124_ (.A(net25),
    .B(_0643_),
    .C(_0651_),
    .Y(_0683_));
 AO21x1_ASAP7_75t_R _2125_ (.A1(net65),
    .A2(_0676_),
    .B(_0683_),
    .Y(_0684_));
 OA222x2_ASAP7_75t_R _2126_ (.A1(_0654_),
    .A2(_0680_),
    .B1(_0682_),
    .B2(_0650_),
    .C1(_0684_),
    .C2(_0663_),
    .Y(net381));
 AND3x1_ASAP7_75t_R _2127_ (.A(net261),
    .B(_0995_),
    .C(_0504_),
    .Y(_0685_));
 AND2x2_ASAP7_75t_R _2128_ (.A(net301),
    .B(_0482_),
    .Y(_0686_));
 OR3x1_ASAP7_75t_R _2129_ (.A(_0513_),
    .B(_0685_),
    .C(_0686_),
    .Y(net382));
 AND3x1_ASAP7_75t_R _2130_ (.A(net262),
    .B(_0995_),
    .C(_0504_),
    .Y(_0687_));
 AO21x1_ASAP7_75t_R _2131_ (.A1(net303),
    .A2(_0507_),
    .B(_0687_),
    .Y(_0688_));
 AND3x1_ASAP7_75t_R _2132_ (.A(net184),
    .B(_0995_),
    .C(_0504_),
    .Y(_0689_));
 AO21x1_ASAP7_75t_R _2133_ (.A1(net225),
    .A2(_0507_),
    .B(_0689_),
    .Y(_0690_));
 AO22x1_ASAP7_75t_R _2134_ (.A1(_0495_),
    .A2(_0688_),
    .B1(_0690_),
    .B2(_0489_),
    .Y(net383));
 AND3x1_ASAP7_75t_R _2135_ (.A(net263),
    .B(_0995_),
    .C(_0504_),
    .Y(_0691_));
 AO21x1_ASAP7_75t_R _2136_ (.A1(net304),
    .A2(_0507_),
    .B(_0691_),
    .Y(_0692_));
 AND3x1_ASAP7_75t_R _2137_ (.A(net185),
    .B(_0995_),
    .C(_0504_),
    .Y(_0693_));
 AO21x1_ASAP7_75t_R _2138_ (.A1(net226),
    .A2(_0507_),
    .B(_0693_),
    .Y(_0694_));
 AO22x1_ASAP7_75t_R _2139_ (.A1(_0495_),
    .A2(_0692_),
    .B1(_0694_),
    .B2(_0489_),
    .Y(net384));
 AND3x1_ASAP7_75t_R _2140_ (.A(net264),
    .B(_0995_),
    .C(_0504_),
    .Y(_0695_));
 AO21x1_ASAP7_75t_R _2141_ (.A1(net305),
    .A2(_0507_),
    .B(_0695_),
    .Y(_0696_));
 AND3x1_ASAP7_75t_R _2142_ (.A(net186),
    .B(_0995_),
    .C(_0504_),
    .Y(_0697_));
 AO21x1_ASAP7_75t_R _2143_ (.A1(net227),
    .A2(_0507_),
    .B(_0697_),
    .Y(_0698_));
 AO22x1_ASAP7_75t_R _2144_ (.A1(_0495_),
    .A2(_0696_),
    .B1(_0698_),
    .B2(_0489_),
    .Y(net385));
 AND3x1_ASAP7_75t_R _2145_ (.A(net187),
    .B(_0671_),
    .C(_0509_),
    .Y(_0699_));
 AO21x1_ASAP7_75t_R _2146_ (.A1(net228),
    .A2(_0655_),
    .B(_0699_),
    .Y(_0700_));
 AND3x1_ASAP7_75t_R _2147_ (.A(net265),
    .B(_0658_),
    .C(_0666_),
    .Y(_0701_));
 AO21x1_ASAP7_75t_R _2148_ (.A1(net306),
    .A2(_0514_),
    .B(_0701_),
    .Y(_0702_));
 AND3x1_ASAP7_75t_R _2149_ (.A(net30),
    .B(_0643_),
    .C(_0651_),
    .Y(_0703_));
 AO21x1_ASAP7_75t_R _2150_ (.A1(net71),
    .A2(_0676_),
    .B(_0703_),
    .Y(_0704_));
 OA222x2_ASAP7_75t_R _2151_ (.A1(_0654_),
    .A2(_0700_),
    .B1(_0702_),
    .B2(_0650_),
    .C1(_0704_),
    .C2(_0663_),
    .Y(net386));
 AND3x1_ASAP7_75t_R _2152_ (.A(net191),
    .B(_0671_),
    .C(_0509_),
    .Y(_0705_));
 AO21x1_ASAP7_75t_R _2153_ (.A1(net192),
    .A2(_0655_),
    .B(_0705_),
    .Y(_0706_));
 AND3x1_ASAP7_75t_R _2154_ (.A(net269),
    .B(_0658_),
    .C(_0666_),
    .Y(_0707_));
 AO21x1_ASAP7_75t_R _2155_ (.A1(net270),
    .A2(_0514_),
    .B(_0707_),
    .Y(_0708_));
 AND3x1_ASAP7_75t_R _2156_ (.A(net34),
    .B(_0643_),
    .C(_0651_),
    .Y(_0709_));
 AO21x1_ASAP7_75t_R _2157_ (.A1(net35),
    .A2(_0676_),
    .B(_0709_),
    .Y(_0710_));
 OA222x2_ASAP7_75t_R _2158_ (.A1(_0654_),
    .A2(_0706_),
    .B1(_0708_),
    .B2(_0650_),
    .C1(_0710_),
    .C2(_0663_),
    .Y(net387));
 AND3x1_ASAP7_75t_R _2159_ (.A(net202),
    .B(_0671_),
    .C(_0509_),
    .Y(_0711_));
 AO21x1_ASAP7_75t_R _2160_ (.A1(net193),
    .A2(_0655_),
    .B(_0711_),
    .Y(_0712_));
 AND3x1_ASAP7_75t_R _2161_ (.A(net280),
    .B(_0658_),
    .C(_0666_),
    .Y(_0713_));
 AO21x1_ASAP7_75t_R _2162_ (.A1(net271),
    .A2(_0514_),
    .B(_0713_),
    .Y(_0714_));
 AND3x1_ASAP7_75t_R _2163_ (.A(net45),
    .B(_0643_),
    .C(_0651_),
    .Y(_0715_));
 AO21x1_ASAP7_75t_R _2164_ (.A1(net36),
    .A2(_0676_),
    .B(_0715_),
    .Y(_0716_));
 OA222x2_ASAP7_75t_R _2165_ (.A1(_0654_),
    .A2(_0712_),
    .B1(_0714_),
    .B2(_0650_),
    .C1(_0716_),
    .C2(_0663_),
    .Y(net388));
 AND3x1_ASAP7_75t_R _2166_ (.A(net213),
    .B(_0671_),
    .C(_0509_),
    .Y(_0717_));
 AO21x1_ASAP7_75t_R _2167_ (.A1(net194),
    .A2(_0655_),
    .B(_0717_),
    .Y(_0718_));
 AND3x1_ASAP7_75t_R _2168_ (.A(net291),
    .B(_0658_),
    .C(_0666_),
    .Y(_0719_));
 AO21x1_ASAP7_75t_R _2169_ (.A1(net272),
    .A2(_0514_),
    .B(_0719_),
    .Y(_0720_));
 AND3x1_ASAP7_75t_R _2170_ (.A(net56),
    .B(_0643_),
    .C(_0651_),
    .Y(_0721_));
 AO21x1_ASAP7_75t_R _2171_ (.A1(net37),
    .A2(_0676_),
    .B(_0721_),
    .Y(_0722_));
 OA222x2_ASAP7_75t_R _2172_ (.A1(_0654_),
    .A2(_0718_),
    .B1(_0720_),
    .B2(_0650_),
    .C1(_0722_),
    .C2(_0663_),
    .Y(net389));
 AND3x1_ASAP7_75t_R _2173_ (.A(net224),
    .B(_0671_),
    .C(_0509_),
    .Y(_0723_));
 AO21x1_ASAP7_75t_R _2174_ (.A1(net195),
    .A2(_0655_),
    .B(_0723_),
    .Y(_0724_));
 AND3x1_ASAP7_75t_R _2175_ (.A(net302),
    .B(_0658_),
    .C(_0666_),
    .Y(_0725_));
 AO21x1_ASAP7_75t_R _2176_ (.A1(net273),
    .A2(_0514_),
    .B(_0725_),
    .Y(_0726_));
 AND3x1_ASAP7_75t_R _2177_ (.A(net67),
    .B(_0994_),
    .C(_0651_),
    .Y(_0727_));
 AO21x1_ASAP7_75t_R _2178_ (.A1(net38),
    .A2(_0676_),
    .B(_0727_),
    .Y(_0728_));
 OA222x2_ASAP7_75t_R _2179_ (.A1(_0654_),
    .A2(_0724_),
    .B1(_0726_),
    .B2(_0650_),
    .C1(_0728_),
    .C2(_0663_),
    .Y(net390));
 AND3x1_ASAP7_75t_R _2180_ (.A(net229),
    .B(_0671_),
    .C(_0509_),
    .Y(_0729_));
 AO21x1_ASAP7_75t_R _2181_ (.A1(net196),
    .A2(_0655_),
    .B(_0729_),
    .Y(_0730_));
 AND3x1_ASAP7_75t_R _2182_ (.A(net307),
    .B(_0658_),
    .C(_0666_),
    .Y(_0731_));
 AO21x1_ASAP7_75t_R _2183_ (.A1(net274),
    .A2(_0514_),
    .B(_0731_),
    .Y(_0732_));
 AND3x1_ASAP7_75t_R _2184_ (.A(net72),
    .B(_0994_),
    .C(_0479_),
    .Y(_0733_));
 AO21x1_ASAP7_75t_R _2185_ (.A1(net39),
    .A2(_0676_),
    .B(_0733_),
    .Y(_0734_));
 OA222x2_ASAP7_75t_R _2186_ (.A1(_0654_),
    .A2(_0730_),
    .B1(_0732_),
    .B2(_0512_),
    .C1(_0734_),
    .C2(_0663_),
    .Y(net391));
 AND3x1_ASAP7_75t_R _2187_ (.A(net230),
    .B(_0671_),
    .C(_0509_),
    .Y(_0735_));
 AO21x1_ASAP7_75t_R _2188_ (.A1(net197),
    .A2(_0502_),
    .B(_0735_),
    .Y(_0736_));
 AND3x1_ASAP7_75t_R _2189_ (.A(net308),
    .B(_0515_),
    .C(_0666_),
    .Y(_0737_));
 AO21x1_ASAP7_75t_R _2190_ (.A1(net275),
    .A2(_0514_),
    .B(_0737_),
    .Y(_0738_));
 AND3x1_ASAP7_75t_R _2191_ (.A(net73),
    .B(_0994_),
    .C(_0479_),
    .Y(_0739_));
 AO21x1_ASAP7_75t_R _2192_ (.A1(net40),
    .A2(_0676_),
    .B(_0739_),
    .Y(_0740_));
 OA222x2_ASAP7_75t_R _2193_ (.A1(_0498_),
    .A2(_0736_),
    .B1(_0738_),
    .B2(_0512_),
    .C1(_0740_),
    .C2(_0486_),
    .Y(net392));
 AND3x1_ASAP7_75t_R _2194_ (.A(net231),
    .B(_0671_),
    .C(_0509_),
    .Y(_0741_));
 AO21x1_ASAP7_75t_R _2195_ (.A1(net198),
    .A2(_0502_),
    .B(_0741_),
    .Y(_0742_));
 AND3x1_ASAP7_75t_R _2196_ (.A(net309),
    .B(_0515_),
    .C(_0516_),
    .Y(_0743_));
 AO21x1_ASAP7_75t_R _2197_ (.A1(net276),
    .A2(_0514_),
    .B(_0743_),
    .Y(_0744_));
 AND3x1_ASAP7_75t_R _2198_ (.A(net74),
    .B(_0994_),
    .C(_0479_),
    .Y(_0745_));
 AO21x1_ASAP7_75t_R _2199_ (.A1(net41),
    .A2(_0676_),
    .B(_0745_),
    .Y(_0746_));
 OA222x2_ASAP7_75t_R _2200_ (.A1(_0498_),
    .A2(_0742_),
    .B1(_0744_),
    .B2(_0512_),
    .C1(_0746_),
    .C2(_0486_),
    .Y(net393));
 BUFx6f_ASAP7_75t_R _2201_ (.A(_1153_),
    .Y(_0747_));
 BUFx6f_ASAP7_75t_R _2202_ (.A(_0747_),
    .Y(_0748_));
 BUFx6f_ASAP7_75t_R _2203_ (.A(_1041_),
    .Y(_0749_));
 BUFx6f_ASAP7_75t_R _2204_ (.A(_0749_),
    .Y(_0750_));
 AND2x2_ASAP7_75t_R _2205_ (.A(net31),
    .B(_0750_),
    .Y(_0751_));
 AO21x1_ASAP7_75t_R _2206_ (.A1(net79),
    .A2(_0748_),
    .B(_0751_),
    .Y(_0752_));
 AND2x2_ASAP7_75t_R _2207_ (.A(net1),
    .B(net435),
    .Y(_0753_));
 AO21x1_ASAP7_75t_R _2208_ (.A1(_1179_),
    .A2(_0752_),
    .B(_0753_),
    .Y(net398));
 AND2x2_ASAP7_75t_R _2209_ (.A(net42),
    .B(_0750_),
    .Y(_0754_));
 AO21x1_ASAP7_75t_R _2210_ (.A1(net80),
    .A2(_0748_),
    .B(_0754_),
    .Y(_0755_));
 AND2x2_ASAP7_75t_R _2211_ (.A(net2),
    .B(net435),
    .Y(_0756_));
 AO21x1_ASAP7_75t_R _2212_ (.A1(_1179_),
    .A2(_0755_),
    .B(_0756_),
    .Y(net399));
 AND2x2_ASAP7_75t_R _2213_ (.A(net43),
    .B(_0750_),
    .Y(_0757_));
 AO21x1_ASAP7_75t_R _2214_ (.A1(net81),
    .A2(_0748_),
    .B(_0757_),
    .Y(_0758_));
 AND2x2_ASAP7_75t_R _2215_ (.A(net3),
    .B(net435),
    .Y(_0759_));
 AO21x1_ASAP7_75t_R _2216_ (.A1(_1179_),
    .A2(_0758_),
    .B(_0759_),
    .Y(net400));
 AND2x2_ASAP7_75t_R _2217_ (.A(net44),
    .B(_0750_),
    .Y(_0760_));
 AO21x1_ASAP7_75t_R _2218_ (.A1(net82),
    .A2(_0748_),
    .B(_0760_),
    .Y(_0761_));
 AND2x2_ASAP7_75t_R _2219_ (.A(net4),
    .B(net435),
    .Y(_0762_));
 AO21x1_ASAP7_75t_R _2220_ (.A1(_1179_),
    .A2(_0761_),
    .B(_0762_),
    .Y(net401));
 AND2x2_ASAP7_75t_R _2221_ (.A(net46),
    .B(_0750_),
    .Y(_0763_));
 AO21x1_ASAP7_75t_R _2222_ (.A1(net83),
    .A2(_0748_),
    .B(_0763_),
    .Y(_0764_));
 AND2x2_ASAP7_75t_R _2223_ (.A(net5),
    .B(net435),
    .Y(_0765_));
 AO21x1_ASAP7_75t_R _2224_ (.A1(_1179_),
    .A2(_0764_),
    .B(_0765_),
    .Y(net402));
 AND2x2_ASAP7_75t_R _2225_ (.A(net47),
    .B(_0750_),
    .Y(_0766_));
 AO21x1_ASAP7_75t_R _2226_ (.A1(net84),
    .A2(_0748_),
    .B(_0766_),
    .Y(_0767_));
 AND2x2_ASAP7_75t_R _2227_ (.A(net6),
    .B(net435),
    .Y(_0768_));
 AO21x1_ASAP7_75t_R _2228_ (.A1(_1179_),
    .A2(_0767_),
    .B(_0768_),
    .Y(net403));
 AND2x2_ASAP7_75t_R _2229_ (.A(net48),
    .B(_0750_),
    .Y(_0769_));
 AO21x1_ASAP7_75t_R _2230_ (.A1(net85),
    .A2(_0748_),
    .B(_0769_),
    .Y(_0770_));
 AND2x2_ASAP7_75t_R _2231_ (.A(net7),
    .B(net435),
    .Y(_0771_));
 AO21x1_ASAP7_75t_R _2232_ (.A1(_1179_),
    .A2(_0770_),
    .B(_0771_),
    .Y(net404));
 AND2x2_ASAP7_75t_R _2233_ (.A(net49),
    .B(_0750_),
    .Y(_0772_));
 AO21x1_ASAP7_75t_R _2234_ (.A1(net86),
    .A2(_0748_),
    .B(_0772_),
    .Y(_0773_));
 AND2x2_ASAP7_75t_R _2235_ (.A(net8),
    .B(net435),
    .Y(_0774_));
 AO21x1_ASAP7_75t_R _2236_ (.A1(_1179_),
    .A2(_0773_),
    .B(_0774_),
    .Y(net405));
 AND2x2_ASAP7_75t_R _2237_ (.A(net50),
    .B(_0750_),
    .Y(_0775_));
 AO21x1_ASAP7_75t_R _2238_ (.A1(net87),
    .A2(_0748_),
    .B(_0775_),
    .Y(_0776_));
 AND2x2_ASAP7_75t_R _2239_ (.A(net9),
    .B(net435),
    .Y(_0777_));
 AO21x1_ASAP7_75t_R _2240_ (.A1(_1179_),
    .A2(_0776_),
    .B(_0777_),
    .Y(net406));
 BUFx6f_ASAP7_75t_R _2241_ (.A(_0989_),
    .Y(_0778_));
 BUFx6f_ASAP7_75t_R _2242_ (.A(_0778_),
    .Y(_0779_));
 AND2x2_ASAP7_75t_R _2243_ (.A(net51),
    .B(_0750_),
    .Y(_0780_));
 AO21x1_ASAP7_75t_R _2244_ (.A1(net88),
    .A2(_0748_),
    .B(_0780_),
    .Y(_0781_));
 BUFx6f_ASAP7_75t_R _2245_ (.A(_0990_),
    .Y(_0782_));
 BUFx6f_ASAP7_75t_R _2246_ (.A(_0782_),
    .Y(_0783_));
 AND2x2_ASAP7_75t_R _2247_ (.A(net10),
    .B(_0783_),
    .Y(_0784_));
 AO21x1_ASAP7_75t_R _2248_ (.A1(_0779_),
    .A2(_0781_),
    .B(_0784_),
    .Y(net407));
 BUFx6f_ASAP7_75t_R _2249_ (.A(_0747_),
    .Y(_0785_));
 BUFx6f_ASAP7_75t_R _2250_ (.A(_0749_),
    .Y(_0786_));
 AND2x2_ASAP7_75t_R _2251_ (.A(net52),
    .B(_0786_),
    .Y(_0787_));
 AO21x1_ASAP7_75t_R _2252_ (.A1(net89),
    .A2(_0785_),
    .B(_0787_),
    .Y(_0788_));
 AND2x2_ASAP7_75t_R _2253_ (.A(net11),
    .B(_0783_),
    .Y(_0789_));
 AO21x1_ASAP7_75t_R _2254_ (.A1(_0779_),
    .A2(_0788_),
    .B(_0789_),
    .Y(net408));
 AND2x2_ASAP7_75t_R _2255_ (.A(net32),
    .B(_0786_),
    .Y(_0790_));
 AO21x1_ASAP7_75t_R _2256_ (.A1(net90),
    .A2(_0785_),
    .B(_0790_),
    .Y(_0791_));
 AND2x2_ASAP7_75t_R _2257_ (.A(net12),
    .B(_0783_),
    .Y(_0792_));
 AO21x1_ASAP7_75t_R _2258_ (.A1(_0779_),
    .A2(_0791_),
    .B(_0792_),
    .Y(net409));
 AND2x2_ASAP7_75t_R _2259_ (.A(net53),
    .B(_0786_),
    .Y(_0793_));
 AO21x1_ASAP7_75t_R _2260_ (.A1(net91),
    .A2(_0785_),
    .B(_0793_),
    .Y(_0794_));
 AND2x2_ASAP7_75t_R _2261_ (.A(net13),
    .B(_0783_),
    .Y(_0795_));
 AO21x1_ASAP7_75t_R _2262_ (.A1(_0779_),
    .A2(_0794_),
    .B(_0795_),
    .Y(net410));
 AND2x2_ASAP7_75t_R _2263_ (.A(net54),
    .B(_0786_),
    .Y(_0796_));
 AO21x1_ASAP7_75t_R _2264_ (.A1(net92),
    .A2(_0785_),
    .B(_0796_),
    .Y(_0797_));
 AND2x2_ASAP7_75t_R _2265_ (.A(net14),
    .B(_0783_),
    .Y(_0798_));
 AO21x1_ASAP7_75t_R _2266_ (.A1(_0779_),
    .A2(_0797_),
    .B(_0798_),
    .Y(net411));
 AND2x2_ASAP7_75t_R _2267_ (.A(net55),
    .B(_0786_),
    .Y(_0799_));
 AO21x1_ASAP7_75t_R _2268_ (.A1(net93),
    .A2(_0785_),
    .B(_0799_),
    .Y(_0800_));
 AND2x2_ASAP7_75t_R _2269_ (.A(net15),
    .B(_0783_),
    .Y(_0801_));
 AO21x1_ASAP7_75t_R _2270_ (.A1(_0779_),
    .A2(_0800_),
    .B(_0801_),
    .Y(net412));
 AND2x2_ASAP7_75t_R _2271_ (.A(net57),
    .B(_0786_),
    .Y(_0802_));
 AO21x1_ASAP7_75t_R _2272_ (.A1(net94),
    .A2(_0785_),
    .B(_0802_),
    .Y(_0803_));
 AND2x2_ASAP7_75t_R _2273_ (.A(net16),
    .B(_0783_),
    .Y(_0804_));
 AO21x1_ASAP7_75t_R _2274_ (.A1(_0779_),
    .A2(_0803_),
    .B(_0804_),
    .Y(net413));
 AND2x2_ASAP7_75t_R _2275_ (.A(net58),
    .B(_0786_),
    .Y(_0805_));
 AO21x1_ASAP7_75t_R _2276_ (.A1(net95),
    .A2(_0785_),
    .B(_0805_),
    .Y(_0806_));
 AND2x2_ASAP7_75t_R _2277_ (.A(net17),
    .B(_0783_),
    .Y(_0807_));
 AO21x1_ASAP7_75t_R _2278_ (.A1(_0779_),
    .A2(_0806_),
    .B(_0807_),
    .Y(net414));
 AND2x2_ASAP7_75t_R _2279_ (.A(net59),
    .B(_0786_),
    .Y(_0808_));
 AO21x1_ASAP7_75t_R _2280_ (.A1(net96),
    .A2(_0785_),
    .B(_0808_),
    .Y(_0809_));
 AND2x2_ASAP7_75t_R _2281_ (.A(net18),
    .B(_0783_),
    .Y(_0810_));
 AO21x1_ASAP7_75t_R _2282_ (.A1(_0779_),
    .A2(_0809_),
    .B(_0810_),
    .Y(net415));
 AND2x2_ASAP7_75t_R _2283_ (.A(net60),
    .B(_0786_),
    .Y(_0811_));
 AO21x1_ASAP7_75t_R _2284_ (.A1(net97),
    .A2(_0785_),
    .B(_0811_),
    .Y(_0812_));
 AND2x2_ASAP7_75t_R _2285_ (.A(net19),
    .B(_0783_),
    .Y(_0813_));
 AO21x1_ASAP7_75t_R _2286_ (.A1(_0779_),
    .A2(_0812_),
    .B(_0813_),
    .Y(net416));
 BUFx6f_ASAP7_75t_R _2287_ (.A(_0778_),
    .Y(_0814_));
 AND2x2_ASAP7_75t_R _2288_ (.A(net61),
    .B(_0786_),
    .Y(_0815_));
 AO21x1_ASAP7_75t_R _2289_ (.A1(net98),
    .A2(_0785_),
    .B(_0815_),
    .Y(_0816_));
 BUFx6f_ASAP7_75t_R _2290_ (.A(_0782_),
    .Y(_0817_));
 AND2x2_ASAP7_75t_R _2291_ (.A(net20),
    .B(_0817_),
    .Y(_0818_));
 AO21x1_ASAP7_75t_R _2292_ (.A1(_0814_),
    .A2(_0816_),
    .B(_0818_),
    .Y(net417));
 BUFx6f_ASAP7_75t_R _2293_ (.A(_0747_),
    .Y(_0819_));
 BUFx6f_ASAP7_75t_R _2294_ (.A(_0749_),
    .Y(_0820_));
 AND2x2_ASAP7_75t_R _2295_ (.A(net62),
    .B(_0820_),
    .Y(_0821_));
 AO21x1_ASAP7_75t_R _2296_ (.A1(net99),
    .A2(_0819_),
    .B(_0821_),
    .Y(_0822_));
 AND2x2_ASAP7_75t_R _2297_ (.A(net21),
    .B(_0817_),
    .Y(_0823_));
 AO21x1_ASAP7_75t_R _2298_ (.A1(_0814_),
    .A2(_0822_),
    .B(_0823_),
    .Y(net418));
 AND2x2_ASAP7_75t_R _2299_ (.A(net63),
    .B(_0820_),
    .Y(_0824_));
 AO21x1_ASAP7_75t_R _2300_ (.A1(net100),
    .A2(_0819_),
    .B(_0824_),
    .Y(_0825_));
 AND2x2_ASAP7_75t_R _2301_ (.A(net22),
    .B(_0817_),
    .Y(_0826_));
 AO21x1_ASAP7_75t_R _2302_ (.A1(_0814_),
    .A2(_0825_),
    .B(_0826_),
    .Y(net419));
 AND2x2_ASAP7_75t_R _2303_ (.A(net33),
    .B(_0820_),
    .Y(_0827_));
 AO21x1_ASAP7_75t_R _2304_ (.A1(net101),
    .A2(_0819_),
    .B(_0827_),
    .Y(_0828_));
 AND2x2_ASAP7_75t_R _2305_ (.A(net23),
    .B(_0817_),
    .Y(_0829_));
 AO21x1_ASAP7_75t_R _2306_ (.A1(_0814_),
    .A2(_0828_),
    .B(_0829_),
    .Y(net420));
 AND2x2_ASAP7_75t_R _2307_ (.A(net64),
    .B(_0820_),
    .Y(_0830_));
 AO21x1_ASAP7_75t_R _2308_ (.A1(net102),
    .A2(_0819_),
    .B(_0830_),
    .Y(_0831_));
 AND2x2_ASAP7_75t_R _2309_ (.A(net24),
    .B(_0817_),
    .Y(_0832_));
 AO21x1_ASAP7_75t_R _2310_ (.A1(_0814_),
    .A2(_0831_),
    .B(_0832_),
    .Y(net421));
 AND2x2_ASAP7_75t_R _2311_ (.A(net65),
    .B(_0820_),
    .Y(_0833_));
 AO21x1_ASAP7_75t_R _2312_ (.A1(net103),
    .A2(_0819_),
    .B(_0833_),
    .Y(_0834_));
 AND2x2_ASAP7_75t_R _2313_ (.A(net25),
    .B(_0817_),
    .Y(_0835_));
 AO21x1_ASAP7_75t_R _2314_ (.A1(_0814_),
    .A2(_0834_),
    .B(_0835_),
    .Y(net422));
 AND2x2_ASAP7_75t_R _2315_ (.A(net66),
    .B(_0820_),
    .Y(_0836_));
 AO21x1_ASAP7_75t_R _2316_ (.A1(net104),
    .A2(_0819_),
    .B(_0836_),
    .Y(_0837_));
 AND2x2_ASAP7_75t_R _2317_ (.A(net26),
    .B(_0817_),
    .Y(_0838_));
 AO21x1_ASAP7_75t_R _2318_ (.A1(_0814_),
    .A2(_0837_),
    .B(_0838_),
    .Y(net423));
 AND2x2_ASAP7_75t_R _2319_ (.A(net68),
    .B(_0820_),
    .Y(_0839_));
 AO21x1_ASAP7_75t_R _2320_ (.A1(net105),
    .A2(_0819_),
    .B(_0839_),
    .Y(_0840_));
 AND2x2_ASAP7_75t_R _2321_ (.A(net27),
    .B(_0817_),
    .Y(_0841_));
 AO21x1_ASAP7_75t_R _2322_ (.A1(_0814_),
    .A2(_0840_),
    .B(_0841_),
    .Y(net424));
 AND2x2_ASAP7_75t_R _2323_ (.A(net69),
    .B(_0820_),
    .Y(_0842_));
 AO21x1_ASAP7_75t_R _2324_ (.A1(net106),
    .A2(_0819_),
    .B(_0842_),
    .Y(_0843_));
 AND2x2_ASAP7_75t_R _2325_ (.A(net28),
    .B(_0817_),
    .Y(_0844_));
 AO21x1_ASAP7_75t_R _2326_ (.A1(_0814_),
    .A2(_0843_),
    .B(_0844_),
    .Y(net425));
 AND2x2_ASAP7_75t_R _2327_ (.A(net70),
    .B(_0820_),
    .Y(_0845_));
 AO21x1_ASAP7_75t_R _2328_ (.A1(net107),
    .A2(_0819_),
    .B(_0845_),
    .Y(_0846_));
 AND2x2_ASAP7_75t_R _2329_ (.A(net29),
    .B(_0817_),
    .Y(_0847_));
 AO21x1_ASAP7_75t_R _2330_ (.A1(_0814_),
    .A2(_0846_),
    .B(_0847_),
    .Y(net426));
 AND2x2_ASAP7_75t_R _2331_ (.A(net71),
    .B(_0820_),
    .Y(_0848_));
 AO21x1_ASAP7_75t_R _2332_ (.A1(net108),
    .A2(_0819_),
    .B(_0848_),
    .Y(_0849_));
 AND2x2_ASAP7_75t_R _2333_ (.A(net30),
    .B(_0782_),
    .Y(_0850_));
 AO21x1_ASAP7_75t_R _2334_ (.A1(_0778_),
    .A2(_0849_),
    .B(_0850_),
    .Y(net427));
 AND2x2_ASAP7_75t_R _2335_ (.A(net35),
    .B(_0749_),
    .Y(_0851_));
 AO21x1_ASAP7_75t_R _2336_ (.A1(net112),
    .A2(_0747_),
    .B(_0851_),
    .Y(_0852_));
 AND2x2_ASAP7_75t_R _2337_ (.A(net34),
    .B(_0782_),
    .Y(_0853_));
 AO21x1_ASAP7_75t_R _2338_ (.A1(_0778_),
    .A2(_0852_),
    .B(_0853_),
    .Y(net428));
 AND2x2_ASAP7_75t_R _2339_ (.A(net36),
    .B(_0749_),
    .Y(_0854_));
 AO21x1_ASAP7_75t_R _2340_ (.A1(net123),
    .A2(_0747_),
    .B(_0854_),
    .Y(_0855_));
 AND2x2_ASAP7_75t_R _2341_ (.A(net45),
    .B(_0782_),
    .Y(_0856_));
 AO21x1_ASAP7_75t_R _2342_ (.A1(_0778_),
    .A2(_0855_),
    .B(_0856_),
    .Y(net429));
 AND2x2_ASAP7_75t_R _2343_ (.A(net37),
    .B(_0749_),
    .Y(_0857_));
 AO21x1_ASAP7_75t_R _2344_ (.A1(net134),
    .A2(_0747_),
    .B(_0857_),
    .Y(_0858_));
 AND2x2_ASAP7_75t_R _2345_ (.A(net56),
    .B(_0782_),
    .Y(_0859_));
 AO21x1_ASAP7_75t_R _2346_ (.A1(_0778_),
    .A2(_0858_),
    .B(_0859_),
    .Y(net430));
 AND2x2_ASAP7_75t_R _2347_ (.A(net38),
    .B(_0749_),
    .Y(_0860_));
 AO21x1_ASAP7_75t_R _2348_ (.A1(net145),
    .A2(_0747_),
    .B(_0860_),
    .Y(_0861_));
 AND2x2_ASAP7_75t_R _2349_ (.A(net67),
    .B(_0782_),
    .Y(_0862_));
 AO21x1_ASAP7_75t_R _2350_ (.A1(_0778_),
    .A2(_0861_),
    .B(_0862_),
    .Y(net431));
 AND2x2_ASAP7_75t_R _2351_ (.A(net39),
    .B(_0749_),
    .Y(_0863_));
 AO21x1_ASAP7_75t_R _2352_ (.A1(net150),
    .A2(_0747_),
    .B(_0863_),
    .Y(_0864_));
 AND2x2_ASAP7_75t_R _2353_ (.A(net72),
    .B(_0782_),
    .Y(_0865_));
 AO21x1_ASAP7_75t_R _2354_ (.A1(_0778_),
    .A2(_0864_),
    .B(_0865_),
    .Y(net432));
 AND2x2_ASAP7_75t_R _2355_ (.A(net40),
    .B(_0749_),
    .Y(_0866_));
 AO21x1_ASAP7_75t_R _2356_ (.A1(net151),
    .A2(_0747_),
    .B(_0866_),
    .Y(_0867_));
 AND2x2_ASAP7_75t_R _2357_ (.A(net73),
    .B(_0782_),
    .Y(_0868_));
 AO21x1_ASAP7_75t_R _2358_ (.A1(_0778_),
    .A2(_0867_),
    .B(_0868_),
    .Y(net433));
 AND2x2_ASAP7_75t_R _2359_ (.A(net41),
    .B(_0749_),
    .Y(_0869_));
 AO21x1_ASAP7_75t_R _2360_ (.A1(net152),
    .A2(_0747_),
    .B(_0869_),
    .Y(_0870_));
 AND2x2_ASAP7_75t_R _2361_ (.A(net74),
    .B(_0782_),
    .Y(_0871_));
 AO21x1_ASAP7_75t_R _2362_ (.A1(_0778_),
    .A2(_0870_),
    .B(_0871_),
    .Y(net434));
 BUFx6f_ASAP7_75t_R _2363_ (.A(_1038_),
    .Y(_0872_));
 AND2x2_ASAP7_75t_R _2364_ (.A(net79),
    .B(_0872_),
    .Y(_0873_));
 AO21x1_ASAP7_75t_R _2365_ (.A1(net109),
    .A2(net477),
    .B(_0873_),
    .Y(net439));
 BUFx6f_ASAP7_75t_R _2366_ (.A(_0872_),
    .Y(_0874_));
 AND2x2_ASAP7_75t_R _2367_ (.A(net120),
    .B(net477),
    .Y(_0875_));
 AO21x1_ASAP7_75t_R _2368_ (.A1(net80),
    .A2(_0874_),
    .B(_0875_),
    .Y(net440));
 AND2x2_ASAP7_75t_R _2369_ (.A(net121),
    .B(net477),
    .Y(_0876_));
 AO21x1_ASAP7_75t_R _2370_ (.A1(net81),
    .A2(_0874_),
    .B(_0876_),
    .Y(net441));
 AND2x2_ASAP7_75t_R _2371_ (.A(net122),
    .B(net477),
    .Y(_0877_));
 AO21x1_ASAP7_75t_R _2372_ (.A1(net82),
    .A2(_0874_),
    .B(_0877_),
    .Y(net442));
 AND2x2_ASAP7_75t_R _2373_ (.A(net124),
    .B(net477),
    .Y(_0878_));
 AO21x1_ASAP7_75t_R _2374_ (.A1(net83),
    .A2(_0874_),
    .B(_0878_),
    .Y(net443));
 AND2x2_ASAP7_75t_R _2375_ (.A(net125),
    .B(net477),
    .Y(_0879_));
 AO21x1_ASAP7_75t_R _2376_ (.A1(net84),
    .A2(_0874_),
    .B(_0879_),
    .Y(net444));
 AND2x2_ASAP7_75t_R _2377_ (.A(net126),
    .B(net477),
    .Y(_0880_));
 AO21x1_ASAP7_75t_R _2378_ (.A1(net85),
    .A2(_0874_),
    .B(_0880_),
    .Y(net445));
 AND2x2_ASAP7_75t_R _2379_ (.A(net127),
    .B(net477),
    .Y(_0881_));
 AO21x1_ASAP7_75t_R _2380_ (.A1(net86),
    .A2(_0874_),
    .B(_0881_),
    .Y(net446));
 AND2x2_ASAP7_75t_R _2381_ (.A(net128),
    .B(net477),
    .Y(_0882_));
 AO21x1_ASAP7_75t_R _2382_ (.A1(net87),
    .A2(_0874_),
    .B(_0882_),
    .Y(net447));
 BUFx6f_ASAP7_75t_R _2383_ (.A(_1039_),
    .Y(_0883_));
 BUFx6f_ASAP7_75t_R _2384_ (.A(_0883_),
    .Y(_0884_));
 AND2x2_ASAP7_75t_R _2385_ (.A(net129),
    .B(_0884_),
    .Y(_0885_));
 AO21x1_ASAP7_75t_R _2386_ (.A1(net88),
    .A2(_0874_),
    .B(_0885_),
    .Y(net448));
 AND2x2_ASAP7_75t_R _2387_ (.A(net130),
    .B(_0884_),
    .Y(_0886_));
 AO21x1_ASAP7_75t_R _2388_ (.A1(net89),
    .A2(_0874_),
    .B(_0886_),
    .Y(net449));
 BUFx6f_ASAP7_75t_R _2389_ (.A(_0872_),
    .Y(_0887_));
 AND2x2_ASAP7_75t_R _2390_ (.A(net110),
    .B(_0884_),
    .Y(_0888_));
 AO21x1_ASAP7_75t_R _2391_ (.A1(net90),
    .A2(_0887_),
    .B(_0888_),
    .Y(net450));
 AND2x2_ASAP7_75t_R _2392_ (.A(net131),
    .B(_0884_),
    .Y(_0889_));
 AO21x1_ASAP7_75t_R _2393_ (.A1(net91),
    .A2(_0887_),
    .B(_0889_),
    .Y(net451));
 AND2x2_ASAP7_75t_R _2394_ (.A(net132),
    .B(_0884_),
    .Y(_0890_));
 AO21x1_ASAP7_75t_R _2395_ (.A1(net92),
    .A2(_0887_),
    .B(_0890_),
    .Y(net452));
 AND2x2_ASAP7_75t_R _2396_ (.A(net133),
    .B(_0884_),
    .Y(_0891_));
 AO21x1_ASAP7_75t_R _2397_ (.A1(net93),
    .A2(_0887_),
    .B(_0891_),
    .Y(net453));
 AND2x2_ASAP7_75t_R _2398_ (.A(net135),
    .B(_0884_),
    .Y(_0892_));
 AO21x1_ASAP7_75t_R _2399_ (.A1(net94),
    .A2(_0887_),
    .B(_0892_),
    .Y(net454));
 AND2x2_ASAP7_75t_R _2400_ (.A(net136),
    .B(_0884_),
    .Y(_0893_));
 AO21x1_ASAP7_75t_R _2401_ (.A1(net95),
    .A2(_0887_),
    .B(_0893_),
    .Y(net455));
 AND2x2_ASAP7_75t_R _2402_ (.A(net137),
    .B(_0884_),
    .Y(_0894_));
 AO21x1_ASAP7_75t_R _2403_ (.A1(net96),
    .A2(_0887_),
    .B(_0894_),
    .Y(net456));
 AND2x2_ASAP7_75t_R _2404_ (.A(net138),
    .B(_0884_),
    .Y(_0895_));
 AO21x1_ASAP7_75t_R _2405_ (.A1(net97),
    .A2(_0887_),
    .B(_0895_),
    .Y(net457));
 BUFx6f_ASAP7_75t_R _2406_ (.A(_0883_),
    .Y(_0896_));
 AND2x2_ASAP7_75t_R _2407_ (.A(net139),
    .B(_0896_),
    .Y(_0897_));
 AO21x1_ASAP7_75t_R _2408_ (.A1(net98),
    .A2(_0887_),
    .B(_0897_),
    .Y(net458));
 AND2x2_ASAP7_75t_R _2409_ (.A(net140),
    .B(_0896_),
    .Y(_0898_));
 AO21x1_ASAP7_75t_R _2410_ (.A1(net99),
    .A2(_0887_),
    .B(_0898_),
    .Y(net459));
 BUFx6f_ASAP7_75t_R _2411_ (.A(_0872_),
    .Y(_0899_));
 AND2x2_ASAP7_75t_R _2412_ (.A(net141),
    .B(_0896_),
    .Y(_0900_));
 AO21x1_ASAP7_75t_R _2413_ (.A1(net100),
    .A2(_0899_),
    .B(_0900_),
    .Y(net460));
 AND2x2_ASAP7_75t_R _2414_ (.A(net111),
    .B(_0896_),
    .Y(_0901_));
 AO21x1_ASAP7_75t_R _2415_ (.A1(net101),
    .A2(_0899_),
    .B(_0901_),
    .Y(net461));
 AND2x2_ASAP7_75t_R _2416_ (.A(net142),
    .B(_0896_),
    .Y(_0902_));
 AO21x1_ASAP7_75t_R _2417_ (.A1(net102),
    .A2(_0899_),
    .B(_0902_),
    .Y(net462));
 AND2x2_ASAP7_75t_R _2418_ (.A(net143),
    .B(_0896_),
    .Y(_0903_));
 AO21x1_ASAP7_75t_R _2419_ (.A1(net103),
    .A2(_0899_),
    .B(_0903_),
    .Y(net463));
 AND2x2_ASAP7_75t_R _2420_ (.A(net144),
    .B(_0896_),
    .Y(_0904_));
 AO21x1_ASAP7_75t_R _2421_ (.A1(net104),
    .A2(_0899_),
    .B(_0904_),
    .Y(net464));
 AND2x2_ASAP7_75t_R _2422_ (.A(net146),
    .B(_0896_),
    .Y(_0905_));
 AO21x1_ASAP7_75t_R _2423_ (.A1(net105),
    .A2(_0899_),
    .B(_0905_),
    .Y(net465));
 AND2x2_ASAP7_75t_R _2424_ (.A(net147),
    .B(_0896_),
    .Y(_0906_));
 AO21x1_ASAP7_75t_R _2425_ (.A1(net106),
    .A2(_0899_),
    .B(_0906_),
    .Y(net466));
 AND2x2_ASAP7_75t_R _2426_ (.A(net148),
    .B(_0896_),
    .Y(_0907_));
 AO21x1_ASAP7_75t_R _2427_ (.A1(net107),
    .A2(_0899_),
    .B(_0907_),
    .Y(net467));
 AND2x2_ASAP7_75t_R _2428_ (.A(net149),
    .B(_0883_),
    .Y(_0908_));
 AO21x1_ASAP7_75t_R _2429_ (.A1(net108),
    .A2(_0899_),
    .B(_0908_),
    .Y(net468));
 AND2x2_ASAP7_75t_R _2430_ (.A(net113),
    .B(_0883_),
    .Y(_0909_));
 AO21x1_ASAP7_75t_R _2431_ (.A1(net112),
    .A2(_0899_),
    .B(_0909_),
    .Y(net469));
 AND2x2_ASAP7_75t_R _2432_ (.A(net114),
    .B(_0883_),
    .Y(_0910_));
 AO21x1_ASAP7_75t_R _2433_ (.A1(net123),
    .A2(_0872_),
    .B(_0910_),
    .Y(net470));
 AND2x2_ASAP7_75t_R _2434_ (.A(net115),
    .B(_0883_),
    .Y(_0911_));
 AO21x1_ASAP7_75t_R _2435_ (.A1(net134),
    .A2(_0872_),
    .B(_0911_),
    .Y(net471));
 AND2x2_ASAP7_75t_R _2436_ (.A(net116),
    .B(_0883_),
    .Y(_0912_));
 AO21x1_ASAP7_75t_R _2437_ (.A1(net145),
    .A2(_0872_),
    .B(_0912_),
    .Y(net472));
 AND2x2_ASAP7_75t_R _2438_ (.A(net117),
    .B(_0883_),
    .Y(_0913_));
 AO21x1_ASAP7_75t_R _2439_ (.A1(net150),
    .A2(_0872_),
    .B(_0913_),
    .Y(net473));
 AND2x2_ASAP7_75t_R _2440_ (.A(net118),
    .B(_0883_),
    .Y(_0914_));
 AO21x1_ASAP7_75t_R _2441_ (.A1(net151),
    .A2(_0872_),
    .B(_0914_),
    .Y(net474));
 AND2x2_ASAP7_75t_R _2442_ (.A(net119),
    .B(_0883_),
    .Y(_0915_));
 AO21x1_ASAP7_75t_R _2443_ (.A1(net152),
    .A2(_0872_),
    .B(_0915_),
    .Y(net475));
 FAx1_ASAP7_75t_R _2444_ (.SN(_0072_),
    .A(_1169_),
    .B(_0071_),
    .CI(_1170_),
    .CON(_0100_));
 FAx1_ASAP7_75t_R _2445_ (.SN(_0101_),
    .A(\credit_pi_route_inst.u1_counters_inst.o_credits[5] ),
    .B(\credit_pi_route_inst.u1_counters_inst.o_credits[6] ),
    .CI(net477),
    .CON(_0013_));
 FAx1_ASAP7_75t_R _2446_ (.SN(_0063_),
    .A(_0062_),
    .B(_1171_),
    .CI(_1172_),
    .CON(_0020_));
 FAx1_ASAP7_75t_R _2447_ (.SN(_0061_),
    .A(_0060_),
    .B(_1173_),
    .CI(_1174_),
    .CON(_0026_));
 FAx1_ASAP7_75t_R _2448_ (.SN(_0067_),
    .A(_0066_),
    .B(_1175_),
    .CI(_1176_),
    .CON(_0033_));
 FAx1_ASAP7_75t_R _2449_ (.SN(_0065_),
    .A(_0064_),
    .B(_1177_),
    .CI(_1178_),
    .CON(_0039_));
 FAx1_ASAP7_75t_R _2450_ (.SN(_0102_),
    .A(\credit_pi_route_inst.u0_counters_inst.o_credits[5] ),
    .B(\credit_pi_route_inst.u0_counters_inst.o_credits[6] ),
    .CI(net436),
    .CON(_0046_));
 FAx1_ASAP7_75t_R _2451_ (.SN(_0069_),
    .A(_1179_),
    .B(_0068_),
    .CI(_1180_),
    .CON(_0103_));
 HAxp5_ASAP7_75t_R _2452_ (.A(net476),
    .B(\credit_pi_route_inst.u1_counters_inst.o_credits[1] ),
    .CON(_0006_),
    .SN(_0004_));
 HAxp5_ASAP7_75t_R _2453_ (.A(net476),
    .B(\credit_pi_route_inst.u1_counters_inst.o_credits[2] ),
    .CON(_0008_),
    .SN(_0005_));
 HAxp5_ASAP7_75t_R _2454_ (.A(net476),
    .B(\credit_pi_route_inst.u1_counters_inst.o_credits[3] ),
    .CON(_0009_),
    .SN(_0007_));
 HAxp5_ASAP7_75t_R _2455_ (.A(\credit_pi_route_inst.u1_counters_inst.o_credits[6] ),
    .B(net477),
    .CON(_0012_),
    .SN(_0010_));
 HAxp5_ASAP7_75t_R _2456_ (.A(\credit_pi_route_inst.u1_counters_inst.o_credits[7] ),
    .B(net477),
    .CON(_0015_),
    .SN(_0011_));
 HAxp5_ASAP7_75t_R _2457_ (.A(\credit_pi_route_inst.u1_counters_inst.o_credits[8] ),
    .B(net477),
    .CON(_0016_),
    .SN(_0014_));
 HAxp5_ASAP7_75t_R _2458_ (.A(\credit_pi_route_inst.l_counters_inst.o_credits[6] ),
    .B(net354),
    .CON(_0019_),
    .SN(_0017_));
 HAxp5_ASAP7_75t_R _2459_ (.A(\credit_pi_route_inst.l_counters_inst.o_credits[7] ),
    .B(net354),
    .CON(_0022_),
    .SN(_0018_));
 HAxp5_ASAP7_75t_R _2460_ (.A(\credit_pi_route_inst.l_counters_inst.o_credits[8] ),
    .B(net354),
    .CON(_0104_),
    .SN(_0021_));
 HAxp5_ASAP7_75t_R _2461_ (.A(\credit_pi_route_inst.l_counters_inst.o_credits[1] ),
    .B(net353),
    .CON(_0025_),
    .SN(_0023_));
 HAxp5_ASAP7_75t_R _2462_ (.A(\credit_pi_route_inst.l_counters_inst.o_credits[2] ),
    .B(net353),
    .CON(_0028_),
    .SN(_0024_));
 HAxp5_ASAP7_75t_R _2463_ (.A(\credit_pi_route_inst.l_counters_inst.o_credits[3] ),
    .B(net353),
    .CON(_0029_),
    .SN(_0027_));
 HAxp5_ASAP7_75t_R _2464_ (.A(\credit_pi_route_inst.r_counters_inst.o_credits[6] ),
    .B(net395),
    .CON(_0032_),
    .SN(_0030_));
 HAxp5_ASAP7_75t_R _2465_ (.A(\credit_pi_route_inst.r_counters_inst.o_credits[7] ),
    .B(net395),
    .CON(_0035_),
    .SN(_0031_));
 HAxp5_ASAP7_75t_R _2466_ (.A(\credit_pi_route_inst.r_counters_inst.o_credits[8] ),
    .B(net395),
    .CON(_0105_),
    .SN(_0034_));
 HAxp5_ASAP7_75t_R _2467_ (.A(\credit_pi_route_inst.r_counters_inst.o_credits[1] ),
    .B(net394),
    .CON(_0038_),
    .SN(_0036_));
 HAxp5_ASAP7_75t_R _2468_ (.A(\credit_pi_route_inst.r_counters_inst.o_credits[2] ),
    .B(net394),
    .CON(_0041_),
    .SN(_0037_));
 HAxp5_ASAP7_75t_R _2469_ (.A(\credit_pi_route_inst.r_counters_inst.o_credits[3] ),
    .B(net394),
    .CON(_0042_),
    .SN(_0040_));
 HAxp5_ASAP7_75t_R _2470_ (.A(\credit_pi_route_inst.u0_counters_inst.o_credits[6] ),
    .B(net436),
    .CON(_0045_),
    .SN(_0043_));
 HAxp5_ASAP7_75t_R _2471_ (.A(\credit_pi_route_inst.u0_counters_inst.o_credits[7] ),
    .B(net436),
    .CON(_0048_),
    .SN(_0044_));
 HAxp5_ASAP7_75t_R _2472_ (.A(\credit_pi_route_inst.u0_counters_inst.o_credits[8] ),
    .B(net436),
    .CON(_0049_),
    .SN(_0047_));
 HAxp5_ASAP7_75t_R _2473_ (.A(net435),
    .B(\credit_pi_route_inst.u0_counters_inst.o_credits[1] ),
    .CON(_0052_),
    .SN(_0050_));
 HAxp5_ASAP7_75t_R _2474_ (.A(net435),
    .B(\credit_pi_route_inst.u0_counters_inst.o_credits[2] ),
    .CON(_0054_),
    .SN(_0051_));
 HAxp5_ASAP7_75t_R _2475_ (.A(net435),
    .B(\credit_pi_route_inst.u0_counters_inst.o_credits[3] ),
    .CON(_0055_),
    .SN(_0053_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.l_counters_inst.o_credits[0]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0106_),
    .QN(_0060_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.l_counters_inst.o_credits[1]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0107_),
    .QN(_1173_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.l_counters_inst.o_credits[2]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0108_),
    .QN(_0096_));
 DFFHQNx1_ASAP7_75t_R \credit_pi_route_inst.l_counters_inst.o_credits[3]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0109_),
    .QN(_0095_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.l_counters_inst.o_credits[4]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0110_),
    .QN(_0094_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.l_counters_inst.o_credits[5]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0111_),
    .QN(_0062_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.l_counters_inst.o_credits[6]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0112_),
    .QN(_1171_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.l_counters_inst.o_credits[7]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0113_),
    .QN(_0093_));
 DFFHQNx1_ASAP7_75t_R \credit_pi_route_inst.l_counters_inst.o_credits[8]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0114_),
    .QN(_0092_));
 DFFHQNx1_ASAP7_75t_R \credit_pi_route_inst.l_counters_inst.o_credits[9]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0115_),
    .QN(_0091_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.r_counters_inst.o_credits[0]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0116_),
    .QN(_0064_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.r_counters_inst.o_credits[1]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0117_),
    .QN(_1177_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.r_counters_inst.o_credits[2]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0118_),
    .QN(_0090_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.r_counters_inst.o_credits[3]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0119_),
    .QN(_0089_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.r_counters_inst.o_credits[4]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0120_),
    .QN(_0088_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.r_counters_inst.o_credits[5]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0121_),
    .QN(_0066_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.r_counters_inst.o_credits[6]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0122_),
    .QN(_1175_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.r_counters_inst.o_credits[7]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0123_),
    .QN(_0087_));
 DFFHQNx1_ASAP7_75t_R \credit_pi_route_inst.r_counters_inst.o_credits[8]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0124_),
    .QN(_0086_));
 DFFHQNx1_ASAP7_75t_R \credit_pi_route_inst.r_counters_inst.o_credits[9]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0125_),
    .QN(_0097_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.state[0]$_DFF_P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0000_),
    .QN(_0098_));
 DFFHQNx1_ASAP7_75t_R \credit_pi_route_inst.state[1]$_DFF_P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0001_),
    .QN(_0056_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.state[2]$_DFF_P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0002_),
    .QN(_0099_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.state[3]$_DFF_P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0003_),
    .QN(_0057_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u0_counters_inst.o_credits[0]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0126_),
    .QN(_0068_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u0_counters_inst.o_credits[1]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0127_),
    .QN(_1180_));
 DFFHQNx1_ASAP7_75t_R \credit_pi_route_inst.u0_counters_inst.o_credits[2]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0128_),
    .QN(_0085_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u0_counters_inst.o_credits[3]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0129_),
    .QN(_0084_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u0_counters_inst.o_credits[4]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0130_),
    .QN(_0058_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u0_counters_inst.o_credits[5]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0131_),
    .QN(_0070_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u0_counters_inst.o_credits[6]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0132_),
    .QN(_0083_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u0_counters_inst.o_credits[7]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0133_),
    .QN(_0082_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u0_counters_inst.o_credits[8]$_SDFFE_PP1P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_0134_),
    .QN(_0081_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u0_counters_inst.o_credits[9]$_SDFFE_PP1P_  (.CLK(clknet_2_2__leaf_clk),
    .D(_0135_),
    .QN(_0080_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u1_counters_inst.o_credits[0]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0136_),
    .QN(_0071_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u1_counters_inst.o_credits[1]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0137_),
    .QN(_1170_));
 DFFHQNx1_ASAP7_75t_R \credit_pi_route_inst.u1_counters_inst.o_credits[2]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0138_),
    .QN(_0079_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u1_counters_inst.o_credits[3]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0139_),
    .QN(_0078_));
 DFFHQNx1_ASAP7_75t_R \credit_pi_route_inst.u1_counters_inst.o_credits[4]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0140_),
    .QN(_0059_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u1_counters_inst.o_credits[5]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0141_),
    .QN(_0073_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u1_counters_inst.o_credits[6]$_SDFFE_PP1P_  (.CLK(clknet_2_0__leaf_clk),
    .D(_0142_),
    .QN(_0077_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u1_counters_inst.o_credits[7]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0143_),
    .QN(_0076_));
 DFFHQNx3_ASAP7_75t_R \credit_pi_route_inst.u1_counters_inst.o_credits[8]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0144_),
    .QN(_0075_));
 DFFHQNx1_ASAP7_75t_R \credit_pi_route_inst.u1_counters_inst.o_credits[9]$_SDFFE_PP1P_  (.CLK(clknet_2_1__leaf_clk),
    .D(_0145_),
    .QN(_0074_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Left_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Left_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Left_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Left_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Left_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Left_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Left_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Left_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Left_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Left_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Left_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Left_133 ();
 BUFx3_ASAP7_75t_R input1 (.A(l_i[0]),
    .Y(net1));
 BUFx3_ASAP7_75t_R input2 (.A(l_i[10]),
    .Y(net2));
 BUFx3_ASAP7_75t_R input3 (.A(l_i[11]),
    .Y(net3));
 BUFx3_ASAP7_75t_R input4 (.A(l_i[12]),
    .Y(net4));
 BUFx3_ASAP7_75t_R input5 (.A(l_i[13]),
    .Y(net5));
 BUFx3_ASAP7_75t_R input6 (.A(l_i[14]),
    .Y(net6));
 BUFx3_ASAP7_75t_R input7 (.A(l_i[15]),
    .Y(net7));
 BUFx3_ASAP7_75t_R input8 (.A(l_i[16]),
    .Y(net8));
 BUFx3_ASAP7_75t_R input9 (.A(l_i[17]),
    .Y(net9));
 BUFx3_ASAP7_75t_R input10 (.A(l_i[18]),
    .Y(net10));
 BUFx3_ASAP7_75t_R input11 (.A(l_i[19]),
    .Y(net11));
 BUFx3_ASAP7_75t_R input12 (.A(l_i[1]),
    .Y(net12));
 BUFx3_ASAP7_75t_R input13 (.A(l_i[20]),
    .Y(net13));
 BUFx3_ASAP7_75t_R input14 (.A(l_i[21]),
    .Y(net14));
 BUFx3_ASAP7_75t_R input15 (.A(l_i[22]),
    .Y(net15));
 BUFx3_ASAP7_75t_R input16 (.A(l_i[23]),
    .Y(net16));
 BUFx3_ASAP7_75t_R input17 (.A(l_i[24]),
    .Y(net17));
 BUFx3_ASAP7_75t_R input18 (.A(l_i[25]),
    .Y(net18));
 BUFx3_ASAP7_75t_R input19 (.A(l_i[26]),
    .Y(net19));
 BUFx3_ASAP7_75t_R input20 (.A(l_i[27]),
    .Y(net20));
 BUFx3_ASAP7_75t_R input21 (.A(l_i[28]),
    .Y(net21));
 BUFx3_ASAP7_75t_R input22 (.A(l_i[29]),
    .Y(net22));
 BUFx3_ASAP7_75t_R input23 (.A(l_i[2]),
    .Y(net23));
 BUFx3_ASAP7_75t_R input24 (.A(l_i[30]),
    .Y(net24));
 BUFx3_ASAP7_75t_R input25 (.A(l_i[31]),
    .Y(net25));
 BUFx3_ASAP7_75t_R input26 (.A(l_i[32]),
    .Y(net26));
 BUFx3_ASAP7_75t_R input27 (.A(l_i[33]),
    .Y(net27));
 BUFx3_ASAP7_75t_R input28 (.A(l_i[34]),
    .Y(net28));
 BUFx3_ASAP7_75t_R input29 (.A(l_i[35]),
    .Y(net29));
 BUFx3_ASAP7_75t_R input30 (.A(l_i[36]),
    .Y(net30));
 BUFx3_ASAP7_75t_R input31 (.A(l_i[37]),
    .Y(net31));
 BUFx3_ASAP7_75t_R input32 (.A(l_i[38]),
    .Y(net32));
 BUFx3_ASAP7_75t_R input33 (.A(l_i[39]),
    .Y(net33));
 BUFx3_ASAP7_75t_R input34 (.A(l_i[3]),
    .Y(net34));
 BUFx3_ASAP7_75t_R input35 (.A(l_i[40]),
    .Y(net35));
 BUFx3_ASAP7_75t_R input36 (.A(l_i[41]),
    .Y(net36));
 BUFx3_ASAP7_75t_R input37 (.A(l_i[42]),
    .Y(net37));
 BUFx3_ASAP7_75t_R input38 (.A(l_i[43]),
    .Y(net38));
 BUFx3_ASAP7_75t_R input39 (.A(l_i[44]),
    .Y(net39));
 BUFx3_ASAP7_75t_R input40 (.A(l_i[45]),
    .Y(net40));
 BUFx3_ASAP7_75t_R input41 (.A(l_i[46]),
    .Y(net41));
 BUFx3_ASAP7_75t_R input42 (.A(l_i[47]),
    .Y(net42));
 BUFx3_ASAP7_75t_R input43 (.A(l_i[48]),
    .Y(net43));
 BUFx3_ASAP7_75t_R input44 (.A(l_i[49]),
    .Y(net44));
 BUFx3_ASAP7_75t_R input45 (.A(l_i[4]),
    .Y(net45));
 BUFx3_ASAP7_75t_R input46 (.A(l_i[50]),
    .Y(net46));
 BUFx3_ASAP7_75t_R input47 (.A(l_i[51]),
    .Y(net47));
 BUFx3_ASAP7_75t_R input48 (.A(l_i[52]),
    .Y(net48));
 BUFx3_ASAP7_75t_R input49 (.A(l_i[53]),
    .Y(net49));
 BUFx3_ASAP7_75t_R input50 (.A(l_i[54]),
    .Y(net50));
 BUFx3_ASAP7_75t_R input51 (.A(l_i[55]),
    .Y(net51));
 BUFx3_ASAP7_75t_R input52 (.A(l_i[56]),
    .Y(net52));
 BUFx3_ASAP7_75t_R input53 (.A(l_i[57]),
    .Y(net53));
 BUFx3_ASAP7_75t_R input54 (.A(l_i[58]),
    .Y(net54));
 BUFx3_ASAP7_75t_R input55 (.A(l_i[59]),
    .Y(net55));
 BUFx3_ASAP7_75t_R input56 (.A(l_i[5]),
    .Y(net56));
 BUFx3_ASAP7_75t_R input57 (.A(l_i[60]),
    .Y(net57));
 BUFx3_ASAP7_75t_R input58 (.A(l_i[61]),
    .Y(net58));
 BUFx3_ASAP7_75t_R input59 (.A(l_i[62]),
    .Y(net59));
 BUFx3_ASAP7_75t_R input60 (.A(l_i[63]),
    .Y(net60));
 BUFx3_ASAP7_75t_R input61 (.A(l_i[64]),
    .Y(net61));
 BUFx3_ASAP7_75t_R input62 (.A(l_i[65]),
    .Y(net62));
 BUFx3_ASAP7_75t_R input63 (.A(l_i[66]),
    .Y(net63));
 BUFx3_ASAP7_75t_R input64 (.A(l_i[67]),
    .Y(net64));
 BUFx3_ASAP7_75t_R input65 (.A(l_i[68]),
    .Y(net65));
 BUFx3_ASAP7_75t_R input66 (.A(l_i[69]),
    .Y(net66));
 BUFx3_ASAP7_75t_R input67 (.A(l_i[6]),
    .Y(net67));
 BUFx3_ASAP7_75t_R input68 (.A(l_i[70]),
    .Y(net68));
 BUFx3_ASAP7_75t_R input69 (.A(l_i[71]),
    .Y(net69));
 BUFx3_ASAP7_75t_R input70 (.A(l_i[72]),
    .Y(net70));
 BUFx3_ASAP7_75t_R input71 (.A(l_i[73]),
    .Y(net71));
 BUFx3_ASAP7_75t_R input72 (.A(l_i[7]),
    .Y(net72));
 BUFx3_ASAP7_75t_R input73 (.A(l_i[8]),
    .Y(net73));
 BUFx3_ASAP7_75t_R input74 (.A(l_i[9]),
    .Y(net74));
 BUFx3_ASAP7_75t_R input75 (.A(l_i_v[0]),
    .Y(net75));
 BUFx3_ASAP7_75t_R input76 (.A(l_i_v[1]),
    .Y(net76));
 BUFx3_ASAP7_75t_R input77 (.A(l_o_credit_gnt[0]),
    .Y(net77));
 BUFx3_ASAP7_75t_R input78 (.A(l_o_credit_gnt[1]),
    .Y(net78));
 BUFx3_ASAP7_75t_R input79 (.A(r_i[0]),
    .Y(net79));
 BUFx3_ASAP7_75t_R input80 (.A(r_i[10]),
    .Y(net80));
 BUFx3_ASAP7_75t_R input81 (.A(r_i[11]),
    .Y(net81));
 BUFx3_ASAP7_75t_R input82 (.A(r_i[12]),
    .Y(net82));
 BUFx3_ASAP7_75t_R input83 (.A(r_i[13]),
    .Y(net83));
 BUFx3_ASAP7_75t_R input84 (.A(r_i[14]),
    .Y(net84));
 BUFx3_ASAP7_75t_R input85 (.A(r_i[15]),
    .Y(net85));
 BUFx3_ASAP7_75t_R input86 (.A(r_i[16]),
    .Y(net86));
 BUFx3_ASAP7_75t_R input87 (.A(r_i[17]),
    .Y(net87));
 BUFx3_ASAP7_75t_R input88 (.A(r_i[18]),
    .Y(net88));
 BUFx3_ASAP7_75t_R input89 (.A(r_i[19]),
    .Y(net89));
 BUFx3_ASAP7_75t_R input90 (.A(r_i[1]),
    .Y(net90));
 BUFx3_ASAP7_75t_R input91 (.A(r_i[20]),
    .Y(net91));
 BUFx3_ASAP7_75t_R input92 (.A(r_i[21]),
    .Y(net92));
 BUFx3_ASAP7_75t_R input93 (.A(r_i[22]),
    .Y(net93));
 BUFx3_ASAP7_75t_R input94 (.A(r_i[23]),
    .Y(net94));
 BUFx3_ASAP7_75t_R input95 (.A(r_i[24]),
    .Y(net95));
 BUFx3_ASAP7_75t_R input96 (.A(r_i[25]),
    .Y(net96));
 BUFx3_ASAP7_75t_R input97 (.A(r_i[26]),
    .Y(net97));
 BUFx3_ASAP7_75t_R input98 (.A(r_i[27]),
    .Y(net98));
 BUFx3_ASAP7_75t_R input99 (.A(r_i[28]),
    .Y(net99));
 BUFx3_ASAP7_75t_R input100 (.A(r_i[29]),
    .Y(net100));
 BUFx3_ASAP7_75t_R input101 (.A(r_i[2]),
    .Y(net101));
 BUFx3_ASAP7_75t_R input102 (.A(r_i[30]),
    .Y(net102));
 BUFx3_ASAP7_75t_R input103 (.A(r_i[31]),
    .Y(net103));
 BUFx3_ASAP7_75t_R input104 (.A(r_i[32]),
    .Y(net104));
 BUFx3_ASAP7_75t_R input105 (.A(r_i[33]),
    .Y(net105));
 BUFx3_ASAP7_75t_R input106 (.A(r_i[34]),
    .Y(net106));
 BUFx3_ASAP7_75t_R input107 (.A(r_i[35]),
    .Y(net107));
 BUFx3_ASAP7_75t_R input108 (.A(r_i[36]),
    .Y(net108));
 BUFx3_ASAP7_75t_R input109 (.A(r_i[37]),
    .Y(net109));
 BUFx3_ASAP7_75t_R input110 (.A(r_i[38]),
    .Y(net110));
 BUFx3_ASAP7_75t_R input111 (.A(r_i[39]),
    .Y(net111));
 BUFx3_ASAP7_75t_R input112 (.A(r_i[3]),
    .Y(net112));
 BUFx3_ASAP7_75t_R input113 (.A(r_i[40]),
    .Y(net113));
 BUFx3_ASAP7_75t_R input114 (.A(r_i[41]),
    .Y(net114));
 BUFx3_ASAP7_75t_R input115 (.A(r_i[42]),
    .Y(net115));
 BUFx3_ASAP7_75t_R input116 (.A(r_i[43]),
    .Y(net116));
 BUFx3_ASAP7_75t_R input117 (.A(r_i[44]),
    .Y(net117));
 BUFx3_ASAP7_75t_R input118 (.A(r_i[45]),
    .Y(net118));
 BUFx3_ASAP7_75t_R input119 (.A(r_i[46]),
    .Y(net119));
 BUFx3_ASAP7_75t_R input120 (.A(r_i[47]),
    .Y(net120));
 BUFx3_ASAP7_75t_R input121 (.A(r_i[48]),
    .Y(net121));
 BUFx3_ASAP7_75t_R input122 (.A(r_i[49]),
    .Y(net122));
 BUFx3_ASAP7_75t_R input123 (.A(r_i[4]),
    .Y(net123));
 BUFx3_ASAP7_75t_R input124 (.A(r_i[50]),
    .Y(net124));
 BUFx3_ASAP7_75t_R input125 (.A(r_i[51]),
    .Y(net125));
 BUFx3_ASAP7_75t_R input126 (.A(r_i[52]),
    .Y(net126));
 BUFx3_ASAP7_75t_R input127 (.A(r_i[53]),
    .Y(net127));
 BUFx3_ASAP7_75t_R input128 (.A(r_i[54]),
    .Y(net128));
 BUFx3_ASAP7_75t_R input129 (.A(r_i[55]),
    .Y(net129));
 BUFx3_ASAP7_75t_R input130 (.A(r_i[56]),
    .Y(net130));
 BUFx3_ASAP7_75t_R input131 (.A(r_i[57]),
    .Y(net131));
 BUFx3_ASAP7_75t_R input132 (.A(r_i[58]),
    .Y(net132));
 BUFx3_ASAP7_75t_R input133 (.A(r_i[59]),
    .Y(net133));
 BUFx3_ASAP7_75t_R input134 (.A(r_i[5]),
    .Y(net134));
 BUFx3_ASAP7_75t_R input135 (.A(r_i[60]),
    .Y(net135));
 BUFx3_ASAP7_75t_R input136 (.A(r_i[61]),
    .Y(net136));
 BUFx3_ASAP7_75t_R input137 (.A(r_i[62]),
    .Y(net137));
 BUFx3_ASAP7_75t_R input138 (.A(r_i[63]),
    .Y(net138));
 BUFx3_ASAP7_75t_R input139 (.A(r_i[64]),
    .Y(net139));
 BUFx3_ASAP7_75t_R input140 (.A(r_i[65]),
    .Y(net140));
 BUFx3_ASAP7_75t_R input141 (.A(r_i[66]),
    .Y(net141));
 BUFx3_ASAP7_75t_R input142 (.A(r_i[67]),
    .Y(net142));
 BUFx3_ASAP7_75t_R input143 (.A(r_i[68]),
    .Y(net143));
 BUFx3_ASAP7_75t_R input144 (.A(r_i[69]),
    .Y(net144));
 BUFx3_ASAP7_75t_R input145 (.A(r_i[6]),
    .Y(net145));
 BUFx3_ASAP7_75t_R input146 (.A(r_i[70]),
    .Y(net146));
 BUFx3_ASAP7_75t_R input147 (.A(r_i[71]),
    .Y(net147));
 BUFx3_ASAP7_75t_R input148 (.A(r_i[72]),
    .Y(net148));
 BUFx3_ASAP7_75t_R input149 (.A(r_i[73]),
    .Y(net149));
 BUFx3_ASAP7_75t_R input150 (.A(r_i[7]),
    .Y(net150));
 BUFx3_ASAP7_75t_R input151 (.A(r_i[8]),
    .Y(net151));
 BUFx3_ASAP7_75t_R input152 (.A(r_i[9]),
    .Y(net152));
 BUFx3_ASAP7_75t_R input153 (.A(r_i_v[0]),
    .Y(net153));
 BUFx3_ASAP7_75t_R input154 (.A(r_i_v[1]),
    .Y(net154));
 BUFx3_ASAP7_75t_R input155 (.A(r_o_credit_gnt[0]),
    .Y(net155));
 BUFx3_ASAP7_75t_R input156 (.A(r_o_credit_gnt[1]),
    .Y(net156));
 BUFx6f_ASAP7_75t_R input157 (.A(rst),
    .Y(net157));
 BUFx3_ASAP7_75t_R input158 (.A(u0_i[0]),
    .Y(net158));
 BUFx3_ASAP7_75t_R input159 (.A(u0_i[10]),
    .Y(net159));
 BUFx3_ASAP7_75t_R input160 (.A(u0_i[11]),
    .Y(net160));
 BUFx3_ASAP7_75t_R input161 (.A(u0_i[12]),
    .Y(net161));
 BUFx3_ASAP7_75t_R input162 (.A(u0_i[13]),
    .Y(net162));
 BUFx3_ASAP7_75t_R input163 (.A(u0_i[14]),
    .Y(net163));
 BUFx3_ASAP7_75t_R input164 (.A(u0_i[15]),
    .Y(net164));
 BUFx3_ASAP7_75t_R input165 (.A(u0_i[16]),
    .Y(net165));
 BUFx3_ASAP7_75t_R input166 (.A(u0_i[17]),
    .Y(net166));
 BUFx3_ASAP7_75t_R input167 (.A(u0_i[18]),
    .Y(net167));
 BUFx3_ASAP7_75t_R input168 (.A(u0_i[19]),
    .Y(net168));
 BUFx3_ASAP7_75t_R input169 (.A(u0_i[1]),
    .Y(net169));
 BUFx3_ASAP7_75t_R input170 (.A(u0_i[20]),
    .Y(net170));
 BUFx3_ASAP7_75t_R input171 (.A(u0_i[21]),
    .Y(net171));
 BUFx3_ASAP7_75t_R input172 (.A(u0_i[22]),
    .Y(net172));
 BUFx3_ASAP7_75t_R input173 (.A(u0_i[23]),
    .Y(net173));
 BUFx3_ASAP7_75t_R input174 (.A(u0_i[24]),
    .Y(net174));
 BUFx3_ASAP7_75t_R input175 (.A(u0_i[25]),
    .Y(net175));
 BUFx3_ASAP7_75t_R input176 (.A(u0_i[26]),
    .Y(net176));
 BUFx3_ASAP7_75t_R input177 (.A(u0_i[27]),
    .Y(net177));
 BUFx3_ASAP7_75t_R input178 (.A(u0_i[28]),
    .Y(net178));
 BUFx3_ASAP7_75t_R input179 (.A(u0_i[29]),
    .Y(net179));
 BUFx3_ASAP7_75t_R input180 (.A(u0_i[2]),
    .Y(net180));
 BUFx3_ASAP7_75t_R input181 (.A(u0_i[30]),
    .Y(net181));
 BUFx3_ASAP7_75t_R input182 (.A(u0_i[31]),
    .Y(net182));
 BUFx3_ASAP7_75t_R input183 (.A(u0_i[32]),
    .Y(net183));
 BUFx3_ASAP7_75t_R input184 (.A(u0_i[33]),
    .Y(net184));
 BUFx3_ASAP7_75t_R input185 (.A(u0_i[34]),
    .Y(net185));
 BUFx3_ASAP7_75t_R input186 (.A(u0_i[35]),
    .Y(net186));
 BUFx3_ASAP7_75t_R input187 (.A(u0_i[36]),
    .Y(net187));
 BUFx3_ASAP7_75t_R input188 (.A(u0_i[37]),
    .Y(net188));
 BUFx3_ASAP7_75t_R input189 (.A(u0_i[38]),
    .Y(net189));
 BUFx3_ASAP7_75t_R input190 (.A(u0_i[39]),
    .Y(net190));
 BUFx3_ASAP7_75t_R input191 (.A(u0_i[3]),
    .Y(net191));
 BUFx3_ASAP7_75t_R input192 (.A(u0_i[40]),
    .Y(net192));
 BUFx3_ASAP7_75t_R input193 (.A(u0_i[41]),
    .Y(net193));
 BUFx3_ASAP7_75t_R input194 (.A(u0_i[42]),
    .Y(net194));
 BUFx3_ASAP7_75t_R input195 (.A(u0_i[43]),
    .Y(net195));
 BUFx3_ASAP7_75t_R input196 (.A(u0_i[44]),
    .Y(net196));
 BUFx3_ASAP7_75t_R input197 (.A(u0_i[45]),
    .Y(net197));
 BUFx3_ASAP7_75t_R input198 (.A(u0_i[46]),
    .Y(net198));
 BUFx3_ASAP7_75t_R input199 (.A(u0_i[47]),
    .Y(net199));
 BUFx3_ASAP7_75t_R input200 (.A(u0_i[48]),
    .Y(net200));
 BUFx3_ASAP7_75t_R input201 (.A(u0_i[49]),
    .Y(net201));
 BUFx3_ASAP7_75t_R input202 (.A(u0_i[4]),
    .Y(net202));
 BUFx3_ASAP7_75t_R input203 (.A(u0_i[50]),
    .Y(net203));
 BUFx3_ASAP7_75t_R input204 (.A(u0_i[51]),
    .Y(net204));
 BUFx3_ASAP7_75t_R input205 (.A(u0_i[52]),
    .Y(net205));
 BUFx3_ASAP7_75t_R input206 (.A(u0_i[53]),
    .Y(net206));
 BUFx3_ASAP7_75t_R input207 (.A(u0_i[54]),
    .Y(net207));
 BUFx3_ASAP7_75t_R input208 (.A(u0_i[55]),
    .Y(net208));
 BUFx3_ASAP7_75t_R input209 (.A(u0_i[56]),
    .Y(net209));
 BUFx3_ASAP7_75t_R input210 (.A(u0_i[57]),
    .Y(net210));
 BUFx3_ASAP7_75t_R input211 (.A(u0_i[58]),
    .Y(net211));
 BUFx3_ASAP7_75t_R input212 (.A(u0_i[59]),
    .Y(net212));
 BUFx3_ASAP7_75t_R input213 (.A(u0_i[5]),
    .Y(net213));
 BUFx3_ASAP7_75t_R input214 (.A(u0_i[60]),
    .Y(net214));
 BUFx3_ASAP7_75t_R input215 (.A(u0_i[61]),
    .Y(net215));
 BUFx3_ASAP7_75t_R input216 (.A(u0_i[62]),
    .Y(net216));
 BUFx3_ASAP7_75t_R input217 (.A(u0_i[63]),
    .Y(net217));
 BUFx3_ASAP7_75t_R input218 (.A(u0_i[64]),
    .Y(net218));
 BUFx3_ASAP7_75t_R input219 (.A(u0_i[65]),
    .Y(net219));
 BUFx3_ASAP7_75t_R input220 (.A(u0_i[66]),
    .Y(net220));
 BUFx3_ASAP7_75t_R input221 (.A(u0_i[67]),
    .Y(net221));
 BUFx3_ASAP7_75t_R input222 (.A(u0_i[68]),
    .Y(net222));
 BUFx3_ASAP7_75t_R input223 (.A(u0_i[69]),
    .Y(net223));
 BUFx3_ASAP7_75t_R input224 (.A(u0_i[6]),
    .Y(net224));
 BUFx3_ASAP7_75t_R input225 (.A(u0_i[70]),
    .Y(net225));
 BUFx3_ASAP7_75t_R input226 (.A(u0_i[71]),
    .Y(net226));
 BUFx3_ASAP7_75t_R input227 (.A(u0_i[72]),
    .Y(net227));
 BUFx3_ASAP7_75t_R input228 (.A(u0_i[73]),
    .Y(net228));
 BUFx3_ASAP7_75t_R input229 (.A(u0_i[7]),
    .Y(net229));
 BUFx3_ASAP7_75t_R input230 (.A(u0_i[8]),
    .Y(net230));
 BUFx3_ASAP7_75t_R input231 (.A(u0_i[9]),
    .Y(net231));
 BUFx3_ASAP7_75t_R input232 (.A(u0_i_v[0]),
    .Y(net232));
 BUFx3_ASAP7_75t_R input233 (.A(u0_i_v[1]),
    .Y(net233));
 BUFx3_ASAP7_75t_R input234 (.A(u0_o_credit_gnt[0]),
    .Y(net234));
 BUFx3_ASAP7_75t_R input235 (.A(u0_o_credit_gnt[1]),
    .Y(net235));
 BUFx3_ASAP7_75t_R input236 (.A(u1_i[0]),
    .Y(net236));
 BUFx3_ASAP7_75t_R input237 (.A(u1_i[10]),
    .Y(net237));
 BUFx3_ASAP7_75t_R input238 (.A(u1_i[11]),
    .Y(net238));
 BUFx3_ASAP7_75t_R input239 (.A(u1_i[12]),
    .Y(net239));
 BUFx3_ASAP7_75t_R input240 (.A(u1_i[13]),
    .Y(net240));
 BUFx3_ASAP7_75t_R input241 (.A(u1_i[14]),
    .Y(net241));
 BUFx3_ASAP7_75t_R input242 (.A(u1_i[15]),
    .Y(net242));
 BUFx3_ASAP7_75t_R input243 (.A(u1_i[16]),
    .Y(net243));
 BUFx3_ASAP7_75t_R input244 (.A(u1_i[17]),
    .Y(net244));
 BUFx3_ASAP7_75t_R input245 (.A(u1_i[18]),
    .Y(net245));
 BUFx3_ASAP7_75t_R input246 (.A(u1_i[19]),
    .Y(net246));
 BUFx3_ASAP7_75t_R input247 (.A(u1_i[1]),
    .Y(net247));
 BUFx3_ASAP7_75t_R input248 (.A(u1_i[20]),
    .Y(net248));
 BUFx3_ASAP7_75t_R input249 (.A(u1_i[21]),
    .Y(net249));
 BUFx3_ASAP7_75t_R input250 (.A(u1_i[22]),
    .Y(net250));
 BUFx3_ASAP7_75t_R input251 (.A(u1_i[23]),
    .Y(net251));
 BUFx3_ASAP7_75t_R input252 (.A(u1_i[24]),
    .Y(net252));
 BUFx3_ASAP7_75t_R input253 (.A(u1_i[25]),
    .Y(net253));
 BUFx3_ASAP7_75t_R input254 (.A(u1_i[26]),
    .Y(net254));
 BUFx3_ASAP7_75t_R input255 (.A(u1_i[27]),
    .Y(net255));
 BUFx3_ASAP7_75t_R input256 (.A(u1_i[28]),
    .Y(net256));
 BUFx3_ASAP7_75t_R input257 (.A(u1_i[29]),
    .Y(net257));
 BUFx3_ASAP7_75t_R input258 (.A(u1_i[2]),
    .Y(net258));
 BUFx3_ASAP7_75t_R input259 (.A(u1_i[30]),
    .Y(net259));
 BUFx3_ASAP7_75t_R input260 (.A(u1_i[31]),
    .Y(net260));
 BUFx3_ASAP7_75t_R input261 (.A(u1_i[32]),
    .Y(net261));
 BUFx3_ASAP7_75t_R input262 (.A(u1_i[33]),
    .Y(net262));
 BUFx3_ASAP7_75t_R input263 (.A(u1_i[34]),
    .Y(net263));
 BUFx3_ASAP7_75t_R input264 (.A(u1_i[35]),
    .Y(net264));
 BUFx3_ASAP7_75t_R input265 (.A(u1_i[36]),
    .Y(net265));
 BUFx3_ASAP7_75t_R input266 (.A(u1_i[37]),
    .Y(net266));
 BUFx3_ASAP7_75t_R input267 (.A(u1_i[38]),
    .Y(net267));
 BUFx3_ASAP7_75t_R input268 (.A(u1_i[39]),
    .Y(net268));
 BUFx3_ASAP7_75t_R input269 (.A(u1_i[3]),
    .Y(net269));
 BUFx3_ASAP7_75t_R input270 (.A(u1_i[40]),
    .Y(net270));
 BUFx3_ASAP7_75t_R input271 (.A(u1_i[41]),
    .Y(net271));
 BUFx3_ASAP7_75t_R input272 (.A(u1_i[42]),
    .Y(net272));
 BUFx3_ASAP7_75t_R input273 (.A(u1_i[43]),
    .Y(net273));
 BUFx3_ASAP7_75t_R input274 (.A(u1_i[44]),
    .Y(net274));
 BUFx3_ASAP7_75t_R input275 (.A(u1_i[45]),
    .Y(net275));
 BUFx3_ASAP7_75t_R input276 (.A(u1_i[46]),
    .Y(net276));
 BUFx3_ASAP7_75t_R input277 (.A(u1_i[47]),
    .Y(net277));
 BUFx3_ASAP7_75t_R input278 (.A(u1_i[48]),
    .Y(net278));
 BUFx3_ASAP7_75t_R input279 (.A(u1_i[49]),
    .Y(net279));
 BUFx3_ASAP7_75t_R input280 (.A(u1_i[4]),
    .Y(net280));
 BUFx3_ASAP7_75t_R input281 (.A(u1_i[50]),
    .Y(net281));
 BUFx3_ASAP7_75t_R input282 (.A(u1_i[51]),
    .Y(net282));
 BUFx3_ASAP7_75t_R input283 (.A(u1_i[52]),
    .Y(net283));
 BUFx3_ASAP7_75t_R input284 (.A(u1_i[53]),
    .Y(net284));
 BUFx3_ASAP7_75t_R input285 (.A(u1_i[54]),
    .Y(net285));
 BUFx3_ASAP7_75t_R input286 (.A(u1_i[55]),
    .Y(net286));
 BUFx3_ASAP7_75t_R input287 (.A(u1_i[56]),
    .Y(net287));
 BUFx3_ASAP7_75t_R input288 (.A(u1_i[57]),
    .Y(net288));
 BUFx3_ASAP7_75t_R input289 (.A(u1_i[58]),
    .Y(net289));
 BUFx3_ASAP7_75t_R input290 (.A(u1_i[59]),
    .Y(net290));
 BUFx3_ASAP7_75t_R input291 (.A(u1_i[5]),
    .Y(net291));
 BUFx3_ASAP7_75t_R input292 (.A(u1_i[60]),
    .Y(net292));
 BUFx3_ASAP7_75t_R input293 (.A(u1_i[61]),
    .Y(net293));
 BUFx3_ASAP7_75t_R input294 (.A(u1_i[62]),
    .Y(net294));
 BUFx3_ASAP7_75t_R input295 (.A(u1_i[63]),
    .Y(net295));
 BUFx3_ASAP7_75t_R input296 (.A(u1_i[64]),
    .Y(net296));
 BUFx3_ASAP7_75t_R input297 (.A(u1_i[65]),
    .Y(net297));
 BUFx3_ASAP7_75t_R input298 (.A(u1_i[66]),
    .Y(net298));
 BUFx3_ASAP7_75t_R input299 (.A(u1_i[67]),
    .Y(net299));
 BUFx3_ASAP7_75t_R input300 (.A(u1_i[68]),
    .Y(net300));
 BUFx3_ASAP7_75t_R input301 (.A(u1_i[69]),
    .Y(net301));
 BUFx3_ASAP7_75t_R input302 (.A(u1_i[6]),
    .Y(net302));
 BUFx3_ASAP7_75t_R input303 (.A(u1_i[70]),
    .Y(net303));
 BUFx3_ASAP7_75t_R input304 (.A(u1_i[71]),
    .Y(net304));
 BUFx3_ASAP7_75t_R input305 (.A(u1_i[72]),
    .Y(net305));
 BUFx3_ASAP7_75t_R input306 (.A(u1_i[73]),
    .Y(net306));
 BUFx3_ASAP7_75t_R input307 (.A(u1_i[7]),
    .Y(net307));
 BUFx3_ASAP7_75t_R input308 (.A(u1_i[8]),
    .Y(net308));
 BUFx3_ASAP7_75t_R input309 (.A(u1_i[9]),
    .Y(net309));
 BUFx3_ASAP7_75t_R input310 (.A(u1_i_v[0]),
    .Y(net310));
 BUFx3_ASAP7_75t_R input311 (.A(u1_i_v[1]),
    .Y(net311));
 BUFx3_ASAP7_75t_R input312 (.A(u1_o_credit_gnt[0]),
    .Y(net312));
 BUFx3_ASAP7_75t_R input313 (.A(u1_o_credit_gnt[1]),
    .Y(net313));
 BUFx3_ASAP7_75t_R output314 (.A(net314),
    .Y(l_i_bp[0]));
 BUFx3_ASAP7_75t_R output315 (.A(net315),
    .Y(l_i_bp[1]));
 BUFx3_ASAP7_75t_R output316 (.A(net316),
    .Y(l_o[0]));
 BUFx3_ASAP7_75t_R output317 (.A(net317),
    .Y(l_o[10]));
 BUFx3_ASAP7_75t_R output318 (.A(net318),
    .Y(l_o[11]));
 BUFx3_ASAP7_75t_R output319 (.A(net319),
    .Y(l_o[12]));
 BUFx3_ASAP7_75t_R output320 (.A(net320),
    .Y(l_o[13]));
 BUFx3_ASAP7_75t_R output321 (.A(net321),
    .Y(l_o[14]));
 BUFx3_ASAP7_75t_R output322 (.A(net322),
    .Y(l_o[15]));
 BUFx3_ASAP7_75t_R output323 (.A(net323),
    .Y(l_o[16]));
 BUFx3_ASAP7_75t_R output324 (.A(net324),
    .Y(l_o[17]));
 BUFx3_ASAP7_75t_R output325 (.A(net325),
    .Y(l_o[18]));
 BUFx3_ASAP7_75t_R output326 (.A(net326),
    .Y(l_o[19]));
 BUFx3_ASAP7_75t_R output327 (.A(net327),
    .Y(l_o[1]));
 BUFx3_ASAP7_75t_R output328 (.A(net328),
    .Y(l_o[20]));
 BUFx3_ASAP7_75t_R output329 (.A(net329),
    .Y(l_o[21]));
 BUFx3_ASAP7_75t_R output330 (.A(net330),
    .Y(l_o[22]));
 BUFx3_ASAP7_75t_R output331 (.A(net331),
    .Y(l_o[23]));
 BUFx3_ASAP7_75t_R output332 (.A(net332),
    .Y(l_o[24]));
 BUFx3_ASAP7_75t_R output333 (.A(net333),
    .Y(l_o[25]));
 BUFx3_ASAP7_75t_R output334 (.A(net334),
    .Y(l_o[26]));
 BUFx3_ASAP7_75t_R output335 (.A(net335),
    .Y(l_o[27]));
 BUFx3_ASAP7_75t_R output336 (.A(net336),
    .Y(l_o[28]));
 BUFx3_ASAP7_75t_R output337 (.A(net337),
    .Y(l_o[29]));
 BUFx3_ASAP7_75t_R output338 (.A(net338),
    .Y(l_o[2]));
 BUFx3_ASAP7_75t_R output339 (.A(net339),
    .Y(l_o[30]));
 BUFx3_ASAP7_75t_R output340 (.A(net340),
    .Y(l_o[31]));
 BUFx3_ASAP7_75t_R output341 (.A(net341),
    .Y(l_o[32]));
 BUFx3_ASAP7_75t_R output342 (.A(net342),
    .Y(l_o[33]));
 BUFx3_ASAP7_75t_R output343 (.A(net343),
    .Y(l_o[34]));
 BUFx3_ASAP7_75t_R output344 (.A(net344),
    .Y(l_o[35]));
 BUFx3_ASAP7_75t_R output345 (.A(net345),
    .Y(l_o[36]));
 BUFx3_ASAP7_75t_R output346 (.A(net346),
    .Y(l_o[3]));
 BUFx3_ASAP7_75t_R output347 (.A(net347),
    .Y(l_o[4]));
 BUFx3_ASAP7_75t_R output348 (.A(net348),
    .Y(l_o[5]));
 BUFx3_ASAP7_75t_R output349 (.A(net349),
    .Y(l_o[6]));
 BUFx3_ASAP7_75t_R output350 (.A(net350),
    .Y(l_o[7]));
 BUFx3_ASAP7_75t_R output351 (.A(net351),
    .Y(l_o[8]));
 BUFx3_ASAP7_75t_R output352 (.A(net352),
    .Y(l_o[9]));
 BUFx3_ASAP7_75t_R output353 (.A(net353),
    .Y(l_o_v[0]));
 BUFx3_ASAP7_75t_R output354 (.A(net354),
    .Y(l_o_v[1]));
 BUFx3_ASAP7_75t_R output355 (.A(net355),
    .Y(r_i_bp[0]));
 BUFx3_ASAP7_75t_R output356 (.A(net356),
    .Y(r_i_bp[1]));
 BUFx3_ASAP7_75t_R output357 (.A(net357),
    .Y(r_o[0]));
 BUFx3_ASAP7_75t_R output358 (.A(net358),
    .Y(r_o[10]));
 BUFx3_ASAP7_75t_R output359 (.A(net359),
    .Y(r_o[11]));
 BUFx3_ASAP7_75t_R output360 (.A(net360),
    .Y(r_o[12]));
 BUFx3_ASAP7_75t_R output361 (.A(net361),
    .Y(r_o[13]));
 BUFx3_ASAP7_75t_R output362 (.A(net362),
    .Y(r_o[14]));
 BUFx3_ASAP7_75t_R output363 (.A(net363),
    .Y(r_o[15]));
 BUFx3_ASAP7_75t_R output364 (.A(net364),
    .Y(r_o[16]));
 BUFx3_ASAP7_75t_R output365 (.A(net365),
    .Y(r_o[17]));
 BUFx3_ASAP7_75t_R output366 (.A(net366),
    .Y(r_o[18]));
 BUFx3_ASAP7_75t_R output367 (.A(net367),
    .Y(r_o[19]));
 BUFx3_ASAP7_75t_R output368 (.A(net368),
    .Y(r_o[1]));
 BUFx3_ASAP7_75t_R output369 (.A(net369),
    .Y(r_o[20]));
 BUFx3_ASAP7_75t_R output370 (.A(net370),
    .Y(r_o[21]));
 BUFx3_ASAP7_75t_R output371 (.A(net371),
    .Y(r_o[22]));
 BUFx3_ASAP7_75t_R output372 (.A(net372),
    .Y(r_o[23]));
 BUFx3_ASAP7_75t_R output373 (.A(net373),
    .Y(r_o[24]));
 BUFx3_ASAP7_75t_R output374 (.A(net374),
    .Y(r_o[25]));
 BUFx3_ASAP7_75t_R output375 (.A(net375),
    .Y(r_o[26]));
 BUFx3_ASAP7_75t_R output376 (.A(net376),
    .Y(r_o[27]));
 BUFx3_ASAP7_75t_R output377 (.A(net377),
    .Y(r_o[28]));
 BUFx3_ASAP7_75t_R output378 (.A(net378),
    .Y(r_o[29]));
 BUFx3_ASAP7_75t_R output379 (.A(net379),
    .Y(r_o[2]));
 BUFx3_ASAP7_75t_R output380 (.A(net380),
    .Y(r_o[30]));
 BUFx3_ASAP7_75t_R output381 (.A(net381),
    .Y(r_o[31]));
 BUFx3_ASAP7_75t_R output382 (.A(net382),
    .Y(r_o[32]));
 BUFx3_ASAP7_75t_R output383 (.A(net383),
    .Y(r_o[33]));
 BUFx3_ASAP7_75t_R output384 (.A(net384),
    .Y(r_o[34]));
 BUFx3_ASAP7_75t_R output385 (.A(net385),
    .Y(r_o[35]));
 BUFx3_ASAP7_75t_R output386 (.A(net386),
    .Y(r_o[36]));
 BUFx3_ASAP7_75t_R output387 (.A(net387),
    .Y(r_o[3]));
 BUFx3_ASAP7_75t_R output388 (.A(net388),
    .Y(r_o[4]));
 BUFx3_ASAP7_75t_R output389 (.A(net389),
    .Y(r_o[5]));
 BUFx3_ASAP7_75t_R output390 (.A(net390),
    .Y(r_o[6]));
 BUFx3_ASAP7_75t_R output391 (.A(net391),
    .Y(r_o[7]));
 BUFx3_ASAP7_75t_R output392 (.A(net392),
    .Y(r_o[8]));
 BUFx3_ASAP7_75t_R output393 (.A(net393),
    .Y(r_o[9]));
 BUFx3_ASAP7_75t_R output394 (.A(net394),
    .Y(r_o_v[0]));
 BUFx3_ASAP7_75t_R output395 (.A(net395),
    .Y(r_o_v[1]));
 BUFx3_ASAP7_75t_R output396 (.A(net396),
    .Y(u0_i_bp[0]));
 BUFx3_ASAP7_75t_R output397 (.A(net397),
    .Y(u0_i_bp[1]));
 BUFx3_ASAP7_75t_R output398 (.A(net398),
    .Y(u0_o[0]));
 BUFx3_ASAP7_75t_R output399 (.A(net399),
    .Y(u0_o[10]));
 BUFx3_ASAP7_75t_R output400 (.A(net400),
    .Y(u0_o[11]));
 BUFx3_ASAP7_75t_R output401 (.A(net401),
    .Y(u0_o[12]));
 BUFx3_ASAP7_75t_R output402 (.A(net402),
    .Y(u0_o[13]));
 BUFx3_ASAP7_75t_R output403 (.A(net403),
    .Y(u0_o[14]));
 BUFx3_ASAP7_75t_R output404 (.A(net404),
    .Y(u0_o[15]));
 BUFx3_ASAP7_75t_R output405 (.A(net405),
    .Y(u0_o[16]));
 BUFx3_ASAP7_75t_R output406 (.A(net406),
    .Y(u0_o[17]));
 BUFx3_ASAP7_75t_R output407 (.A(net407),
    .Y(u0_o[18]));
 BUFx3_ASAP7_75t_R output408 (.A(net408),
    .Y(u0_o[19]));
 BUFx3_ASAP7_75t_R output409 (.A(net409),
    .Y(u0_o[1]));
 BUFx3_ASAP7_75t_R output410 (.A(net410),
    .Y(u0_o[20]));
 BUFx3_ASAP7_75t_R output411 (.A(net411),
    .Y(u0_o[21]));
 BUFx3_ASAP7_75t_R output412 (.A(net412),
    .Y(u0_o[22]));
 BUFx3_ASAP7_75t_R output413 (.A(net413),
    .Y(u0_o[23]));
 BUFx3_ASAP7_75t_R output414 (.A(net414),
    .Y(u0_o[24]));
 BUFx3_ASAP7_75t_R output415 (.A(net415),
    .Y(u0_o[25]));
 BUFx3_ASAP7_75t_R output416 (.A(net416),
    .Y(u0_o[26]));
 BUFx3_ASAP7_75t_R output417 (.A(net417),
    .Y(u0_o[27]));
 BUFx3_ASAP7_75t_R output418 (.A(net418),
    .Y(u0_o[28]));
 BUFx3_ASAP7_75t_R output419 (.A(net419),
    .Y(u0_o[29]));
 BUFx3_ASAP7_75t_R output420 (.A(net420),
    .Y(u0_o[2]));
 BUFx3_ASAP7_75t_R output421 (.A(net421),
    .Y(u0_o[30]));
 BUFx3_ASAP7_75t_R output422 (.A(net422),
    .Y(u0_o[31]));
 BUFx3_ASAP7_75t_R output423 (.A(net423),
    .Y(u0_o[32]));
 BUFx3_ASAP7_75t_R output424 (.A(net424),
    .Y(u0_o[33]));
 BUFx3_ASAP7_75t_R output425 (.A(net425),
    .Y(u0_o[34]));
 BUFx3_ASAP7_75t_R output426 (.A(net426),
    .Y(u0_o[35]));
 BUFx3_ASAP7_75t_R output427 (.A(net427),
    .Y(u0_o[36]));
 BUFx3_ASAP7_75t_R output428 (.A(net428),
    .Y(u0_o[3]));
 BUFx3_ASAP7_75t_R output429 (.A(net429),
    .Y(u0_o[4]));
 BUFx3_ASAP7_75t_R output430 (.A(net430),
    .Y(u0_o[5]));
 BUFx3_ASAP7_75t_R output431 (.A(net431),
    .Y(u0_o[6]));
 BUFx3_ASAP7_75t_R output432 (.A(net432),
    .Y(u0_o[7]));
 BUFx3_ASAP7_75t_R output433 (.A(net433),
    .Y(u0_o[8]));
 BUFx3_ASAP7_75t_R output434 (.A(net434),
    .Y(u0_o[9]));
 BUFx3_ASAP7_75t_R output435 (.A(net435),
    .Y(u0_o_v[0]));
 BUFx3_ASAP7_75t_R output436 (.A(net436),
    .Y(u0_o_v[1]));
 BUFx3_ASAP7_75t_R output437 (.A(net437),
    .Y(u1_i_bp[0]));
 BUFx3_ASAP7_75t_R output438 (.A(net438),
    .Y(u1_i_bp[1]));
 BUFx3_ASAP7_75t_R output439 (.A(net439),
    .Y(u1_o[0]));
 BUFx3_ASAP7_75t_R output440 (.A(net440),
    .Y(u1_o[10]));
 BUFx3_ASAP7_75t_R output441 (.A(net441),
    .Y(u1_o[11]));
 BUFx3_ASAP7_75t_R output442 (.A(net442),
    .Y(u1_o[12]));
 BUFx3_ASAP7_75t_R output443 (.A(net443),
    .Y(u1_o[13]));
 BUFx3_ASAP7_75t_R output444 (.A(net444),
    .Y(u1_o[14]));
 BUFx3_ASAP7_75t_R output445 (.A(net445),
    .Y(u1_o[15]));
 BUFx3_ASAP7_75t_R output446 (.A(net446),
    .Y(u1_o[16]));
 BUFx3_ASAP7_75t_R output447 (.A(net447),
    .Y(u1_o[17]));
 BUFx3_ASAP7_75t_R output448 (.A(net448),
    .Y(u1_o[18]));
 BUFx3_ASAP7_75t_R output449 (.A(net449),
    .Y(u1_o[19]));
 BUFx3_ASAP7_75t_R output450 (.A(net450),
    .Y(u1_o[1]));
 BUFx3_ASAP7_75t_R output451 (.A(net451),
    .Y(u1_o[20]));
 BUFx3_ASAP7_75t_R output452 (.A(net452),
    .Y(u1_o[21]));
 BUFx3_ASAP7_75t_R output453 (.A(net453),
    .Y(u1_o[22]));
 BUFx3_ASAP7_75t_R output454 (.A(net454),
    .Y(u1_o[23]));
 BUFx3_ASAP7_75t_R output455 (.A(net455),
    .Y(u1_o[24]));
 BUFx3_ASAP7_75t_R output456 (.A(net456),
    .Y(u1_o[25]));
 BUFx3_ASAP7_75t_R output457 (.A(net457),
    .Y(u1_o[26]));
 BUFx3_ASAP7_75t_R output458 (.A(net458),
    .Y(u1_o[27]));
 BUFx3_ASAP7_75t_R output459 (.A(net459),
    .Y(u1_o[28]));
 BUFx3_ASAP7_75t_R output460 (.A(net460),
    .Y(u1_o[29]));
 BUFx3_ASAP7_75t_R output461 (.A(net461),
    .Y(u1_o[2]));
 BUFx3_ASAP7_75t_R output462 (.A(net462),
    .Y(u1_o[30]));
 BUFx3_ASAP7_75t_R output463 (.A(net463),
    .Y(u1_o[31]));
 BUFx3_ASAP7_75t_R output464 (.A(net464),
    .Y(u1_o[32]));
 BUFx3_ASAP7_75t_R output465 (.A(net465),
    .Y(u1_o[33]));
 BUFx3_ASAP7_75t_R output466 (.A(net466),
    .Y(u1_o[34]));
 BUFx3_ASAP7_75t_R output467 (.A(net467),
    .Y(u1_o[35]));
 BUFx3_ASAP7_75t_R output468 (.A(net468),
    .Y(u1_o[36]));
 BUFx3_ASAP7_75t_R output469 (.A(net469),
    .Y(u1_o[3]));
 BUFx3_ASAP7_75t_R output470 (.A(net470),
    .Y(u1_o[4]));
 BUFx3_ASAP7_75t_R output471 (.A(net471),
    .Y(u1_o[5]));
 BUFx3_ASAP7_75t_R output472 (.A(net472),
    .Y(u1_o[6]));
 BUFx3_ASAP7_75t_R output473 (.A(net473),
    .Y(u1_o[7]));
 BUFx3_ASAP7_75t_R output474 (.A(net474),
    .Y(u1_o[8]));
 BUFx3_ASAP7_75t_R output475 (.A(net475),
    .Y(u1_o[9]));
 BUFx3_ASAP7_75t_R output476 (.A(net476),
    .Y(u1_o_v[0]));
 BUFx3_ASAP7_75t_R output477 (.A(net477),
    .Y(u1_o_v[1]));
 BUFx4_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_0__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_1__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_2__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_3__leaf_clk));
 BUFx12_ASAP7_75t_R clkload0 (.A(clknet_2_1__leaf_clk));
 BUFx4f_ASAP7_75t_R clkload1 (.A(clknet_2_2__leaf_clk));
 BUFx12_ASAP7_75t_R clkload2 (.A(clknet_2_3__leaf_clk));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 FILLER_ASAP7_75t_R FILLER_0_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_54 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174 ();
 FILLER_ASAP7_75t_R FILLER_0_238 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258 ();
 FILLER_ASAP7_75t_R FILLER_0_264 ();
 DECAPx1_ASAP7_75t_R FILLER_0_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_276 ();
 DECAPx2_ASAP7_75t_R FILLER_0_283 ();
 DECAPx2_ASAP7_75t_R FILLER_0_331 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx2_ASAP7_75t_R FILLER_1_68 ();
 FILLER_ASAP7_75t_R FILLER_1_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_76 ();
 FILLER_ASAP7_75t_R FILLER_1_83 ();
 FILLER_ASAP7_75t_R FILLER_1_88 ();
 FILLER_ASAP7_75t_R FILLER_1_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_113 ();
 FILLER_ASAP7_75t_R FILLER_1_126 ();
 DECAPx2_ASAP7_75t_R FILLER_1_134 ();
 FILLER_ASAP7_75t_R FILLER_1_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_230 ();
 FILLER_ASAP7_75t_R FILLER_1_243 ();
 DECAPx10_ASAP7_75t_R FILLER_1_257 ();
 DECAPx10_ASAP7_75t_R FILLER_1_279 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx6_ASAP7_75t_R FILLER_2_46 ();
 FILLER_ASAP7_75t_R FILLER_2_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_62 ();
 FILLER_ASAP7_75t_R FILLER_2_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_117 ();
 DECAPx2_ASAP7_75t_R FILLER_2_136 ();
 FILLER_ASAP7_75t_R FILLER_2_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_157 ();
 FILLER_ASAP7_75t_R FILLER_2_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_166 ();
 DECAPx2_ASAP7_75t_R FILLER_2_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_197 ();
 DECAPx2_ASAP7_75t_R FILLER_2_204 ();
 FILLER_ASAP7_75t_R FILLER_2_210 ();
 FILLER_ASAP7_75t_R FILLER_2_218 ();
 DECAPx2_ASAP7_75t_R FILLER_2_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_244 ();
 DECAPx10_ASAP7_75t_R FILLER_2_251 ();
 DECAPx4_ASAP7_75t_R FILLER_2_273 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx1_ASAP7_75t_R FILLER_3_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_90 ();
 FILLER_ASAP7_75t_R FILLER_3_116 ();
 DECAPx2_ASAP7_75t_R FILLER_3_140 ();
 FILLER_ASAP7_75t_R FILLER_3_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_167 ();
 DECAPx2_ASAP7_75t_R FILLER_3_174 ();
 DECAPx1_ASAP7_75t_R FILLER_3_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_196 ();
 DECAPx6_ASAP7_75t_R FILLER_3_203 ();
 DECAPx2_ASAP7_75t_R FILLER_3_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_223 ();
 DECAPx10_ASAP7_75t_R FILLER_3_242 ();
 DECAPx10_ASAP7_75t_R FILLER_3_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_286 ();
 DECAPx4_ASAP7_75t_R FILLER_3_293 ();
 FILLER_ASAP7_75t_R FILLER_3_303 ();
 FILLER_ASAP7_75t_R FILLER_3_311 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx2_ASAP7_75t_R FILLER_4_46 ();
 FILLER_ASAP7_75t_R FILLER_4_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_54 ();
 DECAPx10_ASAP7_75t_R FILLER_4_66 ();
 FILLER_ASAP7_75t_R FILLER_4_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_90 ();
 FILLER_ASAP7_75t_R FILLER_4_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_100 ();
 DECAPx10_ASAP7_75t_R FILLER_4_104 ();
 DECAPx10_ASAP7_75t_R FILLER_4_126 ();
 DECAPx10_ASAP7_75t_R FILLER_4_148 ();
 DECAPx10_ASAP7_75t_R FILLER_4_170 ();
 DECAPx10_ASAP7_75t_R FILLER_4_192 ();
 DECAPx10_ASAP7_75t_R FILLER_4_214 ();
 DECAPx10_ASAP7_75t_R FILLER_4_236 ();
 DECAPx10_ASAP7_75t_R FILLER_4_258 ();
 DECAPx2_ASAP7_75t_R FILLER_4_280 ();
 FILLER_ASAP7_75t_R FILLER_4_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_288 ();
 DECAPx2_ASAP7_75t_R FILLER_4_295 ();
 DECAPx2_ASAP7_75t_R FILLER_4_313 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx6_ASAP7_75t_R FILLER_5_24 ();
 DECAPx2_ASAP7_75t_R FILLER_5_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_44 ();
 FILLER_ASAP7_75t_R FILLER_5_65 ();
 DECAPx4_ASAP7_75t_R FILLER_5_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_94 ();
 FILLER_ASAP7_75t_R FILLER_5_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_114 ();
 FILLER_ASAP7_75t_R FILLER_5_121 ();
 DECAPx10_ASAP7_75t_R FILLER_5_129 ();
 DECAPx10_ASAP7_75t_R FILLER_5_151 ();
 DECAPx10_ASAP7_75t_R FILLER_5_173 ();
 DECAPx10_ASAP7_75t_R FILLER_5_195 ();
 DECAPx10_ASAP7_75t_R FILLER_5_217 ();
 DECAPx10_ASAP7_75t_R FILLER_5_239 ();
 DECAPx10_ASAP7_75t_R FILLER_5_261 ();
 DECAPx6_ASAP7_75t_R FILLER_5_283 ();
 FILLER_ASAP7_75t_R FILLER_5_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_324 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx1_ASAP7_75t_R FILLER_6_24 ();
 DECAPx4_ASAP7_75t_R FILLER_6_39 ();
 FILLER_ASAP7_75t_R FILLER_6_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_51 ();
 DECAPx1_ASAP7_75t_R FILLER_6_58 ();
 DECAPx1_ASAP7_75t_R FILLER_6_74 ();
 FILLER_ASAP7_75t_R FILLER_6_100 ();
 DECAPx1_ASAP7_75t_R FILLER_6_114 ();
 DECAPx10_ASAP7_75t_R FILLER_6_146 ();
 DECAPx10_ASAP7_75t_R FILLER_6_168 ();
 DECAPx10_ASAP7_75t_R FILLER_6_190 ();
 DECAPx6_ASAP7_75t_R FILLER_6_212 ();
 DECAPx2_ASAP7_75t_R FILLER_6_232 ();
 DECAPx6_ASAP7_75t_R FILLER_6_244 ();
 FILLER_ASAP7_75t_R FILLER_6_258 ();
 DECAPx10_ASAP7_75t_R FILLER_6_266 ();
 DECAPx6_ASAP7_75t_R FILLER_6_288 ();
 DECAPx1_ASAP7_75t_R FILLER_6_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_306 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_24 ();
 FILLER_ASAP7_75t_R FILLER_7_63 ();
 DECAPx2_ASAP7_75t_R FILLER_7_82 ();
 DECAPx4_ASAP7_75t_R FILLER_7_94 ();
 FILLER_ASAP7_75t_R FILLER_7_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_115 ();
 DECAPx10_ASAP7_75t_R FILLER_7_128 ();
 DECAPx10_ASAP7_75t_R FILLER_7_150 ();
 DECAPx10_ASAP7_75t_R FILLER_7_172 ();
 DECAPx10_ASAP7_75t_R FILLER_7_194 ();
 DECAPx1_ASAP7_75t_R FILLER_7_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_220 ();
 DECAPx2_ASAP7_75t_R FILLER_7_245 ();
 DECAPx1_ASAP7_75t_R FILLER_7_257 ();
 DECAPx1_ASAP7_75t_R FILLER_7_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_277 ();
 DECAPx1_ASAP7_75t_R FILLER_7_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_300 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx1_ASAP7_75t_R FILLER_8_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_28 ();
 DECAPx4_ASAP7_75t_R FILLER_8_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_45 ();
 DECAPx6_ASAP7_75t_R FILLER_8_49 ();
 DECAPx2_ASAP7_75t_R FILLER_8_63 ();
 DECAPx4_ASAP7_75t_R FILLER_8_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_87 ();
 FILLER_ASAP7_75t_R FILLER_8_94 ();
 DECAPx10_ASAP7_75t_R FILLER_8_119 ();
 DECAPx10_ASAP7_75t_R FILLER_8_141 ();
 DECAPx10_ASAP7_75t_R FILLER_8_163 ();
 DECAPx10_ASAP7_75t_R FILLER_8_185 ();
 DECAPx4_ASAP7_75t_R FILLER_8_207 ();
 FILLER_ASAP7_75t_R FILLER_8_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_219 ();
 DECAPx2_ASAP7_75t_R FILLER_8_232 ();
 DECAPx4_ASAP7_75t_R FILLER_8_250 ();
 FILLER_ASAP7_75t_R FILLER_8_260 ();
 DECAPx1_ASAP7_75t_R FILLER_8_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_278 ();
 DECAPx1_ASAP7_75t_R FILLER_8_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_313 ();
 DECAPx1_ASAP7_75t_R FILLER_8_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_336 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx2_ASAP7_75t_R FILLER_9_24 ();
 DECAPx1_ASAP7_75t_R FILLER_9_44 ();
 DECAPx1_ASAP7_75t_R FILLER_9_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_69 ();
 DECAPx2_ASAP7_75t_R FILLER_9_79 ();
 FILLER_ASAP7_75t_R FILLER_9_105 ();
 DECAPx4_ASAP7_75t_R FILLER_9_113 ();
 FILLER_ASAP7_75t_R FILLER_9_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_125 ();
 DECAPx10_ASAP7_75t_R FILLER_9_131 ();
 DECAPx10_ASAP7_75t_R FILLER_9_153 ();
 DECAPx10_ASAP7_75t_R FILLER_9_175 ();
 DECAPx10_ASAP7_75t_R FILLER_9_197 ();
 DECAPx2_ASAP7_75t_R FILLER_9_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_225 ();
 DECAPx1_ASAP7_75t_R FILLER_9_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_273 ();
 FILLER_ASAP7_75t_R FILLER_9_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_294 ();
 DECAPx6_ASAP7_75t_R FILLER_10_2 ();
 FILLER_ASAP7_75t_R FILLER_10_38 ();
 DECAPx2_ASAP7_75t_R FILLER_10_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_66 ();
 DECAPx4_ASAP7_75t_R FILLER_10_78 ();
 FILLER_ASAP7_75t_R FILLER_10_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_10_98 ();
 DECAPx10_ASAP7_75t_R FILLER_10_120 ();
 DECAPx10_ASAP7_75t_R FILLER_10_142 ();
 DECAPx10_ASAP7_75t_R FILLER_10_164 ();
 DECAPx6_ASAP7_75t_R FILLER_10_186 ();
 FILLER_ASAP7_75t_R FILLER_10_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_215 ();
 FILLER_ASAP7_75t_R FILLER_10_222 ();
 DECAPx4_ASAP7_75t_R FILLER_10_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_246 ();
 DECAPx4_ASAP7_75t_R FILLER_10_253 ();
 FILLER_ASAP7_75t_R FILLER_10_263 ();
 DECAPx2_ASAP7_75t_R FILLER_10_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_277 ();
 DECAPx2_ASAP7_75t_R FILLER_10_290 ();
 DECAPx1_ASAP7_75t_R FILLER_10_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_318 ();
 DECAPx10_ASAP7_75t_R FILLER_11_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_37 ();
 FILLER_ASAP7_75t_R FILLER_11_44 ();
 DECAPx2_ASAP7_75t_R FILLER_11_52 ();
 FILLER_ASAP7_75t_R FILLER_11_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_60 ();
 FILLER_ASAP7_75t_R FILLER_11_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_74 ();
 DECAPx4_ASAP7_75t_R FILLER_11_81 ();
 FILLER_ASAP7_75t_R FILLER_11_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_93 ();
 DECAPx2_ASAP7_75t_R FILLER_11_100 ();
 FILLER_ASAP7_75t_R FILLER_11_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_108 ();
 DECAPx1_ASAP7_75t_R FILLER_11_131 ();
 DECAPx10_ASAP7_75t_R FILLER_11_153 ();
 DECAPx10_ASAP7_75t_R FILLER_11_175 ();
 DECAPx1_ASAP7_75t_R FILLER_11_197 ();
 FILLER_ASAP7_75t_R FILLER_11_207 ();
 DECAPx6_ASAP7_75t_R FILLER_11_227 ();
 DECAPx2_ASAP7_75t_R FILLER_11_241 ();
 DECAPx10_ASAP7_75t_R FILLER_11_253 ();
 DECAPx6_ASAP7_75t_R FILLER_11_275 ();
 DECAPx2_ASAP7_75t_R FILLER_11_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_302 ();
 FILLER_ASAP7_75t_R FILLER_11_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_330 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_12_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_46 ();
 FILLER_ASAP7_75t_R FILLER_12_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_61 ();
 DECAPx1_ASAP7_75t_R FILLER_12_65 ();
 DECAPx2_ASAP7_75t_R FILLER_12_81 ();
 DECAPx1_ASAP7_75t_R FILLER_12_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_113 ();
 DECAPx10_ASAP7_75t_R FILLER_12_126 ();
 DECAPx10_ASAP7_75t_R FILLER_12_148 ();
 DECAPx10_ASAP7_75t_R FILLER_12_170 ();
 DECAPx10_ASAP7_75t_R FILLER_12_192 ();
 FILLER_ASAP7_75t_R FILLER_12_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_216 ();
 DECAPx6_ASAP7_75t_R FILLER_12_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_237 ();
 FILLER_ASAP7_75t_R FILLER_12_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_250 ();
 DECAPx1_ASAP7_75t_R FILLER_12_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_261 ();
 DECAPx4_ASAP7_75t_R FILLER_12_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_303 ();
 FILLER_ASAP7_75t_R FILLER_12_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_324 ();
 DECAPx4_ASAP7_75t_R FILLER_13_2 ();
 FILLER_ASAP7_75t_R FILLER_13_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_14 ();
 FILLER_ASAP7_75t_R FILLER_13_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_29 ();
 DECAPx4_ASAP7_75t_R FILLER_13_33 ();
 FILLER_ASAP7_75t_R FILLER_13_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_45 ();
 DECAPx1_ASAP7_75t_R FILLER_13_66 ();
 FILLER_ASAP7_75t_R FILLER_13_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_94 ();
 FILLER_ASAP7_75t_R FILLER_13_107 ();
 DECAPx10_ASAP7_75t_R FILLER_13_126 ();
 DECAPx2_ASAP7_75t_R FILLER_13_148 ();
 FILLER_ASAP7_75t_R FILLER_13_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_156 ();
 DECAPx6_ASAP7_75t_R FILLER_13_163 ();
 DECAPx1_ASAP7_75t_R FILLER_13_183 ();
 DECAPx10_ASAP7_75t_R FILLER_13_193 ();
 FILLER_ASAP7_75t_R FILLER_13_215 ();
 FILLER_ASAP7_75t_R FILLER_13_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_231 ();
 DECAPx1_ASAP7_75t_R FILLER_13_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_258 ();
 DECAPx1_ASAP7_75t_R FILLER_13_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_307 ();
 FILLER_ASAP7_75t_R FILLER_13_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_316 ();
 FILLER_ASAP7_75t_R FILLER_13_329 ();
 DECAPx2_ASAP7_75t_R FILLER_14_2 ();
 FILLER_ASAP7_75t_R FILLER_14_8 ();
 DECAPx10_ASAP7_75t_R FILLER_14_51 ();
 DECAPx6_ASAP7_75t_R FILLER_14_73 ();
 DECAPx2_ASAP7_75t_R FILLER_14_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_93 ();
 DECAPx2_ASAP7_75t_R FILLER_14_111 ();
 FILLER_ASAP7_75t_R FILLER_14_117 ();
 FILLER_ASAP7_75t_R FILLER_14_134 ();
 FILLER_ASAP7_75t_R FILLER_14_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_197 ();
 DECAPx1_ASAP7_75t_R FILLER_14_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_252 ();
 DECAPx1_ASAP7_75t_R FILLER_14_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_300 ();
 FILLER_ASAP7_75t_R FILLER_14_307 ();
 FILLER_ASAP7_75t_R FILLER_14_321 ();
 FILLER_ASAP7_75t_R FILLER_14_335 ();
 DECAPx2_ASAP7_75t_R FILLER_15_2 ();
 FILLER_ASAP7_75t_R FILLER_15_8 ();
 FILLER_ASAP7_75t_R FILLER_15_21 ();
 FILLER_ASAP7_75t_R FILLER_15_29 ();
 DECAPx10_ASAP7_75t_R FILLER_15_67 ();
 DECAPx4_ASAP7_75t_R FILLER_15_89 ();
 FILLER_ASAP7_75t_R FILLER_15_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_101 ();
 DECAPx2_ASAP7_75t_R FILLER_15_141 ();
 FILLER_ASAP7_75t_R FILLER_15_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_149 ();
 FILLER_ASAP7_75t_R FILLER_15_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_180 ();
 DECAPx6_ASAP7_75t_R FILLER_15_196 ();
 DECAPx2_ASAP7_75t_R FILLER_15_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_255 ();
 FILLER_ASAP7_75t_R FILLER_15_262 ();
 DECAPx2_ASAP7_75t_R FILLER_15_276 ();
 FILLER_ASAP7_75t_R FILLER_15_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_304 ();
 FILLER_ASAP7_75t_R FILLER_15_335 ();
 FILLER_ASAP7_75t_R FILLER_16_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_4 ();
 DECAPx6_ASAP7_75t_R FILLER_16_22 ();
 DECAPx1_ASAP7_75t_R FILLER_16_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_40 ();
 DECAPx6_ASAP7_75t_R FILLER_16_47 ();
 FILLER_ASAP7_75t_R FILLER_16_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_63 ();
 DECAPx4_ASAP7_75t_R FILLER_16_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_92 ();
 FILLER_ASAP7_75t_R FILLER_16_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_113 ();
 FILLER_ASAP7_75t_R FILLER_16_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_119 ();
 DECAPx6_ASAP7_75t_R FILLER_16_139 ();
 DECAPx4_ASAP7_75t_R FILLER_16_165 ();
 FILLER_ASAP7_75t_R FILLER_16_175 ();
 DECAPx1_ASAP7_75t_R FILLER_16_183 ();
 DECAPx10_ASAP7_75t_R FILLER_16_199 ();
 DECAPx1_ASAP7_75t_R FILLER_16_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_249 ();
 DECAPx2_ASAP7_75t_R FILLER_16_262 ();
 FILLER_ASAP7_75t_R FILLER_16_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_270 ();
 DECAPx2_ASAP7_75t_R FILLER_16_283 ();
 FILLER_ASAP7_75t_R FILLER_16_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_304 ();
 FILLER_ASAP7_75t_R FILLER_16_329 ();
 DECAPx4_ASAP7_75t_R FILLER_17_2 ();
 DECAPx6_ASAP7_75t_R FILLER_17_18 ();
 FILLER_ASAP7_75t_R FILLER_17_32 ();
 DECAPx2_ASAP7_75t_R FILLER_17_54 ();
 DECAPx2_ASAP7_75t_R FILLER_17_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_100 ();
 DECAPx10_ASAP7_75t_R FILLER_17_124 ();
 DECAPx2_ASAP7_75t_R FILLER_17_146 ();
 FILLER_ASAP7_75t_R FILLER_17_152 ();
 DECAPx10_ASAP7_75t_R FILLER_17_166 ();
 DECAPx2_ASAP7_75t_R FILLER_17_188 ();
 FILLER_ASAP7_75t_R FILLER_17_194 ();
 DECAPx4_ASAP7_75t_R FILLER_17_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_218 ();
 FILLER_ASAP7_75t_R FILLER_17_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_240 ();
 DECAPx6_ASAP7_75t_R FILLER_17_247 ();
 DECAPx1_ASAP7_75t_R FILLER_17_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_265 ();
 DECAPx4_ASAP7_75t_R FILLER_17_272 ();
 FILLER_ASAP7_75t_R FILLER_17_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_307 ();
 DECAPx1_ASAP7_75t_R FILLER_17_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_330 ();
 FILLER_ASAP7_75t_R FILLER_18_2 ();
 DECAPx4_ASAP7_75t_R FILLER_18_27 ();
 FILLER_ASAP7_75t_R FILLER_18_37 ();
 FILLER_ASAP7_75t_R FILLER_18_56 ();
 DECAPx4_ASAP7_75t_R FILLER_18_65 ();
 FILLER_ASAP7_75t_R FILLER_18_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_77 ();
 DECAPx1_ASAP7_75t_R FILLER_18_114 ();
 DECAPx4_ASAP7_75t_R FILLER_18_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_150 ();
 FILLER_ASAP7_75t_R FILLER_18_185 ();
 FILLER_ASAP7_75t_R FILLER_18_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_201 ();
 DECAPx4_ASAP7_75t_R FILLER_18_208 ();
 FILLER_ASAP7_75t_R FILLER_18_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_220 ();
 DECAPx4_ASAP7_75t_R FILLER_18_239 ();
 FILLER_ASAP7_75t_R FILLER_18_249 ();
 FILLER_ASAP7_75t_R FILLER_18_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_259 ();
 FILLER_ASAP7_75t_R FILLER_18_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_316 ();
 FILLER_ASAP7_75t_R FILLER_18_329 ();
 DECAPx1_ASAP7_75t_R FILLER_19_2 ();
 FILLER_ASAP7_75t_R FILLER_19_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_20 ();
 DECAPx2_ASAP7_75t_R FILLER_19_43 ();
 DECAPx4_ASAP7_75t_R FILLER_19_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_81 ();
 DECAPx10_ASAP7_75t_R FILLER_19_95 ();
 DECAPx2_ASAP7_75t_R FILLER_19_117 ();
 FILLER_ASAP7_75t_R FILLER_19_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_125 ();
 DECAPx6_ASAP7_75t_R FILLER_19_143 ();
 DECAPx1_ASAP7_75t_R FILLER_19_157 ();
 DECAPx1_ASAP7_75t_R FILLER_19_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_188 ();
 DECAPx10_ASAP7_75t_R FILLER_19_202 ();
 DECAPx4_ASAP7_75t_R FILLER_19_242 ();
 FILLER_ASAP7_75t_R FILLER_19_252 ();
 DECAPx2_ASAP7_75t_R FILLER_19_282 ();
 FILLER_ASAP7_75t_R FILLER_19_288 ();
 FILLER_ASAP7_75t_R FILLER_19_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_336 ();
 DECAPx2_ASAP7_75t_R FILLER_20_2 ();
 DECAPx4_ASAP7_75t_R FILLER_20_16 ();
 FILLER_ASAP7_75t_R FILLER_20_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_28 ();
 DECAPx6_ASAP7_75t_R FILLER_20_59 ();
 FILLER_ASAP7_75t_R FILLER_20_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_85 ();
 DECAPx6_ASAP7_75t_R FILLER_20_98 ();
 FILLER_ASAP7_75t_R FILLER_20_112 ();
 DECAPx6_ASAP7_75t_R FILLER_20_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_150 ();
 DECAPx4_ASAP7_75t_R FILLER_20_163 ();
 FILLER_ASAP7_75t_R FILLER_20_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_175 ();
 FILLER_ASAP7_75t_R FILLER_20_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_184 ();
 DECAPx1_ASAP7_75t_R FILLER_20_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_195 ();
 DECAPx1_ASAP7_75t_R FILLER_20_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_206 ();
 DECAPx1_ASAP7_75t_R FILLER_20_217 ();
 FILLER_ASAP7_75t_R FILLER_20_227 ();
 DECAPx4_ASAP7_75t_R FILLER_20_245 ();
 FILLER_ASAP7_75t_R FILLER_20_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_257 ();
 DECAPx2_ASAP7_75t_R FILLER_20_276 ();
 DECAPx1_ASAP7_75t_R FILLER_20_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_310 ();
 FILLER_ASAP7_75t_R FILLER_20_335 ();
 DECAPx4_ASAP7_75t_R FILLER_21_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_12 ();
 DECAPx2_ASAP7_75t_R FILLER_21_19 ();
 DECAPx10_ASAP7_75t_R FILLER_21_43 ();
 DECAPx6_ASAP7_75t_R FILLER_21_96 ();
 FILLER_ASAP7_75t_R FILLER_21_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_112 ();
 FILLER_ASAP7_75t_R FILLER_21_119 ();
 DECAPx6_ASAP7_75t_R FILLER_21_136 ();
 DECAPx4_ASAP7_75t_R FILLER_21_162 ();
 FILLER_ASAP7_75t_R FILLER_21_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_193 ();
 DECAPx6_ASAP7_75t_R FILLER_21_206 ();
 DECAPx2_ASAP7_75t_R FILLER_21_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_240 ();
 DECAPx4_ASAP7_75t_R FILLER_21_251 ();
 DECAPx2_ASAP7_75t_R FILLER_21_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_277 ();
 DECAPx1_ASAP7_75t_R FILLER_21_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_318 ();
 DECAPx1_ASAP7_75t_R FILLER_22_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_6 ();
 DECAPx6_ASAP7_75t_R FILLER_22_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_27 ();
 DECAPx2_ASAP7_75t_R FILLER_22_39 ();
 FILLER_ASAP7_75t_R FILLER_22_45 ();
 DECAPx6_ASAP7_75t_R FILLER_22_69 ();
 FILLER_ASAP7_75t_R FILLER_22_83 ();
 DECAPx2_ASAP7_75t_R FILLER_22_91 ();
 FILLER_ASAP7_75t_R FILLER_22_97 ();
 DECAPx6_ASAP7_75t_R FILLER_22_133 ();
 DECAPx1_ASAP7_75t_R FILLER_22_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_183 ();
 FILLER_ASAP7_75t_R FILLER_22_191 ();
 DECAPx2_ASAP7_75t_R FILLER_22_201 ();
 FILLER_ASAP7_75t_R FILLER_22_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_209 ();
 DECAPx10_ASAP7_75t_R FILLER_22_220 ();
 DECAPx10_ASAP7_75t_R FILLER_22_242 ();
 DECAPx6_ASAP7_75t_R FILLER_22_264 ();
 FILLER_ASAP7_75t_R FILLER_22_278 ();
 DECAPx1_ASAP7_75t_R FILLER_22_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_336 ();
 DECAPx2_ASAP7_75t_R FILLER_23_2 ();
 DECAPx2_ASAP7_75t_R FILLER_23_36 ();
 DECAPx4_ASAP7_75t_R FILLER_23_52 ();
 FILLER_ASAP7_75t_R FILLER_23_62 ();
 DECAPx2_ASAP7_75t_R FILLER_23_72 ();
 FILLER_ASAP7_75t_R FILLER_23_78 ();
 DECAPx4_ASAP7_75t_R FILLER_23_96 ();
 FILLER_ASAP7_75t_R FILLER_23_106 ();
 FILLER_ASAP7_75t_R FILLER_23_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_114 ();
 DECAPx6_ASAP7_75t_R FILLER_23_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_135 ();
 DECAPx2_ASAP7_75t_R FILLER_23_146 ();
 DECAPx1_ASAP7_75t_R FILLER_23_164 ();
 DECAPx10_ASAP7_75t_R FILLER_23_190 ();
 FILLER_ASAP7_75t_R FILLER_23_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_214 ();
 DECAPx10_ASAP7_75t_R FILLER_23_235 ();
 DECAPx6_ASAP7_75t_R FILLER_23_257 ();
 DECAPx2_ASAP7_75t_R FILLER_23_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_291 ();
 FILLER_ASAP7_75t_R FILLER_23_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_300 ();
 DECAPx4_ASAP7_75t_R FILLER_24_2 ();
 FILLER_ASAP7_75t_R FILLER_24_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_60 ();
 DECAPx4_ASAP7_75t_R FILLER_24_69 ();
 FILLER_ASAP7_75t_R FILLER_24_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_81 ();
 FILLER_ASAP7_75t_R FILLER_24_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_94 ();
 FILLER_ASAP7_75t_R FILLER_24_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_135 ();
 DECAPx4_ASAP7_75t_R FILLER_24_139 ();
 FILLER_ASAP7_75t_R FILLER_24_149 ();
 DECAPx6_ASAP7_75t_R FILLER_24_163 ();
 DECAPx2_ASAP7_75t_R FILLER_24_177 ();
 FILLER_ASAP7_75t_R FILLER_24_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_189 ();
 DECAPx1_ASAP7_75t_R FILLER_24_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_206 ();
 FILLER_ASAP7_75t_R FILLER_24_213 ();
 DECAPx6_ASAP7_75t_R FILLER_24_225 ();
 DECAPx1_ASAP7_75t_R FILLER_24_239 ();
 FILLER_ASAP7_75t_R FILLER_24_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_261 ();
 DECAPx4_ASAP7_75t_R FILLER_24_272 ();
 FILLER_ASAP7_75t_R FILLER_24_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_301 ();
 DECAPx4_ASAP7_75t_R FILLER_24_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_330 ();
 DECAPx10_ASAP7_75t_R FILLER_25_2 ();
 DECAPx2_ASAP7_75t_R FILLER_25_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_40 ();
 DECAPx4_ASAP7_75t_R FILLER_25_54 ();
 DECAPx1_ASAP7_75t_R FILLER_25_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_82 ();
 DECAPx1_ASAP7_75t_R FILLER_25_86 ();
 DECAPx2_ASAP7_75t_R FILLER_25_106 ();
 FILLER_ASAP7_75t_R FILLER_25_151 ();
 DECAPx6_ASAP7_75t_R FILLER_25_159 ();
 DECAPx2_ASAP7_75t_R FILLER_25_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_199 ();
 FILLER_ASAP7_75t_R FILLER_25_206 ();
 DECAPx1_ASAP7_75t_R FILLER_25_214 ();
 FILLER_ASAP7_75t_R FILLER_25_224 ();
 DECAPx4_ASAP7_75t_R FILLER_25_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_252 ();
 DECAPx6_ASAP7_75t_R FILLER_25_263 ();
 DECAPx2_ASAP7_75t_R FILLER_25_277 ();
 FILLER_ASAP7_75t_R FILLER_25_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_291 ();
 FILLER_ASAP7_75t_R FILLER_25_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_324 ();
 DECAPx10_ASAP7_75t_R FILLER_26_2 ();
 DECAPx4_ASAP7_75t_R FILLER_26_24 ();
 FILLER_ASAP7_75t_R FILLER_26_34 ();
 DECAPx2_ASAP7_75t_R FILLER_26_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_61 ();
 DECAPx2_ASAP7_75t_R FILLER_26_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_74 ();
 FILLER_ASAP7_75t_R FILLER_26_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_101 ();
 FILLER_ASAP7_75t_R FILLER_26_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_120 ();
 DECAPx4_ASAP7_75t_R FILLER_26_145 ();
 FILLER_ASAP7_75t_R FILLER_26_155 ();
 DECAPx2_ASAP7_75t_R FILLER_26_175 ();
 DECAPx4_ASAP7_75t_R FILLER_26_191 ();
 FILLER_ASAP7_75t_R FILLER_26_201 ();
 FILLER_ASAP7_75t_R FILLER_26_209 ();
 DECAPx2_ASAP7_75t_R FILLER_26_229 ();
 DECAPx2_ASAP7_75t_R FILLER_26_255 ();
 FILLER_ASAP7_75t_R FILLER_26_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_263 ();
 DECAPx1_ASAP7_75t_R FILLER_26_280 ();
 DECAPx1_ASAP7_75t_R FILLER_26_290 ();
 DECAPx1_ASAP7_75t_R FILLER_26_300 ();
 FILLER_ASAP7_75t_R FILLER_26_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_330 ();
 FILLER_ASAP7_75t_R FILLER_27_2 ();
 DECAPx2_ASAP7_75t_R FILLER_27_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_22 ();
 DECAPx2_ASAP7_75t_R FILLER_27_57 ();
 DECAPx2_ASAP7_75t_R FILLER_27_75 ();
 DECAPx1_ASAP7_75t_R FILLER_27_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_97 ();
 DECAPx2_ASAP7_75t_R FILLER_27_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_112 ();
 DECAPx2_ASAP7_75t_R FILLER_27_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_129 ();
 DECAPx4_ASAP7_75t_R FILLER_27_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_158 ();
 DECAPx2_ASAP7_75t_R FILLER_27_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_184 ();
 DECAPx10_ASAP7_75t_R FILLER_27_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_217 ();
 DECAPx6_ASAP7_75t_R FILLER_27_248 ();
 DECAPx1_ASAP7_75t_R FILLER_27_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_276 ();
 FILLER_ASAP7_75t_R FILLER_27_323 ();
 FILLER_ASAP7_75t_R FILLER_28_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_4 ();
 DECAPx4_ASAP7_75t_R FILLER_28_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_27 ();
 FILLER_ASAP7_75t_R FILLER_28_38 ();
 DECAPx4_ASAP7_75t_R FILLER_28_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_79 ();
 DECAPx4_ASAP7_75t_R FILLER_28_90 ();
 FILLER_ASAP7_75t_R FILLER_28_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_102 ();
 DECAPx10_ASAP7_75t_R FILLER_28_135 ();
 DECAPx10_ASAP7_75t_R FILLER_28_157 ();
 DECAPx10_ASAP7_75t_R FILLER_28_179 ();
 FILLER_ASAP7_75t_R FILLER_28_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_220 ();
 DECAPx1_ASAP7_75t_R FILLER_28_233 ();
 FILLER_ASAP7_75t_R FILLER_28_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_249 ();
 DECAPx6_ASAP7_75t_R FILLER_28_260 ();
 DECAPx1_ASAP7_75t_R FILLER_28_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_2 ();
 DECAPx2_ASAP7_75t_R FILLER_29_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_15 ();
 FILLER_ASAP7_75t_R FILLER_29_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_30 ();
 DECAPx4_ASAP7_75t_R FILLER_29_37 ();
 DECAPx4_ASAP7_75t_R FILLER_29_60 ();
 FILLER_ASAP7_75t_R FILLER_29_70 ();
 DECAPx4_ASAP7_75t_R FILLER_29_89 ();
 FILLER_ASAP7_75t_R FILLER_29_99 ();
 FILLER_ASAP7_75t_R FILLER_29_117 ();
 DECAPx10_ASAP7_75t_R FILLER_29_133 ();
 DECAPx6_ASAP7_75t_R FILLER_29_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_186 ();
 DECAPx4_ASAP7_75t_R FILLER_29_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_207 ();
 FILLER_ASAP7_75t_R FILLER_29_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_222 ();
 DECAPx10_ASAP7_75t_R FILLER_29_239 ();
 DECAPx6_ASAP7_75t_R FILLER_29_261 ();
 DECAPx1_ASAP7_75t_R FILLER_29_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_296 ();
 DECAPx1_ASAP7_75t_R FILLER_29_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_336 ();
 DECAPx1_ASAP7_75t_R FILLER_30_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_6 ();
 DECAPx2_ASAP7_75t_R FILLER_30_35 ();
 FILLER_ASAP7_75t_R FILLER_30_41 ();
 FILLER_ASAP7_75t_R FILLER_30_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_73 ();
 FILLER_ASAP7_75t_R FILLER_30_119 ();
 DECAPx10_ASAP7_75t_R FILLER_30_128 ();
 DECAPx10_ASAP7_75t_R FILLER_30_150 ();
 DECAPx2_ASAP7_75t_R FILLER_30_172 ();
 FILLER_ASAP7_75t_R FILLER_30_178 ();
 DECAPx2_ASAP7_75t_R FILLER_30_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_222 ();
 DECAPx2_ASAP7_75t_R FILLER_30_235 ();
 FILLER_ASAP7_75t_R FILLER_30_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_243 ();
 FILLER_ASAP7_75t_R FILLER_30_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_256 ();
 DECAPx10_ASAP7_75t_R FILLER_30_267 ();
 DECAPx2_ASAP7_75t_R FILLER_30_289 ();
 FILLER_ASAP7_75t_R FILLER_30_295 ();
 DECAPx1_ASAP7_75t_R FILLER_30_321 ();
 DECAPx2_ASAP7_75t_R FILLER_30_331 ();
 FILLER_ASAP7_75t_R FILLER_31_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_4 ();
 DECAPx1_ASAP7_75t_R FILLER_31_28 ();
 DECAPx10_ASAP7_75t_R FILLER_31_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_78 ();
 DECAPx4_ASAP7_75t_R FILLER_31_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_101 ();
 DECAPx6_ASAP7_75t_R FILLER_31_134 ();
 DECAPx2_ASAP7_75t_R FILLER_31_148 ();
 DECAPx6_ASAP7_75t_R FILLER_31_168 ();
 DECAPx4_ASAP7_75t_R FILLER_31_192 ();
 FILLER_ASAP7_75t_R FILLER_31_202 ();
 DECAPx2_ASAP7_75t_R FILLER_31_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_222 ();
 DECAPx2_ASAP7_75t_R FILLER_31_229 ();
 DECAPx10_ASAP7_75t_R FILLER_31_245 ();
 FILLER_ASAP7_75t_R FILLER_31_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_269 ();
 DECAPx10_ASAP7_75t_R FILLER_31_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_302 ();
 FILLER_ASAP7_75t_R FILLER_32_8 ();
 DECAPx2_ASAP7_75t_R FILLER_32_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_28 ();
 DECAPx6_ASAP7_75t_R FILLER_32_51 ();
 DECAPx2_ASAP7_75t_R FILLER_32_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_71 ();
 FILLER_ASAP7_75t_R FILLER_32_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_128 ();
 DECAPx2_ASAP7_75t_R FILLER_32_139 ();
 FILLER_ASAP7_75t_R FILLER_32_155 ();
 DECAPx2_ASAP7_75t_R FILLER_32_163 ();
 FILLER_ASAP7_75t_R FILLER_32_169 ();
 DECAPx6_ASAP7_75t_R FILLER_32_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_195 ();
 FILLER_ASAP7_75t_R FILLER_32_212 ();
 DECAPx1_ASAP7_75t_R FILLER_32_220 ();
 DECAPx1_ASAP7_75t_R FILLER_32_230 ();
 FILLER_ASAP7_75t_R FILLER_32_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_242 ();
 DECAPx10_ASAP7_75t_R FILLER_32_253 ();
 DECAPx1_ASAP7_75t_R FILLER_32_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_279 ();
 DECAPx1_ASAP7_75t_R FILLER_32_290 ();
 DECAPx2_ASAP7_75t_R FILLER_32_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_324 ();
 DECAPx2_ASAP7_75t_R FILLER_33_2 ();
 DECAPx6_ASAP7_75t_R FILLER_33_44 ();
 DECAPx2_ASAP7_75t_R FILLER_33_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_64 ();
 DECAPx2_ASAP7_75t_R FILLER_33_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_83 ();
 DECAPx4_ASAP7_75t_R FILLER_33_96 ();
 DECAPx1_ASAP7_75t_R FILLER_33_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_119 ();
 DECAPx1_ASAP7_75t_R FILLER_33_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_132 ();
 FILLER_ASAP7_75t_R FILLER_33_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_141 ();
 DECAPx4_ASAP7_75t_R FILLER_33_172 ();
 FILLER_ASAP7_75t_R FILLER_33_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_205 ();
 DECAPx2_ASAP7_75t_R FILLER_33_218 ();
 DECAPx2_ASAP7_75t_R FILLER_33_236 ();
 FILLER_ASAP7_75t_R FILLER_33_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_244 ();
 DECAPx10_ASAP7_75t_R FILLER_33_255 ();
 DECAPx6_ASAP7_75t_R FILLER_33_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_42 ();
 DECAPx4_ASAP7_75t_R FILLER_34_59 ();
 FILLER_ASAP7_75t_R FILLER_34_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_71 ();
 DECAPx10_ASAP7_75t_R FILLER_34_83 ();
 DECAPx6_ASAP7_75t_R FILLER_34_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_119 ();
 FILLER_ASAP7_75t_R FILLER_34_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_142 ();
 DECAPx1_ASAP7_75t_R FILLER_34_155 ();
 DECAPx10_ASAP7_75t_R FILLER_34_169 ();
 DECAPx1_ASAP7_75t_R FILLER_34_191 ();
 DECAPx2_ASAP7_75t_R FILLER_34_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_225 ();
 DECAPx2_ASAP7_75t_R FILLER_34_238 ();
 DECAPx2_ASAP7_75t_R FILLER_34_254 ();
 FILLER_ASAP7_75t_R FILLER_34_260 ();
 DECAPx4_ASAP7_75t_R FILLER_34_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_295 ();
 FILLER_ASAP7_75t_R FILLER_34_308 ();
 FILLER_ASAP7_75t_R FILLER_34_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_22 ();
 DECAPx6_ASAP7_75t_R FILLER_35_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_104 ();
 DECAPx1_ASAP7_75t_R FILLER_35_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_125 ();
 DECAPx1_ASAP7_75t_R FILLER_35_136 ();
 DECAPx6_ASAP7_75t_R FILLER_35_146 ();
 DECAPx6_ASAP7_75t_R FILLER_35_186 ();
 FILLER_ASAP7_75t_R FILLER_35_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_237 ();
 DECAPx10_ASAP7_75t_R FILLER_35_248 ();
 DECAPx2_ASAP7_75t_R FILLER_35_270 ();
 FILLER_ASAP7_75t_R FILLER_35_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_278 ();
 FILLER_ASAP7_75t_R FILLER_35_315 ();
 FILLER_ASAP7_75t_R FILLER_35_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_8 ();
 FILLER_ASAP7_75t_R FILLER_36_18 ();
 FILLER_ASAP7_75t_R FILLER_36_24 ();
 FILLER_ASAP7_75t_R FILLER_36_32 ();
 DECAPx2_ASAP7_75t_R FILLER_36_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_60 ();
 DECAPx1_ASAP7_75t_R FILLER_36_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_71 ();
 FILLER_ASAP7_75t_R FILLER_36_82 ();
 DECAPx2_ASAP7_75t_R FILLER_36_90 ();
 FILLER_ASAP7_75t_R FILLER_36_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_98 ();
 DECAPx2_ASAP7_75t_R FILLER_36_105 ();
 FILLER_ASAP7_75t_R FILLER_36_111 ();
 FILLER_ASAP7_75t_R FILLER_36_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_137 ();
 DECAPx4_ASAP7_75t_R FILLER_36_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_162 ();
 FILLER_ASAP7_75t_R FILLER_36_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_183 ();
 FILLER_ASAP7_75t_R FILLER_36_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_196 ();
 DECAPx2_ASAP7_75t_R FILLER_36_207 ();
 FILLER_ASAP7_75t_R FILLER_36_213 ();
 DECAPx2_ASAP7_75t_R FILLER_36_221 ();
 FILLER_ASAP7_75t_R FILLER_36_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_229 ();
 DECAPx1_ASAP7_75t_R FILLER_36_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_250 ();
 DECAPx1_ASAP7_75t_R FILLER_36_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_281 ();
 DECAPx1_ASAP7_75t_R FILLER_36_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_292 ();
 DECAPx2_ASAP7_75t_R FILLER_37_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_8 ();
 DECAPx2_ASAP7_75t_R FILLER_37_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_37 ();
 DECAPx2_ASAP7_75t_R FILLER_37_56 ();
 FILLER_ASAP7_75t_R FILLER_37_62 ();
 DECAPx4_ASAP7_75t_R FILLER_37_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_80 ();
 FILLER_ASAP7_75t_R FILLER_37_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_89 ();
 DECAPx2_ASAP7_75t_R FILLER_37_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_102 ();
 DECAPx1_ASAP7_75t_R FILLER_37_109 ();
 DECAPx10_ASAP7_75t_R FILLER_37_125 ();
 DECAPx10_ASAP7_75t_R FILLER_37_147 ();
 DECAPx2_ASAP7_75t_R FILLER_37_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_175 ();
 DECAPx6_ASAP7_75t_R FILLER_37_182 ();
 DECAPx1_ASAP7_75t_R FILLER_37_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_200 ();
 DECAPx6_ASAP7_75t_R FILLER_37_221 ();
 FILLER_ASAP7_75t_R FILLER_37_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_237 ();
 DECAPx10_ASAP7_75t_R FILLER_37_248 ();
 FILLER_ASAP7_75t_R FILLER_37_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_305 ();
 DECAPx1_ASAP7_75t_R FILLER_37_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_328 ();
 FILLER_ASAP7_75t_R FILLER_37_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_14 ();
 DECAPx1_ASAP7_75t_R FILLER_38_34 ();
 DECAPx4_ASAP7_75t_R FILLER_38_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_56 ();
 DECAPx6_ASAP7_75t_R FILLER_38_74 ();
 FILLER_ASAP7_75t_R FILLER_38_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_90 ();
 DECAPx1_ASAP7_75t_R FILLER_38_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_109 ();
 FILLER_ASAP7_75t_R FILLER_38_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_126 ();
 DECAPx2_ASAP7_75t_R FILLER_38_134 ();
 FILLER_ASAP7_75t_R FILLER_38_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_142 ();
 DECAPx6_ASAP7_75t_R FILLER_38_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_175 ();
 DECAPx2_ASAP7_75t_R FILLER_38_194 ();
 DECAPx1_ASAP7_75t_R FILLER_38_212 ();
 DECAPx10_ASAP7_75t_R FILLER_38_226 ();
 DECAPx1_ASAP7_75t_R FILLER_38_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_252 ();
 DECAPx4_ASAP7_75t_R FILLER_38_263 ();
 FILLER_ASAP7_75t_R FILLER_38_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_275 ();
 FILLER_ASAP7_75t_R FILLER_38_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_310 ();
 FILLER_ASAP7_75t_R FILLER_38_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_2 ();
 DECAPx2_ASAP7_75t_R FILLER_39_60 ();
 FILLER_ASAP7_75t_R FILLER_39_66 ();
 FILLER_ASAP7_75t_R FILLER_39_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_82 ();
 FILLER_ASAP7_75t_R FILLER_39_100 ();
 DECAPx2_ASAP7_75t_R FILLER_39_105 ();
 DECAPx6_ASAP7_75t_R FILLER_39_159 ();
 DECAPx1_ASAP7_75t_R FILLER_39_173 ();
 DECAPx2_ASAP7_75t_R FILLER_39_189 ();
 FILLER_ASAP7_75t_R FILLER_39_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_256 ();
 DECAPx10_ASAP7_75t_R FILLER_39_267 ();
 DECAPx10_ASAP7_75t_R FILLER_39_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_2 ();
 DECAPx1_ASAP7_75t_R FILLER_40_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_13 ();
 FILLER_ASAP7_75t_R FILLER_40_27 ();
 FILLER_ASAP7_75t_R FILLER_40_40 ();
 DECAPx1_ASAP7_75t_R FILLER_40_70 ();
 DECAPx1_ASAP7_75t_R FILLER_40_86 ();
 DECAPx2_ASAP7_75t_R FILLER_40_97 ();
 FILLER_ASAP7_75t_R FILLER_40_103 ();
 DECAPx2_ASAP7_75t_R FILLER_40_117 ();
 FILLER_ASAP7_75t_R FILLER_40_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_125 ();
 FILLER_ASAP7_75t_R FILLER_40_136 ();
 DECAPx1_ASAP7_75t_R FILLER_40_144 ();
 DECAPx2_ASAP7_75t_R FILLER_40_154 ();
 FILLER_ASAP7_75t_R FILLER_40_160 ();
 DECAPx2_ASAP7_75t_R FILLER_40_168 ();
 DECAPx4_ASAP7_75t_R FILLER_40_184 ();
 DECAPx2_ASAP7_75t_R FILLER_40_226 ();
 DECAPx1_ASAP7_75t_R FILLER_40_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_246 ();
 DECAPx2_ASAP7_75t_R FILLER_40_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_263 ();
 DECAPx4_ASAP7_75t_R FILLER_40_274 ();
 FILLER_ASAP7_75t_R FILLER_40_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_293 ();
 FILLER_ASAP7_75t_R FILLER_40_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_309 ();
 DECAPx2_ASAP7_75t_R FILLER_40_328 ();
 FILLER_ASAP7_75t_R FILLER_40_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_336 ();
 FILLER_ASAP7_75t_R FILLER_41_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_15 ();
 DECAPx2_ASAP7_75t_R FILLER_41_34 ();
 DECAPx6_ASAP7_75t_R FILLER_41_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_73 ();
 FILLER_ASAP7_75t_R FILLER_41_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_92 ();
 FILLER_ASAP7_75t_R FILLER_41_99 ();
 FILLER_ASAP7_75t_R FILLER_41_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_109 ();
 DECAPx10_ASAP7_75t_R FILLER_41_120 ();
 DECAPx6_ASAP7_75t_R FILLER_41_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_156 ();
 DECAPx4_ASAP7_75t_R FILLER_41_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_185 ();
 DECAPx10_ASAP7_75t_R FILLER_41_214 ();
 DECAPx10_ASAP7_75t_R FILLER_41_236 ();
 DECAPx10_ASAP7_75t_R FILLER_41_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_287 ();
 DECAPx4_ASAP7_75t_R FILLER_41_304 ();
 DECAPx1_ASAP7_75t_R FILLER_41_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_330 ();
 DECAPx6_ASAP7_75t_R FILLER_42_2 ();
 DECAPx1_ASAP7_75t_R FILLER_42_16 ();
 DECAPx4_ASAP7_75t_R FILLER_42_32 ();
 FILLER_ASAP7_75t_R FILLER_42_42 ();
 FILLER_ASAP7_75t_R FILLER_42_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_85 ();
 DECAPx10_ASAP7_75t_R FILLER_42_101 ();
 DECAPx6_ASAP7_75t_R FILLER_42_123 ();
 DECAPx1_ASAP7_75t_R FILLER_42_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_141 ();
 DECAPx1_ASAP7_75t_R FILLER_42_152 ();
 FILLER_ASAP7_75t_R FILLER_42_168 ();
 DECAPx10_ASAP7_75t_R FILLER_42_176 ();
 FILLER_ASAP7_75t_R FILLER_42_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_200 ();
 DECAPx1_ASAP7_75t_R FILLER_42_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_215 ();
 DECAPx1_ASAP7_75t_R FILLER_42_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_230 ();
 DECAPx10_ASAP7_75t_R FILLER_42_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_287 ();
 DECAPx4_ASAP7_75t_R FILLER_42_306 ();
 FILLER_ASAP7_75t_R FILLER_42_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_330 ();
 DECAPx1_ASAP7_75t_R FILLER_43_2 ();
 DECAPx4_ASAP7_75t_R FILLER_43_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_22 ();
 DECAPx6_ASAP7_75t_R FILLER_43_35 ();
 FILLER_ASAP7_75t_R FILLER_43_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_51 ();
 DECAPx1_ASAP7_75t_R FILLER_43_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_67 ();
 DECAPx1_ASAP7_75t_R FILLER_43_81 ();
 FILLER_ASAP7_75t_R FILLER_43_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_93 ();
 FILLER_ASAP7_75t_R FILLER_43_103 ();
 FILLER_ASAP7_75t_R FILLER_43_116 ();
 DECAPx6_ASAP7_75t_R FILLER_43_124 ();
 FILLER_ASAP7_75t_R FILLER_43_138 ();
 DECAPx4_ASAP7_75t_R FILLER_43_152 ();
 FILLER_ASAP7_75t_R FILLER_43_162 ();
 DECAPx6_ASAP7_75t_R FILLER_43_170 ();
 DECAPx10_ASAP7_75t_R FILLER_43_196 ();
 DECAPx10_ASAP7_75t_R FILLER_43_218 ();
 DECAPx6_ASAP7_75t_R FILLER_43_240 ();
 FILLER_ASAP7_75t_R FILLER_43_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_256 ();
 DECAPx4_ASAP7_75t_R FILLER_43_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_287 ();
 DECAPx2_ASAP7_75t_R FILLER_43_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_324 ();
 DECAPx4_ASAP7_75t_R FILLER_44_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_12 ();
 DECAPx2_ASAP7_75t_R FILLER_44_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_37 ();
 FILLER_ASAP7_75t_R FILLER_44_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_97 ();
 FILLER_ASAP7_75t_R FILLER_44_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_120 ();
 FILLER_ASAP7_75t_R FILLER_44_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_162 ();
 DECAPx6_ASAP7_75t_R FILLER_44_169 ();
 DECAPx2_ASAP7_75t_R FILLER_44_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_213 ();
 DECAPx10_ASAP7_75t_R FILLER_44_226 ();
 DECAPx10_ASAP7_75t_R FILLER_44_248 ();
 DECAPx6_ASAP7_75t_R FILLER_44_270 ();
 FILLER_ASAP7_75t_R FILLER_44_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_286 ();
 FILLER_ASAP7_75t_R FILLER_44_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_302 ();
 DECAPx1_ASAP7_75t_R FILLER_44_327 ();
 DECAPx2_ASAP7_75t_R FILLER_45_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_20 ();
 DECAPx1_ASAP7_75t_R FILLER_45_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_47 ();
 DECAPx1_ASAP7_75t_R FILLER_45_54 ();
 DECAPx1_ASAP7_75t_R FILLER_45_78 ();
 DECAPx10_ASAP7_75t_R FILLER_45_94 ();
 DECAPx10_ASAP7_75t_R FILLER_45_116 ();
 DECAPx2_ASAP7_75t_R FILLER_45_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_144 ();
 DECAPx2_ASAP7_75t_R FILLER_45_151 ();
 DECAPx6_ASAP7_75t_R FILLER_45_167 ();
 DECAPx4_ASAP7_75t_R FILLER_45_203 ();
 FILLER_ASAP7_75t_R FILLER_45_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_221 ();
 DECAPx6_ASAP7_75t_R FILLER_45_234 ();
 DECAPx1_ASAP7_75t_R FILLER_45_248 ();
 DECAPx10_ASAP7_75t_R FILLER_45_262 ();
 DECAPx2_ASAP7_75t_R FILLER_45_290 ();
 FILLER_ASAP7_75t_R FILLER_45_314 ();
 FILLER_ASAP7_75t_R FILLER_45_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_330 ();
 DECAPx4_ASAP7_75t_R FILLER_46_2 ();
 FILLER_ASAP7_75t_R FILLER_46_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_14 ();
 DECAPx10_ASAP7_75t_R FILLER_46_26 ();
 DECAPx10_ASAP7_75t_R FILLER_46_48 ();
 DECAPx10_ASAP7_75t_R FILLER_46_70 ();
 DECAPx10_ASAP7_75t_R FILLER_46_92 ();
 DECAPx6_ASAP7_75t_R FILLER_46_114 ();
 DECAPx2_ASAP7_75t_R FILLER_46_128 ();
 DECAPx4_ASAP7_75t_R FILLER_46_146 ();
 FILLER_ASAP7_75t_R FILLER_46_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_158 ();
 DECAPx4_ASAP7_75t_R FILLER_46_177 ();
 DECAPx4_ASAP7_75t_R FILLER_46_199 ();
 DECAPx6_ASAP7_75t_R FILLER_46_225 ();
 DECAPx1_ASAP7_75t_R FILLER_46_239 ();
 DECAPx1_ASAP7_75t_R FILLER_46_253 ();
 DECAPx4_ASAP7_75t_R FILLER_46_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_277 ();
 DECAPx2_ASAP7_75t_R FILLER_46_312 ();
 DECAPx2_ASAP7_75t_R FILLER_46_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_336 ();
 DECAPx1_ASAP7_75t_R FILLER_47_17 ();
 DECAPx4_ASAP7_75t_R FILLER_47_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_59 ();
 FILLER_ASAP7_75t_R FILLER_47_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_73 ();
 FILLER_ASAP7_75t_R FILLER_47_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_96 ();
 DECAPx6_ASAP7_75t_R FILLER_47_117 ();
 FILLER_ASAP7_75t_R FILLER_47_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_133 ();
 DECAPx1_ASAP7_75t_R FILLER_47_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_150 ();
 FILLER_ASAP7_75t_R FILLER_47_157 ();
 FILLER_ASAP7_75t_R FILLER_47_165 ();
 DECAPx1_ASAP7_75t_R FILLER_47_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_183 ();
 DECAPx4_ASAP7_75t_R FILLER_47_190 ();
 FILLER_ASAP7_75t_R FILLER_47_200 ();
 DECAPx4_ASAP7_75t_R FILLER_47_208 ();
 FILLER_ASAP7_75t_R FILLER_47_218 ();
 FILLER_ASAP7_75t_R FILLER_47_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_234 ();
 DECAPx6_ASAP7_75t_R FILLER_47_265 ();
 FILLER_ASAP7_75t_R FILLER_47_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_330 ();
 FILLER_ASAP7_75t_R FILLER_48_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_4 ();
 DECAPx1_ASAP7_75t_R FILLER_48_19 ();
 DECAPx2_ASAP7_75t_R FILLER_48_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_93 ();
 DECAPx1_ASAP7_75t_R FILLER_48_100 ();
 DECAPx6_ASAP7_75t_R FILLER_48_107 ();
 FILLER_ASAP7_75t_R FILLER_48_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_148 ();
 DECAPx10_ASAP7_75t_R FILLER_48_155 ();
 DECAPx4_ASAP7_75t_R FILLER_48_177 ();
 FILLER_ASAP7_75t_R FILLER_48_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_195 ();
 DECAPx4_ASAP7_75t_R FILLER_48_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_225 ();
 DECAPx1_ASAP7_75t_R FILLER_48_232 ();
 DECAPx2_ASAP7_75t_R FILLER_48_246 ();
 FILLER_ASAP7_75t_R FILLER_48_252 ();
 DECAPx2_ASAP7_75t_R FILLER_48_264 ();
 FILLER_ASAP7_75t_R FILLER_48_270 ();
 FILLER_ASAP7_75t_R FILLER_48_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_284 ();
 DECAPx1_ASAP7_75t_R FILLER_48_291 ();
 DECAPx1_ASAP7_75t_R FILLER_49_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_25 ();
 DECAPx10_ASAP7_75t_R FILLER_49_38 ();
 DECAPx6_ASAP7_75t_R FILLER_49_60 ();
 FILLER_ASAP7_75t_R FILLER_49_74 ();
 DECAPx4_ASAP7_75t_R FILLER_49_102 ();
 FILLER_ASAP7_75t_R FILLER_49_144 ();
 FILLER_ASAP7_75t_R FILLER_49_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_167 ();
 DECAPx2_ASAP7_75t_R FILLER_49_174 ();
 FILLER_ASAP7_75t_R FILLER_49_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_199 ();
 DECAPx1_ASAP7_75t_R FILLER_49_212 ();
 DECAPx10_ASAP7_75t_R FILLER_49_222 ();
 DECAPx2_ASAP7_75t_R FILLER_49_244 ();
 FILLER_ASAP7_75t_R FILLER_49_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_252 ();
 DECAPx6_ASAP7_75t_R FILLER_49_265 ();
 DECAPx2_ASAP7_75t_R FILLER_49_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_285 ();
 FILLER_ASAP7_75t_R FILLER_49_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_306 ();
 DECAPx1_ASAP7_75t_R FILLER_50_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_6 ();
 FILLER_ASAP7_75t_R FILLER_50_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_25 ();
 DECAPx2_ASAP7_75t_R FILLER_50_41 ();
 DECAPx4_ASAP7_75t_R FILLER_50_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_68 ();
 DECAPx4_ASAP7_75t_R FILLER_50_81 ();
 DECAPx4_ASAP7_75t_R FILLER_50_97 ();
 FILLER_ASAP7_75t_R FILLER_50_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_109 ();
 DECAPx4_ASAP7_75t_R FILLER_50_124 ();
 FILLER_ASAP7_75t_R FILLER_50_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_136 ();
 DECAPx4_ASAP7_75t_R FILLER_50_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_183 ();
 DECAPx1_ASAP7_75t_R FILLER_50_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_194 ();
 DECAPx4_ASAP7_75t_R FILLER_50_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_211 ();
 DECAPx10_ASAP7_75t_R FILLER_50_230 ();
 DECAPx2_ASAP7_75t_R FILLER_50_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_320 ();
 FILLER_ASAP7_75t_R FILLER_50_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_336 ();
 DECAPx1_ASAP7_75t_R FILLER_51_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_6 ();
 DECAPx1_ASAP7_75t_R FILLER_51_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_22 ();
 FILLER_ASAP7_75t_R FILLER_51_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_31 ();
 DECAPx2_ASAP7_75t_R FILLER_51_38 ();
 FILLER_ASAP7_75t_R FILLER_51_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_46 ();
 DECAPx2_ASAP7_75t_R FILLER_51_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_97 ();
 FILLER_ASAP7_75t_R FILLER_51_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_111 ();
 DECAPx4_ASAP7_75t_R FILLER_51_118 ();
 FILLER_ASAP7_75t_R FILLER_51_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_130 ();
 DECAPx1_ASAP7_75t_R FILLER_51_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_159 ();
 DECAPx2_ASAP7_75t_R FILLER_51_172 ();
 FILLER_ASAP7_75t_R FILLER_51_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_180 ();
 DECAPx4_ASAP7_75t_R FILLER_51_199 ();
 FILLER_ASAP7_75t_R FILLER_51_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_211 ();
 DECAPx6_ASAP7_75t_R FILLER_51_234 ();
 FILLER_ASAP7_75t_R FILLER_51_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_250 ();
 FILLER_ASAP7_75t_R FILLER_51_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_330 ();
 DECAPx1_ASAP7_75t_R FILLER_52_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_12 ();
 FILLER_ASAP7_75t_R FILLER_52_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_40 ();
 DECAPx10_ASAP7_75t_R FILLER_52_57 ();
 DECAPx2_ASAP7_75t_R FILLER_52_79 ();
 FILLER_ASAP7_75t_R FILLER_52_85 ();
 DECAPx4_ASAP7_75t_R FILLER_52_129 ();
 FILLER_ASAP7_75t_R FILLER_52_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_148 ();
 FILLER_ASAP7_75t_R FILLER_52_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_169 ();
 FILLER_ASAP7_75t_R FILLER_52_180 ();
 DECAPx2_ASAP7_75t_R FILLER_52_192 ();
 FILLER_ASAP7_75t_R FILLER_52_198 ();
 DECAPx1_ASAP7_75t_R FILLER_52_212 ();
 DECAPx10_ASAP7_75t_R FILLER_52_228 ();
 FILLER_ASAP7_75t_R FILLER_52_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_252 ();
 FILLER_ASAP7_75t_R FILLER_52_259 ();
 FILLER_ASAP7_75t_R FILLER_52_273 ();
 DECAPx1_ASAP7_75t_R FILLER_52_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_285 ();
 FILLER_ASAP7_75t_R FILLER_52_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_330 ();
 DECAPx2_ASAP7_75t_R FILLER_53_2 ();
 FILLER_ASAP7_75t_R FILLER_53_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_10 ();
 FILLER_ASAP7_75t_R FILLER_53_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_20 ();
 DECAPx4_ASAP7_75t_R FILLER_53_58 ();
 FILLER_ASAP7_75t_R FILLER_53_68 ();
 DECAPx4_ASAP7_75t_R FILLER_53_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_98 ();
 DECAPx4_ASAP7_75t_R FILLER_53_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_136 ();
 DECAPx1_ASAP7_75t_R FILLER_53_165 ();
 FILLER_ASAP7_75t_R FILLER_53_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_181 ();
 DECAPx1_ASAP7_75t_R FILLER_53_188 ();
 DECAPx4_ASAP7_75t_R FILLER_53_204 ();
 DECAPx6_ASAP7_75t_R FILLER_53_226 ();
 DECAPx1_ASAP7_75t_R FILLER_53_240 ();
 FILLER_ASAP7_75t_R FILLER_53_268 ();
 DECAPx1_ASAP7_75t_R FILLER_53_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_292 ();
 FILLER_ASAP7_75t_R FILLER_53_323 ();
 DECAPx4_ASAP7_75t_R FILLER_54_2 ();
 FILLER_ASAP7_75t_R FILLER_54_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_14 ();
 DECAPx10_ASAP7_75t_R FILLER_54_35 ();
 DECAPx2_ASAP7_75t_R FILLER_54_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_63 ();
 DECAPx2_ASAP7_75t_R FILLER_54_86 ();
 FILLER_ASAP7_75t_R FILLER_54_92 ();
 DECAPx2_ASAP7_75t_R FILLER_54_100 ();
 DECAPx6_ASAP7_75t_R FILLER_54_120 ();
 DECAPx1_ASAP7_75t_R FILLER_54_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_138 ();
 DECAPx10_ASAP7_75t_R FILLER_54_145 ();
 DECAPx6_ASAP7_75t_R FILLER_54_167 ();
 DECAPx1_ASAP7_75t_R FILLER_54_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_185 ();
 DECAPx10_ASAP7_75t_R FILLER_54_198 ();
 DECAPx6_ASAP7_75t_R FILLER_54_220 ();
 DECAPx1_ASAP7_75t_R FILLER_54_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_238 ();
 FILLER_ASAP7_75t_R FILLER_54_287 ();
 DECAPx6_ASAP7_75t_R FILLER_55_2 ();
 DECAPx1_ASAP7_75t_R FILLER_55_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_20 ();
 DECAPx10_ASAP7_75t_R FILLER_55_55 ();
 DECAPx4_ASAP7_75t_R FILLER_55_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_99 ();
 DECAPx1_ASAP7_75t_R FILLER_55_119 ();
 DECAPx10_ASAP7_75t_R FILLER_55_135 ();
 DECAPx10_ASAP7_75t_R FILLER_55_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_179 ();
 DECAPx6_ASAP7_75t_R FILLER_55_198 ();
 DECAPx2_ASAP7_75t_R FILLER_55_212 ();
 DECAPx1_ASAP7_75t_R FILLER_55_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_228 ();
 DECAPx2_ASAP7_75t_R FILLER_55_241 ();
 FILLER_ASAP7_75t_R FILLER_55_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_280 ();
 FILLER_ASAP7_75t_R FILLER_55_299 ();
 DECAPx10_ASAP7_75t_R FILLER_56_2 ();
 DECAPx10_ASAP7_75t_R FILLER_56_24 ();
 DECAPx10_ASAP7_75t_R FILLER_56_46 ();
 DECAPx2_ASAP7_75t_R FILLER_56_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_74 ();
 DECAPx6_ASAP7_75t_R FILLER_56_97 ();
 DECAPx2_ASAP7_75t_R FILLER_56_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_128 ();
 DECAPx10_ASAP7_75t_R FILLER_56_151 ();
 DECAPx2_ASAP7_75t_R FILLER_56_173 ();
 FILLER_ASAP7_75t_R FILLER_56_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_199 ();
 DECAPx2_ASAP7_75t_R FILLER_56_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_218 ();
 FILLER_ASAP7_75t_R FILLER_56_225 ();
 DECAPx2_ASAP7_75t_R FILLER_56_233 ();
 FILLER_ASAP7_75t_R FILLER_56_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_247 ();
 FILLER_ASAP7_75t_R FILLER_56_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_304 ();
 FILLER_ASAP7_75t_R FILLER_56_335 ();
 DECAPx10_ASAP7_75t_R FILLER_57_2 ();
 DECAPx10_ASAP7_75t_R FILLER_57_24 ();
 DECAPx10_ASAP7_75t_R FILLER_57_46 ();
 DECAPx6_ASAP7_75t_R FILLER_57_68 ();
 FILLER_ASAP7_75t_R FILLER_57_82 ();
 DECAPx1_ASAP7_75t_R FILLER_57_104 ();
 DECAPx1_ASAP7_75t_R FILLER_57_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_115 ();
 FILLER_ASAP7_75t_R FILLER_57_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_190 ();
 FILLER_ASAP7_75t_R FILLER_57_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_199 ();
 FILLER_ASAP7_75t_R FILLER_57_212 ();
 FILLER_ASAP7_75t_R FILLER_57_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_246 ();
 DECAPx2_ASAP7_75t_R FILLER_57_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_291 ();
 FILLER_ASAP7_75t_R FILLER_57_298 ();
 FILLER_ASAP7_75t_R FILLER_57_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_315 ();
 FILLER_ASAP7_75t_R FILLER_57_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_324 ();
 DECAPx10_ASAP7_75t_R FILLER_58_2 ();
 DECAPx10_ASAP7_75t_R FILLER_58_24 ();
 DECAPx10_ASAP7_75t_R FILLER_58_46 ();
 DECAPx10_ASAP7_75t_R FILLER_58_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_102 ();
 DECAPx1_ASAP7_75t_R FILLER_58_129 ();
 FILLER_ASAP7_75t_R FILLER_58_151 ();
 DECAPx10_ASAP7_75t_R FILLER_58_159 ();
 FILLER_ASAP7_75t_R FILLER_58_181 ();
 DECAPx1_ASAP7_75t_R FILLER_58_195 ();
 DECAPx2_ASAP7_75t_R FILLER_58_205 ();
 FILLER_ASAP7_75t_R FILLER_58_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_213 ();
 FILLER_ASAP7_75t_R FILLER_58_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_247 ();
 FILLER_ASAP7_75t_R FILLER_58_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_274 ();
 DECAPx1_ASAP7_75t_R FILLER_58_303 ();
 DECAPx10_ASAP7_75t_R FILLER_59_2 ();
 DECAPx10_ASAP7_75t_R FILLER_59_24 ();
 DECAPx10_ASAP7_75t_R FILLER_59_46 ();
 DECAPx10_ASAP7_75t_R FILLER_59_68 ();
 DECAPx6_ASAP7_75t_R FILLER_59_90 ();
 FILLER_ASAP7_75t_R FILLER_59_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_106 ();
 FILLER_ASAP7_75t_R FILLER_59_116 ();
 DECAPx6_ASAP7_75t_R FILLER_59_125 ();
 DECAPx1_ASAP7_75t_R FILLER_59_139 ();
 DECAPx10_ASAP7_75t_R FILLER_59_149 ();
 DECAPx10_ASAP7_75t_R FILLER_59_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_193 ();
 FILLER_ASAP7_75t_R FILLER_59_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_202 ();
 FILLER_ASAP7_75t_R FILLER_59_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_221 ();
 DECAPx1_ASAP7_75t_R FILLER_59_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_250 ();
 DECAPx1_ASAP7_75t_R FILLER_59_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_291 ();
 DECAPx1_ASAP7_75t_R FILLER_59_298 ();
 DECAPx2_ASAP7_75t_R FILLER_59_308 ();
 DECAPx1_ASAP7_75t_R FILLER_59_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_330 ();
 DECAPx10_ASAP7_75t_R FILLER_60_2 ();
 DECAPx10_ASAP7_75t_R FILLER_60_24 ();
 DECAPx10_ASAP7_75t_R FILLER_60_46 ();
 DECAPx10_ASAP7_75t_R FILLER_60_68 ();
 DECAPx6_ASAP7_75t_R FILLER_60_90 ();
 DECAPx2_ASAP7_75t_R FILLER_60_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_110 ();
 DECAPx6_ASAP7_75t_R FILLER_60_119 ();
 DECAPx1_ASAP7_75t_R FILLER_60_133 ();
 DECAPx10_ASAP7_75t_R FILLER_60_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_165 ();
 DECAPx4_ASAP7_75t_R FILLER_60_172 ();
 FILLER_ASAP7_75t_R FILLER_60_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_184 ();
 DECAPx1_ASAP7_75t_R FILLER_60_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_208 ();
 DECAPx2_ASAP7_75t_R FILLER_60_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_251 ();
 FILLER_ASAP7_75t_R FILLER_60_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_330 ();
 DECAPx10_ASAP7_75t_R FILLER_61_2 ();
 DECAPx10_ASAP7_75t_R FILLER_61_24 ();
 DECAPx10_ASAP7_75t_R FILLER_61_46 ();
 DECAPx10_ASAP7_75t_R FILLER_61_68 ();
 DECAPx10_ASAP7_75t_R FILLER_61_90 ();
 DECAPx10_ASAP7_75t_R FILLER_61_112 ();
 DECAPx2_ASAP7_75t_R FILLER_61_152 ();
 DECAPx1_ASAP7_75t_R FILLER_61_170 ();
 DECAPx2_ASAP7_75t_R FILLER_61_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_202 ();
 FILLER_ASAP7_75t_R FILLER_61_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_217 ();
 FILLER_ASAP7_75t_R FILLER_61_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_230 ();
 DECAPx2_ASAP7_75t_R FILLER_61_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_286 ();
 DECAPx2_ASAP7_75t_R FILLER_61_303 ();
 DECAPx1_ASAP7_75t_R FILLER_61_315 ();
 DECAPx10_ASAP7_75t_R FILLER_62_2 ();
 DECAPx10_ASAP7_75t_R FILLER_62_24 ();
 DECAPx10_ASAP7_75t_R FILLER_62_46 ();
 DECAPx4_ASAP7_75t_R FILLER_62_68 ();
 FILLER_ASAP7_75t_R FILLER_62_78 ();
 DECAPx6_ASAP7_75t_R FILLER_62_86 ();
 FILLER_ASAP7_75t_R FILLER_62_100 ();
 FILLER_ASAP7_75t_R FILLER_62_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_110 ();
 DECAPx2_ASAP7_75t_R FILLER_62_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_123 ();
 DECAPx2_ASAP7_75t_R FILLER_62_148 ();
 FILLER_ASAP7_75t_R FILLER_62_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_156 ();
 FILLER_ASAP7_75t_R FILLER_62_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_165 ();
 FILLER_ASAP7_75t_R FILLER_62_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_174 ();
 DECAPx6_ASAP7_75t_R FILLER_62_187 ();
 DECAPx2_ASAP7_75t_R FILLER_62_207 ();
 FILLER_ASAP7_75t_R FILLER_62_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_259 ();
 FILLER_ASAP7_75t_R FILLER_62_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_274 ();
 DECAPx1_ASAP7_75t_R FILLER_62_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_291 ();
 FILLER_ASAP7_75t_R FILLER_62_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_330 ();
 DECAPx10_ASAP7_75t_R FILLER_63_2 ();
 DECAPx10_ASAP7_75t_R FILLER_63_24 ();
 DECAPx10_ASAP7_75t_R FILLER_63_46 ();
 DECAPx4_ASAP7_75t_R FILLER_63_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_78 ();
 DECAPx6_ASAP7_75t_R FILLER_63_85 ();
 DECAPx1_ASAP7_75t_R FILLER_63_99 ();
 FILLER_ASAP7_75t_R FILLER_63_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_117 ();
 FILLER_ASAP7_75t_R FILLER_63_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_176 ();
 DECAPx2_ASAP7_75t_R FILLER_63_183 ();
 DECAPx2_ASAP7_75t_R FILLER_63_195 ();
 FILLER_ASAP7_75t_R FILLER_63_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_221 ();
 FILLER_ASAP7_75t_R FILLER_63_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_230 ();
 FILLER_ASAP7_75t_R FILLER_63_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_272 ();
 FILLER_ASAP7_75t_R FILLER_63_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_330 ();
 DECAPx10_ASAP7_75t_R FILLER_64_2 ();
 DECAPx10_ASAP7_75t_R FILLER_64_24 ();
 DECAPx10_ASAP7_75t_R FILLER_64_46 ();
 DECAPx1_ASAP7_75t_R FILLER_64_68 ();
 FILLER_ASAP7_75t_R FILLER_64_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_80 ();
 FILLER_ASAP7_75t_R FILLER_64_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_107 ();
 FILLER_ASAP7_75t_R FILLER_64_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_122 ();
 DECAPx1_ASAP7_75t_R FILLER_64_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_139 ();
 FILLER_ASAP7_75t_R FILLER_64_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_191 ();
 DECAPx2_ASAP7_75t_R FILLER_64_198 ();
 FILLER_ASAP7_75t_R FILLER_64_204 ();
 DECAPx1_ASAP7_75t_R FILLER_64_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_324 ();
 DECAPx10_ASAP7_75t_R FILLER_65_2 ();
 DECAPx10_ASAP7_75t_R FILLER_65_24 ();
 DECAPx6_ASAP7_75t_R FILLER_65_46 ();
 FILLER_ASAP7_75t_R FILLER_65_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_336 ();
 DECAPx10_ASAP7_75t_R FILLER_66_2 ();
 DECAPx10_ASAP7_75t_R FILLER_66_24 ();
 DECAPx4_ASAP7_75t_R FILLER_66_46 ();
 FILLER_ASAP7_75t_R FILLER_66_56 ();
 DECAPx1_ASAP7_75t_R FILLER_66_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_81 ();
 FILLER_ASAP7_75t_R FILLER_66_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_108 ();
 DECAPx1_ASAP7_75t_R FILLER_66_115 ();
 DECAPx1_ASAP7_75t_R FILLER_66_131 ();
 FILLER_ASAP7_75t_R FILLER_66_141 ();
 FILLER_ASAP7_75t_R FILLER_66_167 ();
 FILLER_ASAP7_75t_R FILLER_66_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_183 ();
 FILLER_ASAP7_75t_R FILLER_66_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_336 ();
endmodule
