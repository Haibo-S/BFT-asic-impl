module ibex_core (alert_major_o,
    alert_minor_o,
    clk_i,
    core_sleep_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_nm_i,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    hart_id_i,
    instr_addr_o,
    instr_rdata_i,
    irq_fast_i);
 output alert_major_o;
 output alert_minor_o;
 input clk_i;
 output core_sleep_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_nm_i;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 input [31:0] hart_id_i;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [14:0] irq_fast_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire net1975;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire _18110_;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire _18328_;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire _18403_;
 wire _18404_;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire _18412_;
 wire _18413_;
 wire _18414_;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire _18429_;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire _18438_;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire _18454_;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire _18461_;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire _18521_;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire _18609_;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire _18622_;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire _18628_;
 wire _18629_;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire _18652_;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire _18660_;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire _18664_;
 wire _18665_;
 wire _18666_;
 wire _18667_;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire _18686_;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire _18700_;
 wire _18701_;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire _18709_;
 wire _18710_;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire clk_i_regs;
 wire net277;
 wire \alu_adder_result_ex[0] ;
 wire \alu_adder_result_ex[10] ;
 wire \alu_adder_result_ex[11] ;
 wire \alu_adder_result_ex[12] ;
 wire \alu_adder_result_ex[13] ;
 wire \alu_adder_result_ex[14] ;
 wire \alu_adder_result_ex[15] ;
 wire \alu_adder_result_ex[16] ;
 wire \alu_adder_result_ex[17] ;
 wire \alu_adder_result_ex[18] ;
 wire \alu_adder_result_ex[19] ;
 wire \alu_adder_result_ex[1] ;
 wire \alu_adder_result_ex[20] ;
 wire \alu_adder_result_ex[21] ;
 wire \alu_adder_result_ex[22] ;
 wire \alu_adder_result_ex[23] ;
 wire \alu_adder_result_ex[24] ;
 wire \alu_adder_result_ex[25] ;
 wire \alu_adder_result_ex[26] ;
 wire \alu_adder_result_ex[27] ;
 wire \alu_adder_result_ex[28] ;
 wire \alu_adder_result_ex[29] ;
 wire \alu_adder_result_ex[2] ;
 wire \alu_adder_result_ex[30] ;
 wire \alu_adder_result_ex[31] ;
 wire \alu_adder_result_ex[3] ;
 wire \alu_adder_result_ex[4] ;
 wire \alu_adder_result_ex[5] ;
 wire \alu_adder_result_ex[6] ;
 wire \alu_adder_result_ex[7] ;
 wire \alu_adder_result_ex[8] ;
 wire \alu_adder_result_ex[9] ;
 wire clk;
 wire core_busy_d;
 wire \core_clock_gate_i.en_latch ;
 wire net171;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[0] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[1] ;
 wire \cs_registers_i.mhpmcounter[1856] ;
 wire \cs_registers_i.mhpmcounter[1857] ;
 wire \cs_registers_i.pc_id_i[1] ;
 wire \cs_registers_i.pc_id_i[2] ;
 wire \cs_registers_i.pc_if_i[2] ;
 wire \cs_registers_i.priv_mode_id_o[0] ;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ;
 wire \id_stage_i.branch_set_d ;
 wire \id_stage_i.controller_i.exc_req_d ;
 wire \id_stage_i.controller_i.illegal_insn_d ;
 wire \id_stage_i.controller_i.load_err_i ;
 wire \id_stage_i.controller_i.store_err_i ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ;
 wire \if_stage_i.instr_valid_id_d ;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire clknet_0_clk_i;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_leaf_0_clk_i_regs;
 wire clknet_leaf_1_clk_i_regs;
 wire clknet_leaf_2_clk_i_regs;
 wire clknet_leaf_3_clk_i_regs;
 wire clknet_leaf_4_clk_i_regs;
 wire clknet_leaf_5_clk_i_regs;
 wire clknet_leaf_6_clk_i_regs;
 wire clknet_leaf_7_clk_i_regs;
 wire clknet_leaf_8_clk_i_regs;
 wire clknet_leaf_9_clk_i_regs;
 wire clknet_leaf_10_clk_i_regs;
 wire clknet_leaf_11_clk_i_regs;
 wire clknet_leaf_12_clk_i_regs;
 wire clknet_leaf_13_clk_i_regs;
 wire clknet_leaf_14_clk_i_regs;
 wire clknet_leaf_15_clk_i_regs;
 wire clknet_leaf_16_clk_i_regs;
 wire clknet_leaf_17_clk_i_regs;
 wire clknet_leaf_18_clk_i_regs;
 wire clknet_leaf_19_clk_i_regs;
 wire clknet_leaf_20_clk_i_regs;
 wire clknet_leaf_21_clk_i_regs;
 wire clknet_0_clk_i_regs;
 wire clknet_1_0__leaf_clk_i_regs;
 wire clknet_1_1__leaf_clk_i_regs;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire delaynet_0_core_clock;
 wire delaynet_1_core_clock;
 wire delaynet_2_core_clock;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1976;
 wire net1977;

 OA211x2_ASAP7_75t_R _18722_ (.A1(_15597_),
    .A2(_04250_),
    .B(_04316_),
    .C(_15266_),
    .Y(_04317_));
 NAND2x1_ASAP7_75t_R _18723_ (.A(net1958),
    .B(_01205_),
    .Y(_04318_));
 OA211x2_ASAP7_75t_R _18724_ (.A1(_15597_),
    .A2(_04253_),
    .B(_04318_),
    .C(_15274_),
    .Y(_04319_));
 OR3x1_ASAP7_75t_R _18725_ (.A(_15278_),
    .B(_04317_),
    .C(_04319_),
    .Y(_04320_));
 OA211x2_ASAP7_75t_R _18726_ (.A1(_16368_),
    .A2(_04315_),
    .B(_04320_),
    .C(_15312_),
    .Y(_04321_));
 NAND2x1_ASAP7_75t_R _18727_ (.A(_15306_),
    .B(_01202_),
    .Y(_04322_));
 OA211x2_ASAP7_75t_R _18728_ (.A1(_15734_),
    .A2(_04258_),
    .B(_04322_),
    .C(_16948_),
    .Y(_04323_));
 NAND2x1_ASAP7_75t_R _18729_ (.A(_15306_),
    .B(_01201_),
    .Y(_04324_));
 OA211x2_ASAP7_75t_R _18730_ (.A1(_15734_),
    .A2(_04261_),
    .B(_04324_),
    .C(_15294_),
    .Y(_04325_));
 OR3x1_ASAP7_75t_R _18731_ (.A(_15287_),
    .B(_04323_),
    .C(_04325_),
    .Y(_04326_));
 NAND2x1_ASAP7_75t_R _18732_ (.A(_15306_),
    .B(_01210_),
    .Y(_04327_));
 OA211x2_ASAP7_75t_R _18733_ (.A1(_15734_),
    .A2(_04265_),
    .B(_04327_),
    .C(_16948_),
    .Y(_04328_));
 NAND2x1_ASAP7_75t_R _18734_ (.A(_15306_),
    .B(_01209_),
    .Y(_04329_));
 OA211x2_ASAP7_75t_R _18735_ (.A1(_15483_),
    .A2(_04268_),
    .B(_04329_),
    .C(_15294_),
    .Y(_04330_));
 OR3x1_ASAP7_75t_R _18736_ (.A(_15336_),
    .B(_04328_),
    .C(_04330_),
    .Y(_04331_));
 AND3x1_ASAP7_75t_R _18737_ (.A(_15252_),
    .B(_04326_),
    .C(_04331_),
    .Y(_04332_));
 OR3x2_ASAP7_75t_R _18738_ (.A(_15251_),
    .B(_04321_),
    .C(_04332_),
    .Y(_04333_));
 NAND2x1_ASAP7_75t_R _18739_ (.A(_15485_),
    .B(_01218_),
    .Y(_04334_));
 OA211x2_ASAP7_75t_R _18740_ (.A1(_15340_),
    .A2(_04274_),
    .B(_04334_),
    .C(_16948_),
    .Y(_04335_));
 NAND2x1_ASAP7_75t_R _18741_ (.A(_15485_),
    .B(_01217_),
    .Y(_04336_));
 OA211x2_ASAP7_75t_R _18742_ (.A1(_15734_),
    .A2(_04277_),
    .B(_04336_),
    .C(_15294_),
    .Y(_04337_));
 OR3x1_ASAP7_75t_R _18743_ (.A(_15287_),
    .B(_04335_),
    .C(_04337_),
    .Y(_04338_));
 NAND2x1_ASAP7_75t_R _18744_ (.A(_15485_),
    .B(_01226_),
    .Y(_04339_));
 OA211x2_ASAP7_75t_R _18745_ (.A1(_15734_),
    .A2(_04281_),
    .B(_04339_),
    .C(_16948_),
    .Y(_04340_));
 NAND2x1_ASAP7_75t_R _18746_ (.A(_15306_),
    .B(_01225_),
    .Y(_04341_));
 OA211x2_ASAP7_75t_R _18747_ (.A1(_15734_),
    .A2(_04284_),
    .B(_04341_),
    .C(_15294_),
    .Y(_04342_));
 OR3x1_ASAP7_75t_R _18748_ (.A(_15336_),
    .B(_04340_),
    .C(_04342_),
    .Y(_04343_));
 AND3x1_ASAP7_75t_R _18749_ (.A(_15252_),
    .B(_04338_),
    .C(_04343_),
    .Y(_04344_));
 NOR2x1_ASAP7_75t_R _18750_ (.A(_15632_),
    .B(_01223_),
    .Y(_04345_));
 AO21x1_ASAP7_75t_R _18751_ (.A1(_15437_),
    .A2(_04289_),
    .B(_04345_),
    .Y(_04346_));
 NAND2x1_ASAP7_75t_R _18752_ (.A(_15485_),
    .B(_01222_),
    .Y(_04347_));
 OA211x2_ASAP7_75t_R _18753_ (.A1(_16109_),
    .A2(_04292_),
    .B(_04347_),
    .C(_16948_),
    .Y(_04348_));
 AO21x1_ASAP7_75t_R _18754_ (.A1(_16354_),
    .A2(_04346_),
    .B(_04348_),
    .Y(_04349_));
 NAND2x1_ASAP7_75t_R _18755_ (.A(net1968),
    .B(_01214_),
    .Y(_04350_));
 OA211x2_ASAP7_75t_R _18756_ (.A1(_15597_),
    .A2(_04296_),
    .B(_04350_),
    .C(_15266_),
    .Y(_04351_));
 NAND2x1_ASAP7_75t_R _18757_ (.A(net1968),
    .B(_01213_),
    .Y(_04352_));
 OA211x2_ASAP7_75t_R _18758_ (.A1(_15597_),
    .A2(_04299_),
    .B(_04352_),
    .C(_15274_),
    .Y(_04353_));
 OR3x1_ASAP7_75t_R _18759_ (.A(_15254_),
    .B(_04351_),
    .C(_04353_),
    .Y(_04354_));
 OA211x2_ASAP7_75t_R _18760_ (.A1(_15475_),
    .A2(_04349_),
    .B(_04354_),
    .C(_15312_),
    .Y(_04355_));
 OR3x2_ASAP7_75t_R _18761_ (.A(_15316_),
    .B(_04344_),
    .C(_04355_),
    .Y(_04356_));
 AND2x6_ASAP7_75t_R _18762_ (.A(_04333_),
    .B(_04356_),
    .Y(_04357_));
 INVx2_ASAP7_75t_R _18763_ (.A(_04357_),
    .Y(_04358_));
 OA211x2_ASAP7_75t_R _18764_ (.A1(_13837_),
    .A2(_16386_),
    .B(_16389_),
    .C(_15370_),
    .Y(_04359_));
 AOI21x1_ASAP7_75t_R _18765_ (.A1(_15250_),
    .A2(_04358_),
    .B(_04359_),
    .Y(_18684_));
 INVx1_ASAP7_75t_R _18766_ (.A(_18684_),
    .Y(_18682_));
 AND2x2_ASAP7_75t_R _18767_ (.A(_14756_),
    .B(_01769_),
    .Y(_04360_));
 AO21x1_ASAP7_75t_R _18768_ (.A1(_13092_),
    .A2(_01232_),
    .B(_04360_),
    .Y(_04361_));
 OAI22x1_ASAP7_75t_R _18769_ (.A1(_01231_),
    .A2(_13102_),
    .B1(_04361_),
    .B2(_14975_),
    .Y(_04362_));
 INVx2_ASAP7_75t_R _18770_ (.A(_01240_),
    .Y(_04363_));
 NAND2x1_ASAP7_75t_R _18771_ (.A(_13165_),
    .B(_01238_),
    .Y(_04364_));
 OA211x2_ASAP7_75t_R _18772_ (.A1(_13097_),
    .A2(_04363_),
    .B(_04364_),
    .C(_14914_),
    .Y(_04365_));
 INVx2_ASAP7_75t_R _18773_ (.A(_01239_),
    .Y(_04366_));
 NAND2x1_ASAP7_75t_R _18774_ (.A(_14697_),
    .B(_01237_),
    .Y(_04367_));
 OA211x2_ASAP7_75t_R _18775_ (.A1(_14360_),
    .A2(_04366_),
    .B(_04367_),
    .C(_14463_),
    .Y(_04368_));
 OR3x1_ASAP7_75t_R _18776_ (.A(_13105_),
    .B(_04365_),
    .C(_04368_),
    .Y(_04369_));
 OA211x2_ASAP7_75t_R _18777_ (.A1(_13086_),
    .A2(_04362_),
    .B(_04369_),
    .C(_14466_),
    .Y(_04370_));
 INVx2_ASAP7_75t_R _18778_ (.A(_01236_),
    .Y(_04371_));
 NAND2x1_ASAP7_75t_R _18779_ (.A(_14815_),
    .B(_01234_),
    .Y(_04372_));
 OA211x2_ASAP7_75t_R _18780_ (.A1(_14943_),
    .A2(_04371_),
    .B(_04372_),
    .C(_14494_),
    .Y(_04373_));
 INVx1_ASAP7_75t_R _18781_ (.A(_01235_),
    .Y(_04374_));
 NAND2x1_ASAP7_75t_R _18782_ (.A(_13189_),
    .B(_01233_),
    .Y(_04375_));
 OA211x2_ASAP7_75t_R _18783_ (.A1(_14496_),
    .A2(_04374_),
    .B(_04375_),
    .C(_14498_),
    .Y(_04376_));
 OR3x1_ASAP7_75t_R _18784_ (.A(_14489_),
    .B(_04373_),
    .C(_04376_),
    .Y(_04377_));
 INVx2_ASAP7_75t_R _18785_ (.A(_01244_),
    .Y(_04378_));
 NAND2x1_ASAP7_75t_R _18786_ (.A(_14492_),
    .B(_01242_),
    .Y(_04379_));
 OA211x2_ASAP7_75t_R _18787_ (.A1(_14491_),
    .A2(_04378_),
    .B(_04379_),
    .C(_14504_),
    .Y(_04380_));
 INVx2_ASAP7_75t_R _18788_ (.A(_01243_),
    .Y(_04381_));
 NAND2x1_ASAP7_75t_R _18789_ (.A(_13189_),
    .B(_01241_),
    .Y(_04382_));
 OA211x2_ASAP7_75t_R _18790_ (.A1(_14506_),
    .A2(_04381_),
    .B(_04382_),
    .C(_14498_),
    .Y(_04383_));
 OR3x1_ASAP7_75t_R _18791_ (.A(_14929_),
    .B(_04380_),
    .C(_04383_),
    .Y(_04384_));
 AND3x1_ASAP7_75t_R _18792_ (.A(_14488_),
    .B(_04377_),
    .C(_04384_),
    .Y(_04385_));
 OR3x2_ASAP7_75t_R _18793_ (.A(_14447_),
    .B(_04370_),
    .C(_04385_),
    .Y(_04386_));
 INVx1_ASAP7_75t_R _18794_ (.A(_01252_),
    .Y(_04387_));
 NAND2x1_ASAP7_75t_R _18795_ (.A(_14752_),
    .B(_01250_),
    .Y(_04388_));
 OA211x2_ASAP7_75t_R _18796_ (.A1(_14985_),
    .A2(_04387_),
    .B(_04388_),
    .C(_14923_),
    .Y(_04389_));
 INVx1_ASAP7_75t_R _18797_ (.A(_01251_),
    .Y(_04390_));
 NAND2x1_ASAP7_75t_R _18798_ (.A(_14815_),
    .B(_01249_),
    .Y(_04391_));
 OA211x2_ASAP7_75t_R _18799_ (.A1(_14491_),
    .A2(_04390_),
    .B(_04391_),
    .C(_14926_),
    .Y(_04392_));
 OR3x1_ASAP7_75t_R _18800_ (.A(_14489_),
    .B(_04389_),
    .C(_04392_),
    .Y(_04393_));
 INVx1_ASAP7_75t_R _18801_ (.A(_01260_),
    .Y(_04394_));
 NAND2x1_ASAP7_75t_R _18802_ (.A(_14808_),
    .B(_01258_),
    .Y(_04395_));
 OA211x2_ASAP7_75t_R _18803_ (.A1(_14921_),
    .A2(_04394_),
    .B(_04395_),
    .C(_14923_),
    .Y(_04396_));
 INVx1_ASAP7_75t_R _18804_ (.A(_01259_),
    .Y(_04397_));
 NAND2x1_ASAP7_75t_R _18805_ (.A(_14492_),
    .B(_01257_),
    .Y(_04398_));
 OA211x2_ASAP7_75t_R _18806_ (.A1(_14501_),
    .A2(_04397_),
    .B(_04398_),
    .C(_14926_),
    .Y(_04399_));
 OR3x1_ASAP7_75t_R _18807_ (.A(_14929_),
    .B(_04396_),
    .C(_04399_),
    .Y(_04400_));
 AND3x1_ASAP7_75t_R _18808_ (.A(_14488_),
    .B(_04393_),
    .C(_04400_),
    .Y(_04401_));
 INVx2_ASAP7_75t_R _18809_ (.A(_01253_),
    .Y(_04402_));
 NOR2x1_ASAP7_75t_R _18810_ (.A(_14717_),
    .B(_01255_),
    .Y(_04403_));
 AO21x1_ASAP7_75t_R _18811_ (.A1(_14358_),
    .A2(_04402_),
    .B(_04403_),
    .Y(_04404_));
 INVx2_ASAP7_75t_R _18812_ (.A(_01256_),
    .Y(_04405_));
 NAND2x1_ASAP7_75t_R _18813_ (.A(_14367_),
    .B(_01254_),
    .Y(_04406_));
 OA211x2_ASAP7_75t_R _18814_ (.A1(_14366_),
    .A2(_04405_),
    .B(_04406_),
    .C(_14369_),
    .Y(_04407_));
 AO21x1_ASAP7_75t_R _18815_ (.A1(_13187_),
    .A2(_04404_),
    .B(_04407_),
    .Y(_04408_));
 INVx2_ASAP7_75t_R _18816_ (.A(_01248_),
    .Y(_04409_));
 NAND2x1_ASAP7_75t_R _18817_ (.A(_14697_),
    .B(_01246_),
    .Y(_04410_));
 OA211x2_ASAP7_75t_R _18818_ (.A1(_14360_),
    .A2(_04409_),
    .B(_04410_),
    .C(_14914_),
    .Y(_04411_));
 INVx2_ASAP7_75t_R _18819_ (.A(_01247_),
    .Y(_04412_));
 NAND2x1_ASAP7_75t_R _18820_ (.A(_14697_),
    .B(_01245_),
    .Y(_04413_));
 OA211x2_ASAP7_75t_R _18821_ (.A1(_14455_),
    .A2(_04412_),
    .B(_04413_),
    .C(_14463_),
    .Y(_04414_));
 OR3x1_ASAP7_75t_R _18822_ (.A(_13085_),
    .B(_04411_),
    .C(_04414_),
    .Y(_04415_));
 OA211x2_ASAP7_75t_R _18823_ (.A1(_13186_),
    .A2(_04408_),
    .B(_04415_),
    .C(_14466_),
    .Y(_04416_));
 OR3x2_ASAP7_75t_R _18824_ (.A(_14487_),
    .B(_04401_),
    .C(_04416_),
    .Y(_04417_));
 AO21x2_ASAP7_75t_R _18825_ (.A1(_04386_),
    .A2(_04417_),
    .B(_14377_),
    .Y(_04418_));
 BUFx6f_ASAP7_75t_R _18826_ (.A(_01488_),
    .Y(_04419_));
 AND2x2_ASAP7_75t_R _18827_ (.A(_01458_),
    .B(_14381_),
    .Y(_04420_));
 OAI22x1_ASAP7_75t_R _18828_ (.A1(_04419_),
    .A2(_14967_),
    .B1(_14968_),
    .B2(_04420_),
    .Y(_04421_));
 NAND2x2_ASAP7_75t_R _18829_ (.A(_04418_),
    .B(_04421_),
    .Y(_18688_));
 INVx1_ASAP7_75t_R _18830_ (.A(_18688_),
    .Y(_18690_));
 BUFx6f_ASAP7_75t_R _18831_ (.A(_00161_),
    .Y(_04422_));
 OR3x1_ASAP7_75t_R _18832_ (.A(_04422_),
    .B(_14627_),
    .C(_14649_),
    .Y(_04423_));
 OAI21x1_ASAP7_75t_R _18833_ (.A1(_14646_),
    .A2(_18688_),
    .B(_04423_),
    .Y(_18062_));
 AND2x2_ASAP7_75t_R _18834_ (.A(_15437_),
    .B(_01769_),
    .Y(_04424_));
 AO21x1_ASAP7_75t_R _18835_ (.A1(_15436_),
    .A2(_01232_),
    .B(_04424_),
    .Y(_04425_));
 OAI22x1_ASAP7_75t_R _18836_ (.A1(_01231_),
    .A2(_15435_),
    .B1(_04425_),
    .B2(_15296_),
    .Y(_04426_));
 NAND2x1_ASAP7_75t_R _18837_ (.A(_15302_),
    .B(_01238_),
    .Y(_04427_));
 OA211x2_ASAP7_75t_R _18838_ (.A1(_15445_),
    .A2(_04363_),
    .B(_04427_),
    .C(_15443_),
    .Y(_04428_));
 NAND2x1_ASAP7_75t_R _18839_ (.A(_15302_),
    .B(_01237_),
    .Y(_04429_));
 OA211x2_ASAP7_75t_R _18840_ (.A1(_15445_),
    .A2(_04366_),
    .B(_04429_),
    .C(_15309_),
    .Y(_04430_));
 OR3x1_ASAP7_75t_R _18841_ (.A(_15298_),
    .B(_04428_),
    .C(_04430_),
    .Y(_04431_));
 OA211x2_ASAP7_75t_R _18842_ (.A1(_15288_),
    .A2(_04426_),
    .B(_04431_),
    .C(_15360_),
    .Y(_04432_));
 NAND2x1_ASAP7_75t_R _18843_ (.A(_15451_),
    .B(_01234_),
    .Y(_04433_));
 OA211x2_ASAP7_75t_R _18844_ (.A1(_15450_),
    .A2(_04371_),
    .B(_04433_),
    .C(_15323_),
    .Y(_04434_));
 NAND2x1_ASAP7_75t_R _18845_ (.A(_15454_),
    .B(_01233_),
    .Y(_04435_));
 OA211x2_ASAP7_75t_R _18846_ (.A1(_15320_),
    .A2(_04374_),
    .B(_04435_),
    .C(_15275_),
    .Y(_04436_));
 OR3x1_ASAP7_75t_R _18847_ (.A(_15318_),
    .B(_04434_),
    .C(_04436_),
    .Y(_04437_));
 NAND2x1_ASAP7_75t_R _18848_ (.A(_15454_),
    .B(_01242_),
    .Y(_04438_));
 OA211x2_ASAP7_75t_R _18849_ (.A1(_15450_),
    .A2(_04378_),
    .B(_04438_),
    .C(_15323_),
    .Y(_04439_));
 NAND2x1_ASAP7_75t_R _18850_ (.A(_16106_),
    .B(_01241_),
    .Y(_04440_));
 OA211x2_ASAP7_75t_R _18851_ (.A1(_15320_),
    .A2(_04381_),
    .B(_04440_),
    .C(_15275_),
    .Y(_04441_));
 OR3x1_ASAP7_75t_R _18852_ (.A(_15279_),
    .B(_04439_),
    .C(_04441_),
    .Y(_04442_));
 AND3x1_ASAP7_75t_R _18853_ (.A(_15317_),
    .B(_04437_),
    .C(_04442_),
    .Y(_04443_));
 OR3x2_ASAP7_75t_R _18854_ (.A(_15434_),
    .B(_04432_),
    .C(_04443_),
    .Y(_04444_));
 NAND2x1_ASAP7_75t_R _18855_ (.A(_15326_),
    .B(_01250_),
    .Y(_04445_));
 OA211x2_ASAP7_75t_R _18856_ (.A1(_15467_),
    .A2(_04387_),
    .B(_04445_),
    .C(_15349_),
    .Y(_04446_));
 NAND2x1_ASAP7_75t_R _18857_ (.A(_15262_),
    .B(_01249_),
    .Y(_04447_));
 OA211x2_ASAP7_75t_R _18858_ (.A1(_15471_),
    .A2(_04390_),
    .B(_04447_),
    .C(_15456_),
    .Y(_04448_));
 OR3x1_ASAP7_75t_R _18859_ (.A(_15318_),
    .B(_04446_),
    .C(_04448_),
    .Y(_04449_));
 NAND2x1_ASAP7_75t_R _18860_ (.A(_15326_),
    .B(_01258_),
    .Y(_04450_));
 OA211x2_ASAP7_75t_R _18861_ (.A1(_15471_),
    .A2(_04394_),
    .B(_04450_),
    .C(_15349_),
    .Y(_04451_));
 NAND2x1_ASAP7_75t_R _18862_ (.A(_15262_),
    .B(_01257_),
    .Y(_04452_));
 OA211x2_ASAP7_75t_R _18863_ (.A1(_15471_),
    .A2(_04397_),
    .B(_04452_),
    .C(_15456_),
    .Y(_04453_));
 OR3x1_ASAP7_75t_R _18864_ (.A(_15475_),
    .B(_04451_),
    .C(_04453_),
    .Y(_04454_));
 AND3x1_ASAP7_75t_R _18865_ (.A(_15317_),
    .B(_04449_),
    .C(_04454_),
    .Y(_04455_));
 NOR2x1_ASAP7_75t_R _18866_ (.A(_15486_),
    .B(_01255_),
    .Y(_04456_));
 AO21x1_ASAP7_75t_R _18867_ (.A1(_15484_),
    .A2(_04402_),
    .B(_04456_),
    .Y(_04457_));
 NAND2x1_ASAP7_75t_R _18868_ (.A(_15347_),
    .B(_01254_),
    .Y(_04458_));
 OA211x2_ASAP7_75t_R _18869_ (.A1(_15490_),
    .A2(_04405_),
    .B(_04458_),
    .C(_15469_),
    .Y(_04459_));
 AO21x1_ASAP7_75t_R _18870_ (.A1(_15339_),
    .A2(_04457_),
    .B(_04459_),
    .Y(_04460_));
 NAND2x1_ASAP7_75t_R _18871_ (.A(_15354_),
    .B(_01246_),
    .Y(_04461_));
 OA211x2_ASAP7_75t_R _18872_ (.A1(_15441_),
    .A2(_04409_),
    .B(_04461_),
    .C(_15443_),
    .Y(_04462_));
 NAND2x1_ASAP7_75t_R _18873_ (.A(_15354_),
    .B(_01245_),
    .Y(_04463_));
 OA211x2_ASAP7_75t_R _18874_ (.A1(_15441_),
    .A2(_04412_),
    .B(_04463_),
    .C(_15497_),
    .Y(_04464_));
 OR3x1_ASAP7_75t_R _18875_ (.A(_15352_),
    .B(_04462_),
    .C(_04464_),
    .Y(_04465_));
 OA211x2_ASAP7_75t_R _18876_ (.A1(_15482_),
    .A2(_04460_),
    .B(_04465_),
    .C(_15360_),
    .Y(_04466_));
 OR3x2_ASAP7_75t_R _18877_ (.A(_15466_),
    .B(_04455_),
    .C(_04466_),
    .Y(_04467_));
 NAND2x2_ASAP7_75t_R _18878_ (.A(_04444_),
    .B(_04467_),
    .Y(_04468_));
 OA211x2_ASAP7_75t_R _18879_ (.A1(_13909_),
    .A2(_16386_),
    .B(_16389_),
    .C(_15370_),
    .Y(_04469_));
 AOI21x1_ASAP7_75t_R _18880_ (.A1(_15250_),
    .A2(_04468_),
    .B(_04469_),
    .Y(_18689_));
 INVx1_ASAP7_75t_R _18881_ (.A(_18689_),
    .Y(_18687_));
 OA21x2_ASAP7_75t_R _18882_ (.A1(_01230_),
    .A2(_01229_),
    .B(_01262_),
    .Y(_04470_));
 AO21x1_ASAP7_75t_R _18883_ (.A1(_01133_),
    .A2(_01166_),
    .B(_01165_),
    .Y(_04471_));
 OR2x2_ASAP7_75t_R _18884_ (.A(_01197_),
    .B(_01229_),
    .Y(_04472_));
 AO21x1_ASAP7_75t_R _18885_ (.A1(_01198_),
    .A2(_04471_),
    .B(_04472_),
    .Y(_04473_));
 OA21x2_ASAP7_75t_R _18886_ (.A1(_01166_),
    .A2(_01165_),
    .B(_01198_),
    .Y(_04474_));
 AND3x1_ASAP7_75t_R _18887_ (.A(_01134_),
    .B(_04470_),
    .C(_04474_),
    .Y(_04475_));
 AO22x1_ASAP7_75t_R _18888_ (.A1(_04470_),
    .A2(_04473_),
    .B1(_04475_),
    .B2(_01101_),
    .Y(_04476_));
 AND4x1_ASAP7_75t_R _18889_ (.A(_16513_),
    .B(_16504_),
    .C(_16505_),
    .D(_16506_),
    .Y(_04477_));
 OA211x2_ASAP7_75t_R _18890_ (.A1(_16749_),
    .A2(_04477_),
    .B(_04475_),
    .C(_01102_),
    .Y(_04478_));
 OR2x2_ASAP7_75t_R _18891_ (.A(_04476_),
    .B(_04478_),
    .Y(_04479_));
 XNOR2x1_ASAP7_75t_R _18892_ (.B(_04479_),
    .Y(_04480_),
    .A(_01261_));
 INVx5_ASAP7_75t_R _18893_ (.A(_04480_),
    .Y(\alu_adder_result_ex[27] ));
 INVx1_ASAP7_75t_R _18894_ (.A(_01229_),
    .Y(_04481_));
 OA21x2_ASAP7_75t_R _18895_ (.A1(_01134_),
    .A2(_01133_),
    .B(_01166_),
    .Y(_04482_));
 OA21x2_ASAP7_75t_R _18896_ (.A1(_01165_),
    .A2(_04482_),
    .B(_01198_),
    .Y(_04483_));
 OA21x2_ASAP7_75t_R _18897_ (.A1(_01197_),
    .A2(_04483_),
    .B(_01230_),
    .Y(_04484_));
 AND3x1_ASAP7_75t_R _18898_ (.A(_04481_),
    .B(_16759_),
    .C(_04484_),
    .Y(_04485_));
 OA21x2_ASAP7_75t_R _18899_ (.A1(_16756_),
    .A2(_16758_),
    .B(_04485_),
    .Y(_04486_));
 OR3x2_ASAP7_75t_R _18900_ (.A(_01165_),
    .B(_01197_),
    .C(_04242_),
    .Y(_04487_));
 OR2x2_ASAP7_75t_R _18901_ (.A(_04481_),
    .B(_04487_),
    .Y(_04488_));
 NOR3x1_ASAP7_75t_R _18902_ (.A(_16756_),
    .B(_16758_),
    .C(_04488_),
    .Y(_04489_));
 NOR2x1_ASAP7_75t_R _18903_ (.A(_16759_),
    .B(_04487_),
    .Y(_04490_));
 INVx1_ASAP7_75t_R _18904_ (.A(_04484_),
    .Y(_04491_));
 AND3x1_ASAP7_75t_R _18905_ (.A(_04481_),
    .B(_04484_),
    .C(_04487_),
    .Y(_04492_));
 AO21x1_ASAP7_75t_R _18906_ (.A1(_01229_),
    .A2(_04491_),
    .B(_04492_),
    .Y(_04493_));
 AO21x2_ASAP7_75t_R _18907_ (.A1(_01229_),
    .A2(_04490_),
    .B(_04493_),
    .Y(_04494_));
 NOR3x2_ASAP7_75t_R _18908_ (.B(_04489_),
    .C(_04494_),
    .Y(_04495_),
    .A(_04486_));
 INVx5_ASAP7_75t_R _18909_ (.A(_04495_),
    .Y(\alu_adder_result_ex[26] ));
 INVx2_ASAP7_75t_R _18910_ (.A(_01285_),
    .Y(_04496_));
 NOR2x1_ASAP7_75t_R _18911_ (.A(_14717_),
    .B(_01287_),
    .Y(_04497_));
 AO21x1_ASAP7_75t_R _18912_ (.A1(_14358_),
    .A2(_04496_),
    .B(_04497_),
    .Y(_04498_));
 INVx2_ASAP7_75t_R _18913_ (.A(_01288_),
    .Y(_04499_));
 NAND2x1_ASAP7_75t_R _18914_ (.A(_14301_),
    .B(_01286_),
    .Y(_04500_));
 OA211x2_ASAP7_75t_R _18915_ (.A1(_14299_),
    .A2(_04499_),
    .B(_04500_),
    .C(_14369_),
    .Y(_04501_));
 AO21x1_ASAP7_75t_R _18916_ (.A1(_13187_),
    .A2(_04498_),
    .B(_04501_),
    .Y(_04502_));
 INVx2_ASAP7_75t_R _18917_ (.A(_01280_),
    .Y(_04503_));
 NAND2x1_ASAP7_75t_R _18918_ (.A(_14517_),
    .B(_01278_),
    .Y(_04504_));
 OA211x2_ASAP7_75t_R _18919_ (.A1(_14516_),
    .A2(_04503_),
    .B(_04504_),
    .C(_14472_),
    .Y(_04505_));
 INVx2_ASAP7_75t_R _18920_ (.A(_01279_),
    .Y(_04506_));
 NAND2x1_ASAP7_75t_R _18921_ (.A(_14470_),
    .B(_01277_),
    .Y(_04507_));
 OA211x2_ASAP7_75t_R _18922_ (.A1(_13193_),
    .A2(_04506_),
    .B(_04507_),
    .C(_14476_),
    .Y(_04508_));
 OA21x2_ASAP7_75t_R _18923_ (.A1(_04505_),
    .A2(_04508_),
    .B(_14291_),
    .Y(_04509_));
 AO21x1_ASAP7_75t_R _18924_ (.A1(_14448_),
    .A2(_04502_),
    .B(_04509_),
    .Y(_04510_));
 INVx2_ASAP7_75t_R _18925_ (.A(_01284_),
    .Y(_04511_));
 NAND2x1_ASAP7_75t_R _18926_ (.A(_13142_),
    .B(_01282_),
    .Y(_04512_));
 OA211x2_ASAP7_75t_R _18927_ (.A1(_14455_),
    .A2(_04511_),
    .B(_04512_),
    .C(_14458_),
    .Y(_04513_));
 INVx2_ASAP7_75t_R _18928_ (.A(_01283_),
    .Y(_04514_));
 NAND2x1_ASAP7_75t_R _18929_ (.A(_14292_),
    .B(_01281_),
    .Y(_04515_));
 OA211x2_ASAP7_75t_R _18930_ (.A1(_15052_),
    .A2(_04514_),
    .B(_04515_),
    .C(_14463_),
    .Y(_04516_));
 OR3x1_ASAP7_75t_R _18931_ (.A(_13085_),
    .B(_04513_),
    .C(_04516_),
    .Y(_04517_));
 INVx2_ASAP7_75t_R _18932_ (.A(_01292_),
    .Y(_04518_));
 NAND2x1_ASAP7_75t_R _18933_ (.A(_13142_),
    .B(_01290_),
    .Y(_04519_));
 OA211x2_ASAP7_75t_R _18934_ (.A1(_14461_),
    .A2(_04518_),
    .B(_04519_),
    .C(_14458_),
    .Y(_04520_));
 INVx2_ASAP7_75t_R _18935_ (.A(_01291_),
    .Y(_04521_));
 NAND2x1_ASAP7_75t_R _18936_ (.A(_14292_),
    .B(_01289_),
    .Y(_04522_));
 OA211x2_ASAP7_75t_R _18937_ (.A1(_15052_),
    .A2(_04521_),
    .B(_04522_),
    .C(_14463_),
    .Y(_04523_));
 OR3x1_ASAP7_75t_R _18938_ (.A(_14454_),
    .B(_04520_),
    .C(_04523_),
    .Y(_04524_));
 AND3x1_ASAP7_75t_R _18939_ (.A(_14468_),
    .B(_04517_),
    .C(_04524_),
    .Y(_04525_));
 AO21x1_ASAP7_75t_R _18940_ (.A1(_14778_),
    .A2(_04510_),
    .B(_04525_),
    .Y(_04526_));
 AND2x2_ASAP7_75t_R _18941_ (.A(_14678_),
    .B(_01768_),
    .Y(_04527_));
 AO21x1_ASAP7_75t_R _18942_ (.A1(_14285_),
    .A2(_01264_),
    .B(_04527_),
    .Y(_04528_));
 OAI22x1_ASAP7_75t_R _18943_ (.A1(_01263_),
    .A2(_13101_),
    .B1(_04528_),
    .B2(_14710_),
    .Y(_04529_));
 INVx2_ASAP7_75t_R _18944_ (.A(_01272_),
    .Y(_04530_));
 NAND2x1_ASAP7_75t_R _18945_ (.A(_13096_),
    .B(_01270_),
    .Y(_04531_));
 OA211x2_ASAP7_75t_R _18946_ (.A1(_14507_),
    .A2(_04530_),
    .B(_04531_),
    .C(_14762_),
    .Y(_04532_));
 INVx2_ASAP7_75t_R _18947_ (.A(_01271_),
    .Y(_04533_));
 NAND2x1_ASAP7_75t_R _18948_ (.A(_13096_),
    .B(_01269_),
    .Y(_04534_));
 OA211x2_ASAP7_75t_R _18949_ (.A1(_14517_),
    .A2(_04533_),
    .B(_04534_),
    .C(_14765_),
    .Y(_04535_));
 OR3x1_ASAP7_75t_R _18950_ (.A(_13185_),
    .B(_04532_),
    .C(_04535_),
    .Y(_04536_));
 OA211x2_ASAP7_75t_R _18951_ (.A1(_14448_),
    .A2(_04529_),
    .B(_04536_),
    .C(_14466_),
    .Y(_04537_));
 INVx1_ASAP7_75t_R _18952_ (.A(_01268_),
    .Y(_04538_));
 NAND2x1_ASAP7_75t_R _18953_ (.A(_14490_),
    .B(_01266_),
    .Y(_04539_));
 OA211x2_ASAP7_75t_R _18954_ (.A1(_13200_),
    .A2(_04538_),
    .B(_04539_),
    .C(_14740_),
    .Y(_04540_));
 INVx1_ASAP7_75t_R _18955_ (.A(_01267_),
    .Y(_04541_));
 NAND2x1_ASAP7_75t_R _18956_ (.A(_14490_),
    .B(_01265_),
    .Y(_04542_));
 OA211x2_ASAP7_75t_R _18957_ (.A1(_14653_),
    .A2(_04541_),
    .B(_04542_),
    .C(_14743_),
    .Y(_04543_));
 OR3x1_ASAP7_75t_R _18958_ (.A(_14737_),
    .B(_04540_),
    .C(_04543_),
    .Y(_04544_));
 INVx1_ASAP7_75t_R _18959_ (.A(_01276_),
    .Y(_04545_));
 NAND2x1_ASAP7_75t_R _18960_ (.A(_14490_),
    .B(_01274_),
    .Y(_04546_));
 OA211x2_ASAP7_75t_R _18961_ (.A1(_13200_),
    .A2(_04545_),
    .B(_04546_),
    .C(_14740_),
    .Y(_04547_));
 INVx2_ASAP7_75t_R _18962_ (.A(_01275_),
    .Y(_04548_));
 NAND2x1_ASAP7_75t_R _18963_ (.A(_13192_),
    .B(_01273_),
    .Y(_04549_));
 OA211x2_ASAP7_75t_R _18964_ (.A1(_14653_),
    .A2(_04548_),
    .B(_04549_),
    .C(_14732_),
    .Y(_04550_));
 OR3x1_ASAP7_75t_R _18965_ (.A(_14454_),
    .B(_04547_),
    .C(_04550_),
    .Y(_04551_));
 AND3x1_ASAP7_75t_R _18966_ (.A(_14468_),
    .B(_04544_),
    .C(_04551_),
    .Y(_04552_));
 OR3x1_ASAP7_75t_R _18967_ (.A(_14447_),
    .B(_04537_),
    .C(_04552_),
    .Y(_04553_));
 OA21x2_ASAP7_75t_R _18968_ (.A1(_14339_),
    .A2(_04526_),
    .B(_04553_),
    .Y(_04554_));
 AND2x2_ASAP7_75t_R _18969_ (.A(_01457_),
    .B(_14772_),
    .Y(_04555_));
 OAI22x1_ASAP7_75t_R _18970_ (.A1(_01487_),
    .A2(_14967_),
    .B1(_14968_),
    .B2(_04555_),
    .Y(_04556_));
 OA21x2_ASAP7_75t_R _18971_ (.A1(_14709_),
    .A2(_04554_),
    .B(_04556_),
    .Y(_04557_));
 BUFx6f_ASAP7_75t_R _18972_ (.A(_04557_),
    .Y(_18695_));
 INVx2_ASAP7_75t_R _18973_ (.A(_18695_),
    .Y(_18693_));
 BUFx6f_ASAP7_75t_R _18974_ (.A(_00169_),
    .Y(_04558_));
 INVx1_ASAP7_75t_R _18975_ (.A(_04558_),
    .Y(_04559_));
 AND3x1_ASAP7_75t_R _18976_ (.A(_04559_),
    .B(_14625_),
    .C(_14907_),
    .Y(_04560_));
 AO21x1_ASAP7_75t_R _18977_ (.A1(_14903_),
    .A2(_18695_),
    .B(_04560_),
    .Y(_18064_));
 AND2x2_ASAP7_75t_R _18978_ (.A(_15489_),
    .B(_01768_),
    .Y(_04561_));
 AO21x1_ASAP7_75t_R _18979_ (.A1(_15290_),
    .A2(_01264_),
    .B(_04561_),
    .Y(_04562_));
 OAI22x1_ASAP7_75t_R _18980_ (.A1(_01263_),
    .A2(_15289_),
    .B1(_04562_),
    .B2(_15593_),
    .Y(_04563_));
 NAND2x1_ASAP7_75t_R _18981_ (.A(_15306_),
    .B(_01270_),
    .Y(_04564_));
 OA211x2_ASAP7_75t_R _18982_ (.A1(_15354_),
    .A2(_04530_),
    .B(_04564_),
    .C(_16948_),
    .Y(_04565_));
 NAND2x1_ASAP7_75t_R _18983_ (.A(_15306_),
    .B(_01269_),
    .Y(_04566_));
 OA211x2_ASAP7_75t_R _18984_ (.A1(_15354_),
    .A2(_04533_),
    .B(_04566_),
    .C(_15294_),
    .Y(_04567_));
 OR3x1_ASAP7_75t_R _18985_ (.A(_15336_),
    .B(_04565_),
    .C(_04567_),
    .Y(_04568_));
 OA211x2_ASAP7_75t_R _18986_ (.A1(_16368_),
    .A2(_04563_),
    .B(_04568_),
    .C(_15312_),
    .Y(_04569_));
 NAND2x1_ASAP7_75t_R _18987_ (.A(_15259_),
    .B(_01266_),
    .Y(_04570_));
 OA211x2_ASAP7_75t_R _18988_ (.A1(_15262_),
    .A2(_04538_),
    .B(_04570_),
    .C(_15752_),
    .Y(_04571_));
 NAND2x1_ASAP7_75t_R _18989_ (.A(_15342_),
    .B(_01265_),
    .Y(_04572_));
 OA211x2_ASAP7_75t_R _18990_ (.A1(_15451_),
    .A2(_04541_),
    .B(_04572_),
    .C(_15592_),
    .Y(_04573_));
 OR3x1_ASAP7_75t_R _18991_ (.A(_15287_),
    .B(_04571_),
    .C(_04573_),
    .Y(_04574_));
 NAND2x1_ASAP7_75t_R _18992_ (.A(_15342_),
    .B(_01274_),
    .Y(_04575_));
 OA211x2_ASAP7_75t_R _18993_ (.A1(_15270_),
    .A2(_04545_),
    .B(_04575_),
    .C(_15752_),
    .Y(_04576_));
 NAND2x1_ASAP7_75t_R _18994_ (.A(_15342_),
    .B(_01273_),
    .Y(_04577_));
 OA211x2_ASAP7_75t_R _18995_ (.A1(_15451_),
    .A2(_04548_),
    .B(_04577_),
    .C(_15592_),
    .Y(_04578_));
 OR3x1_ASAP7_75t_R _18996_ (.A(_15336_),
    .B(_04576_),
    .C(_04578_),
    .Y(_04579_));
 AND3x1_ASAP7_75t_R _18997_ (.A(_15252_),
    .B(_04574_),
    .C(_04579_),
    .Y(_04580_));
 OR3x2_ASAP7_75t_R _18998_ (.A(_15251_),
    .B(_04569_),
    .C(_04580_),
    .Y(_04581_));
 NAND2x1_ASAP7_75t_R _18999_ (.A(_15259_),
    .B(_01282_),
    .Y(_04582_));
 OA211x2_ASAP7_75t_R _19000_ (.A1(_15262_),
    .A2(_04511_),
    .B(_04582_),
    .C(_15752_),
    .Y(_04583_));
 NAND2x1_ASAP7_75t_R _19001_ (.A(_15259_),
    .B(_01281_),
    .Y(_04584_));
 OA211x2_ASAP7_75t_R _19002_ (.A1(_15270_),
    .A2(_04514_),
    .B(_04584_),
    .C(_15592_),
    .Y(_04585_));
 OR3x1_ASAP7_75t_R _19003_ (.A(_15287_),
    .B(_04583_),
    .C(_04585_),
    .Y(_04586_));
 NAND2x1_ASAP7_75t_R _19004_ (.A(_15259_),
    .B(_01290_),
    .Y(_04587_));
 OA211x2_ASAP7_75t_R _19005_ (.A1(_15262_),
    .A2(_04518_),
    .B(_04587_),
    .C(_15752_),
    .Y(_04588_));
 NAND2x1_ASAP7_75t_R _19006_ (.A(_15342_),
    .B(_01289_),
    .Y(_04589_));
 OA211x2_ASAP7_75t_R _19007_ (.A1(_15270_),
    .A2(_04521_),
    .B(_04589_),
    .C(_15592_),
    .Y(_04590_));
 OR3x1_ASAP7_75t_R _19008_ (.A(_15336_),
    .B(_04588_),
    .C(_04590_),
    .Y(_04591_));
 AND3x1_ASAP7_75t_R _19009_ (.A(_15253_),
    .B(_04586_),
    .C(_04591_),
    .Y(_04592_));
 NOR2x1_ASAP7_75t_R _19010_ (.A(_15483_),
    .B(_01287_),
    .Y(_04593_));
 AO21x1_ASAP7_75t_R _19011_ (.A1(_15445_),
    .A2(_04496_),
    .B(_04593_),
    .Y(_04594_));
 NAND2x1_ASAP7_75t_R _19012_ (.A(_15259_),
    .B(_01286_),
    .Y(_04595_));
 OA211x2_ASAP7_75t_R _19013_ (.A1(_15347_),
    .A2(_04499_),
    .B(_04595_),
    .C(_15752_),
    .Y(_04596_));
 AO21x1_ASAP7_75t_R _19014_ (.A1(_15593_),
    .A2(_04594_),
    .B(_04596_),
    .Y(_04597_));
 NAND2x1_ASAP7_75t_R _19015_ (.A(net1971),
    .B(_01278_),
    .Y(_04598_));
 OA211x2_ASAP7_75t_R _19016_ (.A1(_15302_),
    .A2(_04503_),
    .B(_04598_),
    .C(_16948_),
    .Y(_04599_));
 NAND2x1_ASAP7_75t_R _19017_ (.A(net1971),
    .B(_01277_),
    .Y(_04600_));
 OA211x2_ASAP7_75t_R _19018_ (.A1(_15302_),
    .A2(_04506_),
    .B(_04600_),
    .C(_15274_),
    .Y(_04601_));
 OR3x1_ASAP7_75t_R _19019_ (.A(_15287_),
    .B(_04599_),
    .C(_04601_),
    .Y(_04602_));
 OA211x2_ASAP7_75t_R _19020_ (.A1(_15596_),
    .A2(_04597_),
    .B(_04602_),
    .C(_15312_),
    .Y(_04603_));
 OR3x2_ASAP7_75t_R _19021_ (.A(_15316_),
    .B(_04592_),
    .C(_04603_),
    .Y(_04604_));
 AND2x6_ASAP7_75t_R _19022_ (.A(_04581_),
    .B(_04604_),
    .Y(_04605_));
 INVx2_ASAP7_75t_R _19023_ (.A(_04605_),
    .Y(_04606_));
 OA211x2_ASAP7_75t_R _19024_ (.A1(_01513_),
    .A2(_15364_),
    .B(_16388_),
    .C(_15370_),
    .Y(_04607_));
 AOI21x1_ASAP7_75t_R _19025_ (.A1(_15250_),
    .A2(_04606_),
    .B(_04607_),
    .Y(_18694_));
 INVx1_ASAP7_75t_R _19026_ (.A(_18694_),
    .Y(_18692_));
 AND2x2_ASAP7_75t_R _19027_ (.A(_14717_),
    .B(_01767_),
    .Y(_04608_));
 AO21x1_ASAP7_75t_R _19028_ (.A1(_14286_),
    .A2(_01296_),
    .B(_04608_),
    .Y(_04609_));
 OAI22x1_ASAP7_75t_R _19029_ (.A1(_01295_),
    .A2(_14284_),
    .B1(_04609_),
    .B2(_13090_),
    .Y(_04610_));
 INVx1_ASAP7_75t_R _19030_ (.A(_01304_),
    .Y(_04611_));
 NAND2x1_ASAP7_75t_R _19031_ (.A(_14507_),
    .B(_01302_),
    .Y(_04612_));
 OA211x2_ASAP7_75t_R _19032_ (.A1(_14516_),
    .A2(_04611_),
    .B(_04612_),
    .C(_14472_),
    .Y(_04613_));
 INVx1_ASAP7_75t_R _19033_ (.A(_01303_),
    .Y(_04614_));
 NAND2x1_ASAP7_75t_R _19034_ (.A(_14517_),
    .B(_01301_),
    .Y(_04615_));
 OA211x2_ASAP7_75t_R _19035_ (.A1(_13193_),
    .A2(_04614_),
    .B(_04615_),
    .C(_14476_),
    .Y(_04616_));
 OR3x1_ASAP7_75t_R _19036_ (.A(_14353_),
    .B(_04613_),
    .C(_04616_),
    .Y(_04617_));
 OA211x2_ASAP7_75t_R _19037_ (.A1(_13086_),
    .A2(_04610_),
    .B(_04617_),
    .C(_14852_),
    .Y(_04618_));
 INVx1_ASAP7_75t_R _19038_ (.A(_01300_),
    .Y(_04619_));
 NAND2x1_ASAP7_75t_R _19039_ (.A(_13200_),
    .B(_01298_),
    .Y(_04620_));
 OA211x2_ASAP7_75t_R _19040_ (.A1(_13197_),
    .A2(_04619_),
    .B(_04620_),
    .C(_14856_),
    .Y(_04621_));
 INVx1_ASAP7_75t_R _19041_ (.A(_01299_),
    .Y(_04622_));
 NAND2x1_ASAP7_75t_R _19042_ (.A(_14858_),
    .B(_01297_),
    .Y(_04623_));
 OA211x2_ASAP7_75t_R _19043_ (.A1(_14854_),
    .A2(_04622_),
    .B(_04623_),
    .C(_14874_),
    .Y(_04624_));
 OR3x1_ASAP7_75t_R _19044_ (.A(_15117_),
    .B(_04621_),
    .C(_04624_),
    .Y(_04625_));
 INVx1_ASAP7_75t_R _19045_ (.A(_01308_),
    .Y(_04626_));
 NAND2x1_ASAP7_75t_R _19046_ (.A(_14653_),
    .B(_01306_),
    .Y(_04627_));
 OA211x2_ASAP7_75t_R _19047_ (.A1(_13197_),
    .A2(_04626_),
    .B(_04627_),
    .C(_14856_),
    .Y(_04628_));
 INVx1_ASAP7_75t_R _19048_ (.A(_01307_),
    .Y(_04629_));
 NAND2x1_ASAP7_75t_R _19049_ (.A(_14858_),
    .B(_01305_),
    .Y(_04630_));
 OA211x2_ASAP7_75t_R _19050_ (.A1(_14854_),
    .A2(_04629_),
    .B(_04630_),
    .C(_14874_),
    .Y(_04631_));
 OR3x1_ASAP7_75t_R _19051_ (.A(_14877_),
    .B(_04628_),
    .C(_04631_),
    .Y(_04632_));
 AND3x1_ASAP7_75t_R _19052_ (.A(_14340_),
    .B(_04625_),
    .C(_04632_),
    .Y(_04633_));
 OR3x1_ASAP7_75t_R _19053_ (.A(_13082_),
    .B(_04618_),
    .C(_04633_),
    .Y(_04634_));
 INVx2_ASAP7_75t_R _19054_ (.A(_01316_),
    .Y(_04635_));
 NAND2x1_ASAP7_75t_R _19055_ (.A(_13200_),
    .B(_01314_),
    .Y(_04636_));
 OA211x2_ASAP7_75t_R _19056_ (.A1(_13197_),
    .A2(_04635_),
    .B(_04636_),
    .C(_14856_),
    .Y(_04637_));
 INVx2_ASAP7_75t_R _19057_ (.A(_01315_),
    .Y(_04638_));
 NAND2x1_ASAP7_75t_R _19058_ (.A(_14858_),
    .B(_01313_),
    .Y(_04639_));
 OA211x2_ASAP7_75t_R _19059_ (.A1(_14854_),
    .A2(_04638_),
    .B(_04639_),
    .C(_14874_),
    .Y(_04640_));
 OR3x1_ASAP7_75t_R _19060_ (.A(_15117_),
    .B(_04637_),
    .C(_04640_),
    .Y(_04641_));
 INVx2_ASAP7_75t_R _19061_ (.A(_01324_),
    .Y(_04642_));
 NAND2x1_ASAP7_75t_R _19062_ (.A(_14653_),
    .B(_01322_),
    .Y(_04643_));
 OA211x2_ASAP7_75t_R _19063_ (.A1(_14854_),
    .A2(_04642_),
    .B(_04643_),
    .C(_14856_),
    .Y(_04644_));
 INVx2_ASAP7_75t_R _19064_ (.A(_01323_),
    .Y(_04645_));
 NAND2x1_ASAP7_75t_R _19065_ (.A(_14858_),
    .B(_01321_),
    .Y(_04646_));
 OA211x2_ASAP7_75t_R _19066_ (.A1(_14854_),
    .A2(_04645_),
    .B(_04646_),
    .C(_14874_),
    .Y(_04647_));
 OR3x1_ASAP7_75t_R _19067_ (.A(_14877_),
    .B(_04644_),
    .C(_04647_),
    .Y(_04648_));
 AND3x1_ASAP7_75t_R _19068_ (.A(_13129_),
    .B(_04641_),
    .C(_04648_),
    .Y(_04649_));
 INVx2_ASAP7_75t_R _19069_ (.A(_01317_),
    .Y(_04650_));
 NOR2x1_ASAP7_75t_R _19070_ (.A(_14943_),
    .B(_01319_),
    .Y(_04651_));
 AO21x1_ASAP7_75t_R _19071_ (.A1(_13190_),
    .A2(_04650_),
    .B(_04651_),
    .Y(_04652_));
 INVx2_ASAP7_75t_R _19072_ (.A(_01320_),
    .Y(_04653_));
 NAND2x1_ASAP7_75t_R _19073_ (.A(_14888_),
    .B(_01318_),
    .Y(_04654_));
 OA211x2_ASAP7_75t_R _19074_ (.A1(_14886_),
    .A2(_04653_),
    .B(_04654_),
    .C(_14652_),
    .Y(_04655_));
 AO21x1_ASAP7_75t_R _19075_ (.A1(_14975_),
    .A2(_04652_),
    .B(_04655_),
    .Y(_04656_));
 INVx2_ASAP7_75t_R _19076_ (.A(_01312_),
    .Y(_04657_));
 NAND2x1_ASAP7_75t_R _19077_ (.A(_14310_),
    .B(_01310_),
    .Y(_04658_));
 OA211x2_ASAP7_75t_R _19078_ (.A1(_14474_),
    .A2(_04657_),
    .B(_04658_),
    .C(_13115_),
    .Y(_04659_));
 INVx2_ASAP7_75t_R _19079_ (.A(_01311_),
    .Y(_04660_));
 NAND2x1_ASAP7_75t_R _19080_ (.A(_14317_),
    .B(_01309_),
    .Y(_04661_));
 OA211x2_ASAP7_75t_R _19081_ (.A1(_13107_),
    .A2(_04660_),
    .B(_04661_),
    .C(_14476_),
    .Y(_04662_));
 OR3x1_ASAP7_75t_R _19082_ (.A(_14469_),
    .B(_04659_),
    .C(_04662_),
    .Y(_04663_));
 OA211x2_ASAP7_75t_R _19083_ (.A1(_14354_),
    .A2(_04656_),
    .B(_04663_),
    .C(_14852_),
    .Y(_04664_));
 OR3x2_ASAP7_75t_R _19084_ (.A(_13164_),
    .B(_04649_),
    .C(_04664_),
    .Y(_04665_));
 AO21x2_ASAP7_75t_R _19085_ (.A1(_04634_),
    .A2(_04665_),
    .B(_14377_),
    .Y(_04666_));
 BUFx6f_ASAP7_75t_R _19086_ (.A(_01486_),
    .Y(_04667_));
 AND2x2_ASAP7_75t_R _19087_ (.A(_01456_),
    .B(_14381_),
    .Y(_04668_));
 OAI22x1_ASAP7_75t_R _19088_ (.A1(_04667_),
    .A2(_14967_),
    .B1(_14968_),
    .B2(_04668_),
    .Y(_04669_));
 NAND2x2_ASAP7_75t_R _19089_ (.A(_04666_),
    .B(_04669_),
    .Y(_18698_));
 INVx1_ASAP7_75t_R _19090_ (.A(_18698_),
    .Y(_18700_));
 BUFx6f_ASAP7_75t_R _19091_ (.A(_00176_),
    .Y(_04670_));
 INVx1_ASAP7_75t_R _19092_ (.A(_04670_),
    .Y(_04671_));
 AND3x1_ASAP7_75t_R _19093_ (.A(_04671_),
    .B(_14625_),
    .C(_14906_),
    .Y(_04672_));
 AO21x1_ASAP7_75t_R _19094_ (.A1(_14903_),
    .A2(_18700_),
    .B(_04672_),
    .Y(_18066_));
 AND2x2_ASAP7_75t_R _19095_ (.A(_15325_),
    .B(_01767_),
    .Y(_04673_));
 AO21x1_ASAP7_75t_R _19096_ (.A1(_15436_),
    .A2(_01296_),
    .B(_04673_),
    .Y(_04674_));
 OAI22x1_ASAP7_75t_R _19097_ (.A1(_01295_),
    .A2(_15435_),
    .B1(_04674_),
    .B2(_15594_),
    .Y(_04675_));
 NAND2x1_ASAP7_75t_R _19098_ (.A(_15347_),
    .B(_01302_),
    .Y(_04676_));
 OA211x2_ASAP7_75t_R _19099_ (.A1(_15490_),
    .A2(_04611_),
    .B(_04676_),
    .C(_15469_),
    .Y(_04677_));
 NAND2x1_ASAP7_75t_R _19100_ (.A(_15321_),
    .B(_01301_),
    .Y(_04678_));
 OA211x2_ASAP7_75t_R _19101_ (.A1(_15490_),
    .A2(_04614_),
    .B(_04678_),
    .C(_15338_),
    .Y(_04679_));
 OR3x1_ASAP7_75t_R _19102_ (.A(_15475_),
    .B(_04677_),
    .C(_04679_),
    .Y(_04680_));
 OA211x2_ASAP7_75t_R _19103_ (.A1(_15588_),
    .A2(_04675_),
    .B(_04680_),
    .C(_15360_),
    .Y(_04681_));
 NAND2x1_ASAP7_75t_R _19104_ (.A(_15353_),
    .B(_01298_),
    .Y(_04682_));
 OA211x2_ASAP7_75t_R _19105_ (.A1(_15341_),
    .A2(_04619_),
    .B(_04682_),
    .C(_15600_),
    .Y(_04683_));
 NAND2x1_ASAP7_75t_R _19106_ (.A(_15300_),
    .B(_01297_),
    .Y(_04684_));
 OA211x2_ASAP7_75t_R _19107_ (.A1(_15341_),
    .A2(_04622_),
    .B(_04684_),
    .C(_15295_),
    .Y(_04685_));
 OR3x1_ASAP7_75t_R _19108_ (.A(_16368_),
    .B(_04683_),
    .C(_04685_),
    .Y(_04686_));
 NAND2x1_ASAP7_75t_R _19109_ (.A(_15300_),
    .B(_01306_),
    .Y(_04687_));
 OA211x2_ASAP7_75t_R _19110_ (.A1(_15341_),
    .A2(_04626_),
    .B(_04687_),
    .C(_15600_),
    .Y(_04688_));
 NAND2x1_ASAP7_75t_R _19111_ (.A(_15307_),
    .B(_01305_),
    .Y(_04689_));
 OA211x2_ASAP7_75t_R _19112_ (.A1(_15633_),
    .A2(_04629_),
    .B(_04689_),
    .C(_15295_),
    .Y(_04690_));
 OR3x1_ASAP7_75t_R _19113_ (.A(_15596_),
    .B(_04688_),
    .C(_04690_),
    .Y(_04691_));
 AND3x1_ASAP7_75t_R _19114_ (.A(_16218_),
    .B(_04686_),
    .C(_04691_),
    .Y(_04692_));
 OR3x2_ASAP7_75t_R _19115_ (.A(_15434_),
    .B(_04681_),
    .C(_04692_),
    .Y(_04693_));
 NAND2x1_ASAP7_75t_R _19116_ (.A(_15353_),
    .B(_01314_),
    .Y(_04694_));
 OA211x2_ASAP7_75t_R _19117_ (.A1(_15484_),
    .A2(_04635_),
    .B(_04694_),
    .C(_15600_),
    .Y(_04695_));
 NAND2x1_ASAP7_75t_R _19118_ (.A(_15353_),
    .B(_01313_),
    .Y(_04696_));
 OA211x2_ASAP7_75t_R _19119_ (.A1(_15341_),
    .A2(_04638_),
    .B(_04696_),
    .C(_15295_),
    .Y(_04697_));
 OR3x1_ASAP7_75t_R _19120_ (.A(_16368_),
    .B(_04695_),
    .C(_04697_),
    .Y(_04698_));
 NAND2x1_ASAP7_75t_R _19121_ (.A(_15353_),
    .B(_01322_),
    .Y(_04699_));
 OA211x2_ASAP7_75t_R _19122_ (.A1(_15341_),
    .A2(_04642_),
    .B(_04699_),
    .C(_15600_),
    .Y(_04700_));
 NAND2x1_ASAP7_75t_R _19123_ (.A(_15300_),
    .B(_01321_),
    .Y(_04701_));
 OA211x2_ASAP7_75t_R _19124_ (.A1(_15341_),
    .A2(_04645_),
    .B(_04701_),
    .C(_15295_),
    .Y(_04702_));
 OR3x1_ASAP7_75t_R _19125_ (.A(_15596_),
    .B(_04700_),
    .C(_04702_),
    .Y(_04703_));
 AND3x1_ASAP7_75t_R _19126_ (.A(_16218_),
    .B(_04698_),
    .C(_04703_),
    .Y(_04704_));
 NOR2x1_ASAP7_75t_R _19127_ (.A(_15598_),
    .B(_01319_),
    .Y(_04705_));
 AO21x1_ASAP7_75t_R _19128_ (.A1(_16333_),
    .A2(_04650_),
    .B(_04705_),
    .Y(_04706_));
 NAND2x1_ASAP7_75t_R _19129_ (.A(_15445_),
    .B(_01318_),
    .Y(_04707_));
 OA211x2_ASAP7_75t_R _19130_ (.A1(_15484_),
    .A2(_04653_),
    .B(_04707_),
    .C(_15600_),
    .Y(_04708_));
 AO21x1_ASAP7_75t_R _19131_ (.A1(_15296_),
    .A2(_04706_),
    .B(_04708_),
    .Y(_04709_));
 NAND2x1_ASAP7_75t_R _19132_ (.A(_15321_),
    .B(_01310_),
    .Y(_04710_));
 OA211x2_ASAP7_75t_R _19133_ (.A1(_15490_),
    .A2(_04657_),
    .B(_04710_),
    .C(_15469_),
    .Y(_04711_));
 NAND2x1_ASAP7_75t_R _19134_ (.A(_15321_),
    .B(_01309_),
    .Y(_04712_));
 OA211x2_ASAP7_75t_R _19135_ (.A1(_15490_),
    .A2(_04660_),
    .B(_04712_),
    .C(_15338_),
    .Y(_04713_));
 OR3x1_ASAP7_75t_R _19136_ (.A(_16368_),
    .B(_04711_),
    .C(_04713_),
    .Y(_04714_));
 OA211x2_ASAP7_75t_R _19137_ (.A1(_15482_),
    .A2(_04709_),
    .B(_04714_),
    .C(_15360_),
    .Y(_04715_));
 OR3x2_ASAP7_75t_R _19138_ (.A(_15466_),
    .B(_04704_),
    .C(_04715_),
    .Y(_04716_));
 AND2x6_ASAP7_75t_R _19139_ (.A(_04693_),
    .B(_04716_),
    .Y(_04717_));
 INVx2_ASAP7_75t_R _19140_ (.A(_04717_),
    .Y(_04718_));
 OA211x2_ASAP7_75t_R _19141_ (.A1(_01512_),
    .A2(_16386_),
    .B(_16389_),
    .C(_15503_),
    .Y(_04719_));
 AOI21x1_ASAP7_75t_R _19142_ (.A1(_14090_),
    .A2(_04718_),
    .B(_04719_),
    .Y(_18699_));
 INVx1_ASAP7_75t_R _19143_ (.A(_18699_),
    .Y(_18697_));
 OA31x2_ASAP7_75t_R _19144_ (.A1(_01261_),
    .A2(_04476_),
    .A3(_04478_),
    .B1(_01294_),
    .Y(_04720_));
 OA21x2_ASAP7_75t_R _19145_ (.A1(_01293_),
    .A2(_04720_),
    .B(_01326_),
    .Y(_04721_));
 XNOR2x1_ASAP7_75t_R _19146_ (.B(_04721_),
    .Y(_04722_),
    .A(_01325_));
 INVx6_ASAP7_75t_R _19147_ (.A(_04722_),
    .Y(\alu_adder_result_ex[29] ));
 OR3x2_ASAP7_75t_R _19148_ (.A(_01229_),
    .B(_01261_),
    .C(_04487_),
    .Y(_04723_));
 OA21x2_ASAP7_75t_R _19149_ (.A1(_01165_),
    .A2(_04244_),
    .B(_01198_),
    .Y(_04724_));
 OA21x2_ASAP7_75t_R _19150_ (.A1(_01197_),
    .A2(_04724_),
    .B(_01230_),
    .Y(_04725_));
 OA21x2_ASAP7_75t_R _19151_ (.A1(_01229_),
    .A2(_04725_),
    .B(_01262_),
    .Y(_04726_));
 OA21x2_ASAP7_75t_R _19152_ (.A1(_01261_),
    .A2(_04726_),
    .B(_01294_),
    .Y(_04727_));
 OA31x2_ASAP7_75t_R _19153_ (.A1(_16756_),
    .A2(_16758_),
    .A3(_04723_),
    .B1(_04727_),
    .Y(_04728_));
 XNOR2x1_ASAP7_75t_R _19154_ (.B(_04728_),
    .Y(_04729_),
    .A(_01293_));
 INVx4_ASAP7_75t_R _19155_ (.A(_04729_),
    .Y(\alu_adder_result_ex[28] ));
 AND2x2_ASAP7_75t_R _19156_ (.A(_14717_),
    .B(_01766_),
    .Y(_04730_));
 AO21x1_ASAP7_75t_R _19157_ (.A1(_13092_),
    .A2(_01328_),
    .B(_04730_),
    .Y(_04731_));
 OAI22x1_ASAP7_75t_R _19158_ (.A1(_01327_),
    .A2(_13102_),
    .B1(_04731_),
    .B2(_13090_),
    .Y(_04732_));
 INVx1_ASAP7_75t_R _19159_ (.A(_01336_),
    .Y(_04733_));
 NAND2x1_ASAP7_75t_R _19160_ (.A(_14317_),
    .B(_01334_),
    .Y(_04734_));
 OA211x2_ASAP7_75t_R _19161_ (.A1(_14474_),
    .A2(_04733_),
    .B(_04734_),
    .C(_13115_),
    .Y(_04735_));
 INVx1_ASAP7_75t_R _19162_ (.A(_01335_),
    .Y(_04736_));
 NAND2x1_ASAP7_75t_R _19163_ (.A(_13110_),
    .B(_01333_),
    .Y(_04737_));
 OA211x2_ASAP7_75t_R _19164_ (.A1(_13107_),
    .A2(_04736_),
    .B(_04737_),
    .C(_14476_),
    .Y(_04738_));
 OR3x1_ASAP7_75t_R _19165_ (.A(_13105_),
    .B(_04735_),
    .C(_04738_),
    .Y(_04739_));
 OA211x2_ASAP7_75t_R _19166_ (.A1(_13086_),
    .A2(_04732_),
    .B(_04739_),
    .C(_13125_),
    .Y(_04740_));
 INVx1_ASAP7_75t_R _19167_ (.A(_01332_),
    .Y(_04741_));
 NAND2x1_ASAP7_75t_R _19168_ (.A(_13168_),
    .B(_01330_),
    .Y(_04742_));
 OA211x2_ASAP7_75t_R _19169_ (.A1(_13166_),
    .A2(_04741_),
    .B(_04742_),
    .C(_14856_),
    .Y(_04743_));
 INVx2_ASAP7_75t_R _19170_ (.A(_01331_),
    .Y(_04744_));
 NAND2x1_ASAP7_75t_R _19171_ (.A(_13137_),
    .B(_01329_),
    .Y(_04745_));
 OA211x2_ASAP7_75t_R _19172_ (.A1(_13133_),
    .A2(_04744_),
    .B(_04745_),
    .C(_13174_),
    .Y(_04746_));
 OR3x1_ASAP7_75t_R _19173_ (.A(_13131_),
    .B(_04743_),
    .C(_04746_),
    .Y(_04747_));
 INVx1_ASAP7_75t_R _19174_ (.A(_01340_),
    .Y(_04748_));
 NAND2x1_ASAP7_75t_R _19175_ (.A(_13168_),
    .B(_01338_),
    .Y(_04749_));
 OA211x2_ASAP7_75t_R _19176_ (.A1(_13166_),
    .A2(_04748_),
    .B(_04749_),
    .C(_13140_),
    .Y(_04750_));
 INVx1_ASAP7_75t_R _19177_ (.A(_01339_),
    .Y(_04751_));
 NAND2x1_ASAP7_75t_R _19178_ (.A(_13137_),
    .B(_01337_),
    .Y(_04752_));
 OA211x2_ASAP7_75t_R _19179_ (.A1(_13133_),
    .A2(_04751_),
    .B(_04752_),
    .C(_13174_),
    .Y(_04753_));
 OR3x1_ASAP7_75t_R _19180_ (.A(_13153_),
    .B(_04750_),
    .C(_04753_),
    .Y(_04754_));
 AND3x1_ASAP7_75t_R _19181_ (.A(_13129_),
    .B(_04747_),
    .C(_04754_),
    .Y(_04755_));
 OR3x2_ASAP7_75t_R _19182_ (.A(_13082_),
    .B(_04740_),
    .C(_04755_),
    .Y(_04756_));
 INVx1_ASAP7_75t_R _19183_ (.A(_01348_),
    .Y(_04757_));
 NAND2x1_ASAP7_75t_R _19184_ (.A(_13168_),
    .B(_01346_),
    .Y(_04758_));
 OA211x2_ASAP7_75t_R _19185_ (.A1(_13166_),
    .A2(_04757_),
    .B(_04758_),
    .C(_14856_),
    .Y(_04759_));
 INVx1_ASAP7_75t_R _19186_ (.A(_01347_),
    .Y(_04760_));
 NAND2x1_ASAP7_75t_R _19187_ (.A(_13137_),
    .B(_01345_),
    .Y(_04761_));
 OA211x2_ASAP7_75t_R _19188_ (.A1(_13133_),
    .A2(_04760_),
    .B(_04761_),
    .C(_13174_),
    .Y(_04762_));
 OR3x1_ASAP7_75t_R _19189_ (.A(_13131_),
    .B(_04759_),
    .C(_04762_),
    .Y(_04763_));
 INVx1_ASAP7_75t_R _19190_ (.A(_01356_),
    .Y(_04764_));
 NAND2x1_ASAP7_75t_R _19191_ (.A(_13168_),
    .B(_01354_),
    .Y(_04765_));
 OA211x2_ASAP7_75t_R _19192_ (.A1(_13166_),
    .A2(_04764_),
    .B(_04765_),
    .C(_13140_),
    .Y(_04766_));
 INVx1_ASAP7_75t_R _19193_ (.A(_01355_),
    .Y(_04767_));
 NAND2x1_ASAP7_75t_R _19194_ (.A(_13137_),
    .B(_01353_),
    .Y(_04768_));
 OA211x2_ASAP7_75t_R _19195_ (.A1(_13143_),
    .A2(_04767_),
    .B(_04768_),
    .C(_13174_),
    .Y(_04769_));
 OR3x1_ASAP7_75t_R _19196_ (.A(_13153_),
    .B(_04766_),
    .C(_04769_),
    .Y(_04770_));
 AND3x1_ASAP7_75t_R _19197_ (.A(_13129_),
    .B(_04763_),
    .C(_04770_),
    .Y(_04771_));
 INVx2_ASAP7_75t_R _19198_ (.A(_01349_),
    .Y(_04772_));
 NOR2x1_ASAP7_75t_R _19199_ (.A(_14516_),
    .B(_01351_),
    .Y(_04773_));
 AO21x1_ASAP7_75t_R _19200_ (.A1(_13190_),
    .A2(_04772_),
    .B(_04773_),
    .Y(_04774_));
 INVx2_ASAP7_75t_R _19201_ (.A(_01352_),
    .Y(_04775_));
 NAND2x1_ASAP7_75t_R _19202_ (.A(_14738_),
    .B(_01350_),
    .Y(_04776_));
 OA211x2_ASAP7_75t_R _19203_ (.A1(_13197_),
    .A2(_04775_),
    .B(_04776_),
    .C(_13202_),
    .Y(_04777_));
 AO21x1_ASAP7_75t_R _19204_ (.A1(_13187_),
    .A2(_04774_),
    .B(_04777_),
    .Y(_04778_));
 INVx1_ASAP7_75t_R _19205_ (.A(_01344_),
    .Y(_04779_));
 NAND2x1_ASAP7_75t_R _19206_ (.A(_15675_),
    .B(_01342_),
    .Y(_04780_));
 OA211x2_ASAP7_75t_R _19207_ (.A1(_13107_),
    .A2(_04779_),
    .B(_04780_),
    .C(_13115_),
    .Y(_04781_));
 INVx1_ASAP7_75t_R _19208_ (.A(_01343_),
    .Y(_04782_));
 NAND2x1_ASAP7_75t_R _19209_ (.A(_13118_),
    .B(_01341_),
    .Y(_04783_));
 OA211x2_ASAP7_75t_R _19210_ (.A1(_13206_),
    .A2(_04782_),
    .B(_04783_),
    .C(_13120_),
    .Y(_04784_));
 OR3x1_ASAP7_75t_R _19211_ (.A(_13085_),
    .B(_04781_),
    .C(_04784_),
    .Y(_04785_));
 OA211x2_ASAP7_75t_R _19212_ (.A1(_13186_),
    .A2(_04778_),
    .B(_04785_),
    .C(_13125_),
    .Y(_04786_));
 OR3x2_ASAP7_75t_R _19213_ (.A(_13164_),
    .B(_04771_),
    .C(_04786_),
    .Y(_04787_));
 AO21x2_ASAP7_75t_R _19214_ (.A1(_04756_),
    .A2(_04787_),
    .B(_13267_),
    .Y(_04788_));
 AND2x2_ASAP7_75t_R _19215_ (.A(_01454_),
    .B(_14381_),
    .Y(_04789_));
 OAI22x1_ASAP7_75t_R _19216_ (.A1(_01485_),
    .A2(_14967_),
    .B1(_14968_),
    .B2(_04789_),
    .Y(_04790_));
 NAND2x2_ASAP7_75t_R _19217_ (.A(_04788_),
    .B(_04790_),
    .Y(_18703_));
 INVx1_ASAP7_75t_R _19218_ (.A(_18703_),
    .Y(_18705_));
 BUFx6f_ASAP7_75t_R _19219_ (.A(_00181_),
    .Y(_04791_));
 OR3x1_ASAP7_75t_R _19220_ (.A(_04791_),
    .B(_14627_),
    .C(_14649_),
    .Y(_04792_));
 OAI21x1_ASAP7_75t_R _19221_ (.A1(_14646_),
    .A2(_18703_),
    .B(_04792_),
    .Y(_18068_));
 AND2x2_ASAP7_75t_R _19222_ (.A(_15347_),
    .B(_01766_),
    .Y(_04793_));
 AO21x1_ASAP7_75t_R _19223_ (.A1(_15290_),
    .A2(_01328_),
    .B(_04793_),
    .Y(_04794_));
 OAI22x1_ASAP7_75t_R _19224_ (.A1(_01327_),
    .A2(_15289_),
    .B1(_04794_),
    .B2(_15339_),
    .Y(_04795_));
 NAND2x1_ASAP7_75t_R _19225_ (.A(_15597_),
    .B(_01334_),
    .Y(_04796_));
 OA211x2_ASAP7_75t_R _19226_ (.A1(_15437_),
    .A2(_04733_),
    .B(_04796_),
    .C(_15304_),
    .Y(_04797_));
 NAND2x1_ASAP7_75t_R _19227_ (.A(_15319_),
    .B(_01333_),
    .Y(_04798_));
 OA211x2_ASAP7_75t_R _19228_ (.A1(_15437_),
    .A2(_04736_),
    .B(_04798_),
    .C(_15592_),
    .Y(_04799_));
 OR3x1_ASAP7_75t_R _19229_ (.A(_15336_),
    .B(_04797_),
    .C(_04799_),
    .Y(_04800_));
 OA211x2_ASAP7_75t_R _19230_ (.A1(_15288_),
    .A2(_04795_),
    .B(_04800_),
    .C(_15313_),
    .Y(_04801_));
 NAND2x1_ASAP7_75t_R _19231_ (.A(_15734_),
    .B(_01330_),
    .Y(_04802_));
 OA211x2_ASAP7_75t_R _19232_ (.A1(_15486_),
    .A2(_04741_),
    .B(_04802_),
    .C(_15443_),
    .Y(_04803_));
 NAND2x1_ASAP7_75t_R _19233_ (.A(_15483_),
    .B(_01329_),
    .Y(_04804_));
 OA211x2_ASAP7_75t_R _19234_ (.A1(_15589_),
    .A2(_04744_),
    .B(_04804_),
    .C(_15497_),
    .Y(_04805_));
 OR3x1_ASAP7_75t_R _19235_ (.A(_15255_),
    .B(_04803_),
    .C(_04805_),
    .Y(_04806_));
 NAND2x1_ASAP7_75t_R _19236_ (.A(_15483_),
    .B(_01338_),
    .Y(_04807_));
 OA211x2_ASAP7_75t_R _19237_ (.A1(_15486_),
    .A2(_04748_),
    .B(_04807_),
    .C(_15443_),
    .Y(_04808_));
 NAND2x1_ASAP7_75t_R _19238_ (.A(_15483_),
    .B(_01337_),
    .Y(_04809_));
 OA211x2_ASAP7_75t_R _19239_ (.A1(_15589_),
    .A2(_04751_),
    .B(_04809_),
    .C(_15497_),
    .Y(_04810_));
 OR3x1_ASAP7_75t_R _19240_ (.A(_15298_),
    .B(_04808_),
    .C(_04810_),
    .Y(_04811_));
 AND3x1_ASAP7_75t_R _19241_ (.A(_15253_),
    .B(_04806_),
    .C(_04811_),
    .Y(_04812_));
 OR3x2_ASAP7_75t_R _19242_ (.A(_15251_),
    .B(_04801_),
    .C(_04812_),
    .Y(_04813_));
 NAND2x1_ASAP7_75t_R _19243_ (.A(_15618_),
    .B(_01346_),
    .Y(_04814_));
 OA211x2_ASAP7_75t_R _19244_ (.A1(_15622_),
    .A2(_04757_),
    .B(_04814_),
    .C(_15620_),
    .Y(_04815_));
 NAND2x1_ASAP7_75t_R _19245_ (.A(_15340_),
    .B(_01345_),
    .Y(_04816_));
 OA211x2_ASAP7_75t_R _19246_ (.A1(_15622_),
    .A2(_04760_),
    .B(_04816_),
    .C(_15283_),
    .Y(_04817_));
 OR3x1_ASAP7_75t_R _19247_ (.A(_15255_),
    .B(_04815_),
    .C(_04817_),
    .Y(_04818_));
 NAND2x1_ASAP7_75t_R _19248_ (.A(_15340_),
    .B(_01354_),
    .Y(_04819_));
 OA211x2_ASAP7_75t_R _19249_ (.A1(_15622_),
    .A2(_04764_),
    .B(_04819_),
    .C(_15620_),
    .Y(_04820_));
 NAND2x1_ASAP7_75t_R _19250_ (.A(_15340_),
    .B(_01353_),
    .Y(_04821_));
 OA211x2_ASAP7_75t_R _19251_ (.A1(_15343_),
    .A2(_04767_),
    .B(_04821_),
    .C(_15283_),
    .Y(_04822_));
 OR3x1_ASAP7_75t_R _19252_ (.A(_15279_),
    .B(_04820_),
    .C(_04822_),
    .Y(_04823_));
 AND3x1_ASAP7_75t_R _19253_ (.A(_15253_),
    .B(_04818_),
    .C(_04823_),
    .Y(_04824_));
 NOR2x1_ASAP7_75t_R _19254_ (.A(_15353_),
    .B(_01351_),
    .Y(_04825_));
 AO21x1_ASAP7_75t_R _19255_ (.A1(_15633_),
    .A2(_04772_),
    .B(_04825_),
    .Y(_04826_));
 NAND2x1_ASAP7_75t_R _19256_ (.A(_16106_),
    .B(_01350_),
    .Y(_04827_));
 OA211x2_ASAP7_75t_R _19257_ (.A1(_15325_),
    .A2(_04775_),
    .B(_04827_),
    .C(_15267_),
    .Y(_04828_));
 AO21x1_ASAP7_75t_R _19258_ (.A1(_15339_),
    .A2(_04826_),
    .B(_04828_),
    .Y(_04829_));
 NAND2x1_ASAP7_75t_R _19259_ (.A(_15597_),
    .B(_01342_),
    .Y(_04830_));
 OA211x2_ASAP7_75t_R _19260_ (.A1(_15307_),
    .A2(_04779_),
    .B(_04830_),
    .C(_15304_),
    .Y(_04831_));
 NAND2x1_ASAP7_75t_R _19261_ (.A(_15597_),
    .B(_01341_),
    .Y(_04832_));
 OA211x2_ASAP7_75t_R _19262_ (.A1(_15437_),
    .A2(_04782_),
    .B(_04832_),
    .C(_15592_),
    .Y(_04833_));
 OR3x1_ASAP7_75t_R _19263_ (.A(_15352_),
    .B(_04831_),
    .C(_04833_),
    .Y(_04834_));
 OA211x2_ASAP7_75t_R _19264_ (.A1(_15337_),
    .A2(_04829_),
    .B(_04834_),
    .C(_15313_),
    .Y(_04835_));
 OR3x2_ASAP7_75t_R _19265_ (.A(_15316_),
    .B(_04824_),
    .C(_04835_),
    .Y(_04836_));
 NAND2x2_ASAP7_75t_R _19266_ (.A(_04813_),
    .B(_04836_),
    .Y(_04837_));
 OA211x2_ASAP7_75t_R _19267_ (.A1(_14122_),
    .A2(_16386_),
    .B(_16389_),
    .C(_15370_),
    .Y(_04838_));
 AOI21x1_ASAP7_75t_R _19268_ (.A1(_15250_),
    .A2(_04837_),
    .B(_04838_),
    .Y(_18704_));
 INVx1_ASAP7_75t_R _19269_ (.A(_18704_),
    .Y(_18702_));
 BUFx6f_ASAP7_75t_R _19270_ (.A(_00343_),
    .Y(_04839_));
 INVx2_ASAP7_75t_R _19271_ (.A(_01387_),
    .Y(_04840_));
 NAND2x1_ASAP7_75t_R _19272_ (.A(_13093_),
    .B(_01385_),
    .Y(_04841_));
 OA211x2_ASAP7_75t_R _19273_ (.A1(_04839_),
    .A2(_04840_),
    .B(_04841_),
    .C(_13087_),
    .Y(_04842_));
 INVx2_ASAP7_75t_R _19274_ (.A(_01388_),
    .Y(_04843_));
 NAND2x1_ASAP7_75t_R _19275_ (.A(_13093_),
    .B(_01386_),
    .Y(_04844_));
 OA211x2_ASAP7_75t_R _19276_ (.A1(_04839_),
    .A2(_04843_),
    .B(_04844_),
    .C(_13113_),
    .Y(_04845_));
 OA21x2_ASAP7_75t_R _19277_ (.A1(_04842_),
    .A2(_04845_),
    .B(_13084_),
    .Y(_04846_));
 AND2x2_ASAP7_75t_R _19278_ (.A(_13113_),
    .B(_00341_),
    .Y(_04847_));
 INVx2_ASAP7_75t_R _19279_ (.A(_01380_),
    .Y(_04848_));
 NAND2x1_ASAP7_75t_R _19280_ (.A(_13093_),
    .B(_01378_),
    .Y(_04849_));
 OA21x2_ASAP7_75t_R _19281_ (.A1(_04839_),
    .A2(_04848_),
    .B(_04849_),
    .Y(_04850_));
 INVx2_ASAP7_75t_R _19282_ (.A(_01377_),
    .Y(_04851_));
 NOR2x1_ASAP7_75t_R _19283_ (.A(_04839_),
    .B(_01379_),
    .Y(_04852_));
 AO21x1_ASAP7_75t_R _19284_ (.A1(_04839_),
    .A2(_04851_),
    .B(_04852_),
    .Y(_04853_));
 OR2x2_ASAP7_75t_R _19285_ (.A(_13123_),
    .B(_00340_),
    .Y(_04854_));
 AO221x1_ASAP7_75t_R _19286_ (.A1(_04847_),
    .A2(_04850_),
    .B1(_04853_),
    .B2(_14091_),
    .C(_04854_),
    .Y(_04855_));
 INVx1_ASAP7_75t_R _19287_ (.A(_01376_),
    .Y(_04856_));
 NAND2x1_ASAP7_75t_R _19288_ (.A(_13093_),
    .B(_01374_),
    .Y(_04857_));
 OA211x2_ASAP7_75t_R _19289_ (.A1(_13093_),
    .A2(_04856_),
    .B(_04857_),
    .C(_13112_),
    .Y(_04858_));
 INVx1_ASAP7_75t_R _19290_ (.A(_01375_),
    .Y(_04859_));
 NAND2x1_ASAP7_75t_R _19291_ (.A(_13093_),
    .B(_01373_),
    .Y(_04860_));
 OA211x2_ASAP7_75t_R _19292_ (.A1(_13093_),
    .A2(_04859_),
    .B(_04860_),
    .C(_00344_),
    .Y(_04861_));
 OR5x1_ASAP7_75t_R _19293_ (.A(_13127_),
    .B(_13083_),
    .C(_13163_),
    .D(_04858_),
    .E(_04861_),
    .Y(_04862_));
 INVx2_ASAP7_75t_R _19294_ (.A(_01372_),
    .Y(_04863_));
 NAND2x1_ASAP7_75t_R _19295_ (.A(_00342_),
    .B(_01368_),
    .Y(_04864_));
 OA211x2_ASAP7_75t_R _19296_ (.A1(_13123_),
    .A2(_04863_),
    .B(_04864_),
    .C(_13112_),
    .Y(_04865_));
 INVx2_ASAP7_75t_R _19297_ (.A(_01371_),
    .Y(_04866_));
 NAND2x1_ASAP7_75t_R _19298_ (.A(_00342_),
    .B(_01367_),
    .Y(_04867_));
 OA211x2_ASAP7_75t_R _19299_ (.A1(_13123_),
    .A2(_04866_),
    .B(_04867_),
    .C(_00344_),
    .Y(_04868_));
 OR5x1_ASAP7_75t_R _19300_ (.A(_13094_),
    .B(_00341_),
    .C(_13081_),
    .D(_04865_),
    .E(_04868_),
    .Y(_04869_));
 OA211x2_ASAP7_75t_R _19301_ (.A1(_04846_),
    .A2(_04855_),
    .B(_04862_),
    .C(_04869_),
    .Y(_04870_));
 INVx1_ASAP7_75t_R _19302_ (.A(_01369_),
    .Y(_04871_));
 NAND2x1_ASAP7_75t_R _19303_ (.A(_13123_),
    .B(_01365_),
    .Y(_04872_));
 OA211x2_ASAP7_75t_R _19304_ (.A1(_13123_),
    .A2(_04871_),
    .B(_04872_),
    .C(_13087_),
    .Y(_04873_));
 INVx1_ASAP7_75t_R _19305_ (.A(_01370_),
    .Y(_04874_));
 NAND2x1_ASAP7_75t_R _19306_ (.A(_00342_),
    .B(_01366_),
    .Y(_04875_));
 OA211x2_ASAP7_75t_R _19307_ (.A1(_13123_),
    .A2(_04874_),
    .B(_04875_),
    .C(_13113_),
    .Y(_04876_));
 OR4x1_ASAP7_75t_R _19308_ (.A(_13091_),
    .B(_13081_),
    .C(_04873_),
    .D(_04876_),
    .Y(_04877_));
 INVx2_ASAP7_75t_R _19309_ (.A(_01383_),
    .Y(_04878_));
 NAND2x1_ASAP7_75t_R _19310_ (.A(_13093_),
    .B(_01381_),
    .Y(_04879_));
 OA211x2_ASAP7_75t_R _19311_ (.A1(_04839_),
    .A2(_04878_),
    .B(_04879_),
    .C(_00344_),
    .Y(_04880_));
 INVx2_ASAP7_75t_R _19312_ (.A(_01384_),
    .Y(_04881_));
 NAND2x1_ASAP7_75t_R _19313_ (.A(_13093_),
    .B(_01382_),
    .Y(_04882_));
 OA211x2_ASAP7_75t_R _19314_ (.A1(_04839_),
    .A2(_04881_),
    .B(_04882_),
    .C(_13112_),
    .Y(_04883_));
 OR4x1_ASAP7_75t_R _19315_ (.A(_13127_),
    .B(_13163_),
    .C(_04880_),
    .D(_04883_),
    .Y(_04884_));
 AO21x2_ASAP7_75t_R _19316_ (.A1(_04877_),
    .A2(_04884_),
    .B(_13104_),
    .Y(_04885_));
 INVx1_ASAP7_75t_R _19317_ (.A(_01364_),
    .Y(_04886_));
 NAND2x1_ASAP7_75t_R _19318_ (.A(_04839_),
    .B(_01362_),
    .Y(_04887_));
 OA211x2_ASAP7_75t_R _19319_ (.A1(_13094_),
    .A2(_04886_),
    .B(_04887_),
    .C(_13113_),
    .Y(_04888_));
 INVx1_ASAP7_75t_R _19320_ (.A(_01363_),
    .Y(_04889_));
 NAND2x1_ASAP7_75t_R _19321_ (.A(_04839_),
    .B(_01361_),
    .Y(_04890_));
 OA211x2_ASAP7_75t_R _19322_ (.A1(_13094_),
    .A2(_04889_),
    .B(_04890_),
    .C(_13087_),
    .Y(_04891_));
 OR3x1_ASAP7_75t_R _19323_ (.A(_13123_),
    .B(_04888_),
    .C(_04891_),
    .Y(_04892_));
 INVx1_ASAP7_75t_R _19324_ (.A(_01359_),
    .Y(_04893_));
 INVx2_ASAP7_75t_R _19325_ (.A(_01360_),
    .Y(_04894_));
 NAND2x1_ASAP7_75t_R _19326_ (.A(_04839_),
    .B(_01765_),
    .Y(_04895_));
 OA21x2_ASAP7_75t_R _19327_ (.A1(_13094_),
    .A2(_04894_),
    .B(_04895_),
    .Y(_04896_));
 AO221x1_ASAP7_75t_R _19328_ (.A1(_04893_),
    .A2(_14449_),
    .B1(_04896_),
    .B2(_13113_),
    .C(_13127_),
    .Y(_04897_));
 NAND2x1_ASAP7_75t_R _19329_ (.A(_00341_),
    .B(_13163_),
    .Y(_04898_));
 AO21x2_ASAP7_75t_R _19330_ (.A1(_04892_),
    .A2(_04897_),
    .B(_04898_),
    .Y(_04899_));
 NAND3x2_ASAP7_75t_R _19331_ (.B(_04885_),
    .C(_04899_),
    .Y(_04900_),
    .A(_04870_));
 AND2x2_ASAP7_75t_R _19332_ (.A(_13279_),
    .B(_13284_),
    .Y(_04901_));
 OR4x1_ASAP7_75t_R _19333_ (.A(_01484_),
    .B(_13285_),
    .C(_13272_),
    .D(_13291_),
    .Y(_04902_));
 OA21x2_ASAP7_75t_R _19334_ (.A1(_04901_),
    .A2(_04902_),
    .B(_13259_),
    .Y(_04903_));
 NAND2x1_ASAP7_75t_R _19335_ (.A(_13252_),
    .B(_13266_),
    .Y(_04904_));
 AND2x2_ASAP7_75t_R _19336_ (.A(_01453_),
    .B(_14380_),
    .Y(_04905_));
 AOI221x1_ASAP7_75t_R _19337_ (.A1(_14446_),
    .A2(_04900_),
    .B1(_04903_),
    .B2(_04904_),
    .C(_04905_),
    .Y(_18072_));
 INVx3_ASAP7_75t_R _19338_ (.A(_18072_),
    .Y(_18070_));
 NAND2x1_ASAP7_75t_R _19339_ (.A(_13753_),
    .B(_01385_),
    .Y(_04906_));
 OA21x2_ASAP7_75t_R _19340_ (.A1(_13738_),
    .A2(_04840_),
    .B(_04906_),
    .Y(_04907_));
 NAND2x1_ASAP7_75t_R _19341_ (.A(_13695_),
    .B(_01386_),
    .Y(_04908_));
 OA211x2_ASAP7_75t_R _19342_ (.A1(_13734_),
    .A2(_04843_),
    .B(_13889_),
    .C(_04908_),
    .Y(_04909_));
 AO21x1_ASAP7_75t_R _19343_ (.A1(_13895_),
    .A2(_04907_),
    .B(_04909_),
    .Y(_04910_));
 NAND2x1_ASAP7_75t_R _19344_ (.A(_13725_),
    .B(_01370_),
    .Y(_04911_));
 OA21x2_ASAP7_75t_R _19345_ (.A1(_13936_),
    .A2(_04863_),
    .B(_04911_),
    .Y(_04912_));
 NAND2x1_ASAP7_75t_R _19346_ (.A(_13695_),
    .B(_01369_),
    .Y(_04913_));
 OA211x2_ASAP7_75t_R _19347_ (.A1(_13734_),
    .A2(_04866_),
    .B(_13903_),
    .C(_04913_),
    .Y(_04914_));
 AO21x1_ASAP7_75t_R _19348_ (.A1(_13900_),
    .A2(_04912_),
    .B(_04914_),
    .Y(_04915_));
 OA211x2_ASAP7_75t_R _19349_ (.A1(_04910_),
    .A2(_04915_),
    .B(_13669_),
    .C(_13688_),
    .Y(_04916_));
 INVx1_ASAP7_75t_R _19350_ (.A(_01368_),
    .Y(_04917_));
 NAND2x1_ASAP7_75t_R _19351_ (.A(_13518_),
    .B(_01366_),
    .Y(_04918_));
 OA211x2_ASAP7_75t_R _19352_ (.A1(_13348_),
    .A2(_04917_),
    .B(_04918_),
    .C(_13369_),
    .Y(_04919_));
 INVx1_ASAP7_75t_R _19353_ (.A(_01367_),
    .Y(_04920_));
 NAND2x1_ASAP7_75t_R _19354_ (.A(_13518_),
    .B(_01365_),
    .Y(_04921_));
 OA211x2_ASAP7_75t_R _19355_ (.A1(_13348_),
    .A2(_04920_),
    .B(_04921_),
    .C(_13322_),
    .Y(_04922_));
 OR3x1_ASAP7_75t_R _19356_ (.A(_13461_),
    .B(_04919_),
    .C(_04922_),
    .Y(_04923_));
 NAND2x1_ASAP7_75t_R _19357_ (.A(_13518_),
    .B(_01382_),
    .Y(_04924_));
 OA211x2_ASAP7_75t_R _19358_ (.A1(_13348_),
    .A2(_04881_),
    .B(_04924_),
    .C(_13369_),
    .Y(_04925_));
 NAND2x1_ASAP7_75t_R _19359_ (.A(_13518_),
    .B(_01381_),
    .Y(_04926_));
 OA211x2_ASAP7_75t_R _19360_ (.A1(_13348_),
    .A2(_04878_),
    .B(_04926_),
    .C(_13322_),
    .Y(_04927_));
 OR3x1_ASAP7_75t_R _19361_ (.A(_13305_),
    .B(_04925_),
    .C(_04927_),
    .Y(_04928_));
 AND4x1_ASAP7_75t_R _19362_ (.A(_13814_),
    .B(_13688_),
    .C(_04923_),
    .D(_04928_),
    .Y(_04929_));
 NOR2x1_ASAP7_75t_R _19363_ (.A(_13725_),
    .B(_01379_),
    .Y(_04930_));
 AO21x1_ASAP7_75t_R _19364_ (.A1(_13738_),
    .A2(_04851_),
    .B(_04930_),
    .Y(_04931_));
 NAND2x1_ASAP7_75t_R _19365_ (.A(_13339_),
    .B(_01378_),
    .Y(_04932_));
 OA211x2_ASAP7_75t_R _19366_ (.A1(_13773_),
    .A2(_04848_),
    .B(_13637_),
    .C(_04932_),
    .Y(_04933_));
 AO21x1_ASAP7_75t_R _19367_ (.A1(_13632_),
    .A2(_04931_),
    .B(_04933_),
    .Y(_04934_));
 NAND2x1_ASAP7_75t_R _19368_ (.A(_13746_),
    .B(_01373_),
    .Y(_04935_));
 NAND2x1_ASAP7_75t_R _19369_ (.A(_13314_),
    .B(_01375_),
    .Y(_04936_));
 NAND2x1_ASAP7_75t_R _19370_ (.A(_13746_),
    .B(_01374_),
    .Y(_04937_));
 NAND2x1_ASAP7_75t_R _19371_ (.A(_13314_),
    .B(_01376_),
    .Y(_04938_));
 AO33x2_ASAP7_75t_R _19372_ (.A1(_13646_),
    .A2(_04935_),
    .A3(_04936_),
    .B1(_04937_),
    .B2(_04938_),
    .B3(_13641_),
    .Y(_04939_));
 OA211x2_ASAP7_75t_R _19373_ (.A1(_04934_),
    .A2(_04939_),
    .B(_13724_),
    .C(_13764_),
    .Y(_04940_));
 NAND2x1_ASAP7_75t_R _19374_ (.A(_13339_),
    .B(_01765_),
    .Y(_04941_));
 OA211x2_ASAP7_75t_R _19375_ (.A1(_13773_),
    .A2(_04894_),
    .B(_04941_),
    .C(_13346_),
    .Y(_04942_));
 AO21x1_ASAP7_75t_R _19376_ (.A1(_04893_),
    .A2(_13476_),
    .B(_04942_),
    .Y(_04943_));
 NAND2x1_ASAP7_75t_R _19377_ (.A(_13518_),
    .B(_01362_),
    .Y(_04944_));
 OA211x2_ASAP7_75t_R _19378_ (.A1(_13348_),
    .A2(_04886_),
    .B(_04944_),
    .C(_13369_),
    .Y(_04945_));
 NAND2x1_ASAP7_75t_R _19379_ (.A(_13378_),
    .B(_01361_),
    .Y(_04946_));
 OA211x2_ASAP7_75t_R _19380_ (.A1(_13701_),
    .A2(_04889_),
    .B(_04946_),
    .C(_13322_),
    .Y(_04947_));
 OR3x1_ASAP7_75t_R _19381_ (.A(_13814_),
    .B(_04945_),
    .C(_04947_),
    .Y(_04948_));
 OA211x2_ASAP7_75t_R _19382_ (.A1(_13669_),
    .A2(_04943_),
    .B(_04948_),
    .C(_13374_),
    .Y(_04949_));
 OR4x1_ASAP7_75t_R _19383_ (.A(_04916_),
    .B(_04929_),
    .C(_04940_),
    .D(_04949_),
    .Y(_04950_));
 AND4x1_ASAP7_75t_R _19384_ (.A(_15367_),
    .B(_13260_),
    .C(_13426_),
    .D(_13833_),
    .Y(_04951_));
 AO21x1_ASAP7_75t_R _19385_ (.A1(_13302_),
    .A2(_04950_),
    .B(_04951_),
    .Y(_04952_));
 BUFx3_ASAP7_75t_R _19386_ (.A(_04952_),
    .Y(_18071_));
 INVx1_ASAP7_75t_R _19387_ (.A(_18071_),
    .Y(_18069_));
 OR2x6_ASAP7_75t_R _19388_ (.A(_01293_),
    .B(_01325_),
    .Y(_04953_));
 OA21x2_ASAP7_75t_R _19389_ (.A1(_01326_),
    .A2(_01325_),
    .B(_01358_),
    .Y(_04954_));
 OA21x2_ASAP7_75t_R _19390_ (.A1(_04720_),
    .A2(_04953_),
    .B(_04954_),
    .Y(_04955_));
 OA21x2_ASAP7_75t_R _19391_ (.A1(_01357_),
    .A2(_04955_),
    .B(_02223_),
    .Y(_04956_));
 XNOR2x2_ASAP7_75t_R _19392_ (.A(_18070_),
    .B(_18071_),
    .Y(_04957_));
 XNOR2x2_ASAP7_75t_R _19393_ (.A(_15241_),
    .B(_04957_),
    .Y(_04958_));
 BUFx6f_ASAP7_75t_R _19394_ (.A(_00029_),
    .Y(_04959_));
 INVx2_ASAP7_75t_R _19395_ (.A(_04959_),
    .Y(_04960_));
 AND2x2_ASAP7_75t_R _19396_ (.A(_04960_),
    .B(_14641_),
    .Y(_04961_));
 AND3x4_ASAP7_75t_R _19397_ (.A(_04870_),
    .B(_04885_),
    .C(_04899_),
    .Y(_04962_));
 BUFx12f_ASAP7_75t_R _19398_ (.A(_04950_),
    .Y(_04963_));
 AOI22x1_ASAP7_75t_R _19399_ (.A1(_14639_),
    .A2(_04959_),
    .B1(_01732_),
    .B2(_14641_),
    .Y(_04964_));
 OA221x2_ASAP7_75t_R _19400_ (.A1(_14633_),
    .A2(_04962_),
    .B1(_04963_),
    .B2(_14642_),
    .C(_04964_),
    .Y(_04965_));
 OA211x2_ASAP7_75t_R _19401_ (.A1(net1953),
    .A2(_18071_),
    .B(_04961_),
    .C(_04965_),
    .Y(_04966_));
 AO221x1_ASAP7_75t_R _19402_ (.A1(_04960_),
    .A2(_14641_),
    .B1(_04963_),
    .B2(_13969_),
    .C(_04951_),
    .Y(_04967_));
 OAI22x1_ASAP7_75t_R _19403_ (.A1(_04961_),
    .A2(_04965_),
    .B1(_04967_),
    .B2(_15241_),
    .Y(_04968_));
 OA21x2_ASAP7_75t_R _19404_ (.A1(_04966_),
    .A2(_04968_),
    .B(_15234_),
    .Y(_04969_));
 AO21x1_ASAP7_75t_R _19405_ (.A1(_14620_),
    .A2(_04958_),
    .B(_04969_),
    .Y(_04970_));
 XOR2x2_ASAP7_75t_R _19406_ (.A(_04956_),
    .B(_04970_),
    .Y(_04971_));
 INVx6_ASAP7_75t_R _19407_ (.A(_04971_),
    .Y(\alu_adder_result_ex[31] ));
 INVx2_ASAP7_75t_R _19408_ (.A(_01357_),
    .Y(_04972_));
 OR2x2_ASAP7_75t_R _19409_ (.A(_04972_),
    .B(_04953_),
    .Y(_04973_));
 OR2x2_ASAP7_75t_R _19410_ (.A(_04723_),
    .B(_04973_),
    .Y(_04974_));
 NOR3x1_ASAP7_75t_R _19411_ (.A(_16756_),
    .B(_16758_),
    .C(_04974_),
    .Y(_04975_));
 AND2x2_ASAP7_75t_R _19412_ (.A(_04972_),
    .B(_04954_),
    .Y(_04976_));
 OA211x2_ASAP7_75t_R _19413_ (.A1(_16756_),
    .A2(_16758_),
    .B(_04727_),
    .C(_04976_),
    .Y(_04977_));
 NAND3x1_ASAP7_75t_R _19414_ (.A(_04972_),
    .B(_04954_),
    .C(_04953_),
    .Y(_04978_));
 OAI21x1_ASAP7_75t_R _19415_ (.A1(_04972_),
    .A2(_04954_),
    .B(_04978_),
    .Y(_04979_));
 NOR2x1_ASAP7_75t_R _19416_ (.A(_04727_),
    .B(_04973_),
    .Y(_04980_));
 AND3x1_ASAP7_75t_R _19417_ (.A(_04727_),
    .B(_04723_),
    .C(_04976_),
    .Y(_04981_));
 OR3x2_ASAP7_75t_R _19418_ (.A(_04979_),
    .B(_04980_),
    .C(_04981_),
    .Y(_04982_));
 NOR3x2_ASAP7_75t_R _19419_ (.B(_04977_),
    .C(_04982_),
    .Y(_04983_),
    .A(_04975_));
 INVx4_ASAP7_75t_R _19420_ (.A(_04983_),
    .Y(\alu_adder_result_ex[30] ));
 INVx2_ASAP7_75t_R _19421_ (.A(_02062_),
    .Y(\cs_registers_i.priv_mode_id_o[0] ));
 AO21x1_ASAP7_75t_R _19422_ (.A1(_14538_),
    .A2(_14582_),
    .B(_14581_),
    .Y(_04984_));
 OR3x1_ASAP7_75t_R _19423_ (.A(_14560_),
    .B(_14563_),
    .C(_04984_),
    .Y(_04985_));
 AND3x4_ASAP7_75t_R _19424_ (.A(_14126_),
    .B(_14140_),
    .C(_04985_),
    .Y(_04986_));
 AND2x6_ASAP7_75t_R _19425_ (.A(_04986_),
    .B(_14115_),
    .Y(_04987_));
 INVx1_ASAP7_75t_R _19426_ (.A(_02231_),
    .Y(_04988_));
 OAI21x1_ASAP7_75t_R _19427_ (.A1(_04988_),
    .A2(_02230_),
    .B(_02229_),
    .Y(_04989_));
 OA21x2_ASAP7_75t_R _19428_ (.A1(_01392_),
    .A2(_02230_),
    .B(_04989_),
    .Y(_04990_));
 BUFx6f_ASAP7_75t_R _19429_ (.A(_00758_),
    .Y(_04991_));
 AO21x1_ASAP7_75t_R _19430_ (.A1(_13613_),
    .A2(_13690_),
    .B(_14142_),
    .Y(_04992_));
 BUFx6f_ASAP7_75t_R _19431_ (.A(_04992_),
    .Y(_04993_));
 AND2x4_ASAP7_75t_R _19432_ (.A(_13839_),
    .B(_14107_),
    .Y(_04994_));
 NAND2x1_ASAP7_75t_R _19433_ (.A(_14202_),
    .B(_04994_),
    .Y(_04995_));
 NAND2x2_ASAP7_75t_R _19434_ (.A(_13995_),
    .B(_14024_),
    .Y(_04996_));
 AOI22x1_ASAP7_75t_R _19435_ (.A1(_14028_),
    .A2(_14035_),
    .B1(_14042_),
    .B2(_14043_),
    .Y(_04997_));
 OR3x1_ASAP7_75t_R _19436_ (.A(_13389_),
    .B(_14048_),
    .C(_14055_),
    .Y(_04998_));
 AOI22x1_ASAP7_75t_R _19437_ (.A1(_13840_),
    .A2(_14063_),
    .B1(_14070_),
    .B2(_13856_),
    .Y(_04999_));
 OA22x2_ASAP7_75t_R _19438_ (.A1(_13716_),
    .A2(_14078_),
    .B1(_14085_),
    .B2(_14086_),
    .Y(_05000_));
 AND4x1_ASAP7_75t_R _19439_ (.A(_04997_),
    .B(_04998_),
    .C(_04999_),
    .D(_05000_),
    .Y(_05001_));
 AOI211x1_ASAP7_75t_R _19440_ (.A1(_13764_),
    .A2(_14159_),
    .B(_14188_),
    .C(_14200_),
    .Y(_05002_));
 OR4x1_ASAP7_75t_R _19441_ (.A(_13763_),
    .B(_04996_),
    .C(_05001_),
    .D(_05002_),
    .Y(_05003_));
 NAND2x1_ASAP7_75t_R _19442_ (.A(_04995_),
    .B(_05003_),
    .Y(_05004_));
 AND2x6_ASAP7_75t_R _19443_ (.A(_14115_),
    .B(_14141_),
    .Y(_05005_));
 BUFx6f_ASAP7_75t_R _19444_ (.A(_05005_),
    .Y(_05006_));
 OR2x6_ASAP7_75t_R _19445_ (.A(_13302_),
    .B(_14270_),
    .Y(_05007_));
 NAND2x2_ASAP7_75t_R _19446_ (.A(_13969_),
    .B(_14260_),
    .Y(_05008_));
 AND4x1_ASAP7_75t_R _19447_ (.A(_18578_),
    .B(_05006_),
    .C(_05007_),
    .D(_05008_),
    .Y(_05009_));
 AND4x1_ASAP7_75t_R _19448_ (.A(_13813_),
    .B(_13861_),
    .C(_13926_),
    .D(_13927_),
    .Y(_05010_));
 AND3x1_ASAP7_75t_R _19449_ (.A(_13328_),
    .B(_13863_),
    .C(_13930_),
    .Y(_05011_));
 OA21x2_ASAP7_75t_R _19450_ (.A1(_05010_),
    .A2(_05011_),
    .B(_13434_),
    .Y(_05012_));
 OA211x2_ASAP7_75t_R _19451_ (.A1(_13920_),
    .A2(_13923_),
    .B(_14191_),
    .C(_13855_),
    .Y(_05013_));
 OR3x2_ASAP7_75t_R _19452_ (.A(_13306_),
    .B(_05012_),
    .C(_05013_),
    .Y(_05014_));
 OA211x2_ASAP7_75t_R _19453_ (.A1(_13913_),
    .A2(_13916_),
    .B(_14191_),
    .C(_13848_),
    .Y(_05015_));
 OR3x1_ASAP7_75t_R _19454_ (.A(_13328_),
    .B(_13872_),
    .C(_13935_),
    .Y(_05016_));
 OR3x1_ASAP7_75t_R _19455_ (.A(_13813_),
    .B(_13869_),
    .C(_13933_),
    .Y(_05017_));
 AOI21x1_ASAP7_75t_R _19456_ (.A1(_05016_),
    .A2(_05017_),
    .B(_14191_),
    .Y(_05018_));
 OR3x1_ASAP7_75t_R _19457_ (.A(_13764_),
    .B(_05015_),
    .C(_05018_),
    .Y(_05019_));
 AND4x1_ASAP7_75t_R _19458_ (.A(_13688_),
    .B(_13969_),
    .C(_05014_),
    .D(_05019_),
    .Y(_05020_));
 AO211x2_ASAP7_75t_R _19459_ (.A1(_13943_),
    .A2(_13950_),
    .B(_13880_),
    .C(_13887_),
    .Y(_05021_));
 OR5x1_ASAP7_75t_R _19460_ (.A(_13814_),
    .B(_13896_),
    .C(_13905_),
    .D(_13958_),
    .E(_13965_),
    .Y(_05022_));
 OAI21x1_ASAP7_75t_R _19461_ (.A1(_13669_),
    .A2(_05021_),
    .B(_05022_),
    .Y(_05023_));
 AO33x2_ASAP7_75t_R _19462_ (.A1(_13837_),
    .A2(_13910_),
    .A3(_13839_),
    .B1(_05023_),
    .B2(_13302_),
    .B3(_13724_),
    .Y(_05024_));
 OA21x2_ASAP7_75t_R _19463_ (.A1(_05020_),
    .A2(_05024_),
    .B(_13768_),
    .Y(_05025_));
 AND5x1_ASAP7_75t_R _19464_ (.A(_04991_),
    .B(_04993_),
    .C(_05004_),
    .D(_05009_),
    .E(_05025_),
    .Y(_05026_));
 NOR2x1_ASAP7_75t_R _19465_ (.A(_04990_),
    .B(_05026_),
    .Y(_05027_));
 AOI21x1_ASAP7_75t_R _19466_ (.A1(_13541_),
    .A2(_13768_),
    .B(_13448_),
    .Y(_05028_));
 AO32x1_ASAP7_75t_R _19467_ (.A1(_14191_),
    .A2(_13407_),
    .A3(_13855_),
    .B1(_13848_),
    .B2(_13840_),
    .Y(_05029_));
 NOR3x1_ASAP7_75t_R _19468_ (.A(_13858_),
    .B(_13865_),
    .C(_13873_),
    .Y(_05030_));
 NOR3x1_ASAP7_75t_R _19469_ (.A(_13389_),
    .B(_13880_),
    .C(_13887_),
    .Y(_05031_));
 NOR3x1_ASAP7_75t_R _19470_ (.A(_13513_),
    .B(_13896_),
    .C(_13905_),
    .Y(_05032_));
 OR4x1_ASAP7_75t_R _19471_ (.A(_05029_),
    .B(_05030_),
    .C(_05031_),
    .D(_05032_),
    .Y(_05033_));
 AO32x1_ASAP7_75t_R _19472_ (.A1(_14191_),
    .A2(_13407_),
    .A3(_13924_),
    .B1(_13917_),
    .B2(_13840_),
    .Y(_05034_));
 NOR3x1_ASAP7_75t_R _19473_ (.A(_13858_),
    .B(_13931_),
    .C(_13938_),
    .Y(_05035_));
 AND3x1_ASAP7_75t_R _19474_ (.A(_13310_),
    .B(_13943_),
    .C(_13950_),
    .Y(_05036_));
 OA21x2_ASAP7_75t_R _19475_ (.A1(_13958_),
    .A2(_13965_),
    .B(_13694_),
    .Y(_05037_));
 OR4x1_ASAP7_75t_R _19476_ (.A(_05034_),
    .B(_05035_),
    .C(_05036_),
    .D(_05037_),
    .Y(_05038_));
 OAI22x1_ASAP7_75t_R _19477_ (.A1(_13375_),
    .A2(_13777_),
    .B1(_13784_),
    .B2(_13386_),
    .Y(_05039_));
 AO32x1_ASAP7_75t_R _19478_ (.A1(_13814_),
    .A2(_13374_),
    .A3(_13788_),
    .B1(_13795_),
    .B2(_13666_),
    .Y(_05040_));
 AO211x2_ASAP7_75t_R _19479_ (.A1(_13808_),
    .A2(_13812_),
    .B(_13821_),
    .C(_13828_),
    .Y(_05041_));
 OA31x2_ASAP7_75t_R _19480_ (.A1(_05039_),
    .A2(_05040_),
    .A3(_05041_),
    .B1(_13301_),
    .Y(_05042_));
 OA21x2_ASAP7_75t_R _19481_ (.A1(_16387_),
    .A2(_14098_),
    .B(_13763_),
    .Y(_05043_));
 AO31x2_ASAP7_75t_R _19482_ (.A1(_05033_),
    .A2(_05038_),
    .A3(_05042_),
    .B(_05043_),
    .Y(_05044_));
 AND3x1_ASAP7_75t_R _19483_ (.A(_13614_),
    .B(_13690_),
    .C(_05044_),
    .Y(_05045_));
 AND5x1_ASAP7_75t_R _19484_ (.A(_13447_),
    .B(_13541_),
    .C(_13691_),
    .D(_05005_),
    .E(_05044_),
    .Y(_05046_));
 AO21x1_ASAP7_75t_R _19485_ (.A1(_05028_),
    .A2(_05045_),
    .B(_05046_),
    .Y(_05047_));
 AO31x2_ASAP7_75t_R _19486_ (.A1(_13785_),
    .A2(_13796_),
    .A3(_13829_),
    .B(_13763_),
    .Y(_05048_));
 OAI21x1_ASAP7_75t_R _19487_ (.A1(_16387_),
    .A2(_14098_),
    .B(_13763_),
    .Y(_05049_));
 OA31x2_ASAP7_75t_R _19488_ (.A1(_13908_),
    .A2(_13968_),
    .A3(_05048_),
    .B1(_05049_),
    .Y(_05050_));
 NAND2x1_ASAP7_75t_R _19489_ (.A(_05006_),
    .B(_05050_),
    .Y(_05051_));
 NAND3x1_ASAP7_75t_R _19490_ (.A(_13447_),
    .B(_13541_),
    .C(_13691_),
    .Y(_05052_));
 AO211x2_ASAP7_75t_R _19491_ (.A1(_13447_),
    .A2(_13541_),
    .B(_13691_),
    .C(_13768_),
    .Y(_05053_));
 OR2x6_ASAP7_75t_R _19492_ (.A(_13447_),
    .B(_13541_),
    .Y(_05054_));
 AND5x1_ASAP7_75t_R _19493_ (.A(_13614_),
    .B(_05051_),
    .C(_05052_),
    .D(_05053_),
    .E(_05054_),
    .Y(_05055_));
 OR4x1_ASAP7_75t_R _19494_ (.A(_13447_),
    .B(_13541_),
    .C(_13690_),
    .D(_05050_),
    .Y(_05056_));
 OAI21x1_ASAP7_75t_R _19495_ (.A1(_13614_),
    .A2(_05050_),
    .B(_05056_),
    .Y(_05057_));
 OR4x1_ASAP7_75t_R _19496_ (.A(_14143_),
    .B(_05047_),
    .C(_05055_),
    .D(_05057_),
    .Y(_05058_));
 AO221x1_ASAP7_75t_R _19497_ (.A1(_13980_),
    .A2(_13984_),
    .B1(_13991_),
    .B2(_13666_),
    .C(_13994_),
    .Y(_05059_));
 NOR3x1_ASAP7_75t_R _19498_ (.A(_13417_),
    .B(_13998_),
    .C(_14001_),
    .Y(_05060_));
 NOR3x1_ASAP7_75t_R _19499_ (.A(_13544_),
    .B(_14005_),
    .C(_14008_),
    .Y(_05061_));
 NOR3x1_ASAP7_75t_R _19500_ (.A(_13375_),
    .B(_14012_),
    .C(_14015_),
    .Y(_05062_));
 NOR3x1_ASAP7_75t_R _19501_ (.A(_13386_),
    .B(_14019_),
    .C(_14022_),
    .Y(_05063_));
 OR4x1_ASAP7_75t_R _19502_ (.A(_05060_),
    .B(_05061_),
    .C(_05062_),
    .D(_05063_),
    .Y(_05064_));
 OR3x1_ASAP7_75t_R _19503_ (.A(_13763_),
    .B(_05059_),
    .C(_05064_),
    .Y(_05065_));
 OR5x1_ASAP7_75t_R _19504_ (.A(_14202_),
    .B(_01512_),
    .C(_01513_),
    .D(_13302_),
    .E(_16387_),
    .Y(_05066_));
 OA31x2_ASAP7_75t_R _19505_ (.A1(_05065_),
    .A2(_05001_),
    .A3(_14201_),
    .B1(_05066_),
    .Y(_05067_));
 OR3x2_ASAP7_75t_R _19506_ (.A(_14143_),
    .B(_18610_),
    .C(_05067_),
    .Y(_05068_));
 INVx4_ASAP7_75t_R _19507_ (.A(_05068_),
    .Y(_05069_));
 AND2x4_ASAP7_75t_R _19508_ (.A(_05058_),
    .B(_05069_),
    .Y(_05070_));
 BUFx6f_ASAP7_75t_R _19509_ (.A(_05006_),
    .Y(_05071_));
 AND3x4_ASAP7_75t_R _19510_ (.A(_13449_),
    .B(_13543_),
    .C(_05071_),
    .Y(_05072_));
 AND2x4_ASAP7_75t_R _19511_ (.A(_18575_),
    .B(_18580_),
    .Y(_05073_));
 AND2x2_ASAP7_75t_R _19512_ (.A(_18563_),
    .B(_14142_),
    .Y(_05074_));
 OA21x2_ASAP7_75t_R _19513_ (.A1(_13614_),
    .A2(_13769_),
    .B(_18580_),
    .Y(_05075_));
 NOR2x2_ASAP7_75t_R _19514_ (.A(_13447_),
    .B(_13541_),
    .Y(_05076_));
 OA21x2_ASAP7_75t_R _19515_ (.A1(_05074_),
    .A2(_05075_),
    .B(_05076_),
    .Y(_05077_));
 AOI21x1_ASAP7_75t_R _19516_ (.A1(_05072_),
    .A2(_05073_),
    .B(_05077_),
    .Y(_05078_));
 OR2x6_ASAP7_75t_R _19517_ (.A(_05020_),
    .B(_05024_),
    .Y(_05079_));
 AO32x2_ASAP7_75t_R _19518_ (.A1(_14025_),
    .A2(_14089_),
    .A3(_05002_),
    .B1(_04994_),
    .B2(_14122_),
    .Y(_05080_));
 BUFx6f_ASAP7_75t_R _19519_ (.A(_05080_),
    .Y(_05081_));
 AND5x2_ASAP7_75t_R _19520_ (.A(_18568_),
    .B(_05071_),
    .C(_18608_),
    .D(_05079_),
    .E(_05081_),
    .Y(_05082_));
 INVx1_ASAP7_75t_R _19521_ (.A(_05082_),
    .Y(_05083_));
 NAND2x1_ASAP7_75t_R _19522_ (.A(_13614_),
    .B(_13769_),
    .Y(_05084_));
 OR3x1_ASAP7_75t_R _19523_ (.A(_13542_),
    .B(_13614_),
    .C(_14142_),
    .Y(_05085_));
 NAND2x1_ASAP7_75t_R _19524_ (.A(_13451_),
    .B(_18570_),
    .Y(_05086_));
 AO21x1_ASAP7_75t_R _19525_ (.A1(_05084_),
    .A2(_05085_),
    .B(_05086_),
    .Y(_05087_));
 AOI21x1_ASAP7_75t_R _19526_ (.A1(_13969_),
    .A2(_13684_),
    .B(_13689_),
    .Y(_05088_));
 AO21x1_ASAP7_75t_R _19527_ (.A1(_05088_),
    .A2(_05071_),
    .B(_13451_),
    .Y(_05089_));
 OA21x2_ASAP7_75t_R _19528_ (.A1(_13448_),
    .A2(_13769_),
    .B(_13542_),
    .Y(_05090_));
 AOI211x1_ASAP7_75t_R _19529_ (.A1(_13614_),
    .A2(_18570_),
    .B(_18573_),
    .C(_13542_),
    .Y(_05091_));
 AOI22x1_ASAP7_75t_R _19530_ (.A1(_05089_),
    .A2(_05090_),
    .B1(_05091_),
    .B2(_13449_),
    .Y(_05092_));
 NOR2x1_ASAP7_75t_R _19531_ (.A(_05020_),
    .B(_05024_),
    .Y(_05093_));
 OR5x1_ASAP7_75t_R _19532_ (.A(_18578_),
    .B(_14143_),
    .C(_18610_),
    .D(_05093_),
    .E(_05067_),
    .Y(_05094_));
 AO21x2_ASAP7_75t_R _19533_ (.A1(_05087_),
    .A2(_05092_),
    .B(_05094_),
    .Y(_05095_));
 OAI21x1_ASAP7_75t_R _19534_ (.A1(_05078_),
    .A2(_05083_),
    .B(_05095_),
    .Y(_05096_));
 AO211x2_ASAP7_75t_R _19535_ (.A1(_13447_),
    .A2(_13541_),
    .B(_13612_),
    .C(_13691_),
    .Y(_05097_));
 AO21x1_ASAP7_75t_R _19536_ (.A1(_05071_),
    .A2(_05097_),
    .B(_13768_),
    .Y(_05098_));
 NAND2x1_ASAP7_75t_R _19537_ (.A(_13837_),
    .B(_13909_),
    .Y(_05099_));
 NAND2x1_ASAP7_75t_R _19538_ (.A(_05033_),
    .B(_05038_),
    .Y(_05100_));
 AOI22x1_ASAP7_75t_R _19539_ (.A1(_13839_),
    .A2(_05099_),
    .B1(_05100_),
    .B2(_13969_),
    .Y(_05101_));
 AND4x1_ASAP7_75t_R _19540_ (.A(_05009_),
    .B(_05081_),
    .C(_05098_),
    .D(_05101_),
    .Y(_05102_));
 AND2x2_ASAP7_75t_R _19541_ (.A(_05079_),
    .B(_05080_),
    .Y(_05103_));
 OA21x2_ASAP7_75t_R _19542_ (.A1(_13612_),
    .A2(_13691_),
    .B(_05006_),
    .Y(_05104_));
 NAND2x1_ASAP7_75t_R _19543_ (.A(_13769_),
    .B(_05104_),
    .Y(_05105_));
 XNOR2x2_ASAP7_75t_R _19544_ (.A(_13612_),
    .B(_18570_),
    .Y(_05106_));
 AND3x4_ASAP7_75t_R _19545_ (.A(_13448_),
    .B(_13542_),
    .C(_18570_),
    .Y(_05107_));
 AOI21x1_ASAP7_75t_R _19546_ (.A1(_05076_),
    .A2(_05106_),
    .B(_05107_),
    .Y(_05108_));
 OA211x2_ASAP7_75t_R _19547_ (.A1(_05020_),
    .A2(_05024_),
    .B(_13768_),
    .C(_05005_),
    .Y(_05109_));
 AND4x1_ASAP7_75t_R _19548_ (.A(_13836_),
    .B(_18608_),
    .C(_05109_),
    .D(_05080_),
    .Y(_05110_));
 AO32x2_ASAP7_75t_R _19549_ (.A1(_05009_),
    .A2(_05103_),
    .A3(_05105_),
    .B1(_05108_),
    .B2(_05110_),
    .Y(_05111_));
 AND2x6_ASAP7_75t_R _19550_ (.A(_13769_),
    .B(_05080_),
    .Y(_05112_));
 AND4x1_ASAP7_75t_R _19551_ (.A(_05005_),
    .B(_05007_),
    .C(_05008_),
    .D(_05044_),
    .Y(_05113_));
 AND2x6_ASAP7_75t_R _19552_ (.A(_05112_),
    .B(_05113_),
    .Y(_05114_));
 AO21x1_ASAP7_75t_R _19553_ (.A1(_14025_),
    .A2(_14089_),
    .B(_04994_),
    .Y(_05115_));
 AND3x1_ASAP7_75t_R _19554_ (.A(_13768_),
    .B(_05006_),
    .C(_05115_),
    .Y(_05116_));
 NAND2x1_ASAP7_75t_R _19555_ (.A(_14201_),
    .B(_14260_),
    .Y(_05117_));
 OR4x1_ASAP7_75t_R _19556_ (.A(_14122_),
    .B(_13969_),
    .C(_16387_),
    .D(_14270_),
    .Y(_05118_));
 OAI21x1_ASAP7_75t_R _19557_ (.A1(_13763_),
    .A2(_05117_),
    .B(_05118_),
    .Y(_05119_));
 AND3x4_ASAP7_75t_R _19558_ (.A(_05044_),
    .B(_05116_),
    .C(_05119_),
    .Y(_05120_));
 AND2x6_ASAP7_75t_R _19559_ (.A(_13612_),
    .B(_13690_),
    .Y(_05121_));
 AND3x1_ASAP7_75t_R _19560_ (.A(_05006_),
    .B(_05076_),
    .C(_05121_),
    .Y(_05122_));
 BUFx6f_ASAP7_75t_R _19561_ (.A(_05122_),
    .Y(_05123_));
 OA21x2_ASAP7_75t_R _19562_ (.A1(_05114_),
    .A2(_05120_),
    .B(_05123_),
    .Y(_05124_));
 OR3x1_ASAP7_75t_R _19563_ (.A(_05102_),
    .B(_05111_),
    .C(_05124_),
    .Y(_05125_));
 AND3x1_ASAP7_75t_R _19564_ (.A(_18552_),
    .B(_18588_),
    .C(_05004_),
    .Y(_05126_));
 AND3x4_ASAP7_75t_R _19565_ (.A(_05005_),
    .B(_05007_),
    .C(_05008_),
    .Y(_05127_));
 AND3x4_ASAP7_75t_R _19566_ (.A(_13769_),
    .B(_13836_),
    .C(_18583_),
    .Y(_05128_));
 AND2x2_ASAP7_75t_R _19567_ (.A(_05127_),
    .B(_05128_),
    .Y(_05129_));
 AND2x6_ASAP7_75t_R _19568_ (.A(_13543_),
    .B(_05071_),
    .Y(_05130_));
 AND2x6_ASAP7_75t_R _19569_ (.A(_18590_),
    .B(_05080_),
    .Y(_05131_));
 AND3x1_ASAP7_75t_R _19570_ (.A(_05127_),
    .B(_05128_),
    .C(_05131_),
    .Y(_05132_));
 BUFx6f_ASAP7_75t_R _19571_ (.A(_05132_),
    .Y(_05133_));
 AND4x1_ASAP7_75t_R _19572_ (.A(_18578_),
    .B(_18610_),
    .C(_05109_),
    .D(_05004_),
    .Y(_05134_));
 AOI221x1_ASAP7_75t_R _19573_ (.A1(_05126_),
    .A2(_05129_),
    .B1(_05130_),
    .B2(_05133_),
    .C(_05134_),
    .Y(_05135_));
 NOR3x2_ASAP7_75t_R _19574_ (.B(_13542_),
    .C(_14142_),
    .Y(_05136_),
    .A(_13446_));
 AND3x4_ASAP7_75t_R _19575_ (.A(_05112_),
    .B(_05113_),
    .C(_05136_),
    .Y(_05137_));
 OAI21x1_ASAP7_75t_R _19576_ (.A1(_13448_),
    .A2(_13542_),
    .B(_05006_),
    .Y(_05138_));
 AND5x1_ASAP7_75t_R _19577_ (.A(_18575_),
    .B(_05009_),
    .C(_05081_),
    .D(_05101_),
    .E(_05138_),
    .Y(_05139_));
 OAI21x1_ASAP7_75t_R _19578_ (.A1(_05137_),
    .A2(_05139_),
    .B(_04993_),
    .Y(_05140_));
 OAI21x1_ASAP7_75t_R _19579_ (.A1(_05104_),
    .A2(_05135_),
    .B(_05140_),
    .Y(_05141_));
 NOR2x2_ASAP7_75t_R _19580_ (.A(_13542_),
    .B(_18568_),
    .Y(_05142_));
 AO33x2_ASAP7_75t_R _19581_ (.A1(_13614_),
    .A2(_05112_),
    .A3(_05113_),
    .B1(_05128_),
    .B2(_05131_),
    .B3(_05127_),
    .Y(_05143_));
 AO31x2_ASAP7_75t_R _19582_ (.A1(_05127_),
    .A2(_05128_),
    .A3(_05131_),
    .B(_18563_),
    .Y(_05144_));
 AO31x2_ASAP7_75t_R _19583_ (.A1(_13448_),
    .A2(_05112_),
    .A3(_05113_),
    .B(_18565_),
    .Y(_05145_));
 AO22x2_ASAP7_75t_R _19584_ (.A1(_13451_),
    .A2(_05143_),
    .B1(_05144_),
    .B2(_05145_),
    .Y(_05146_));
 AND2x2_ASAP7_75t_R _19585_ (.A(_05142_),
    .B(_05146_),
    .Y(_05147_));
 OR5x2_ASAP7_75t_R _19586_ (.A(_05070_),
    .B(_05096_),
    .C(_05125_),
    .D(_05141_),
    .E(_05147_),
    .Y(_05148_));
 AO21x2_ASAP7_75t_R _19587_ (.A1(_05027_),
    .A2(_05148_),
    .B(_14388_),
    .Y(_05149_));
 INVx1_ASAP7_75t_R _19588_ (.A(_02228_),
    .Y(_05150_));
 INVx1_ASAP7_75t_R _19589_ (.A(_05119_),
    .Y(_05151_));
 INVx2_ASAP7_75t_R _19590_ (.A(_01539_),
    .Y(_05152_));
 INVx3_ASAP7_75t_R _19591_ (.A(_01762_),
    .Y(_05153_));
 BUFx6f_ASAP7_75t_R _19592_ (.A(_01763_),
    .Y(_05154_));
 INVx2_ASAP7_75t_R _19593_ (.A(_01761_),
    .Y(_05155_));
 NAND2x1_ASAP7_75t_R _19594_ (.A(_01760_),
    .B(_05155_),
    .Y(_05156_));
 OR3x2_ASAP7_75t_R _19595_ (.A(_05153_),
    .B(_05154_),
    .C(_05156_),
    .Y(_05157_));
 BUFx12f_ASAP7_75t_R _19596_ (.A(_05157_),
    .Y(_05158_));
 OR3x2_ASAP7_75t_R _19597_ (.A(_13233_),
    .B(_05152_),
    .C(_05158_),
    .Y(_05159_));
 OR4x1_ASAP7_75t_R _19598_ (.A(_05150_),
    .B(_14388_),
    .C(_05151_),
    .D(_05159_),
    .Y(_05160_));
 AND3x1_ASAP7_75t_R _19599_ (.A(_04987_),
    .B(_05149_),
    .C(_05160_),
    .Y(_05161_));
 NOR2x1_ASAP7_75t_R _19600_ (.A(_13233_),
    .B(_05161_),
    .Y(_05162_));
 AND3x1_ASAP7_75t_R _19601_ (.A(_13234_),
    .B(_13228_),
    .C(_13265_),
    .Y(_05163_));
 BUFx6f_ASAP7_75t_R _19602_ (.A(_05163_),
    .Y(_05164_));
 AND3x4_ASAP7_75t_R _19603_ (.A(_14105_),
    .B(_14108_),
    .C(_05164_),
    .Y(_05165_));
 NAND2x1_ASAP7_75t_R _19604_ (.A(_14110_),
    .B(_05164_),
    .Y(_05166_));
 NAND3x1_ASAP7_75t_R _19605_ (.A(_14106_),
    .B(_14108_),
    .C(_05164_),
    .Y(_05167_));
 OAI21x1_ASAP7_75t_R _19606_ (.A1(_01833_),
    .A2(_05166_),
    .B(_05167_),
    .Y(_05168_));
 OA21x2_ASAP7_75t_R _19607_ (.A1(_18080_),
    .A2(_02062_),
    .B(_05168_),
    .Y(_05169_));
 AO21x1_ASAP7_75t_R _19608_ (.A1(_04991_),
    .A2(_05165_),
    .B(_05169_),
    .Y(_05170_));
 INVx3_ASAP7_75t_R _19609_ (.A(_01760_),
    .Y(_05171_));
 BUFx6f_ASAP7_75t_R _19610_ (.A(_01761_),
    .Y(_05172_));
 INVx3_ASAP7_75t_R _19611_ (.A(_01763_),
    .Y(_05173_));
 OR4x1_ASAP7_75t_R _19612_ (.A(_05171_),
    .B(_05172_),
    .C(_01762_),
    .D(_05173_),
    .Y(_05174_));
 OA21x2_ASAP7_75t_R _19613_ (.A1(_05162_),
    .A2(_05170_),
    .B(_05174_),
    .Y(\id_stage_i.controller_i.illegal_insn_d ));
 NAND2x1_ASAP7_75t_R _19614_ (.A(_14103_),
    .B(_05164_),
    .Y(_05175_));
 AND4x1_ASAP7_75t_R _19615_ (.A(_01539_),
    .B(_04987_),
    .C(_05160_),
    .D(_05175_),
    .Y(_05176_));
 AOI21x1_ASAP7_75t_R _19616_ (.A1(_05149_),
    .A2(_05176_),
    .B(_13233_),
    .Y(_05177_));
 OA21x2_ASAP7_75t_R _19617_ (.A1(_05170_),
    .A2(_05177_),
    .B(_05174_),
    .Y(\id_stage_i.controller_i.exc_req_d ));
 BUFx6f_ASAP7_75t_R _19618_ (.A(_01393_),
    .Y(_05178_));
 BUFx6f_ASAP7_75t_R _19619_ (.A(_05178_),
    .Y(_05179_));
 BUFx6f_ASAP7_75t_R _19620_ (.A(_01443_),
    .Y(_05180_));
 AND4x1_ASAP7_75t_R _19621_ (.A(_00375_),
    .B(net80),
    .C(_05180_),
    .D(_01444_),
    .Y(_05181_));
 INVx1_ASAP7_75t_R _19622_ (.A(net25),
    .Y(_05182_));
 NAND2x1_ASAP7_75t_R _19623_ (.A(_05182_),
    .B(_01442_),
    .Y(_05183_));
 NAND2x1_ASAP7_75t_R _19624_ (.A(_05181_),
    .B(_05183_),
    .Y(_05184_));
 NOR2x1_ASAP7_75t_R _19625_ (.A(_05179_),
    .B(_05184_),
    .Y(\id_stage_i.controller_i.store_err_i ));
 AND3x1_ASAP7_75t_R _19626_ (.A(_05179_),
    .B(_05181_),
    .C(_05183_),
    .Y(\id_stage_i.controller_i.load_err_i ));
 INVx1_ASAP7_75t_R _19627_ (.A(_01395_),
    .Y(_05185_));
 BUFx6f_ASAP7_75t_R _19628_ (.A(_00026_),
    .Y(_05186_));
 BUFx6f_ASAP7_75t_R _19629_ (.A(_00027_),
    .Y(_05187_));
 AND4x1_ASAP7_75t_R _19630_ (.A(_05185_),
    .B(_01394_),
    .C(_05186_),
    .D(_05187_),
    .Y(_05188_));
 AND2x6_ASAP7_75t_R _19631_ (.A(_01760_),
    .B(_05155_),
    .Y(_05189_));
 AND3x4_ASAP7_75t_R _19632_ (.A(_01762_),
    .B(_05173_),
    .C(_05189_),
    .Y(_05190_));
 AND3x4_ASAP7_75t_R _19633_ (.A(_13234_),
    .B(_01539_),
    .C(_05190_),
    .Y(_05191_));
 AND3x4_ASAP7_75t_R _19634_ (.A(_04986_),
    .B(_14115_),
    .C(_05191_),
    .Y(_05192_));
 BUFx12f_ASAP7_75t_R _19635_ (.A(_05192_),
    .Y(_05193_));
 AND2x6_ASAP7_75t_R _19636_ (.A(_14541_),
    .B(_14623_),
    .Y(_05194_));
 AND2x6_ASAP7_75t_R _19637_ (.A(_05193_),
    .B(_05194_),
    .Y(_05195_));
 BUFx6f_ASAP7_75t_R _19638_ (.A(_05195_),
    .Y(_05196_));
 BUFx6f_ASAP7_75t_R _19639_ (.A(_01798_),
    .Y(_05197_));
 BUFx6f_ASAP7_75t_R _19640_ (.A(_05197_),
    .Y(_05198_));
 AO21x1_ASAP7_75t_R _19641_ (.A1(_05188_),
    .A2(_05196_),
    .B(_05198_),
    .Y(_05199_));
 INVx5_ASAP7_75t_R _19642_ (.A(_02193_),
    .Y(_05200_));
 NAND2x2_ASAP7_75t_R _19643_ (.A(_05200_),
    .B(_05195_),
    .Y(_05201_));
 BUFx6f_ASAP7_75t_R _19644_ (.A(_05201_),
    .Y(_05202_));
 NAND2x1_ASAP7_75t_R _19645_ (.A(_05199_),
    .B(_05202_),
    .Y(_00005_));
 BUFx12f_ASAP7_75t_R _19646_ (.A(_14634_),
    .Y(_05203_));
 BUFx6f_ASAP7_75t_R _19647_ (.A(_05195_),
    .Y(_05204_));
 NAND2x2_ASAP7_75t_R _19648_ (.A(_05193_),
    .B(_05194_),
    .Y(_05205_));
 BUFx6f_ASAP7_75t_R _19649_ (.A(_05205_),
    .Y(_05206_));
 INVx2_ASAP7_75t_R _19650_ (.A(\alu_adder_result_ex[6] ),
    .Y(_05207_));
 BUFx6f_ASAP7_75t_R _19651_ (.A(_18708_),
    .Y(_05208_));
 INVx4_ASAP7_75t_R _19652_ (.A(_05208_),
    .Y(_05209_));
 OA21x2_ASAP7_75t_R _19653_ (.A1(_15033_),
    .A2(_15034_),
    .B(_15035_),
    .Y(_05210_));
 OA21x2_ASAP7_75t_R _19654_ (.A1(_15029_),
    .A2(_05210_),
    .B(_00768_),
    .Y(_05211_));
 XNOR2x1_ASAP7_75t_R _19655_ (.B(_05211_),
    .Y(_05212_),
    .A(_00767_));
 OA21x2_ASAP7_75t_R _19656_ (.A1(_00761_),
    .A2(_15033_),
    .B(_00764_),
    .Y(_05213_));
 XNOR2x1_ASAP7_75t_R _19657_ (.B(_05213_),
    .Y(_05214_),
    .A(_00763_));
 AND4x1_ASAP7_75t_R _19658_ (.A(_05209_),
    .B(_15040_),
    .C(_05212_),
    .D(_05214_),
    .Y(_05215_));
 AND4x1_ASAP7_75t_R _19659_ (.A(_15166_),
    .B(_15518_),
    .C(_16515_),
    .D(_05215_),
    .Y(_05216_));
 AND5x1_ASAP7_75t_R _19660_ (.A(_15240_),
    .B(_15764_),
    .C(_16004_),
    .D(_16253_),
    .E(_05216_),
    .Y(_05217_));
 OA21x2_ASAP7_75t_R _19661_ (.A1(_14621_),
    .A2(_15044_),
    .B(_15042_),
    .Y(_05218_));
 XNOR2x1_ASAP7_75t_R _19662_ (.B(_05218_),
    .Y(_05219_),
    .A(_00761_));
 AND5x1_ASAP7_75t_R _19663_ (.A(_05207_),
    .B(_16753_),
    .C(_04480_),
    .D(_05217_),
    .E(_05219_),
    .Y(_05220_));
 OA211x2_ASAP7_75t_R _19664_ (.A1(_15241_),
    .A2(_15170_),
    .B(_15172_),
    .C(_00766_),
    .Y(_05221_));
 INVx1_ASAP7_75t_R _19665_ (.A(_15170_),
    .Y(_05222_));
 INVx1_ASAP7_75t_R _19666_ (.A(_15172_),
    .Y(_05223_));
 NAND2x1_ASAP7_75t_R _19667_ (.A(_00766_),
    .B(_15029_),
    .Y(_05224_));
 AO211x2_ASAP7_75t_R _19668_ (.A1(_14632_),
    .A2(_05222_),
    .B(_05223_),
    .C(_05224_),
    .Y(_05225_));
 OAI21x1_ASAP7_75t_R _19669_ (.A1(_15029_),
    .A2(_05221_),
    .B(_05225_),
    .Y(_05226_));
 AND4x1_ASAP7_75t_R _19670_ (.A(_15248_),
    .B(_15524_),
    .C(_15772_),
    .D(_05226_),
    .Y(_05227_));
 AND3x1_ASAP7_75t_R _19671_ (.A(_15179_),
    .B(_16995_),
    .C(_04722_),
    .Y(_05228_));
 AND4x1_ASAP7_75t_R _19672_ (.A(_16267_),
    .B(_05220_),
    .C(_05227_),
    .D(_05228_),
    .Y(_05229_));
 AND4x1_ASAP7_75t_R _19673_ (.A(_16019_),
    .B(_16528_),
    .C(_16761_),
    .D(_04495_),
    .Y(_05230_));
 NAND2x1_ASAP7_75t_R _19674_ (.A(_05229_),
    .B(_05230_),
    .Y(_05231_));
 OR4x1_ASAP7_75t_R _19675_ (.A(\alu_adder_result_ex[24] ),
    .B(\alu_adder_result_ex[28] ),
    .C(\alu_adder_result_ex[31] ),
    .D(\alu_adder_result_ex[30] ),
    .Y(_05232_));
 NOR2x1_ASAP7_75t_R _19676_ (.A(_05231_),
    .B(_05232_),
    .Y(_05233_));
 OR3x1_ASAP7_75t_R _19677_ (.A(_02192_),
    .B(_05206_),
    .C(_05233_),
    .Y(_05234_));
 OAI21x1_ASAP7_75t_R _19678_ (.A1(_05203_),
    .A2(_05204_),
    .B(_05234_),
    .Y(_00004_));
 AND2x6_ASAP7_75t_R _19679_ (.A(_14534_),
    .B(_14624_),
    .Y(_05235_));
 NAND2x2_ASAP7_75t_R _19680_ (.A(_05193_),
    .B(_05235_),
    .Y(_05236_));
 BUFx12f_ASAP7_75t_R _19681_ (.A(_01397_),
    .Y(_05237_));
 AO21x1_ASAP7_75t_R _19682_ (.A1(_14119_),
    .A2(_14624_),
    .B(_02194_),
    .Y(_05238_));
 AND4x1_ASAP7_75t_R _19683_ (.A(_05237_),
    .B(_05193_),
    .C(_05235_),
    .D(_05238_),
    .Y(_05239_));
 AOI21x1_ASAP7_75t_R _19684_ (.A1(_02197_),
    .A2(_05236_),
    .B(_05239_),
    .Y(_00000_));
 AND2x4_ASAP7_75t_R _19685_ (.A(_14533_),
    .B(_15234_),
    .Y(_05240_));
 BUFx6f_ASAP7_75t_R _19686_ (.A(_05240_),
    .Y(_05241_));
 BUFx6f_ASAP7_75t_R _19687_ (.A(_05241_),
    .Y(_05242_));
 OR3x2_ASAP7_75t_R _19688_ (.A(_02194_),
    .B(_13228_),
    .C(_14620_),
    .Y(_05243_));
 BUFx6f_ASAP7_75t_R _19689_ (.A(_05243_),
    .Y(_05244_));
 AND3x1_ASAP7_75t_R _19690_ (.A(_05193_),
    .B(_05242_),
    .C(_05244_),
    .Y(_05245_));
 AOI21x1_ASAP7_75t_R _19691_ (.A1(_05237_),
    .A2(_05236_),
    .B(_05245_),
    .Y(_00001_));
 INVx3_ASAP7_75t_R _19692_ (.A(_02198_),
    .Y(_05246_));
 BUFx6f_ASAP7_75t_R _19693_ (.A(_05246_),
    .Y(_05247_));
 INVx2_ASAP7_75t_R _19694_ (.A(_01798_),
    .Y(_05248_));
 BUFx6f_ASAP7_75t_R _19695_ (.A(_05248_),
    .Y(_05249_));
 AND3x1_ASAP7_75t_R _19696_ (.A(_05249_),
    .B(_05188_),
    .C(_05196_),
    .Y(_05250_));
 AO21x1_ASAP7_75t_R _19697_ (.A1(_05247_),
    .A2(_05206_),
    .B(_05250_),
    .Y(_00002_));
 INVx1_ASAP7_75t_R _19698_ (.A(_05233_),
    .Y(_05251_));
 BUFx6f_ASAP7_75t_R _19699_ (.A(_14636_),
    .Y(_05252_));
 OA211x2_ASAP7_75t_R _19700_ (.A1(_02192_),
    .A2(_05251_),
    .B(_05196_),
    .C(_05252_),
    .Y(_05253_));
 AOI21x1_ASAP7_75t_R _19701_ (.A1(_02199_),
    .A2(_05206_),
    .B(_05253_),
    .Y(_00003_));
 INVx1_ASAP7_75t_R _19702_ (.A(_00748_),
    .Y(\cs_registers_i.mhpmcounter[1856] ));
 INVx2_ASAP7_75t_R _19703_ (.A(_00747_),
    .Y(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ));
 INVx3_ASAP7_75t_R _19704_ (.A(_05219_),
    .Y(\alu_adder_result_ex[2] ));
 INVx3_ASAP7_75t_R _19705_ (.A(_05214_),
    .Y(\alu_adder_result_ex[3] ));
 INVx3_ASAP7_75t_R _19706_ (.A(_05226_),
    .Y(\alu_adder_result_ex[4] ));
 INVx3_ASAP7_75t_R _19707_ (.A(_05212_),
    .Y(\alu_adder_result_ex[5] ));
 INVx1_ASAP7_75t_R _19708_ (.A(_18084_),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ));
 BUFx6f_ASAP7_75t_R _19709_ (.A(_18083_),
    .Y(_05254_));
 INVx3_ASAP7_75t_R _19710_ (.A(_05254_),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ));
 BUFx12f_ASAP7_75t_R _19711_ (.A(\alu_adder_result_ex[0] ),
    .Y(_05255_));
 INVx2_ASAP7_75t_R _19712_ (.A(_05255_),
    .Y(_16999_));
 BUFx6f_ASAP7_75t_R _19713_ (.A(_05244_),
    .Y(_05256_));
 AND2x6_ASAP7_75t_R _19714_ (.A(_05237_),
    .B(_02195_),
    .Y(_05257_));
 BUFx6f_ASAP7_75t_R _19715_ (.A(_05257_),
    .Y(_05258_));
 AND2x6_ASAP7_75t_R _19716_ (.A(_05238_),
    .B(_05258_),
    .Y(_05259_));
 BUFx6f_ASAP7_75t_R _19717_ (.A(_05259_),
    .Y(_05260_));
 OAI22x1_ASAP7_75t_R _19718_ (.A1(_00062_),
    .A2(_05256_),
    .B1(_05260_),
    .B2(_15836_),
    .Y(_18089_));
 INVx2_ASAP7_75t_R _19719_ (.A(_15884_),
    .Y(_05261_));
 NAND2x2_ASAP7_75t_R _19720_ (.A(_05237_),
    .B(_02195_),
    .Y(_05262_));
 AND2x2_ASAP7_75t_R _19721_ (.A(_13420_),
    .B(_05257_),
    .Y(_05263_));
 AO21x1_ASAP7_75t_R _19722_ (.A1(_05261_),
    .A2(_05262_),
    .B(_05263_),
    .Y(_05264_));
 BUFx6f_ASAP7_75t_R _19723_ (.A(_05264_),
    .Y(_05265_));
 NAND2x2_ASAP7_75t_R _19724_ (.A(_05237_),
    .B(_02194_),
    .Y(_05266_));
 BUFx6f_ASAP7_75t_R _19725_ (.A(_05266_),
    .Y(_05267_));
 AND2x6_ASAP7_75t_R _19726_ (.A(_05237_),
    .B(_02194_),
    .Y(_05268_));
 AND3x1_ASAP7_75t_R _19727_ (.A(_14416_),
    .B(_14443_),
    .C(_05268_),
    .Y(_05269_));
 AO21x2_ASAP7_75t_R _19728_ (.A1(_15831_),
    .A2(_05267_),
    .B(_05269_),
    .Y(_05270_));
 BUFx6f_ASAP7_75t_R _19729_ (.A(_05270_),
    .Y(_05271_));
 AND2x2_ASAP7_75t_R _19730_ (.A(_05265_),
    .B(_05271_),
    .Y(_18090_));
 OA22x2_ASAP7_75t_R _19731_ (.A1(_00097_),
    .A2(_05256_),
    .B1(_05260_),
    .B2(_15947_),
    .Y(_17001_));
 OA22x2_ASAP7_75t_R _19732_ (.A1(_00100_),
    .A2(_05256_),
    .B1(_05260_),
    .B2(_16083_),
    .Y(_17005_));
 AND3x1_ASAP7_75t_R _19733_ (.A(_16105_),
    .B(_16130_),
    .C(_05262_),
    .Y(_05272_));
 AO21x2_ASAP7_75t_R _19734_ (.A1(_13601_),
    .A2(_05258_),
    .B(_05272_),
    .Y(_05273_));
 BUFx6f_ASAP7_75t_R _19735_ (.A(_05273_),
    .Y(_05274_));
 AND2x2_ASAP7_75t_R _19736_ (.A(_05271_),
    .B(_05274_),
    .Y(_17007_));
 BUFx6f_ASAP7_75t_R _19737_ (.A(_05244_),
    .Y(_05275_));
 OA22x2_ASAP7_75t_R _19738_ (.A1(_00104_),
    .A2(_05275_),
    .B1(_05260_),
    .B2(_16195_),
    .Y(_17014_));
 OA22x2_ASAP7_75t_R _19739_ (.A1(_00109_),
    .A2(_05275_),
    .B1(_05260_),
    .B2(_16329_),
    .Y(_17020_));
 AND3x4_ASAP7_75t_R _19740_ (.A(_14677_),
    .B(_14702_),
    .C(_05268_),
    .Y(_05276_));
 AO21x2_ASAP7_75t_R _19741_ (.A1(_16078_),
    .A2(_05267_),
    .B(_05276_),
    .Y(_05277_));
 AND2x2_ASAP7_75t_R _19742_ (.A(_05274_),
    .B(_05277_),
    .Y(_17025_));
 AND3x1_ASAP7_75t_R _19743_ (.A(_16217_),
    .B(_16241_),
    .C(_05262_),
    .Y(_05278_));
 AO21x2_ASAP7_75t_R _19744_ (.A1(_13684_),
    .A2(_05258_),
    .B(_05278_),
    .Y(_05279_));
 BUFx12f_ASAP7_75t_R _19745_ (.A(_05279_),
    .Y(_05280_));
 AND2x6_ASAP7_75t_R _19746_ (.A(_15912_),
    .B(_15943_),
    .Y(_05281_));
 AND3x4_ASAP7_75t_R _19747_ (.A(_14486_),
    .B(_14527_),
    .C(_05268_),
    .Y(_05282_));
 AO21x2_ASAP7_75t_R _19748_ (.A1(_05281_),
    .A2(_05267_),
    .B(_05282_),
    .Y(_05283_));
 BUFx12f_ASAP7_75t_R _19749_ (.A(_05283_),
    .Y(_05284_));
 AND2x4_ASAP7_75t_R _19750_ (.A(_05280_),
    .B(_05284_),
    .Y(_17024_));
 BUFx6f_ASAP7_75t_R _19751_ (.A(_05262_),
    .Y(_05285_));
 AND2x2_ASAP7_75t_R _19752_ (.A(_13762_),
    .B(_05257_),
    .Y(_05286_));
 AO21x2_ASAP7_75t_R _19753_ (.A1(_16384_),
    .A2(_05285_),
    .B(_05286_),
    .Y(_05287_));
 BUFx6f_ASAP7_75t_R _19754_ (.A(_05287_),
    .Y(_05288_));
 AND2x2_ASAP7_75t_R _19755_ (.A(_05271_),
    .B(_05288_),
    .Y(_17023_));
 OA22x2_ASAP7_75t_R _19756_ (.A1(_00114_),
    .A2(_05275_),
    .B1(_05260_),
    .B2(_00115_),
    .Y(_17036_));
 OA22x2_ASAP7_75t_R _19757_ (.A1(_00121_),
    .A2(_05275_),
    .B1(_05260_),
    .B2(_16591_),
    .Y(_17048_));
 BUFx6f_ASAP7_75t_R _19758_ (.A(_05268_),
    .Y(_05289_));
 AND3x1_ASAP7_75t_R _19759_ (.A(_16294_),
    .B(_16325_),
    .C(_05266_),
    .Y(_05290_));
 AO21x2_ASAP7_75t_R _19760_ (.A1(_14835_),
    .A2(_05289_),
    .B(_05290_),
    .Y(_05291_));
 AND2x2_ASAP7_75t_R _19761_ (.A(_05274_),
    .B(_05291_),
    .Y(_17053_));
 AND3x1_ASAP7_75t_R _19762_ (.A(_16159_),
    .B(_16190_),
    .C(_05266_),
    .Y(_05292_));
 AO21x2_ASAP7_75t_R _19763_ (.A1(_14770_),
    .A2(_05289_),
    .B(_05292_),
    .Y(_05293_));
 BUFx6f_ASAP7_75t_R _19764_ (.A(_05293_),
    .Y(_05294_));
 AND2x4_ASAP7_75t_R _19765_ (.A(_05280_),
    .B(_05294_),
    .Y(_17052_));
 AND2x2_ASAP7_75t_R _19766_ (.A(_05277_),
    .B(_05288_),
    .Y(_17051_));
 OA22x2_ASAP7_75t_R _19767_ (.A1(_00128_),
    .A2(_05275_),
    .B1(_05260_),
    .B2(_16701_),
    .Y(_17066_));
 AND2x6_ASAP7_75t_R _19768_ (.A(_16417_),
    .B(_16448_),
    .Y(_05295_));
 AND3x1_ASAP7_75t_R _19769_ (.A(_14869_),
    .B(_14898_),
    .C(_05289_),
    .Y(_05296_));
 AO21x2_ASAP7_75t_R _19770_ (.A1(_05295_),
    .A2(_05267_),
    .B(_05296_),
    .Y(_05297_));
 AND2x2_ASAP7_75t_R _19771_ (.A(_05274_),
    .B(_05297_),
    .Y(_17071_));
 AND2x4_ASAP7_75t_R _19772_ (.A(_05280_),
    .B(_05291_),
    .Y(_17070_));
 AND2x2_ASAP7_75t_R _19773_ (.A(_05288_),
    .B(_05294_),
    .Y(_17069_));
 BUFx12f_ASAP7_75t_R _19774_ (.A(_05277_),
    .Y(_05298_));
 AND2x2_ASAP7_75t_R _19775_ (.A(_13830_),
    .B(_05257_),
    .Y(_05299_));
 AO21x2_ASAP7_75t_R _19776_ (.A1(_16498_),
    .A2(_05285_),
    .B(_05299_),
    .Y(_05300_));
 BUFx6f_ASAP7_75t_R _19777_ (.A(_05300_),
    .Y(_05301_));
 BUFx12f_ASAP7_75t_R _19778_ (.A(_05301_),
    .Y(_05302_));
 NAND2x1_ASAP7_75t_R _19779_ (.A(_05298_),
    .B(_05302_),
    .Y(_17078_));
 OA22x2_ASAP7_75t_R _19780_ (.A1(_00135_),
    .A2(_05275_),
    .B1(_05260_),
    .B2(_16823_),
    .Y(_17094_));
 AND2x6_ASAP7_75t_R _19781_ (.A(_14936_),
    .B(_14964_),
    .Y(_05303_));
 AND3x1_ASAP7_75t_R _19782_ (.A(_16555_),
    .B(_16586_),
    .C(_05266_),
    .Y(_05304_));
 AO21x2_ASAP7_75t_R _19783_ (.A1(_05303_),
    .A2(_05289_),
    .B(_05304_),
    .Y(_05305_));
 BUFx12f_ASAP7_75t_R _19784_ (.A(_05305_),
    .Y(_05306_));
 AND2x2_ASAP7_75t_R _19785_ (.A(_05274_),
    .B(_05306_),
    .Y(_17099_));
 AND2x4_ASAP7_75t_R _19786_ (.A(_05280_),
    .B(_05297_),
    .Y(_17098_));
 AND2x2_ASAP7_75t_R _19787_ (.A(_05288_),
    .B(_05291_),
    .Y(_17097_));
 BUFx12f_ASAP7_75t_R _19788_ (.A(_05294_),
    .Y(_05307_));
 NAND2x1_ASAP7_75t_R _19789_ (.A(_05307_),
    .B(_05302_),
    .Y(_17106_));
 OA22x2_ASAP7_75t_R _19790_ (.A1(_00144_),
    .A2(_05275_),
    .B1(_05260_),
    .B2(_16935_),
    .Y(_17116_));
 AND2x6_ASAP7_75t_R _19791_ (.A(_16665_),
    .B(_16696_),
    .Y(_05308_));
 AND3x1_ASAP7_75t_R _19792_ (.A(_14998_),
    .B(_15023_),
    .C(_05289_),
    .Y(_05309_));
 AO21x2_ASAP7_75t_R _19793_ (.A1(_05308_),
    .A2(_05267_),
    .B(_05309_),
    .Y(_05310_));
 AND2x2_ASAP7_75t_R _19794_ (.A(_05274_),
    .B(_05310_),
    .Y(_17121_));
 AND2x4_ASAP7_75t_R _19795_ (.A(_05280_),
    .B(_05305_),
    .Y(_17120_));
 AND2x2_ASAP7_75t_R _19796_ (.A(_05288_),
    .B(_05297_),
    .Y(_17119_));
 BUFx12f_ASAP7_75t_R _19797_ (.A(_05291_),
    .Y(_05311_));
 NAND2x1_ASAP7_75t_R _19798_ (.A(_05311_),
    .B(_05302_),
    .Y(_17127_));
 OA22x2_ASAP7_75t_R _19799_ (.A1(_00152_),
    .A2(_05275_),
    .B1(_05259_),
    .B2(_04310_),
    .Y(_17143_));
 AND3x1_ASAP7_75t_R _19800_ (.A(_16788_),
    .B(_16819_),
    .C(_05266_),
    .Y(_05312_));
 AO21x2_ASAP7_75t_R _19801_ (.A1(_15098_),
    .A2(_05289_),
    .B(_05312_),
    .Y(_05313_));
 AND2x2_ASAP7_75t_R _19802_ (.A(_05274_),
    .B(_05313_),
    .Y(_17148_));
 AND2x4_ASAP7_75t_R _19803_ (.A(_05280_),
    .B(_05310_),
    .Y(_17147_));
 AND2x2_ASAP7_75t_R _19804_ (.A(_05288_),
    .B(_05305_),
    .Y(_17146_));
 BUFx12f_ASAP7_75t_R _19805_ (.A(_05297_),
    .Y(_05314_));
 NAND2x1_ASAP7_75t_R _19806_ (.A(_05314_),
    .B(_05302_),
    .Y(_17153_));
 AND3x1_ASAP7_75t_R _19807_ (.A(_13995_),
    .B(_14024_),
    .C(_05257_),
    .Y(_05315_));
 AO21x1_ASAP7_75t_R _19808_ (.A1(_16870_),
    .A2(_05285_),
    .B(_05315_),
    .Y(_05316_));
 BUFx6f_ASAP7_75t_R _19809_ (.A(_05316_),
    .Y(_05317_));
 BUFx6f_ASAP7_75t_R _19810_ (.A(_05317_),
    .Y(_05318_));
 NAND2x1_ASAP7_75t_R _19811_ (.A(_05298_),
    .B(_05318_),
    .Y(_17163_));
 OA22x2_ASAP7_75t_R _19812_ (.A1(_00160_),
    .A2(_05275_),
    .B1(_05259_),
    .B2(_04422_),
    .Y(_17172_));
 AND3x1_ASAP7_75t_R _19813_ (.A(_15132_),
    .B(_15156_),
    .C(_05289_),
    .Y(_05319_));
 AO21x2_ASAP7_75t_R _19814_ (.A1(_16931_),
    .A2(_05267_),
    .B(_05319_),
    .Y(_05320_));
 AND2x2_ASAP7_75t_R _19815_ (.A(_05274_),
    .B(_05320_),
    .Y(_17177_));
 AND2x4_ASAP7_75t_R _19816_ (.A(_05280_),
    .B(_05313_),
    .Y(_17176_));
 AND2x2_ASAP7_75t_R _19817_ (.A(_05288_),
    .B(_05310_),
    .Y(_17175_));
 NAND2x1_ASAP7_75t_R _19818_ (.A(_05302_),
    .B(_05306_),
    .Y(_17183_));
 NAND2x1_ASAP7_75t_R _19819_ (.A(_05307_),
    .B(_05318_),
    .Y(_17193_));
 AND3x1_ASAP7_75t_R _19820_ (.A(_04444_),
    .B(_04467_),
    .C(_05285_),
    .Y(_05321_));
 AO21x2_ASAP7_75t_R _19821_ (.A1(_14260_),
    .A2(_05258_),
    .B(_05321_),
    .Y(_05322_));
 BUFx6f_ASAP7_75t_R _19822_ (.A(_05322_),
    .Y(_05323_));
 AND2x4_ASAP7_75t_R _19823_ (.A(_05271_),
    .B(_05323_),
    .Y(_17195_));
 OA22x2_ASAP7_75t_R _19824_ (.A1(_00168_),
    .A2(_05275_),
    .B1(_05259_),
    .B2(_04558_),
    .Y(_17210_));
 AND2x6_ASAP7_75t_R _19825_ (.A(_15204_),
    .B(_15227_),
    .Y(_05324_));
 AND3x1_ASAP7_75t_R _19826_ (.A(_04273_),
    .B(_04304_),
    .C(_05266_),
    .Y(_05325_));
 AO21x2_ASAP7_75t_R _19827_ (.A1(_05324_),
    .A2(_05289_),
    .B(_05325_),
    .Y(_05326_));
 AND2x2_ASAP7_75t_R _19828_ (.A(_05273_),
    .B(_05326_),
    .Y(_17215_));
 AND2x4_ASAP7_75t_R _19829_ (.A(_05279_),
    .B(_05320_),
    .Y(_17214_));
 AND2x2_ASAP7_75t_R _19830_ (.A(_05287_),
    .B(_05313_),
    .Y(_17213_));
 BUFx12f_ASAP7_75t_R _19831_ (.A(_05310_),
    .Y(_05327_));
 NAND2x1_ASAP7_75t_R _19832_ (.A(_05302_),
    .B(_05327_),
    .Y(_17221_));
 NAND2x1_ASAP7_75t_R _19833_ (.A(_05311_),
    .B(_05318_),
    .Y(_17230_));
 OA22x2_ASAP7_75t_R _19834_ (.A1(_00175_),
    .A2(_05244_),
    .B1(_05259_),
    .B2(_04670_),
    .Y(_17242_));
 AND2x6_ASAP7_75t_R _19835_ (.A(_14338_),
    .B(_14376_),
    .Y(_05328_));
 AND3x1_ASAP7_75t_R _19836_ (.A(_04386_),
    .B(_04417_),
    .C(_05266_),
    .Y(_05329_));
 AO21x2_ASAP7_75t_R _19837_ (.A1(_05328_),
    .A2(_05289_),
    .B(_05329_),
    .Y(_05330_));
 AND2x2_ASAP7_75t_R _19838_ (.A(_05273_),
    .B(_05330_),
    .Y(_17247_));
 AND2x4_ASAP7_75t_R _19839_ (.A(_05279_),
    .B(_05326_),
    .Y(_17246_));
 AND2x2_ASAP7_75t_R _19840_ (.A(_05287_),
    .B(_05320_),
    .Y(_17245_));
 BUFx12f_ASAP7_75t_R _19841_ (.A(_05313_),
    .Y(_05331_));
 NAND2x1_ASAP7_75t_R _19842_ (.A(_05302_),
    .B(_05331_),
    .Y(_17253_));
 NAND2x1_ASAP7_75t_R _19843_ (.A(_05314_),
    .B(_05318_),
    .Y(_17262_));
 AND2x2_ASAP7_75t_R _19844_ (.A(_05277_),
    .B(_05323_),
    .Y(_17267_));
 AND3x1_ASAP7_75t_R _19845_ (.A(_15315_),
    .B(_15362_),
    .C(_05258_),
    .Y(_05332_));
 AO21x2_ASAP7_75t_R _19846_ (.A1(_04605_),
    .A2(_05285_),
    .B(_05332_),
    .Y(_05333_));
 BUFx6f_ASAP7_75t_R _19847_ (.A(_05333_),
    .Y(_05334_));
 AND2x4_ASAP7_75t_R _19848_ (.A(_05283_),
    .B(_05334_),
    .Y(_17266_));
 AND3x1_ASAP7_75t_R _19849_ (.A(_15465_),
    .B(_15501_),
    .C(_05257_),
    .Y(_05335_));
 AO21x2_ASAP7_75t_R _19850_ (.A1(_04717_),
    .A2(_05285_),
    .B(_05335_),
    .Y(_05336_));
 BUFx6f_ASAP7_75t_R _19851_ (.A(_05336_),
    .Y(_05337_));
 AND2x2_ASAP7_75t_R _19852_ (.A(_05271_),
    .B(_05337_),
    .Y(_17265_));
 OA22x2_ASAP7_75t_R _19853_ (.A1(_00180_),
    .A2(_05244_),
    .B1(_05259_),
    .B2(_04791_),
    .Y(_17280_));
 AND3x1_ASAP7_75t_R _19854_ (.A(_13162_),
    .B(_13216_),
    .C(_05268_),
    .Y(_05338_));
 AO21x1_ASAP7_75t_R _19855_ (.A1(_04554_),
    .A2(_05267_),
    .B(_05338_),
    .Y(_05339_));
 BUFx6f_ASAP7_75t_R _19856_ (.A(_05339_),
    .Y(_05340_));
 BUFx12f_ASAP7_75t_R _19857_ (.A(_05340_),
    .Y(_05341_));
 NAND2x1_ASAP7_75t_R _19858_ (.A(_05274_),
    .B(_05341_),
    .Y(_17285_));
 BUFx12f_ASAP7_75t_R _19859_ (.A(_05320_),
    .Y(_05342_));
 NAND2x1_ASAP7_75t_R _19860_ (.A(_05302_),
    .B(_05342_),
    .Y(_17292_));
 NAND2x1_ASAP7_75t_R _19861_ (.A(_05306_),
    .B(_05318_),
    .Y(_17302_));
 AND2x2_ASAP7_75t_R _19862_ (.A(_05294_),
    .B(_05323_),
    .Y(_17307_));
 AND2x4_ASAP7_75t_R _19863_ (.A(_05277_),
    .B(_05334_),
    .Y(_17306_));
 AND2x2_ASAP7_75t_R _19864_ (.A(_05283_),
    .B(_05337_),
    .Y(_17305_));
 OA22x2_ASAP7_75t_R _19865_ (.A1(_00187_),
    .A2(_05244_),
    .B1(_05259_),
    .B2(_04959_),
    .Y(_17326_));
 AND2x6_ASAP7_75t_R _19866_ (.A(_04634_),
    .B(_04665_),
    .Y(_05343_));
 AND3x1_ASAP7_75t_R _19867_ (.A(_15398_),
    .B(_15429_),
    .C(_05289_),
    .Y(_05344_));
 AO21x2_ASAP7_75t_R _19868_ (.A1(_05343_),
    .A2(_05267_),
    .B(_05344_),
    .Y(_05345_));
 AND2x2_ASAP7_75t_R _19869_ (.A(_05273_),
    .B(_05345_),
    .Y(_17331_));
 AND2x4_ASAP7_75t_R _19870_ (.A(_05279_),
    .B(_05340_),
    .Y(_17330_));
 AND2x2_ASAP7_75t_R _19871_ (.A(_05287_),
    .B(_05330_),
    .Y(_17329_));
 BUFx12f_ASAP7_75t_R _19872_ (.A(_05326_),
    .Y(_05346_));
 NAND2x1_ASAP7_75t_R _19873_ (.A(_05302_),
    .B(_05346_),
    .Y(_17337_));
 NAND2x1_ASAP7_75t_R _19874_ (.A(_05327_),
    .B(_05318_),
    .Y(_17346_));
 AND2x2_ASAP7_75t_R _19875_ (.A(_05291_),
    .B(_05323_),
    .Y(_17351_));
 AND2x4_ASAP7_75t_R _19876_ (.A(_05294_),
    .B(_05334_),
    .Y(_17350_));
 AND2x2_ASAP7_75t_R _19877_ (.A(_05277_),
    .B(_05337_),
    .Y(_17349_));
 AND2x2_ASAP7_75t_R _19878_ (.A(_13837_),
    .B(_14552_),
    .Y(_05347_));
 AO21x2_ASAP7_75t_R _19879_ (.A1(_14272_),
    .A2(_13422_),
    .B(_05347_),
    .Y(_05348_));
 AND3x1_ASAP7_75t_R _19880_ (.A(_15234_),
    .B(_04962_),
    .C(_05348_),
    .Y(_05349_));
 BUFx6f_ASAP7_75t_R _19881_ (.A(_05349_),
    .Y(_05350_));
 AND2x6_ASAP7_75t_R _19882_ (.A(_05266_),
    .B(_05350_),
    .Y(_05351_));
 AND2x6_ASAP7_75t_R _19883_ (.A(_05265_),
    .B(_05351_),
    .Y(_17365_));
 AND3x4_ASAP7_75t_R _19884_ (.A(_15674_),
    .B(_15706_),
    .C(_05268_),
    .Y(_05352_));
 AO21x2_ASAP7_75t_R _19885_ (.A1(_04962_),
    .A2(_05267_),
    .B(_05352_),
    .Y(_05353_));
 AND3x4_ASAP7_75t_R _19886_ (.A(_13495_),
    .B(_13512_),
    .C(_13530_),
    .Y(_05354_));
 NOR2x1_ASAP7_75t_R _19887_ (.A(_15995_),
    .B(_05257_),
    .Y(_05355_));
 AO21x1_ASAP7_75t_R _19888_ (.A1(_05354_),
    .A2(_05257_),
    .B(_05355_),
    .Y(_05356_));
 BUFx6f_ASAP7_75t_R _19889_ (.A(_05356_),
    .Y(_05357_));
 AND2x2_ASAP7_75t_R _19890_ (.A(_05353_),
    .B(_05357_),
    .Y(_17370_));
 AND2x6_ASAP7_75t_R _19891_ (.A(_04756_),
    .B(_04787_),
    .Y(_05358_));
 AND3x1_ASAP7_75t_R _19892_ (.A(_15551_),
    .B(_15582_),
    .C(_05268_),
    .Y(_05359_));
 AO21x2_ASAP7_75t_R _19893_ (.A1(_05358_),
    .A2(_05267_),
    .B(_05359_),
    .Y(_05360_));
 BUFx12f_ASAP7_75t_R _19894_ (.A(_05360_),
    .Y(_05361_));
 AND2x4_ASAP7_75t_R _19895_ (.A(_05273_),
    .B(_05361_),
    .Y(_17369_));
 AND2x2_ASAP7_75t_R _19896_ (.A(_05279_),
    .B(_05345_),
    .Y(_17368_));
 NAND2x1_ASAP7_75t_R _19897_ (.A(_05288_),
    .B(_05341_),
    .Y(_17377_));
 AND3x1_ASAP7_75t_R _19898_ (.A(_16723_),
    .B(_16746_),
    .C(_05262_),
    .Y(_05362_));
 AO21x2_ASAP7_75t_R _19899_ (.A1(_13968_),
    .A2(_05258_),
    .B(_05362_),
    .Y(_05363_));
 BUFx6f_ASAP7_75t_R _19900_ (.A(_05363_),
    .Y(_05364_));
 BUFx12f_ASAP7_75t_R _19901_ (.A(_05364_),
    .Y(_05365_));
 NAND2x1_ASAP7_75t_R _19902_ (.A(_05342_),
    .B(_05365_),
    .Y(_17387_));
 AND2x2_ASAP7_75t_R _19903_ (.A(_14201_),
    .B(_05257_),
    .Y(_05366_));
 AO21x1_ASAP7_75t_R _19904_ (.A1(_04357_),
    .A2(_05285_),
    .B(_05366_),
    .Y(_05367_));
 BUFx6f_ASAP7_75t_R _19905_ (.A(_05367_),
    .Y(_05368_));
 AND2x2_ASAP7_75t_R _19906_ (.A(_05305_),
    .B(_05368_),
    .Y(_17392_));
 AND2x4_ASAP7_75t_R _19907_ (.A(_05297_),
    .B(_05323_),
    .Y(_17391_));
 AND2x2_ASAP7_75t_R _19908_ (.A(_05291_),
    .B(_05334_),
    .Y(_17390_));
 NAND2x1_ASAP7_75t_R _19909_ (.A(_05307_),
    .B(_05337_),
    .Y(_17402_));
 OAI22x1_ASAP7_75t_R _19910_ (.A1(_05237_),
    .A2(_00205_),
    .B1(_05256_),
    .B2(_15947_),
    .Y(_17422_));
 AND2x6_ASAP7_75t_R _19911_ (.A(_05351_),
    .B(_05357_),
    .Y(_17421_));
 BUFx12f_ASAP7_75t_R _19912_ (.A(_05353_),
    .Y(_05369_));
 AND2x2_ASAP7_75t_R _19913_ (.A(_05273_),
    .B(_05369_),
    .Y(_17425_));
 AND2x4_ASAP7_75t_R _19914_ (.A(_05279_),
    .B(_05360_),
    .Y(_17424_));
 AND2x2_ASAP7_75t_R _19915_ (.A(_05287_),
    .B(_05345_),
    .Y(_17423_));
 NAND2x1_ASAP7_75t_R _19916_ (.A(_05302_),
    .B(_05341_),
    .Y(_17433_));
 NAND2x1_ASAP7_75t_R _19917_ (.A(_05318_),
    .B(_05342_),
    .Y(_17443_));
 AND2x2_ASAP7_75t_R _19918_ (.A(_05305_),
    .B(_05323_),
    .Y(_17448_));
 AND2x4_ASAP7_75t_R _19919_ (.A(_05297_),
    .B(_05334_),
    .Y(_17447_));
 AND2x2_ASAP7_75t_R _19920_ (.A(_05291_),
    .B(_05337_),
    .Y(_17446_));
 OR2x2_ASAP7_75t_R _19921_ (.A(net1946),
    .B(_05285_),
    .Y(_05370_));
 OAI21x1_ASAP7_75t_R _19922_ (.A1(_04837_),
    .A2(_05258_),
    .B(_05370_),
    .Y(_05371_));
 BUFx12f_ASAP7_75t_R _19923_ (.A(_05371_),
    .Y(_05372_));
 NAND2x1_ASAP7_75t_R _19924_ (.A(_05307_),
    .B(_05372_),
    .Y(_17457_));
 BUFx6f_ASAP7_75t_R _19925_ (.A(_05244_),
    .Y(_05373_));
 INVx1_ASAP7_75t_R _19926_ (.A(_05348_),
    .Y(_05374_));
 OR4x1_ASAP7_75t_R _19927_ (.A(_05237_),
    .B(_00205_),
    .C(_14620_),
    .D(_05374_),
    .Y(_05375_));
 BUFx6f_ASAP7_75t_R _19928_ (.A(_05375_),
    .Y(_05376_));
 BUFx12f_ASAP7_75t_R _19929_ (.A(_05376_),
    .Y(_05377_));
 OAI21x1_ASAP7_75t_R _19930_ (.A1(_16083_),
    .A2(_05373_),
    .B(_05377_),
    .Y(_17467_));
 BUFx12f_ASAP7_75t_R _19931_ (.A(_05351_),
    .Y(_05378_));
 AND2x6_ASAP7_75t_R _19932_ (.A(_05273_),
    .B(_05378_),
    .Y(_17470_));
 AND2x4_ASAP7_75t_R _19933_ (.A(_05279_),
    .B(_05369_),
    .Y(_17469_));
 AND2x2_ASAP7_75t_R _19934_ (.A(_05287_),
    .B(_05360_),
    .Y(_17468_));
 BUFx12f_ASAP7_75t_R _19935_ (.A(_05345_),
    .Y(_05379_));
 NAND2x1_ASAP7_75t_R _19936_ (.A(_05301_),
    .B(_05379_),
    .Y(_17478_));
 NAND2x1_ASAP7_75t_R _19937_ (.A(_05318_),
    .B(_05346_),
    .Y(_17488_));
 AND2x2_ASAP7_75t_R _19938_ (.A(_05310_),
    .B(_05323_),
    .Y(_17493_));
 AND2x4_ASAP7_75t_R _19939_ (.A(_05305_),
    .B(_05334_),
    .Y(_17492_));
 AND2x2_ASAP7_75t_R _19940_ (.A(_05297_),
    .B(_05337_),
    .Y(_17491_));
 NAND2x1_ASAP7_75t_R _19941_ (.A(_05311_),
    .B(_05372_),
    .Y(_17502_));
 OAI21x1_ASAP7_75t_R _19942_ (.A1(_16195_),
    .A2(_05373_),
    .B(_05377_),
    .Y(_17512_));
 AND2x4_ASAP7_75t_R _19943_ (.A(_05279_),
    .B(_05378_),
    .Y(_17515_));
 AND2x4_ASAP7_75t_R _19944_ (.A(_05287_),
    .B(_05369_),
    .Y(_17514_));
 NAND2x1_ASAP7_75t_R _19945_ (.A(_05301_),
    .B(_05361_),
    .Y(_17523_));
 BUFx12f_ASAP7_75t_R _19946_ (.A(_05330_),
    .Y(_05380_));
 NAND2x1_ASAP7_75t_R _19947_ (.A(_05318_),
    .B(_05380_),
    .Y(_17533_));
 AND2x2_ASAP7_75t_R _19948_ (.A(_05313_),
    .B(_05323_),
    .Y(_17538_));
 AND2x4_ASAP7_75t_R _19949_ (.A(_05310_),
    .B(_05334_),
    .Y(_17537_));
 AND2x2_ASAP7_75t_R _19950_ (.A(_05305_),
    .B(_05337_),
    .Y(_17536_));
 NAND2x1_ASAP7_75t_R _19951_ (.A(_05314_),
    .B(_05372_),
    .Y(_17547_));
 OAI21x1_ASAP7_75t_R _19952_ (.A1(_16329_),
    .A2(_05373_),
    .B(_05377_),
    .Y(_17558_));
 AND2x2_ASAP7_75t_R _19953_ (.A(_05287_),
    .B(_05378_),
    .Y(_17560_));
 NAND2x1_ASAP7_75t_R _19954_ (.A(_05301_),
    .B(_05369_),
    .Y(_17567_));
 NAND2x1_ASAP7_75t_R _19955_ (.A(_05317_),
    .B(_05341_),
    .Y(_17578_));
 AND2x2_ASAP7_75t_R _19956_ (.A(_05320_),
    .B(_05323_),
    .Y(_17583_));
 AND2x4_ASAP7_75t_R _19957_ (.A(_05313_),
    .B(_05334_),
    .Y(_17582_));
 AND2x2_ASAP7_75t_R _19958_ (.A(_05310_),
    .B(_05337_),
    .Y(_17581_));
 NAND2x1_ASAP7_75t_R _19959_ (.A(_05306_),
    .B(_05372_),
    .Y(_17592_));
 OAI21x1_ASAP7_75t_R _19960_ (.A1(_00115_),
    .A2(_05373_),
    .B(_05377_),
    .Y(_17603_));
 AND2x6_ASAP7_75t_R _19961_ (.A(_05301_),
    .B(_05378_),
    .Y(_17610_));
 AND3x1_ASAP7_75t_R _19962_ (.A(_16613_),
    .B(_16636_),
    .C(_05262_),
    .Y(_05381_));
 AO21x2_ASAP7_75t_R _19963_ (.A1(_13908_),
    .A2(_05258_),
    .B(_05381_),
    .Y(_05382_));
 BUFx6f_ASAP7_75t_R _19964_ (.A(_05382_),
    .Y(_05383_));
 AND2x4_ASAP7_75t_R _19965_ (.A(_05353_),
    .B(_05383_),
    .Y(_17609_));
 AND2x2_ASAP7_75t_R _19966_ (.A(_05360_),
    .B(_05364_),
    .Y(_17608_));
 NAND2x1_ASAP7_75t_R _19967_ (.A(_05317_),
    .B(_05379_),
    .Y(_17620_));
 AND2x2_ASAP7_75t_R _19968_ (.A(_05322_),
    .B(_05326_),
    .Y(_17625_));
 AND2x4_ASAP7_75t_R _19969_ (.A(_05320_),
    .B(_05334_),
    .Y(_17624_));
 AND2x2_ASAP7_75t_R _19970_ (.A(_05313_),
    .B(_05337_),
    .Y(_17623_));
 NAND2x1_ASAP7_75t_R _19971_ (.A(_05327_),
    .B(_05372_),
    .Y(_17634_));
 OAI21x1_ASAP7_75t_R _19972_ (.A1(_16591_),
    .A2(_05373_),
    .B(_05377_),
    .Y(_17645_));
 AND2x4_ASAP7_75t_R _19973_ (.A(_05378_),
    .B(_05383_),
    .Y(_17652_));
 AND2x4_ASAP7_75t_R _19974_ (.A(_05353_),
    .B(_05364_),
    .Y(_17651_));
 NAND2x1_ASAP7_75t_R _19975_ (.A(_05317_),
    .B(_05361_),
    .Y(_17661_));
 AND2x2_ASAP7_75t_R _19976_ (.A(_05322_),
    .B(_05330_),
    .Y(_17666_));
 AND2x4_ASAP7_75t_R _19977_ (.A(_05326_),
    .B(_05334_),
    .Y(_17665_));
 AND2x2_ASAP7_75t_R _19978_ (.A(_05320_),
    .B(_05337_),
    .Y(_17664_));
 NAND2x1_ASAP7_75t_R _19979_ (.A(_05331_),
    .B(_05372_),
    .Y(_17675_));
 OAI21x1_ASAP7_75t_R _19980_ (.A1(_16701_),
    .A2(_05373_),
    .B(_05377_),
    .Y(_17686_));
 AND2x2_ASAP7_75t_R _19981_ (.A(_05351_),
    .B(_05364_),
    .Y(_17692_));
 NAND2x1_ASAP7_75t_R _19982_ (.A(_05317_),
    .B(_05369_),
    .Y(_17702_));
 AND2x2_ASAP7_75t_R _19983_ (.A(_05322_),
    .B(_05340_),
    .Y(_17707_));
 AND2x4_ASAP7_75t_R _19984_ (.A(_05330_),
    .B(_05333_),
    .Y(_17706_));
 AND2x2_ASAP7_75t_R _19985_ (.A(_05326_),
    .B(_05336_),
    .Y(_17705_));
 NAND2x1_ASAP7_75t_R _19986_ (.A(_05342_),
    .B(_05372_),
    .Y(_17716_));
 OAI21x1_ASAP7_75t_R _19987_ (.A1(_16823_),
    .A2(_05373_),
    .B(_05377_),
    .Y(_17727_));
 AND2x6_ASAP7_75t_R _19988_ (.A(_05317_),
    .B(_05378_),
    .Y(_17742_));
 AND2x2_ASAP7_75t_R _19989_ (.A(_14089_),
    .B(_05257_),
    .Y(_05384_));
 AO21x1_ASAP7_75t_R _19990_ (.A1(_16983_),
    .A2(_05285_),
    .B(_05384_),
    .Y(_05385_));
 BUFx6f_ASAP7_75t_R _19991_ (.A(_05385_),
    .Y(_05386_));
 AND2x4_ASAP7_75t_R _19992_ (.A(_05353_),
    .B(_05386_),
    .Y(_17741_));
 AND2x2_ASAP7_75t_R _19993_ (.A(_05360_),
    .B(_05368_),
    .Y(_17740_));
 AND2x2_ASAP7_75t_R _19994_ (.A(_05322_),
    .B(_05345_),
    .Y(_17745_));
 AND2x4_ASAP7_75t_R _19995_ (.A(_05333_),
    .B(_05340_),
    .Y(_17744_));
 AND2x2_ASAP7_75t_R _19996_ (.A(_05330_),
    .B(_05336_),
    .Y(_17743_));
 NAND2x1_ASAP7_75t_R _19997_ (.A(_05346_),
    .B(_05372_),
    .Y(_17756_));
 OAI21x1_ASAP7_75t_R _19998_ (.A1(_16935_),
    .A2(_05373_),
    .B(_05377_),
    .Y(_17767_));
 AND2x4_ASAP7_75t_R _19999_ (.A(_05351_),
    .B(_05386_),
    .Y(_17776_));
 AND2x4_ASAP7_75t_R _20000_ (.A(_05353_),
    .B(_05368_),
    .Y(_17775_));
 AND2x2_ASAP7_75t_R _20001_ (.A(_05322_),
    .B(_05360_),
    .Y(_17779_));
 AND2x4_ASAP7_75t_R _20002_ (.A(_05333_),
    .B(_05345_),
    .Y(_17778_));
 AND2x2_ASAP7_75t_R _20003_ (.A(_05336_),
    .B(_05340_),
    .Y(_17777_));
 NAND2x1_ASAP7_75t_R _20004_ (.A(_05380_),
    .B(_05372_),
    .Y(_17792_));
 OAI21x1_ASAP7_75t_R _20005_ (.A1(_04310_),
    .A2(_05373_),
    .B(_05377_),
    .Y(_17803_));
 AND2x2_ASAP7_75t_R _20006_ (.A(_05351_),
    .B(_05368_),
    .Y(_17812_));
 AND2x2_ASAP7_75t_R _20007_ (.A(_05322_),
    .B(_05369_),
    .Y(_17815_));
 AND2x4_ASAP7_75t_R _20008_ (.A(_05333_),
    .B(_05360_),
    .Y(_17814_));
 AND2x2_ASAP7_75t_R _20009_ (.A(_05336_),
    .B(_05345_),
    .Y(_17813_));
 NAND2x1_ASAP7_75t_R _20010_ (.A(_05341_),
    .B(_05372_),
    .Y(_17827_));
 OAI21x1_ASAP7_75t_R _20011_ (.A1(_04422_),
    .A2(_05373_),
    .B(_05377_),
    .Y(_17838_));
 AND2x6_ASAP7_75t_R _20012_ (.A(_05322_),
    .B(_05378_),
    .Y(_17849_));
 AND2x4_ASAP7_75t_R _20013_ (.A(_05333_),
    .B(_05369_),
    .Y(_17848_));
 AND2x2_ASAP7_75t_R _20014_ (.A(_05336_),
    .B(_05360_),
    .Y(_17847_));
 NAND2x1_ASAP7_75t_R _20015_ (.A(_05379_),
    .B(_05371_),
    .Y(_17859_));
 OAI21x1_ASAP7_75t_R _20016_ (.A1(_04558_),
    .A2(_05256_),
    .B(_05376_),
    .Y(_17870_));
 AND2x4_ASAP7_75t_R _20017_ (.A(_05333_),
    .B(_05378_),
    .Y(_17880_));
 AND2x2_ASAP7_75t_R _20018_ (.A(_05336_),
    .B(_05353_),
    .Y(_17879_));
 NAND2x1_ASAP7_75t_R _20019_ (.A(_05361_),
    .B(_05371_),
    .Y(_17889_));
 OAI21x1_ASAP7_75t_R _20020_ (.A1(_04670_),
    .A2(_05256_),
    .B(_05376_),
    .Y(_17900_));
 AND2x4_ASAP7_75t_R _20021_ (.A(_05336_),
    .B(_05378_),
    .Y(_17907_));
 NAND2x1_ASAP7_75t_R _20022_ (.A(_05369_),
    .B(_05371_),
    .Y(_17917_));
 OAI21x1_ASAP7_75t_R _20023_ (.A1(_04791_),
    .A2(_05256_),
    .B(_05376_),
    .Y(_17928_));
 AND2x6_ASAP7_75t_R _20024_ (.A(_05351_),
    .B(_05371_),
    .Y(_17942_));
 NAND2x1_ASAP7_75t_R _20025_ (.A(_15759_),
    .B(_05258_),
    .Y(_05387_));
 OA21x2_ASAP7_75t_R _20026_ (.A1(_04963_),
    .A2(_05258_),
    .B(_05387_),
    .Y(_05388_));
 BUFx12f_ASAP7_75t_R _20027_ (.A(_05388_),
    .Y(_05389_));
 AND2x4_ASAP7_75t_R _20028_ (.A(_05353_),
    .B(_05389_),
    .Y(_17941_));
 AO21x2_ASAP7_75t_R _20029_ (.A1(_13262_),
    .A2(_14272_),
    .B(_05347_),
    .Y(_05390_));
 AND3x4_ASAP7_75t_R _20030_ (.A(_15234_),
    .B(_04963_),
    .C(_05390_),
    .Y(_05391_));
 NAND2x2_ASAP7_75t_R _20031_ (.A(_05285_),
    .B(_05391_),
    .Y(_05392_));
 BUFx6f_ASAP7_75t_R _20032_ (.A(_05392_),
    .Y(_05393_));
 NOR2x1_ASAP7_75t_R _20033_ (.A(_05361_),
    .B(_05393_),
    .Y(_17940_));
 OAI21x1_ASAP7_75t_R _20034_ (.A1(_04959_),
    .A2(_05256_),
    .B(_05376_),
    .Y(_17953_));
 AND2x6_ASAP7_75t_R _20035_ (.A(_05351_),
    .B(_05389_),
    .Y(_17967_));
 NOR2x1_ASAP7_75t_R _20036_ (.A(_05369_),
    .B(_05393_),
    .Y(_17966_));
 OAI21x1_ASAP7_75t_R _20037_ (.A1(_01728_),
    .A2(_05256_),
    .B(_05376_),
    .Y(_17979_));
 NOR2x1_ASAP7_75t_R _20038_ (.A(_05378_),
    .B(_05393_),
    .Y(_17989_));
 INVx5_ASAP7_75t_R _20039_ (.A(net1962),
    .Y(_17736_));
 AO21x1_ASAP7_75t_R _20040_ (.A1(_13441_),
    .A2(_13423_),
    .B(_13424_),
    .Y(_05394_));
 INVx1_ASAP7_75t_R _20041_ (.A(_05394_),
    .Y(_05395_));
 AND3x1_ASAP7_75t_R _20042_ (.A(_13235_),
    .B(_05191_),
    .C(_05395_),
    .Y(_05396_));
 INVx1_ASAP7_75t_R _20043_ (.A(_01764_),
    .Y(_05397_));
 AO31x2_ASAP7_75t_R _20044_ (.A1(_04986_),
    .A2(_14115_),
    .A3(_05396_),
    .B(_05397_),
    .Y(_05398_));
 OR2x2_ASAP7_75t_R _20045_ (.A(_13233_),
    .B(_01539_),
    .Y(_05399_));
 BUFx6f_ASAP7_75t_R _20046_ (.A(_05399_),
    .Y(_05400_));
 AND2x2_ASAP7_75t_R _20047_ (.A(_05190_),
    .B(_05400_),
    .Y(_05401_));
 AND2x6_ASAP7_75t_R _20048_ (.A(_05172_),
    .B(_01762_),
    .Y(_05402_));
 INVx2_ASAP7_75t_R _20049_ (.A(_01398_),
    .Y(_05403_));
 BUFx6f_ASAP7_75t_R _20050_ (.A(_01760_),
    .Y(_05404_));
 OR4x1_ASAP7_75t_R _20051_ (.A(net81),
    .B(_05403_),
    .C(_05404_),
    .D(_05173_),
    .Y(_05405_));
 AND3x4_ASAP7_75t_R _20052_ (.A(_05153_),
    .B(_01763_),
    .C(_05189_),
    .Y(_05406_));
 AND3x4_ASAP7_75t_R _20053_ (.A(_01758_),
    .B(_01759_),
    .C(_02200_),
    .Y(_05407_));
 INVx1_ASAP7_75t_R _20054_ (.A(_05407_),
    .Y(_05408_));
 AO21x2_ASAP7_75t_R _20055_ (.A1(_14109_),
    .A2(_05164_),
    .B(_05408_),
    .Y(_05409_));
 NAND3x1_ASAP7_75t_R _20056_ (.A(_14098_),
    .B(_14101_),
    .C(_14102_),
    .Y(_05410_));
 NAND2x1_ASAP7_75t_R _20057_ (.A(_01391_),
    .B(_05400_),
    .Y(_05411_));
 OR5x2_ASAP7_75t_R _20058_ (.A(_13233_),
    .B(_14119_),
    .C(_14275_),
    .D(_05410_),
    .E(_05411_),
    .Y(_05412_));
 NAND2x1_ASAP7_75t_R _20059_ (.A(_18080_),
    .B(_02062_),
    .Y(_05413_));
 OR3x1_ASAP7_75t_R _20060_ (.A(_18080_),
    .B(_02057_),
    .C(_02062_),
    .Y(_05414_));
 OA21x2_ASAP7_75t_R _20061_ (.A1(_02059_),
    .A2(_05413_),
    .B(_05414_),
    .Y(_05415_));
 AND2x4_ASAP7_75t_R _20062_ (.A(_00758_),
    .B(_05415_),
    .Y(_05416_));
 OR4x1_ASAP7_75t_R _20063_ (.A(_14191_),
    .B(_05407_),
    .C(_05412_),
    .D(_05416_),
    .Y(_05417_));
 INVx1_ASAP7_75t_R _20064_ (.A(net156),
    .Y(_05418_));
 NOR2x1_ASAP7_75t_R _20065_ (.A(_05418_),
    .B(_01919_),
    .Y(_05419_));
 INVx1_ASAP7_75t_R _20066_ (.A(_01911_),
    .Y(_05420_));
 INVx2_ASAP7_75t_R _20067_ (.A(_01912_),
    .Y(_05421_));
 AO22x1_ASAP7_75t_R _20068_ (.A1(net161),
    .A2(_05420_),
    .B1(_05421_),
    .B2(net160),
    .Y(_05422_));
 INVx1_ASAP7_75t_R _20069_ (.A(net163),
    .Y(_05423_));
 INVx2_ASAP7_75t_R _20070_ (.A(net162),
    .Y(_05424_));
 OAI22x1_ASAP7_75t_R _20071_ (.A1(_05423_),
    .A2(_01909_),
    .B1(_01910_),
    .B2(_05424_),
    .Y(_05425_));
 INVx1_ASAP7_75t_R _20072_ (.A(net159),
    .Y(_05426_));
 INVx2_ASAP7_75t_R _20073_ (.A(net158),
    .Y(_05427_));
 OAI22x1_ASAP7_75t_R _20074_ (.A1(_05426_),
    .A2(_01913_),
    .B1(_01914_),
    .B2(_05427_),
    .Y(_05428_));
 INVx1_ASAP7_75t_R _20075_ (.A(net157),
    .Y(_05429_));
 INVx1_ASAP7_75t_R _20076_ (.A(net151),
    .Y(_05430_));
 OAI22x1_ASAP7_75t_R _20077_ (.A1(_05429_),
    .A2(_01915_),
    .B1(_01924_),
    .B2(_05430_),
    .Y(_05431_));
 OR4x1_ASAP7_75t_R _20078_ (.A(_05422_),
    .B(_05425_),
    .C(_05428_),
    .D(_05431_),
    .Y(_05432_));
 INVx1_ASAP7_75t_R _20079_ (.A(_01920_),
    .Y(_05433_));
 INVx1_ASAP7_75t_R _20080_ (.A(_01921_),
    .Y(_05434_));
 AO22x2_ASAP7_75t_R _20081_ (.A1(net155),
    .A2(_05433_),
    .B1(_05434_),
    .B2(net154),
    .Y(_05435_));
 INVx1_ASAP7_75t_R _20082_ (.A(_01922_),
    .Y(_05436_));
 INVx1_ASAP7_75t_R _20083_ (.A(_01923_),
    .Y(_05437_));
 AO22x2_ASAP7_75t_R _20084_ (.A1(net153),
    .A2(_05436_),
    .B1(_05437_),
    .B2(net152),
    .Y(_05438_));
 INVx1_ASAP7_75t_R _20085_ (.A(_01907_),
    .Y(_05439_));
 INVx1_ASAP7_75t_R _20086_ (.A(_01908_),
    .Y(_05440_));
 AO22x2_ASAP7_75t_R _20087_ (.A1(net165),
    .A2(_05439_),
    .B1(_05440_),
    .B2(net164),
    .Y(_05441_));
 OR3x2_ASAP7_75t_R _20088_ (.A(_05435_),
    .B(_05438_),
    .C(_05441_),
    .Y(_05442_));
 INVx1_ASAP7_75t_R _20089_ (.A(net167),
    .Y(_05443_));
 INVx2_ASAP7_75t_R _20090_ (.A(net150),
    .Y(_05444_));
 OAI22x1_ASAP7_75t_R _20091_ (.A1(_05443_),
    .A2(_01916_),
    .B1(_01918_),
    .B2(_05444_),
    .Y(_05445_));
 INVx1_ASAP7_75t_R _20092_ (.A(_01917_),
    .Y(_05446_));
 AO21x1_ASAP7_75t_R _20093_ (.A1(net168),
    .A2(_05446_),
    .B(net166),
    .Y(_05447_));
 OR2x6_ASAP7_75t_R _20094_ (.A(_05445_),
    .B(_05447_),
    .Y(_05448_));
 OR4x1_ASAP7_75t_R _20095_ (.A(_05419_),
    .B(_05432_),
    .C(_05442_),
    .D(_05448_),
    .Y(_05449_));
 INVx1_ASAP7_75t_R _20096_ (.A(_00759_),
    .Y(_05450_));
 OA211x2_ASAP7_75t_R _20097_ (.A1(net166),
    .A2(_05450_),
    .B(_00334_),
    .C(_00758_),
    .Y(_05451_));
 NOR2x1_ASAP7_75t_R _20098_ (.A(_01762_),
    .B(_05154_),
    .Y(_05452_));
 AND3x4_ASAP7_75t_R _20099_ (.A(_05189_),
    .B(_05451_),
    .C(_05452_),
    .Y(_05453_));
 AO32x1_ASAP7_75t_R _20100_ (.A1(_05406_),
    .A2(_05409_),
    .A3(_05417_),
    .B1(_05449_),
    .B2(_05453_),
    .Y(_05454_));
 AO21x1_ASAP7_75t_R _20101_ (.A1(_05402_),
    .A2(_05405_),
    .B(_05454_),
    .Y(_05455_));
 AOI21x1_ASAP7_75t_R _20102_ (.A1(_05398_),
    .A2(_05401_),
    .B(_05455_),
    .Y(_05456_));
 BUFx12f_ASAP7_75t_R _20103_ (.A(_05456_),
    .Y(_05457_));
 BUFx12f_ASAP7_75t_R _20104_ (.A(_05457_),
    .Y(_05458_));
 BUFx12f_ASAP7_75t_R _20105_ (.A(_05458_),
    .Y(_05459_));
 BUFx12f_ASAP7_75t_R _20106_ (.A(_00260_),
    .Y(_05460_));
 BUFx6f_ASAP7_75t_R _20107_ (.A(_05460_),
    .Y(_05461_));
 AOI21x1_ASAP7_75t_R _20108_ (.A1(_01724_),
    .A2(_05459_),
    .B(_05461_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ));
 AO21x2_ASAP7_75t_R _20109_ (.A1(_05398_),
    .A2(_05401_),
    .B(_05455_),
    .Y(_05462_));
 BUFx12f_ASAP7_75t_R _20110_ (.A(_05462_),
    .Y(_05463_));
 BUFx12f_ASAP7_75t_R _20111_ (.A(_05463_),
    .Y(_05464_));
 BUFx12f_ASAP7_75t_R _20112_ (.A(_05464_),
    .Y(_05465_));
 BUFx12f_ASAP7_75t_R _20113_ (.A(_05465_),
    .Y(_05466_));
 BUFx6f_ASAP7_75t_R _20114_ (.A(_05466_),
    .Y(_05467_));
 INVx1_ASAP7_75t_R _20115_ (.A(_14106_),
    .Y(_05468_));
 AND3x1_ASAP7_75t_R _20116_ (.A(_05468_),
    .B(_05406_),
    .C(_05407_),
    .Y(_05469_));
 NAND2x2_ASAP7_75t_R _20117_ (.A(_05165_),
    .B(_05469_),
    .Y(_05470_));
 BUFx6f_ASAP7_75t_R _20118_ (.A(_05470_),
    .Y(_05471_));
 AND2x2_ASAP7_75t_R _20119_ (.A(_05404_),
    .B(_05173_),
    .Y(_05472_));
 AND2x4_ASAP7_75t_R _20120_ (.A(_05171_),
    .B(_05402_),
    .Y(_05473_));
 AOI21x1_ASAP7_75t_R _20121_ (.A1(_05155_),
    .A2(_05472_),
    .B(_05473_),
    .Y(_05474_));
 AO21x2_ASAP7_75t_R _20122_ (.A1(_05167_),
    .A2(_05407_),
    .B(_05174_),
    .Y(_05475_));
 AND3x4_ASAP7_75t_R _20123_ (.A(_05471_),
    .B(_05474_),
    .C(_05475_),
    .Y(_05476_));
 BUFx6f_ASAP7_75t_R _20124_ (.A(_05158_),
    .Y(_05477_));
 NAND2x2_ASAP7_75t_R _20125_ (.A(_05449_),
    .B(_05453_),
    .Y(_05478_));
 NAND2x1_ASAP7_75t_R _20126_ (.A(net154),
    .B(_05434_),
    .Y(_05479_));
 NAND2x1_ASAP7_75t_R _20127_ (.A(net152),
    .B(_05437_),
    .Y(_05480_));
 NAND2x1_ASAP7_75t_R _20128_ (.A(net164),
    .B(_05440_),
    .Y(_05481_));
 INVx1_ASAP7_75t_R _20129_ (.A(_01909_),
    .Y(_05482_));
 INVx1_ASAP7_75t_R _20130_ (.A(net160),
    .Y(_05483_));
 INVx1_ASAP7_75t_R _20131_ (.A(_01913_),
    .Y(_05484_));
 INVx1_ASAP7_75t_R _20132_ (.A(_01915_),
    .Y(_05485_));
 OA211x2_ASAP7_75t_R _20133_ (.A1(_05427_),
    .A2(_01914_),
    .B(_05485_),
    .C(net157),
    .Y(_05486_));
 AO21x1_ASAP7_75t_R _20134_ (.A1(net159),
    .A2(_05484_),
    .B(_05486_),
    .Y(_05487_));
 OA21x2_ASAP7_75t_R _20135_ (.A1(_05483_),
    .A2(_01912_),
    .B(_05487_),
    .Y(_05488_));
 AO21x1_ASAP7_75t_R _20136_ (.A1(net161),
    .A2(_05420_),
    .B(_05488_),
    .Y(_05489_));
 OA21x2_ASAP7_75t_R _20137_ (.A1(_05424_),
    .A2(_01910_),
    .B(_05489_),
    .Y(_05490_));
 AO21x1_ASAP7_75t_R _20138_ (.A1(net163),
    .A2(_05482_),
    .B(_05490_),
    .Y(_05491_));
 AO22x1_ASAP7_75t_R _20139_ (.A1(net165),
    .A2(_05439_),
    .B1(_05481_),
    .B2(_05491_),
    .Y(_05492_));
 AO22x1_ASAP7_75t_R _20140_ (.A1(net153),
    .A2(_05436_),
    .B1(_05480_),
    .B2(_05492_),
    .Y(_05493_));
 AOI22x1_ASAP7_75t_R _20141_ (.A1(net155),
    .A2(_05433_),
    .B1(_05479_),
    .B2(_05493_),
    .Y(_05494_));
 NAND2x1_ASAP7_75t_R _20142_ (.A(net166),
    .B(_00334_),
    .Y(_05495_));
 OR3x2_ASAP7_75t_R _20143_ (.A(_05419_),
    .B(_05432_),
    .C(_05442_),
    .Y(_05496_));
 OA211x2_ASAP7_75t_R _20144_ (.A1(_05419_),
    .A2(_05494_),
    .B(_05495_),
    .C(_05496_),
    .Y(_05497_));
 OR2x6_ASAP7_75t_R _20145_ (.A(_05478_),
    .B(_05497_),
    .Y(_05498_));
 BUFx6f_ASAP7_75t_R _20146_ (.A(_05471_),
    .Y(_05499_));
 BUFx6f_ASAP7_75t_R _20147_ (.A(_05499_),
    .Y(_05500_));
 OR3x2_ASAP7_75t_R _20148_ (.A(_05174_),
    .B(_05167_),
    .C(_05408_),
    .Y(_05501_));
 BUFx6f_ASAP7_75t_R _20149_ (.A(_05501_),
    .Y(_05502_));
 BUFx6f_ASAP7_75t_R _20150_ (.A(_05502_),
    .Y(_05503_));
 BUFx6f_ASAP7_75t_R _20151_ (.A(_05503_),
    .Y(_05504_));
 OA22x2_ASAP7_75t_R _20152_ (.A1(_02032_),
    .A2(_05500_),
    .B1(_05504_),
    .B2(_01934_),
    .Y(_05505_));
 OA211x2_ASAP7_75t_R _20153_ (.A1(_05477_),
    .A2(_05219_),
    .B(_05498_),
    .C(_05505_),
    .Y(_05506_));
 OR3x2_ASAP7_75t_R _20154_ (.A(_05458_),
    .B(_05476_),
    .C(_05506_),
    .Y(_05507_));
 OA21x2_ASAP7_75t_R _20155_ (.A1(_01703_),
    .A2(_05467_),
    .B(_05507_),
    .Y(_05508_));
 INVx1_ASAP7_75t_R _20156_ (.A(_05508_),
    .Y(_18716_));
 OR2x6_ASAP7_75t_R _20157_ (.A(_05174_),
    .B(_05407_),
    .Y(_05509_));
 OA222x2_ASAP7_75t_R _20158_ (.A1(_05158_),
    .A2(_05214_),
    .B1(_05470_),
    .B2(_01399_),
    .C1(_04991_),
    .C2(_05509_),
    .Y(_05510_));
 INVx1_ASAP7_75t_R _20159_ (.A(_05441_),
    .Y(_05511_));
 AOI22x1_ASAP7_75t_R _20160_ (.A1(net161),
    .A2(_05420_),
    .B1(_05421_),
    .B2(net160),
    .Y(_05512_));
 AO21x1_ASAP7_75t_R _20161_ (.A1(_05512_),
    .A2(_05428_),
    .B(_05425_),
    .Y(_05513_));
 AOI21x1_ASAP7_75t_R _20162_ (.A1(_05511_),
    .A2(_05513_),
    .B(_05438_),
    .Y(_05514_));
 AO21x1_ASAP7_75t_R _20163_ (.A1(net166),
    .A2(_00334_),
    .B(_05419_),
    .Y(_05515_));
 INVx1_ASAP7_75t_R _20164_ (.A(_05515_),
    .Y(_05516_));
 OA211x2_ASAP7_75t_R _20165_ (.A1(_05435_),
    .A2(_05514_),
    .B(_05516_),
    .C(_05496_),
    .Y(_05517_));
 OR2x2_ASAP7_75t_R _20166_ (.A(_05478_),
    .B(_05517_),
    .Y(_05518_));
 OA21x2_ASAP7_75t_R _20167_ (.A1(_01931_),
    .A2(_05502_),
    .B(_05518_),
    .Y(_05519_));
 AO21x2_ASAP7_75t_R _20168_ (.A1(_05510_),
    .A2(_05519_),
    .B(_05456_),
    .Y(_05520_));
 OA21x2_ASAP7_75t_R _20169_ (.A1(_01700_),
    .A2(_05463_),
    .B(_05520_),
    .Y(_05521_));
 INVx1_ASAP7_75t_R _20170_ (.A(_05521_),
    .Y(_18719_));
 BUFx12f_ASAP7_75t_R _20171_ (.A(_00750_),
    .Y(_05522_));
 INVx3_ASAP7_75t_R _20172_ (.A(_05522_),
    .Y(_05523_));
 BUFx6f_ASAP7_75t_R _20173_ (.A(_05523_),
    .Y(_05524_));
 BUFx6f_ASAP7_75t_R _20174_ (.A(_05524_),
    .Y(_05525_));
 BUFx6f_ASAP7_75t_R _20175_ (.A(_05525_),
    .Y(_05526_));
 BUFx6f_ASAP7_75t_R _20176_ (.A(_00263_),
    .Y(_05527_));
 AND2x2_ASAP7_75t_R _20177_ (.A(_05527_),
    .B(net124),
    .Y(_05528_));
 NOR2x1_ASAP7_75t_R _20178_ (.A(_05527_),
    .B(_01656_),
    .Y(_05529_));
 INVx1_ASAP7_75t_R _20179_ (.A(_01657_),
    .Y(_05530_));
 AOI22x1_ASAP7_75t_R _20180_ (.A1(net125),
    .A2(_05528_),
    .B1(_05529_),
    .B2(_05530_),
    .Y(_05531_));
 INVx3_ASAP7_75t_R _20181_ (.A(_05527_),
    .Y(_05532_));
 INVx2_ASAP7_75t_R _20182_ (.A(net115),
    .Y(_05533_));
 AND2x2_ASAP7_75t_R _20183_ (.A(_05527_),
    .B(_05533_),
    .Y(_05534_));
 AO21x2_ASAP7_75t_R _20184_ (.A1(_05532_),
    .A2(_01693_),
    .B(_05534_),
    .Y(_05535_));
 AND2x6_ASAP7_75t_R _20185_ (.A(_05531_),
    .B(_05535_),
    .Y(_05536_));
 BUFx6f_ASAP7_75t_R _20186_ (.A(_05532_),
    .Y(_05537_));
 OA211x2_ASAP7_75t_R _20187_ (.A1(_01653_),
    .A2(_01664_),
    .B(_01693_),
    .C(_05537_),
    .Y(_05538_));
 BUFx6f_ASAP7_75t_R _20188_ (.A(_05527_),
    .Y(_05539_));
 AND3x1_ASAP7_75t_R _20189_ (.A(_05539_),
    .B(net117),
    .C(net128),
    .Y(_05540_));
 INVx1_ASAP7_75t_R _20190_ (.A(_05540_),
    .Y(_05541_));
 BUFx6f_ASAP7_75t_R _20191_ (.A(_05522_),
    .Y(_05542_));
 BUFx6f_ASAP7_75t_R _20192_ (.A(_05542_),
    .Y(_05543_));
 BUFx6f_ASAP7_75t_R _20193_ (.A(_05543_),
    .Y(_05544_));
 OA211x2_ASAP7_75t_R _20194_ (.A1(_05534_),
    .A2(_05538_),
    .B(_05541_),
    .C(_05544_),
    .Y(_05545_));
 AOI21x1_ASAP7_75t_R _20195_ (.A1(_05526_),
    .A2(_05536_),
    .B(_05545_),
    .Y(_18551_));
 INVx1_ASAP7_75t_R _20196_ (.A(_18551_),
    .Y(_17999_));
 INVx1_ASAP7_75t_R _20197_ (.A(net170),
    .Y(_05546_));
 NOR2x2_ASAP7_75t_R _20198_ (.A(_05496_),
    .B(_05448_),
    .Y(_05547_));
 INVx2_ASAP7_75t_R _20199_ (.A(net81),
    .Y(_05548_));
 AND2x2_ASAP7_75t_R _20200_ (.A(_05548_),
    .B(_02190_),
    .Y(_05549_));
 AO21x2_ASAP7_75t_R _20201_ (.A1(_05547_),
    .A2(_05549_),
    .B(_01797_),
    .Y(net171));
 NAND2x1_ASAP7_75t_R _20202_ (.A(_05546_),
    .B(net171),
    .Y(_00006_));
 INVx1_ASAP7_75t_R _20203_ (.A(_02329_),
    .Y(_18718_));
 INVx2_ASAP7_75t_R _20204_ (.A(_17997_),
    .Y(\cs_registers_i.pc_if_i[2] ));
 BUFx6f_ASAP7_75t_R _20205_ (.A(_05265_),
    .Y(_05550_));
 NAND2x1_ASAP7_75t_R _20206_ (.A(_05550_),
    .B(_05284_),
    .Y(_17000_));
 BUFx6f_ASAP7_75t_R _20207_ (.A(_05357_),
    .Y(_05551_));
 NAND2x1_ASAP7_75t_R _20208_ (.A(_05284_),
    .B(_05551_),
    .Y(_17003_));
 NAND2x1_ASAP7_75t_R _20209_ (.A(_05298_),
    .B(_05551_),
    .Y(_17012_));
 NAND2x1_ASAP7_75t_R _20210_ (.A(_05307_),
    .B(_05551_),
    .Y(_17018_));
 NAND2x1_ASAP7_75t_R _20211_ (.A(_05311_),
    .B(_05551_),
    .Y(_17034_));
 NAND2x1_ASAP7_75t_R _20212_ (.A(_05284_),
    .B(_05288_),
    .Y(_17039_));
 NAND2x1_ASAP7_75t_R _20213_ (.A(_05314_),
    .B(_05551_),
    .Y(_17046_));
 NAND2x1_ASAP7_75t_R _20214_ (.A(_05306_),
    .B(_05551_),
    .Y(_17064_));
 NAND2x1_ASAP7_75t_R _20215_ (.A(_05271_),
    .B(_05365_),
    .Y(_17076_));
 NAND2x1_ASAP7_75t_R _20216_ (.A(_05327_),
    .B(_05551_),
    .Y(_17092_));
 NAND2x1_ASAP7_75t_R _20217_ (.A(_05284_),
    .B(_05365_),
    .Y(_17104_));
 NAND2x1_ASAP7_75t_R _20218_ (.A(_05331_),
    .B(_05551_),
    .Y(_17114_));
 NAND2x1_ASAP7_75t_R _20219_ (.A(_05298_),
    .B(_05365_),
    .Y(_17125_));
 NAND2x1_ASAP7_75t_R _20220_ (.A(_05342_),
    .B(_05551_),
    .Y(_17141_));
 BUFx12f_ASAP7_75t_R _20221_ (.A(_05383_),
    .Y(_05552_));
 NAND2x1_ASAP7_75t_R _20222_ (.A(_05311_),
    .B(_05552_),
    .Y(_17152_));
 BUFx6f_ASAP7_75t_R _20223_ (.A(_05368_),
    .Y(_05553_));
 NAND2x1_ASAP7_75t_R _20224_ (.A(_05271_),
    .B(_05553_),
    .Y(_17161_));
 NAND2x1_ASAP7_75t_R _20225_ (.A(_05346_),
    .B(_05551_),
    .Y(_17170_));
 NAND2x1_ASAP7_75t_R _20226_ (.A(_05311_),
    .B(_05365_),
    .Y(_17181_));
 NAND2x1_ASAP7_75t_R _20227_ (.A(_05284_),
    .B(_05553_),
    .Y(_17191_));
 NAND2x1_ASAP7_75t_R _20228_ (.A(_05380_),
    .B(_05357_),
    .Y(_17208_));
 NAND2x1_ASAP7_75t_R _20229_ (.A(_05314_),
    .B(_05365_),
    .Y(_17219_));
 NAND2x1_ASAP7_75t_R _20230_ (.A(_05298_),
    .B(_05553_),
    .Y(_17228_));
 NAND2x1_ASAP7_75t_R _20231_ (.A(_05341_),
    .B(_05357_),
    .Y(_17240_));
 NAND2x1_ASAP7_75t_R _20232_ (.A(_05306_),
    .B(_05365_),
    .Y(_17251_));
 NAND2x1_ASAP7_75t_R _20233_ (.A(_05307_),
    .B(_05553_),
    .Y(_17260_));
 NAND2x1_ASAP7_75t_R _20234_ (.A(_05379_),
    .B(_05357_),
    .Y(_17278_));
 NAND2x1_ASAP7_75t_R _20235_ (.A(_05288_),
    .B(_05346_),
    .Y(_17283_));
 NAND2x1_ASAP7_75t_R _20236_ (.A(_05327_),
    .B(_05365_),
    .Y(_17290_));
 NAND2x1_ASAP7_75t_R _20237_ (.A(_05311_),
    .B(_05553_),
    .Y(_17300_));
 NAND2x1_ASAP7_75t_R _20238_ (.A(_05357_),
    .B(_05361_),
    .Y(_17324_));
 NAND2x1_ASAP7_75t_R _20239_ (.A(_05331_),
    .B(_05365_),
    .Y(_17335_));
 NAND2x1_ASAP7_75t_R _20240_ (.A(_05314_),
    .B(_05553_),
    .Y(_17344_));
 NAND2x1_ASAP7_75t_R _20241_ (.A(_05346_),
    .B(_05552_),
    .Y(_17375_));
 BUFx6f_ASAP7_75t_R _20242_ (.A(_05386_),
    .Y(_05554_));
 NAND2x1_ASAP7_75t_R _20243_ (.A(_05327_),
    .B(_05554_),
    .Y(_17385_));
 BUFx6f_ASAP7_75t_R _20244_ (.A(_05389_),
    .Y(_05555_));
 NAND2x1_ASAP7_75t_R _20245_ (.A(_05284_),
    .B(_05555_),
    .Y(_17400_));
 OR2x2_ASAP7_75t_R _20246_ (.A(_05270_),
    .B(_05393_),
    .Y(_17407_));
 NAND2x1_ASAP7_75t_R _20247_ (.A(_05346_),
    .B(_05365_),
    .Y(_17431_));
 NAND2x1_ASAP7_75t_R _20248_ (.A(_05327_),
    .B(_05553_),
    .Y(_17441_));
 OR2x2_ASAP7_75t_R _20249_ (.A(_05283_),
    .B(_05393_),
    .Y(_17455_));
 NAND2x1_ASAP7_75t_R _20250_ (.A(_05380_),
    .B(_05364_),
    .Y(_17476_));
 NAND2x1_ASAP7_75t_R _20251_ (.A(_05331_),
    .B(_05553_),
    .Y(_17486_));
 OR2x2_ASAP7_75t_R _20252_ (.A(_05277_),
    .B(_05393_),
    .Y(_17500_));
 NAND2x1_ASAP7_75t_R _20253_ (.A(_05341_),
    .B(_05364_),
    .Y(_17521_));
 NAND2x1_ASAP7_75t_R _20254_ (.A(_05342_),
    .B(_05553_),
    .Y(_17531_));
 OR2x2_ASAP7_75t_R _20255_ (.A(_05294_),
    .B(_05393_),
    .Y(_17545_));
 NAND2x1_ASAP7_75t_R _20256_ (.A(_05379_),
    .B(_05364_),
    .Y(_17565_));
 NAND2x1_ASAP7_75t_R _20257_ (.A(_05346_),
    .B(_05553_),
    .Y(_17576_));
 OR2x2_ASAP7_75t_R _20258_ (.A(_05291_),
    .B(_05393_),
    .Y(_17590_));
 NAND2x1_ASAP7_75t_R _20259_ (.A(_05380_),
    .B(_05368_),
    .Y(_17618_));
 OR2x2_ASAP7_75t_R _20260_ (.A(_05297_),
    .B(_05393_),
    .Y(_17632_));
 NAND2x1_ASAP7_75t_R _20261_ (.A(_05341_),
    .B(_05368_),
    .Y(_17659_));
 OR2x2_ASAP7_75t_R _20262_ (.A(_05305_),
    .B(_05392_),
    .Y(_17673_));
 NAND2x1_ASAP7_75t_R _20263_ (.A(_05379_),
    .B(_05368_),
    .Y(_17700_));
 OR2x2_ASAP7_75t_R _20264_ (.A(_05310_),
    .B(_05392_),
    .Y(_17714_));
 OR2x2_ASAP7_75t_R _20265_ (.A(_05313_),
    .B(_05392_),
    .Y(_17754_));
 OR2x2_ASAP7_75t_R _20266_ (.A(_05320_),
    .B(_05392_),
    .Y(_17790_));
 OR2x2_ASAP7_75t_R _20267_ (.A(_05326_),
    .B(_05392_),
    .Y(_17825_));
 OR2x2_ASAP7_75t_R _20268_ (.A(_05330_),
    .B(_05392_),
    .Y(_17857_));
 OR2x2_ASAP7_75t_R _20269_ (.A(_05340_),
    .B(_05392_),
    .Y(_17887_));
 OR2x2_ASAP7_75t_R _20270_ (.A(_05345_),
    .B(_05392_),
    .Y(_17915_));
 NAND2x1_ASAP7_75t_R _20271_ (.A(_05550_),
    .B(_05298_),
    .Y(_17004_));
 NAND2x1_ASAP7_75t_R _20272_ (.A(_05550_),
    .B(_05307_),
    .Y(_17013_));
 NAND2x1_ASAP7_75t_R _20273_ (.A(_05550_),
    .B(_05311_),
    .Y(_17019_));
 NAND2x1_ASAP7_75t_R _20274_ (.A(_05550_),
    .B(_05314_),
    .Y(_17035_));
 NAND2x1_ASAP7_75t_R _20275_ (.A(_05298_),
    .B(_05280_),
    .Y(_17040_));
 NAND2x1_ASAP7_75t_R _20276_ (.A(_05550_),
    .B(_05306_),
    .Y(_17047_));
 NAND2x1_ASAP7_75t_R _20277_ (.A(_05550_),
    .B(_05327_),
    .Y(_17065_));
 NAND2x1_ASAP7_75t_R _20278_ (.A(_05284_),
    .B(_05552_),
    .Y(_17077_));
 NAND2x1_ASAP7_75t_R _20279_ (.A(_05550_),
    .B(_05331_),
    .Y(_17093_));
 NAND2x1_ASAP7_75t_R _20280_ (.A(_05298_),
    .B(_05552_),
    .Y(_17105_));
 NAND2x1_ASAP7_75t_R _20281_ (.A(_05550_),
    .B(_05342_),
    .Y(_17115_));
 NAND2x1_ASAP7_75t_R _20282_ (.A(_05307_),
    .B(_05552_),
    .Y(_17126_));
 NAND2x1_ASAP7_75t_R _20283_ (.A(_05550_),
    .B(_05346_),
    .Y(_17142_));
 NAND2x1_ASAP7_75t_R _20284_ (.A(_05284_),
    .B(_05554_),
    .Y(_17162_));
 NAND2x1_ASAP7_75t_R _20285_ (.A(_05265_),
    .B(_05380_),
    .Y(_17171_));
 NAND2x1_ASAP7_75t_R _20286_ (.A(_05314_),
    .B(_05552_),
    .Y(_17182_));
 NAND2x1_ASAP7_75t_R _20287_ (.A(_05298_),
    .B(_05554_),
    .Y(_17192_));
 NAND2x1_ASAP7_75t_R _20288_ (.A(_05265_),
    .B(_05341_),
    .Y(_17209_));
 NAND2x1_ASAP7_75t_R _20289_ (.A(_05306_),
    .B(_05552_),
    .Y(_17220_));
 NAND2x1_ASAP7_75t_R _20290_ (.A(_05307_),
    .B(_05554_),
    .Y(_17229_));
 NAND2x1_ASAP7_75t_R _20291_ (.A(_05265_),
    .B(_05379_),
    .Y(_17241_));
 NAND2x1_ASAP7_75t_R _20292_ (.A(_05327_),
    .B(_05552_),
    .Y(_17252_));
 NAND2x1_ASAP7_75t_R _20293_ (.A(_05311_),
    .B(_05554_),
    .Y(_17261_));
 NAND2x1_ASAP7_75t_R _20294_ (.A(_05265_),
    .B(_05361_),
    .Y(_17279_));
 NAND2x1_ASAP7_75t_R _20295_ (.A(_05280_),
    .B(_05380_),
    .Y(_17284_));
 NAND2x1_ASAP7_75t_R _20296_ (.A(_05331_),
    .B(_05552_),
    .Y(_17291_));
 NAND2x1_ASAP7_75t_R _20297_ (.A(_05314_),
    .B(_05554_),
    .Y(_17301_));
 NAND2x1_ASAP7_75t_R _20298_ (.A(_05265_),
    .B(_05369_),
    .Y(_17325_));
 NAND2x1_ASAP7_75t_R _20299_ (.A(_05342_),
    .B(_05552_),
    .Y(_17336_));
 NAND2x1_ASAP7_75t_R _20300_ (.A(_05306_),
    .B(_05554_),
    .Y(_17345_));
 NAND2x1_ASAP7_75t_R _20301_ (.A(_05301_),
    .B(_05380_),
    .Y(_17376_));
 NAND2x1_ASAP7_75t_R _20302_ (.A(_05331_),
    .B(_05318_),
    .Y(_17386_));
 NAND2x1_ASAP7_75t_R _20303_ (.A(_05298_),
    .B(_05371_),
    .Y(_17401_));
 NAND2x1_ASAP7_75t_R _20304_ (.A(_05380_),
    .B(_05383_),
    .Y(_17432_));
 NAND2x1_ASAP7_75t_R _20305_ (.A(_05331_),
    .B(_05554_),
    .Y(_17442_));
 NAND2x1_ASAP7_75t_R _20306_ (.A(_05277_),
    .B(_05555_),
    .Y(_17456_));
 NAND2x1_ASAP7_75t_R _20307_ (.A(_05341_),
    .B(_05383_),
    .Y(_17477_));
 NAND2x1_ASAP7_75t_R _20308_ (.A(_05342_),
    .B(_05554_),
    .Y(_17487_));
 NAND2x1_ASAP7_75t_R _20309_ (.A(_05294_),
    .B(_05555_),
    .Y(_17501_));
 NAND2x1_ASAP7_75t_R _20310_ (.A(_05379_),
    .B(_05383_),
    .Y(_17522_));
 NAND2x1_ASAP7_75t_R _20311_ (.A(_05346_),
    .B(_05554_),
    .Y(_17532_));
 NAND2x1_ASAP7_75t_R _20312_ (.A(_05311_),
    .B(_05555_),
    .Y(_17546_));
 NAND2x1_ASAP7_75t_R _20313_ (.A(_05361_),
    .B(_05383_),
    .Y(_17566_));
 NAND2x1_ASAP7_75t_R _20314_ (.A(_05380_),
    .B(_05386_),
    .Y(_17577_));
 NAND2x1_ASAP7_75t_R _20315_ (.A(_05314_),
    .B(_05555_),
    .Y(_17591_));
 NAND2x1_ASAP7_75t_R _20316_ (.A(_05340_),
    .B(_05386_),
    .Y(_17619_));
 NAND2x1_ASAP7_75t_R _20317_ (.A(_05306_),
    .B(_05555_),
    .Y(_17633_));
 NAND2x1_ASAP7_75t_R _20318_ (.A(_05379_),
    .B(_05386_),
    .Y(_17660_));
 NAND2x1_ASAP7_75t_R _20319_ (.A(_05327_),
    .B(_05555_),
    .Y(_17674_));
 NAND2x1_ASAP7_75t_R _20320_ (.A(_05361_),
    .B(_05386_),
    .Y(_17701_));
 NAND2x1_ASAP7_75t_R _20321_ (.A(_05331_),
    .B(_05555_),
    .Y(_17715_));
 NAND2x1_ASAP7_75t_R _20322_ (.A(_05342_),
    .B(_05555_),
    .Y(_17755_));
 NAND2x1_ASAP7_75t_R _20323_ (.A(_05326_),
    .B(_05555_),
    .Y(_17791_));
 NAND2x1_ASAP7_75t_R _20324_ (.A(_05330_),
    .B(_05389_),
    .Y(_17826_));
 NAND2x1_ASAP7_75t_R _20325_ (.A(_05340_),
    .B(_05389_),
    .Y(_17858_));
 NAND2x1_ASAP7_75t_R _20326_ (.A(_05379_),
    .B(_05389_),
    .Y(_17888_));
 NAND2x1_ASAP7_75t_R _20327_ (.A(_05361_),
    .B(_05389_),
    .Y(_17916_));
 NAND2x1_ASAP7_75t_R _20328_ (.A(_05526_),
    .B(_05536_),
    .Y(_17998_));
 NAND2x1_ASAP7_75t_R _20329_ (.A(_05271_),
    .B(_05357_),
    .Y(_17002_));
 NAND2x1_ASAP7_75t_R _20330_ (.A(_05274_),
    .B(_05307_),
    .Y(_17041_));
 NAND2x1_ASAP7_75t_R _20331_ (.A(_05294_),
    .B(_05364_),
    .Y(_17154_));
 INVx2_ASAP7_75t_R _20332_ (.A(_05354_),
    .Y(_05556_));
 AND3x4_ASAP7_75t_R _20333_ (.A(_14636_),
    .B(_14633_),
    .C(_14628_),
    .Y(_05557_));
 BUFx6f_ASAP7_75t_R _20334_ (.A(_05557_),
    .Y(_05558_));
 BUFx6f_ASAP7_75t_R _20335_ (.A(_14639_),
    .Y(_05559_));
 AO222x2_ASAP7_75t_R _20336_ (.A1(_05559_),
    .A2(_00097_),
    .B1(_01745_),
    .B2(_14906_),
    .C1(_14528_),
    .C2(_14640_),
    .Y(_05560_));
 AO21x1_ASAP7_75t_R _20337_ (.A1(_05556_),
    .A2(_05558_),
    .B(_05560_),
    .Y(_05561_));
 OR2x2_ASAP7_75t_R _20338_ (.A(_18559_),
    .B(_14632_),
    .Y(_05562_));
 OA21x2_ASAP7_75t_R _20339_ (.A1(_18552_),
    .A2(_14621_),
    .B(_05562_),
    .Y(_05563_));
 AO21x1_ASAP7_75t_R _20340_ (.A1(_15236_),
    .A2(_05561_),
    .B(_05563_),
    .Y(_18009_));
 BUFx6f_ASAP7_75t_R _20341_ (.A(_14621_),
    .Y(_05564_));
 BUFx3_ASAP7_75t_R _20342_ (.A(_14632_),
    .Y(_05565_));
 BUFx6f_ASAP7_75t_R _20343_ (.A(_14636_),
    .Y(_05566_));
 INVx1_ASAP7_75t_R _20344_ (.A(_00100_),
    .Y(_05567_));
 INVx1_ASAP7_75t_R _20345_ (.A(_01734_),
    .Y(_05568_));
 OA222x2_ASAP7_75t_R _20346_ (.A1(_05566_),
    .A2(_05567_),
    .B1(_05568_),
    .B2(_14629_),
    .C1(_14642_),
    .C2(_13601_),
    .Y(_05569_));
 OAI21x1_ASAP7_75t_R _20347_ (.A1(_05203_),
    .A2(_14703_),
    .B(_05569_),
    .Y(_05570_));
 AO22x1_ASAP7_75t_R _20348_ (.A1(_18565_),
    .A2(_05565_),
    .B1(_14625_),
    .B2(_05570_),
    .Y(_05571_));
 AO21x1_ASAP7_75t_R _20349_ (.A1(_18563_),
    .A2(_05564_),
    .B(_05571_),
    .Y(_18011_));
 INVx2_ASAP7_75t_R _20350_ (.A(_13684_),
    .Y(_05572_));
 BUFx6f_ASAP7_75t_R _20351_ (.A(_14639_),
    .Y(_05573_));
 NOR2x1_ASAP7_75t_R _20352_ (.A(_14633_),
    .B(_14770_),
    .Y(_05574_));
 AO221x1_ASAP7_75t_R _20353_ (.A1(_05573_),
    .A2(_00104_),
    .B1(_01731_),
    .B2(_14906_),
    .C(_05574_),
    .Y(_05575_));
 AO21x1_ASAP7_75t_R _20354_ (.A1(_05572_),
    .A2(_05558_),
    .B(_05575_),
    .Y(_05576_));
 AO22x1_ASAP7_75t_R _20355_ (.A1(_18570_),
    .A2(_05565_),
    .B1(_14625_),
    .B2(_05576_),
    .Y(_05577_));
 AO21x1_ASAP7_75t_R _20356_ (.A1(_18568_),
    .A2(_05564_),
    .B(_05577_),
    .Y(_18013_));
 INVx2_ASAP7_75t_R _20357_ (.A(_13762_),
    .Y(_05578_));
 NOR2x1_ASAP7_75t_R _20358_ (.A(_14633_),
    .B(_14835_),
    .Y(_05579_));
 AO221x1_ASAP7_75t_R _20359_ (.A1(_05573_),
    .A2(_00109_),
    .B1(_01730_),
    .B2(_14906_),
    .C(_05579_),
    .Y(_05580_));
 AO21x1_ASAP7_75t_R _20360_ (.A1(_05578_),
    .A2(_05558_),
    .B(_05580_),
    .Y(_05581_));
 AO22x1_ASAP7_75t_R _20361_ (.A1(_18575_),
    .A2(_05565_),
    .B1(_14625_),
    .B2(_05581_),
    .Y(_05582_));
 AO21x1_ASAP7_75t_R _20362_ (.A1(_18573_),
    .A2(_05564_),
    .B(_05582_),
    .Y(_18015_));
 AND2x6_ASAP7_75t_R _20363_ (.A(_14869_),
    .B(_14898_),
    .Y(_05583_));
 INVx1_ASAP7_75t_R _20364_ (.A(_01729_),
    .Y(_05584_));
 OA222x2_ASAP7_75t_R _20365_ (.A1(_05566_),
    .A2(_14904_),
    .B1(_05584_),
    .B2(_14628_),
    .C1(_14642_),
    .C2(_13830_),
    .Y(_05585_));
 OAI21x1_ASAP7_75t_R _20366_ (.A1(_05203_),
    .A2(_05583_),
    .B(_05585_),
    .Y(_05586_));
 AO22x1_ASAP7_75t_R _20367_ (.A1(_18580_),
    .A2(_05565_),
    .B1(_14625_),
    .B2(_05586_),
    .Y(_05587_));
 AO21x1_ASAP7_75t_R _20368_ (.A1(_18578_),
    .A2(_05564_),
    .B(_05587_),
    .Y(_18017_));
 BUFx6f_ASAP7_75t_R _20369_ (.A(_14624_),
    .Y(_05588_));
 BUFx6f_ASAP7_75t_R _20370_ (.A(_14642_),
    .Y(_05589_));
 INVx1_ASAP7_75t_R _20371_ (.A(_01727_),
    .Y(_05590_));
 OA222x2_ASAP7_75t_R _20372_ (.A1(_05566_),
    .A2(_14971_),
    .B1(_05590_),
    .B2(_14628_),
    .C1(_05303_),
    .C2(_14634_),
    .Y(_05591_));
 OAI21x1_ASAP7_75t_R _20373_ (.A1(_13908_),
    .A2(_05589_),
    .B(_05591_),
    .Y(_05592_));
 AO22x1_ASAP7_75t_R _20374_ (.A1(_18585_),
    .A2(_14632_),
    .B1(_05588_),
    .B2(_05592_),
    .Y(_05593_));
 AO21x1_ASAP7_75t_R _20375_ (.A1(_18583_),
    .A2(_05564_),
    .B(_05593_),
    .Y(_18019_));
 INVx1_ASAP7_75t_R _20376_ (.A(_01726_),
    .Y(_05594_));
 AND2x6_ASAP7_75t_R _20377_ (.A(_14998_),
    .B(_15023_),
    .Y(_05595_));
 OA222x2_ASAP7_75t_R _20378_ (.A1(_05566_),
    .A2(_15027_),
    .B1(_05594_),
    .B2(_14628_),
    .C1(_05595_),
    .C2(_14634_),
    .Y(_05596_));
 OAI21x1_ASAP7_75t_R _20379_ (.A1(_13968_),
    .A2(_05589_),
    .B(_05596_),
    .Y(_05597_));
 AO22x1_ASAP7_75t_R _20380_ (.A1(_18590_),
    .A2(_14632_),
    .B1(_05588_),
    .B2(_05597_),
    .Y(_05598_));
 AO21x1_ASAP7_75t_R _20381_ (.A1(_18588_),
    .A2(_05564_),
    .B(_05598_),
    .Y(_18021_));
 BUFx6f_ASAP7_75t_R _20382_ (.A(_14632_),
    .Y(_05599_));
 BUFx6f_ASAP7_75t_R _20383_ (.A(_14634_),
    .Y(_05600_));
 NOR2x1_ASAP7_75t_R _20384_ (.A(_05600_),
    .B(_15098_),
    .Y(_05601_));
 AO222x2_ASAP7_75t_R _20385_ (.A1(_05573_),
    .A2(_00135_),
    .B1(_01725_),
    .B2(_14905_),
    .C1(_05557_),
    .C2(_04996_),
    .Y(_05602_));
 OA21x2_ASAP7_75t_R _20386_ (.A1(_05601_),
    .A2(_05602_),
    .B(_15236_),
    .Y(_05603_));
 AO21x1_ASAP7_75t_R _20387_ (.A1(_18595_),
    .A2(_05599_),
    .B(_05603_),
    .Y(_05604_));
 AO21x1_ASAP7_75t_R _20388_ (.A1(_18593_),
    .A2(_05564_),
    .B(_05604_),
    .Y(_18023_));
 AND2x6_ASAP7_75t_R _20389_ (.A(_15132_),
    .B(_15156_),
    .Y(_05605_));
 AOI22x1_ASAP7_75t_R _20390_ (.A1(_05559_),
    .A2(_00144_),
    .B1(_02201_),
    .B2(_14906_),
    .Y(_05606_));
 OA21x2_ASAP7_75t_R _20391_ (.A1(_14089_),
    .A2(_05589_),
    .B(_05606_),
    .Y(_05607_));
 OAI21x1_ASAP7_75t_R _20392_ (.A1(_05203_),
    .A2(_05605_),
    .B(_05607_),
    .Y(_05608_));
 AO22x1_ASAP7_75t_R _20393_ (.A1(_18600_),
    .A2(_14632_),
    .B1(_05588_),
    .B2(_05608_),
    .Y(_05609_));
 AO21x1_ASAP7_75t_R _20394_ (.A1(_18598_),
    .A2(_05564_),
    .B(_05609_),
    .Y(_18025_));
 NOR2x1_ASAP7_75t_R _20395_ (.A(_05600_),
    .B(_05324_),
    .Y(_05610_));
 AO222x2_ASAP7_75t_R _20396_ (.A1(_05573_),
    .A2(_00152_),
    .B1(_01755_),
    .B2(_14905_),
    .C1(_05557_),
    .C2(_05002_),
    .Y(_05611_));
 OA21x2_ASAP7_75t_R _20397_ (.A1(_05610_),
    .A2(_05611_),
    .B(_15235_),
    .Y(_05612_));
 AO21x1_ASAP7_75t_R _20398_ (.A1(_18605_),
    .A2(_05599_),
    .B(_05612_),
    .Y(_05613_));
 AO21x1_ASAP7_75t_R _20399_ (.A1(_18603_),
    .A2(_05564_),
    .B(_05613_),
    .Y(_18027_));
 INVx1_ASAP7_75t_R _20400_ (.A(_01754_),
    .Y(_05614_));
 OA222x2_ASAP7_75t_R _20401_ (.A1(_05566_),
    .A2(_15232_),
    .B1(_05614_),
    .B2(_14628_),
    .C1(_14642_),
    .C2(_14260_),
    .Y(_05615_));
 OAI21x1_ASAP7_75t_R _20402_ (.A1(_05600_),
    .A2(_05328_),
    .B(_05615_),
    .Y(_05616_));
 AO32x1_ASAP7_75t_R _20403_ (.A1(_05007_),
    .A2(_05008_),
    .A3(_14632_),
    .B1(_14624_),
    .B2(_05616_),
    .Y(_05617_));
 AO21x1_ASAP7_75t_R _20404_ (.A1(_18608_),
    .A2(_05564_),
    .B(_05617_),
    .Y(_18029_));
 NAND2x2_ASAP7_75t_R _20405_ (.A(_13162_),
    .B(_13216_),
    .Y(_05618_));
 AO222x2_ASAP7_75t_R _20406_ (.A1(_05573_),
    .A2(_00168_),
    .B1(_01753_),
    .B2(_14905_),
    .C1(_05557_),
    .C2(_15363_),
    .Y(_05619_));
 AO21x1_ASAP7_75t_R _20407_ (.A1(_14640_),
    .A2(_05618_),
    .B(_05619_),
    .Y(_05620_));
 AO22x1_ASAP7_75t_R _20408_ (.A1(_05599_),
    .A2(_18612_),
    .B1(_05620_),
    .B2(_05588_),
    .Y(_05621_));
 AO21x1_ASAP7_75t_R _20409_ (.A1(_16998_),
    .A2(_18614_),
    .B(_05621_),
    .Y(_18031_));
 BUFx6f_ASAP7_75t_R _20410_ (.A(_14639_),
    .Y(_05622_));
 AO222x2_ASAP7_75t_R _20411_ (.A1(_05622_),
    .A2(_00175_),
    .B1(_01752_),
    .B2(_14906_),
    .C1(_05558_),
    .C2(_15502_),
    .Y(_05623_));
 AND2x6_ASAP7_75t_R _20412_ (.A(_15398_),
    .B(_15429_),
    .Y(_05624_));
 NOR2x1_ASAP7_75t_R _20413_ (.A(_05600_),
    .B(_05624_),
    .Y(_05625_));
 OA21x2_ASAP7_75t_R _20414_ (.A1(_05623_),
    .A2(_05625_),
    .B(_15235_),
    .Y(_05626_));
 AO21x1_ASAP7_75t_R _20415_ (.A1(_05599_),
    .A2(_18617_),
    .B(_05626_),
    .Y(_05627_));
 AO21x1_ASAP7_75t_R _20416_ (.A1(_16998_),
    .A2(_18619_),
    .B(_05627_),
    .Y(_18033_));
 AO222x2_ASAP7_75t_R _20417_ (.A1(_05573_),
    .A2(_00180_),
    .B1(_01751_),
    .B2(_14905_),
    .C1(_05557_),
    .C2(_15646_),
    .Y(_05628_));
 AO21x1_ASAP7_75t_R _20418_ (.A1(_14640_),
    .A2(_15583_),
    .B(_05628_),
    .Y(_05629_));
 AO22x1_ASAP7_75t_R _20419_ (.A1(_05565_),
    .A2(_18622_),
    .B1(_05629_),
    .B2(_05588_),
    .Y(_05630_));
 AO21x1_ASAP7_75t_R _20420_ (.A1(_16998_),
    .A2(_18624_),
    .B(_05630_),
    .Y(_18035_));
 NOR2x1_ASAP7_75t_R _20421_ (.A(_14634_),
    .B(_15707_),
    .Y(_05631_));
 AO221x1_ASAP7_75t_R _20422_ (.A1(_05622_),
    .A2(_00187_),
    .B1(_01750_),
    .B2(_14906_),
    .C(_05631_),
    .Y(_05632_));
 AO21x1_ASAP7_75t_R _20423_ (.A1(_05558_),
    .A2(_15759_),
    .B(_05632_),
    .Y(_05633_));
 AO22x1_ASAP7_75t_R _20424_ (.A1(_05565_),
    .A2(_18627_),
    .B1(_05633_),
    .B2(_05588_),
    .Y(_05634_));
 AO21x1_ASAP7_75t_R _20425_ (.A1(_16998_),
    .A2(_18629_),
    .B(_05634_),
    .Y(_18037_));
 BUFx6f_ASAP7_75t_R _20426_ (.A(_14636_),
    .Y(_05635_));
 INVx1_ASAP7_75t_R _20427_ (.A(_15836_),
    .Y(_05636_));
 INVx1_ASAP7_75t_R _20428_ (.A(_01749_),
    .Y(_05637_));
 OA222x2_ASAP7_75t_R _20429_ (.A1(_05635_),
    .A2(_05636_),
    .B1(_05637_),
    .B2(_14629_),
    .C1(_15831_),
    .C2(_14634_),
    .Y(_05638_));
 OA21x2_ASAP7_75t_R _20430_ (.A1(_05589_),
    .A2(_05261_),
    .B(_05638_),
    .Y(_05639_));
 OAI22x1_ASAP7_75t_R _20431_ (.A1(_15241_),
    .A2(_18634_),
    .B1(_05639_),
    .B2(_14648_),
    .Y(_05640_));
 AO21x1_ASAP7_75t_R _20432_ (.A1(_16998_),
    .A2(_18634_),
    .B(_05640_),
    .Y(_18039_));
 AO222x2_ASAP7_75t_R _20433_ (.A1(_05622_),
    .A2(_15947_),
    .B1(_01748_),
    .B2(_14906_),
    .C1(_05558_),
    .C2(_15995_),
    .Y(_05641_));
 NOR2x1_ASAP7_75t_R _20434_ (.A(_05600_),
    .B(_05281_),
    .Y(_05642_));
 OA21x2_ASAP7_75t_R _20435_ (.A1(_05641_),
    .A2(_05642_),
    .B(_15235_),
    .Y(_05643_));
 AO21x1_ASAP7_75t_R _20436_ (.A1(_05599_),
    .A2(_18637_),
    .B(_05643_),
    .Y(_05644_));
 AO21x1_ASAP7_75t_R _20437_ (.A1(_16998_),
    .A2(_18639_),
    .B(_05644_),
    .Y(_18041_));
 AO222x2_ASAP7_75t_R _20438_ (.A1(_05622_),
    .A2(_16083_),
    .B1(_01747_),
    .B2(_14906_),
    .C1(_05558_),
    .C2(_16131_),
    .Y(_05645_));
 NOR2x1_ASAP7_75t_R _20439_ (.A(_05600_),
    .B(_16078_),
    .Y(_05646_));
 OA21x2_ASAP7_75t_R _20440_ (.A1(_05645_),
    .A2(_05646_),
    .B(_15235_),
    .Y(_05647_));
 AO21x1_ASAP7_75t_R _20441_ (.A1(_05599_),
    .A2(_18642_),
    .B(_05647_),
    .Y(_05648_));
 AO21x1_ASAP7_75t_R _20442_ (.A1(_16998_),
    .A2(_18644_),
    .B(_05648_),
    .Y(_18043_));
 AO222x2_ASAP7_75t_R _20443_ (.A1(_05622_),
    .A2(_16195_),
    .B1(_01746_),
    .B2(_14905_),
    .C1(_05558_),
    .C2(_16242_),
    .Y(_05649_));
 AND2x4_ASAP7_75t_R _20444_ (.A(_16159_),
    .B(_16190_),
    .Y(_05650_));
 NOR2x1_ASAP7_75t_R _20445_ (.A(_05600_),
    .B(_05650_),
    .Y(_05651_));
 OA21x2_ASAP7_75t_R _20446_ (.A1(_05649_),
    .A2(_05651_),
    .B(_15235_),
    .Y(_05652_));
 AO21x1_ASAP7_75t_R _20447_ (.A1(_05599_),
    .A2(_18647_),
    .B(_05652_),
    .Y(_05653_));
 AO21x1_ASAP7_75t_R _20448_ (.A1(_16998_),
    .A2(_18649_),
    .B(_05653_),
    .Y(_18045_));
 AND2x6_ASAP7_75t_R _20449_ (.A(_16294_),
    .B(_16325_),
    .Y(_05654_));
 INVx1_ASAP7_75t_R _20450_ (.A(_01744_),
    .Y(_05655_));
 OA222x2_ASAP7_75t_R _20451_ (.A1(_05635_),
    .A2(_16330_),
    .B1(_05655_),
    .B2(_14629_),
    .C1(_05589_),
    .C2(_16384_),
    .Y(_05656_));
 OA21x2_ASAP7_75t_R _20452_ (.A1(_05203_),
    .A2(_05654_),
    .B(_05656_),
    .Y(_05657_));
 OAI22x1_ASAP7_75t_R _20453_ (.A1(_15241_),
    .A2(_18654_),
    .B1(_05657_),
    .B2(_14648_),
    .Y(_05658_));
 AO21x1_ASAP7_75t_R _20454_ (.A1(_16998_),
    .A2(_18654_),
    .B(_05658_),
    .Y(_18047_));
 BUFx6f_ASAP7_75t_R _20455_ (.A(_14621_),
    .Y(_05659_));
 INVx1_ASAP7_75t_R _20456_ (.A(_01743_),
    .Y(_05660_));
 OA222x2_ASAP7_75t_R _20457_ (.A1(_05635_),
    .A2(_16452_),
    .B1(_05660_),
    .B2(_14629_),
    .C1(_05589_),
    .C2(_16498_),
    .Y(_05661_));
 OA21x2_ASAP7_75t_R _20458_ (.A1(_05203_),
    .A2(_05295_),
    .B(_05661_),
    .Y(_05662_));
 OAI22x1_ASAP7_75t_R _20459_ (.A1(_15241_),
    .A2(_18659_),
    .B1(_05662_),
    .B2(_14648_),
    .Y(_05663_));
 AO21x1_ASAP7_75t_R _20460_ (.A1(_05659_),
    .A2(_18659_),
    .B(_05663_),
    .Y(_18049_));
 AO222x2_ASAP7_75t_R _20461_ (.A1(_05573_),
    .A2(_16591_),
    .B1(_01742_),
    .B2(_14905_),
    .C1(_05558_),
    .C2(_16637_),
    .Y(_05664_));
 NOR2x1_ASAP7_75t_R _20462_ (.A(_05600_),
    .B(_16587_),
    .Y(_05665_));
 OA21x2_ASAP7_75t_R _20463_ (.A1(_05664_),
    .A2(_05665_),
    .B(_15235_),
    .Y(_05666_));
 AO21x1_ASAP7_75t_R _20464_ (.A1(_05599_),
    .A2(_18662_),
    .B(_05666_),
    .Y(_05667_));
 AO21x1_ASAP7_75t_R _20465_ (.A1(_05659_),
    .A2(_18664_),
    .B(_05667_),
    .Y(_18051_));
 AO222x2_ASAP7_75t_R _20466_ (.A1(_05573_),
    .A2(_16701_),
    .B1(_01741_),
    .B2(_14905_),
    .C1(_05558_),
    .C2(_16747_),
    .Y(_05668_));
 NOR2x1_ASAP7_75t_R _20467_ (.A(_14634_),
    .B(_05308_),
    .Y(_05669_));
 OA21x2_ASAP7_75t_R _20468_ (.A1(_05668_),
    .A2(_05669_),
    .B(_15235_),
    .Y(_05670_));
 AO21x1_ASAP7_75t_R _20469_ (.A1(_05599_),
    .A2(_18667_),
    .B(_05670_),
    .Y(_05671_));
 AO21x1_ASAP7_75t_R _20470_ (.A1(_05659_),
    .A2(_18669_),
    .B(_05671_),
    .Y(_18053_));
 AND2x6_ASAP7_75t_R _20471_ (.A(_16788_),
    .B(_16819_),
    .Y(_05672_));
 INVx1_ASAP7_75t_R _20472_ (.A(_01740_),
    .Y(_05673_));
 OA222x2_ASAP7_75t_R _20473_ (.A1(_05635_),
    .A2(_16824_),
    .B1(_05673_),
    .B2(_14629_),
    .C1(_05589_),
    .C2(_16870_),
    .Y(_05674_));
 OA21x2_ASAP7_75t_R _20474_ (.A1(_05600_),
    .A2(_05672_),
    .B(_05674_),
    .Y(_05675_));
 OAI22x1_ASAP7_75t_R _20475_ (.A1(_15241_),
    .A2(_18674_),
    .B1(_05675_),
    .B2(_14648_),
    .Y(_05676_));
 AO21x1_ASAP7_75t_R _20476_ (.A1(_05659_),
    .A2(_18674_),
    .B(_05676_),
    .Y(_18055_));
 INVx1_ASAP7_75t_R _20477_ (.A(_01739_),
    .Y(_05677_));
 OA222x2_ASAP7_75t_R _20478_ (.A1(_05635_),
    .A2(_16936_),
    .B1(_05677_),
    .B2(_14629_),
    .C1(_05589_),
    .C2(_16983_),
    .Y(_05678_));
 OAI21x1_ASAP7_75t_R _20479_ (.A1(_05203_),
    .A2(_16931_),
    .B(_05678_),
    .Y(_05679_));
 AO22x1_ASAP7_75t_R _20480_ (.A1(_05565_),
    .A2(_18677_),
    .B1(_05679_),
    .B2(_05588_),
    .Y(_05680_));
 AO21x1_ASAP7_75t_R _20481_ (.A1(_05659_),
    .A2(_18679_),
    .B(_05680_),
    .Y(_18057_));
 INVx1_ASAP7_75t_R _20482_ (.A(_01738_),
    .Y(_05681_));
 OA222x2_ASAP7_75t_R _20483_ (.A1(_05635_),
    .A2(_04311_),
    .B1(_05681_),
    .B2(_14629_),
    .C1(_05589_),
    .C2(_04357_),
    .Y(_05682_));
 OAI21x1_ASAP7_75t_R _20484_ (.A1(_05203_),
    .A2(_04305_),
    .B(_05682_),
    .Y(_05683_));
 AO22x1_ASAP7_75t_R _20485_ (.A1(_05565_),
    .A2(_18682_),
    .B1(_05683_),
    .B2(_05588_),
    .Y(_05684_));
 AO21x1_ASAP7_75t_R _20486_ (.A1(_05659_),
    .A2(_18684_),
    .B(_05684_),
    .Y(_18059_));
 NAND2x2_ASAP7_75t_R _20487_ (.A(_04386_),
    .B(_04417_),
    .Y(_05685_));
 AO222x2_ASAP7_75t_R _20488_ (.A1(_05573_),
    .A2(_04422_),
    .B1(_01737_),
    .B2(_14905_),
    .C1(_05557_),
    .C2(_04468_),
    .Y(_05686_));
 AO21x1_ASAP7_75t_R _20489_ (.A1(_14640_),
    .A2(_05685_),
    .B(_05686_),
    .Y(_05687_));
 AO22x1_ASAP7_75t_R _20490_ (.A1(_05565_),
    .A2(_18687_),
    .B1(_05687_),
    .B2(_05588_),
    .Y(_05688_));
 AO21x1_ASAP7_75t_R _20491_ (.A1(_05659_),
    .A2(_18689_),
    .B(_05688_),
    .Y(_18061_));
 INVx1_ASAP7_75t_R _20492_ (.A(_01736_),
    .Y(_05689_));
 OA222x2_ASAP7_75t_R _20493_ (.A1(_05635_),
    .A2(_04559_),
    .B1(_05689_),
    .B2(_14629_),
    .C1(_14642_),
    .C2(_04605_),
    .Y(_05690_));
 OAI21x1_ASAP7_75t_R _20494_ (.A1(_05203_),
    .A2(_04554_),
    .B(_05690_),
    .Y(_05691_));
 AO22x1_ASAP7_75t_R _20495_ (.A1(_05565_),
    .A2(_18692_),
    .B1(_05691_),
    .B2(_05588_),
    .Y(_05692_));
 AO21x1_ASAP7_75t_R _20496_ (.A1(_05659_),
    .A2(_18694_),
    .B(_05692_),
    .Y(_18063_));
 INVx1_ASAP7_75t_R _20497_ (.A(_01735_),
    .Y(_05693_));
 OA222x2_ASAP7_75t_R _20498_ (.A1(_05635_),
    .A2(_04671_),
    .B1(_05693_),
    .B2(_14629_),
    .C1(_05589_),
    .C2(_04717_),
    .Y(_05694_));
 OA21x2_ASAP7_75t_R _20499_ (.A1(_05600_),
    .A2(_05343_),
    .B(_05694_),
    .Y(_05695_));
 OAI22x1_ASAP7_75t_R _20500_ (.A1(_15241_),
    .A2(_18699_),
    .B1(_05695_),
    .B2(_14648_),
    .Y(_05696_));
 AO21x1_ASAP7_75t_R _20501_ (.A1(_05659_),
    .A2(_18699_),
    .B(_05696_),
    .Y(_18065_));
 AO222x2_ASAP7_75t_R _20502_ (.A1(_05573_),
    .A2(_04791_),
    .B1(_01733_),
    .B2(_14905_),
    .C1(_05557_),
    .C2(_04837_),
    .Y(_05697_));
 NOR2x1_ASAP7_75t_R _20503_ (.A(_14634_),
    .B(_05358_),
    .Y(_05698_));
 OA21x2_ASAP7_75t_R _20504_ (.A1(_05697_),
    .A2(_05698_),
    .B(_15235_),
    .Y(_05699_));
 AO21x1_ASAP7_75t_R _20505_ (.A1(_05599_),
    .A2(_18702_),
    .B(_05699_),
    .Y(_05700_));
 AO21x1_ASAP7_75t_R _20506_ (.A1(_05659_),
    .A2(_18704_),
    .B(_05700_),
    .Y(_18067_));
 AND2x2_ASAP7_75t_R _20507_ (.A(_05271_),
    .B(_05280_),
    .Y(_18097_));
 AND2x2_ASAP7_75t_R _20508_ (.A(_05271_),
    .B(_05301_),
    .Y(_18113_));
 AND2x2_ASAP7_75t_R _20509_ (.A(_05270_),
    .B(_05383_),
    .Y(_18124_));
 AND2x4_ASAP7_75t_R _20510_ (.A(_05270_),
    .B(_05317_),
    .Y(_18146_));
 INVx1_ASAP7_75t_R _20511_ (.A(_00139_),
    .Y(_17087_));
 AND2x2_ASAP7_75t_R _20512_ (.A(_05270_),
    .B(_05386_),
    .Y(_18158_));
 INVx1_ASAP7_75t_R _20513_ (.A(_00162_),
    .Y(_17198_));
 AND2x4_ASAP7_75t_R _20514_ (.A(_05270_),
    .B(_05333_),
    .Y(_18199_));
 INVx1_ASAP7_75t_R _20515_ (.A(_00170_),
    .Y(_17206_));
 AND2x2_ASAP7_75t_R _20516_ (.A(_05270_),
    .B(_05371_),
    .Y(_18242_));
 AND2x2_ASAP7_75t_R _20517_ (.A(_05270_),
    .B(_05389_),
    .Y(_18263_));
 INVx1_ASAP7_75t_R _20518_ (.A(_00193_),
    .Y(_17322_));
 INVx1_ASAP7_75t_R _20519_ (.A(_05393_),
    .Y(_17366_));
 INVx1_ASAP7_75t_R _20520_ (.A(_00198_),
    .Y(_17363_));
 INVx1_ASAP7_75t_R _20521_ (.A(_00201_),
    .Y(_17406_));
 INVx1_ASAP7_75t_R _20522_ (.A(_00202_),
    .Y(_17419_));
 INVx1_ASAP7_75t_R _20523_ (.A(_00206_),
    .Y(_17507_));
 INVx1_ASAP7_75t_R _20524_ (.A(_17690_),
    .Y(_17646_));
 INVx1_ASAP7_75t_R _20525_ (.A(_00221_),
    .Y(_17721_));
 INVx1_ASAP7_75t_R _20526_ (.A(_00224_),
    .Y(_17761_));
 INVx1_ASAP7_75t_R _20527_ (.A(_00227_),
    .Y(_17797_));
 INVx1_ASAP7_75t_R _20528_ (.A(_17806_),
    .Y(_17768_));
 INVx1_ASAP7_75t_R _20529_ (.A(_00230_),
    .Y(_17832_));
 INVx1_ASAP7_75t_R _20530_ (.A(_17841_),
    .Y(_17804_));
 INVx1_ASAP7_75t_R _20531_ (.A(_17873_),
    .Y(_17839_));
 INVx1_ASAP7_75t_R _20532_ (.A(_17902_),
    .Y(_17871_));
 INVx2_ASAP7_75t_R _20533_ (.A(_00248_),
    .Y(_17990_));
 INVx1_ASAP7_75t_R _20534_ (.A(_00251_),
    .Y(_17993_));
 BUFx6f_ASAP7_75t_R _20535_ (.A(_05071_),
    .Y(_05701_));
 BUFx6f_ASAP7_75t_R _20536_ (.A(_05701_),
    .Y(_05702_));
 NAND2x1_ASAP7_75t_R _20537_ (.A(_18593_),
    .B(_05702_),
    .Y(_18082_));
 AND2x2_ASAP7_75t_R _20538_ (.A(_05273_),
    .B(_05284_),
    .Y(_18098_));
 AND2x2_ASAP7_75t_R _20539_ (.A(_05283_),
    .B(_05301_),
    .Y(_18125_));
 AND2x2_ASAP7_75t_R _20540_ (.A(_05283_),
    .B(_05317_),
    .Y(_18159_));
 INVx1_ASAP7_75t_R _20541_ (.A(_00157_),
    .Y(_18176_));
 AND2x2_ASAP7_75t_R _20542_ (.A(_05283_),
    .B(_05323_),
    .Y(_18200_));
 INVx1_ASAP7_75t_R _20543_ (.A(_00177_),
    .Y(_18227_));
 INVx1_ASAP7_75t_R _20544_ (.A(_00184_),
    .Y(_17323_));
 AND2x2_ASAP7_75t_R _20545_ (.A(_05283_),
    .B(_05371_),
    .Y(_18264_));
 INVx1_ASAP7_75t_R _20546_ (.A(_00190_),
    .Y(_18266_));
 INVx1_ASAP7_75t_R _20547_ (.A(_00192_),
    .Y(_17364_));
 OAI22x1_ASAP7_75t_R _20548_ (.A1(_05237_),
    .A2(_01728_),
    .B1(_05256_),
    .B2(_15836_),
    .Y(_17367_));
 INVx1_ASAP7_75t_R _20549_ (.A(_00196_),
    .Y(_17352_));
 INVx1_ASAP7_75t_R _20550_ (.A(_00197_),
    .Y(_17420_));
 INVx1_ASAP7_75t_R _20551_ (.A(_17772_),
    .Y(_17769_));
 INVx1_ASAP7_75t_R _20552_ (.A(_17774_),
    .Y(_17770_));
 INVx1_ASAP7_75t_R _20553_ (.A(_17807_),
    .Y(_17805_));
 INVx1_ASAP7_75t_R _20554_ (.A(_17842_),
    .Y(_17840_));
 INVx1_ASAP7_75t_R _20555_ (.A(_17874_),
    .Y(_17872_));
 INVx8_ASAP7_75t_R _20556_ (.A(_17564_),
    .Y(_17561_));
 INVx4_ASAP7_75t_R _20557_ (.A(_05460_),
    .Y(_05703_));
 BUFx6f_ASAP7_75t_R _20558_ (.A(_01762_),
    .Y(_05704_));
 NAND2x1_ASAP7_75t_R _20559_ (.A(_05172_),
    .B(_05704_),
    .Y(_05705_));
 AND2x4_ASAP7_75t_R _20560_ (.A(_05404_),
    .B(_05154_),
    .Y(_05706_));
 OR2x6_ASAP7_75t_R _20561_ (.A(_05705_),
    .B(_05706_),
    .Y(_05707_));
 INVx5_ASAP7_75t_R _20562_ (.A(_02205_),
    .Y(_05708_));
 INVx2_ASAP7_75t_R _20563_ (.A(_02206_),
    .Y(_05709_));
 BUFx6f_ASAP7_75t_R _20564_ (.A(_00262_),
    .Y(_05710_));
 INVx5_ASAP7_75t_R _20565_ (.A(_05710_),
    .Y(_05711_));
 BUFx6f_ASAP7_75t_R _20566_ (.A(_05711_),
    .Y(_05712_));
 OA21x2_ASAP7_75t_R _20567_ (.A1(_05708_),
    .A2(_05709_),
    .B(_05712_),
    .Y(_05713_));
 INVx1_ASAP7_75t_R _20568_ (.A(_00261_),
    .Y(_05714_));
 AO221x1_ASAP7_75t_R _20569_ (.A1(_05156_),
    .A2(_05707_),
    .B1(_05713_),
    .B2(_05457_),
    .C(_05714_),
    .Y(_05715_));
 OR2x6_ASAP7_75t_R _20570_ (.A(_05703_),
    .B(_05715_),
    .Y(_05716_));
 INVx2_ASAP7_75t_R _20571_ (.A(_05716_),
    .Y(_05717_));
 BUFx12f_ASAP7_75t_R _20572_ (.A(_05717_),
    .Y(_18717_));
 AND3x1_ASAP7_75t_R _20573_ (.A(_02197_),
    .B(_05193_),
    .C(_05235_),
    .Y(_05718_));
 AOI21x1_ASAP7_75t_R _20574_ (.A1(_02195_),
    .A2(_05236_),
    .B(_05718_),
    .Y(_02333_));
 AND3x1_ASAP7_75t_R _20575_ (.A(_02195_),
    .B(_05193_),
    .C(_05242_),
    .Y(_05719_));
 AOI21x1_ASAP7_75t_R _20576_ (.A1(_02194_),
    .A2(_05236_),
    .B(_05719_),
    .Y(_02334_));
 AND2x4_ASAP7_75t_R _20577_ (.A(_13262_),
    .B(_15234_),
    .Y(_05720_));
 BUFx6f_ASAP7_75t_R _20578_ (.A(_05720_),
    .Y(_05721_));
 BUFx6f_ASAP7_75t_R _20579_ (.A(_05721_),
    .Y(_05722_));
 AO21x1_ASAP7_75t_R _20580_ (.A1(_05193_),
    .A2(_05722_),
    .B(_05559_),
    .Y(_05723_));
 OA21x2_ASAP7_75t_R _20581_ (.A1(_05247_),
    .A2(_05206_),
    .B(_05723_),
    .Y(_02335_));
 BUFx6f_ASAP7_75t_R _20582_ (.A(_05200_),
    .Y(_05724_));
 NAND2x1_ASAP7_75t_R _20583_ (.A(_05203_),
    .B(_05204_),
    .Y(_05725_));
 OA21x2_ASAP7_75t_R _20584_ (.A1(_05724_),
    .A2(_05204_),
    .B(_05725_),
    .Y(_02336_));
 AND3x1_ASAP7_75t_R _20585_ (.A(_02199_),
    .B(_05193_),
    .C(_05722_),
    .Y(_05726_));
 AOI21x1_ASAP7_75t_R _20586_ (.A1(_02192_),
    .A2(_05206_),
    .B(_05726_),
    .Y(_02337_));
 INVx1_ASAP7_75t_R _20587_ (.A(_02191_),
    .Y(_05727_));
 BUFx6f_ASAP7_75t_R _20588_ (.A(_01444_),
    .Y(_05728_));
 INVx1_ASAP7_75t_R _20589_ (.A(_05728_),
    .Y(_05729_));
 NOR2x2_ASAP7_75t_R _20590_ (.A(_14265_),
    .B(_14134_),
    .Y(_05730_));
 AND5x2_ASAP7_75t_R _20591_ (.A(_00375_),
    .B(_13235_),
    .C(_05730_),
    .D(_04987_),
    .E(_05191_),
    .Y(_05731_));
 AND3x1_ASAP7_75t_R _20592_ (.A(_05180_),
    .B(_05728_),
    .C(_05731_),
    .Y(_05732_));
 AO21x1_ASAP7_75t_R _20593_ (.A1(_00375_),
    .A2(_05729_),
    .B(_05732_),
    .Y(_05733_));
 NAND2x1_ASAP7_75t_R _20594_ (.A(net26),
    .B(_05733_),
    .Y(_05734_));
 BUFx6f_ASAP7_75t_R _20595_ (.A(_05734_),
    .Y(_05735_));
 INVx2_ASAP7_75t_R _20596_ (.A(_05734_),
    .Y(_05736_));
 AND3x1_ASAP7_75t_R _20597_ (.A(_14602_),
    .B(_05730_),
    .C(_05736_),
    .Y(_05737_));
 AO21x1_ASAP7_75t_R _20598_ (.A1(_05727_),
    .A2(_05735_),
    .B(_05737_),
    .Y(_02338_));
 INVx2_ASAP7_75t_R _20599_ (.A(_02196_),
    .Y(_05738_));
 OR3x2_ASAP7_75t_R _20600_ (.A(_14274_),
    .B(_14117_),
    .C(_14135_),
    .Y(_05739_));
 NOR2x1_ASAP7_75t_R _20601_ (.A(_05735_),
    .B(_05739_),
    .Y(_05740_));
 AO21x1_ASAP7_75t_R _20602_ (.A1(_05738_),
    .A2(_05735_),
    .B(_05740_),
    .Y(_02339_));
 AO211x2_ASAP7_75t_R _20603_ (.A1(_14261_),
    .A2(_14271_),
    .B(_18580_),
    .C(_14144_),
    .Y(_05741_));
 AO221x1_ASAP7_75t_R _20604_ (.A1(_13839_),
    .A2(_05099_),
    .B1(_05100_),
    .B2(_13969_),
    .C(_05067_),
    .Y(_05742_));
 OA21x2_ASAP7_75t_R _20605_ (.A1(_13449_),
    .A2(_13543_),
    .B(_05701_),
    .Y(_05743_));
 BUFx6f_ASAP7_75t_R _20606_ (.A(_05743_),
    .Y(_05744_));
 OR5x2_ASAP7_75t_R _20607_ (.A(_18573_),
    .B(_05104_),
    .C(_05741_),
    .D(_05742_),
    .E(_05744_),
    .Y(_05745_));
 BUFx6f_ASAP7_75t_R _20608_ (.A(_05745_),
    .Y(_05746_));
 BUFx6f_ASAP7_75t_R _20609_ (.A(_05746_),
    .Y(_05747_));
 AND5x2_ASAP7_75t_R _20610_ (.A(_02228_),
    .B(_05702_),
    .C(_05027_),
    .D(_05151_),
    .E(_05191_),
    .Y(_05748_));
 NAND2x2_ASAP7_75t_R _20611_ (.A(_05148_),
    .B(_05748_),
    .Y(_05749_));
 BUFx6f_ASAP7_75t_R _20612_ (.A(_01396_),
    .Y(_05750_));
 OA21x2_ASAP7_75t_R _20613_ (.A1(_05747_),
    .A2(_05749_),
    .B(_05750_),
    .Y(_05751_));
 OR3x2_ASAP7_75t_R _20614_ (.A(_18563_),
    .B(_18568_),
    .C(_18573_),
    .Y(_05752_));
 OAI21x1_ASAP7_75t_R _20615_ (.A1(_05054_),
    .A2(_05752_),
    .B(_05702_),
    .Y(_05753_));
 BUFx6f_ASAP7_75t_R _20616_ (.A(_05070_),
    .Y(_05754_));
 AO21x1_ASAP7_75t_R _20617_ (.A1(_18575_),
    .A2(_18580_),
    .B(_14144_),
    .Y(_05755_));
 AO32x2_ASAP7_75t_R _20618_ (.A1(_18575_),
    .A2(_18580_),
    .A3(_05072_),
    .B1(_05076_),
    .B2(_05755_),
    .Y(_05756_));
 AND2x2_ASAP7_75t_R _20619_ (.A(_13449_),
    .B(_13543_),
    .Y(_05757_));
 NOR3x1_ASAP7_75t_R _20620_ (.A(_13449_),
    .B(_13543_),
    .C(_18565_),
    .Y(_05758_));
 AND2x2_ASAP7_75t_R _20621_ (.A(_18570_),
    .B(_05701_),
    .Y(_05759_));
 OAI21x1_ASAP7_75t_R _20622_ (.A1(_05757_),
    .A2(_05758_),
    .B(_05759_),
    .Y(_05760_));
 AOI22x1_ASAP7_75t_R _20623_ (.A1(_05082_),
    .A2(_05756_),
    .B1(_05760_),
    .B2(_05110_),
    .Y(_05761_));
 NAND2x2_ASAP7_75t_R _20624_ (.A(_05095_),
    .B(_05761_),
    .Y(_05762_));
 BUFx6f_ASAP7_75t_R _20625_ (.A(_05762_),
    .Y(_05763_));
 INVx2_ASAP7_75t_R _20626_ (.A(_02164_),
    .Y(_05764_));
 AO221x1_ASAP7_75t_R _20627_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .A2(_05754_),
    .B1(_05763_),
    .B2(_05764_),
    .C(_05102_),
    .Y(_05765_));
 AND3x4_ASAP7_75t_R _20628_ (.A(_13451_),
    .B(_18559_),
    .C(_05701_),
    .Y(_05766_));
 NAND2x2_ASAP7_75t_R _20629_ (.A(_05701_),
    .B(_05752_),
    .Y(_05767_));
 AND2x6_ASAP7_75t_R _20630_ (.A(_05766_),
    .B(_05767_),
    .Y(_05768_));
 NAND2x2_ASAP7_75t_R _20631_ (.A(_05058_),
    .B(_05069_),
    .Y(_05769_));
 INVx2_ASAP7_75t_R _20632_ (.A(_05763_),
    .Y(_05770_));
 OAI22x1_ASAP7_75t_R _20633_ (.A1(_00748_),
    .A2(_05769_),
    .B1(_05770_),
    .B2(_02101_),
    .Y(_05771_));
 INVx1_ASAP7_75t_R _20634_ (.A(net83),
    .Y(_05772_));
 NAND2x2_ASAP7_75t_R _20635_ (.A(_05123_),
    .B(_05120_),
    .Y(_05773_));
 BUFx6f_ASAP7_75t_R _20636_ (.A(_05773_),
    .Y(_05774_));
 AND2x6_ASAP7_75t_R _20637_ (.A(_13614_),
    .B(_18570_),
    .Y(_05775_));
 AO21x1_ASAP7_75t_R _20638_ (.A1(_05775_),
    .A2(_05076_),
    .B(_14144_),
    .Y(_05776_));
 BUFx6f_ASAP7_75t_R _20639_ (.A(_05776_),
    .Y(_05777_));
 NAND2x2_ASAP7_75t_R _20640_ (.A(_05133_),
    .B(_05777_),
    .Y(_05778_));
 BUFx6f_ASAP7_75t_R _20641_ (.A(_05778_),
    .Y(_05779_));
 AND2x6_ASAP7_75t_R _20642_ (.A(_04993_),
    .B(_05072_),
    .Y(_05780_));
 NAND2x2_ASAP7_75t_R _20643_ (.A(_05134_),
    .B(_05780_),
    .Y(_05781_));
 BUFx6f_ASAP7_75t_R _20644_ (.A(_05781_),
    .Y(_05782_));
 OA222x2_ASAP7_75t_R _20645_ (.A1(_05772_),
    .A2(_05774_),
    .B1(_05779_),
    .B2(_01906_),
    .C1(_05782_),
    .C2(_01994_),
    .Y(_05783_));
 NAND2x2_ASAP7_75t_R _20646_ (.A(_05133_),
    .B(_05780_),
    .Y(_05784_));
 BUFx6f_ASAP7_75t_R _20647_ (.A(_05784_),
    .Y(_05785_));
 NAND2x2_ASAP7_75t_R _20648_ (.A(_05121_),
    .B(_05137_),
    .Y(_05786_));
 OA21x2_ASAP7_75t_R _20649_ (.A1(_01831_),
    .A2(_05785_),
    .B(_05786_),
    .Y(_05787_));
 OA211x2_ASAP7_75t_R _20650_ (.A1(_05750_),
    .A2(_05747_),
    .B(_05783_),
    .C(_05787_),
    .Y(_05788_));
 NAND3x2_ASAP7_75t_R _20651_ (.B(_05136_),
    .C(_05133_),
    .Y(_05789_),
    .A(_05775_));
 BUFx6f_ASAP7_75t_R _20652_ (.A(_05789_),
    .Y(_05790_));
 BUFx6f_ASAP7_75t_R _20653_ (.A(_05790_),
    .Y(_05791_));
 NAND2x1_ASAP7_75t_R _20654_ (.A(_18573_),
    .B(_05071_),
    .Y(_05792_));
 AND2x2_ASAP7_75t_R _20655_ (.A(_04995_),
    .B(_05003_),
    .Y(_05793_));
 OR5x2_ASAP7_75t_R _20656_ (.A(_18580_),
    .B(_18608_),
    .C(_05093_),
    .D(_05792_),
    .E(_05793_),
    .Y(_05794_));
 NAND2x1_ASAP7_75t_R _20657_ (.A(_18565_),
    .B(_18570_),
    .Y(_05795_));
 OA21x2_ASAP7_75t_R _20658_ (.A1(_05795_),
    .A2(_05054_),
    .B(_05702_),
    .Y(_05796_));
 OR3x1_ASAP7_75t_R _20659_ (.A(_02061_),
    .B(_05794_),
    .C(_05796_),
    .Y(_05797_));
 NAND2x2_ASAP7_75t_R _20660_ (.A(_13451_),
    .B(_05130_),
    .Y(_05798_));
 OR3x2_ASAP7_75t_R _20661_ (.A(_05104_),
    .B(_05794_),
    .C(_05798_),
    .Y(_05799_));
 BUFx6f_ASAP7_75t_R _20662_ (.A(_05799_),
    .Y(_05800_));
 NAND3x2_ASAP7_75t_R _20663_ (.B(_05133_),
    .C(_05766_),
    .Y(_05801_),
    .A(_04993_));
 OA22x2_ASAP7_75t_R _20664_ (.A1(_02026_),
    .A2(_05800_),
    .B1(_05801_),
    .B2(_01962_),
    .Y(_05802_));
 OA211x2_ASAP7_75t_R _20665_ (.A1(_01956_),
    .A2(_05791_),
    .B(_05797_),
    .C(_05802_),
    .Y(_05803_));
 NAND2x1_ASAP7_75t_R _20666_ (.A(_05788_),
    .B(_05803_),
    .Y(_05804_));
 AO221x1_ASAP7_75t_R _20667_ (.A1(_05753_),
    .A2(_05765_),
    .B1(_05768_),
    .B2(_05771_),
    .C(_05804_),
    .Y(_05805_));
 BUFx6f_ASAP7_75t_R _20668_ (.A(_02225_),
    .Y(_05806_));
 AND3x1_ASAP7_75t_R _20669_ (.A(_14280_),
    .B(_14390_),
    .C(_14444_),
    .Y(_05807_));
 AO21x1_ASAP7_75t_R _20670_ (.A1(_02227_),
    .A2(_18556_),
    .B(_05807_),
    .Y(_05808_));
 NAND2x1_ASAP7_75t_R _20671_ (.A(_05806_),
    .B(_05808_),
    .Y(_05809_));
 OA21x2_ASAP7_75t_R _20672_ (.A1(_18554_),
    .A2(_05805_),
    .B(_05809_),
    .Y(_05810_));
 BUFx12f_ASAP7_75t_R _20673_ (.A(_05810_),
    .Y(_05811_));
 NOR3x1_ASAP7_75t_R _20674_ (.A(_05747_),
    .B(_05749_),
    .C(_05811_),
    .Y(_05812_));
 NOR2x1_ASAP7_75t_R _20675_ (.A(_05751_),
    .B(_05812_),
    .Y(_02340_));
 OA21x2_ASAP7_75t_R _20676_ (.A1(_05747_),
    .A2(_05749_),
    .B(_02189_),
    .Y(_05813_));
 BUFx12f_ASAP7_75t_R _20677_ (.A(_05767_),
    .Y(_05814_));
 BUFx6f_ASAP7_75t_R _20678_ (.A(_05130_),
    .Y(_05815_));
 BUFx6f_ASAP7_75t_R _20679_ (.A(_05815_),
    .Y(_05816_));
 INVx1_ASAP7_75t_R _20680_ (.A(_02104_),
    .Y(_05817_));
 INVx1_ASAP7_75t_R _20681_ (.A(_02099_),
    .Y(_05818_));
 AO221x1_ASAP7_75t_R _20682_ (.A1(_05817_),
    .A2(_05070_),
    .B1(_05762_),
    .B2(_05818_),
    .C(_05102_),
    .Y(_05819_));
 INVx1_ASAP7_75t_R _20683_ (.A(_02167_),
    .Y(_05820_));
 BUFx6f_ASAP7_75t_R _20684_ (.A(_05058_),
    .Y(_05821_));
 BUFx3_ASAP7_75t_R _20685_ (.A(_05069_),
    .Y(_05822_));
 BUFx6f_ASAP7_75t_R _20686_ (.A(_02162_),
    .Y(_05823_));
 INVx1_ASAP7_75t_R _20687_ (.A(_05823_),
    .Y(_05824_));
 AO32x1_ASAP7_75t_R _20688_ (.A1(_05820_),
    .A2(_05821_),
    .A3(_05822_),
    .B1(_05762_),
    .B2(_05824_),
    .Y(_05825_));
 BUFx6f_ASAP7_75t_R _20689_ (.A(_05138_),
    .Y(_05826_));
 BUFx6f_ASAP7_75t_R _20690_ (.A(_05826_),
    .Y(_05827_));
 AO32x1_ASAP7_75t_R _20691_ (.A1(_18553_),
    .A2(_05816_),
    .A3(_05819_),
    .B1(_05825_),
    .B2(_05827_),
    .Y(_05828_));
 BUFx6f_ASAP7_75t_R _20692_ (.A(_13451_),
    .Y(_05829_));
 OR5x2_ASAP7_75t_R _20693_ (.A(_05829_),
    .B(_18559_),
    .C(_14144_),
    .D(_05795_),
    .E(_05794_),
    .Y(_05830_));
 BUFx6f_ASAP7_75t_R _20694_ (.A(_05830_),
    .Y(_05831_));
 OA22x2_ASAP7_75t_R _20695_ (.A1(_01934_),
    .A2(_05790_),
    .B1(_05831_),
    .B2(_02032_),
    .Y(_05832_));
 AND3x1_ASAP7_75t_R _20696_ (.A(_05403_),
    .B(_05134_),
    .C(_05777_),
    .Y(_05833_));
 AOI21x1_ASAP7_75t_R _20697_ (.A1(_05775_),
    .A2(_05137_),
    .B(_05833_),
    .Y(_05834_));
 INVx1_ASAP7_75t_R _20698_ (.A(net105),
    .Y(_05835_));
 BUFx6f_ASAP7_75t_R _20699_ (.A(_05778_),
    .Y(_05836_));
 BUFx6f_ASAP7_75t_R _20700_ (.A(_05781_),
    .Y(_05837_));
 OA222x2_ASAP7_75t_R _20701_ (.A1(_05835_),
    .A2(_05774_),
    .B1(_05836_),
    .B2(_01884_),
    .C1(_05837_),
    .C2(_01972_),
    .Y(_05838_));
 BUFx6f_ASAP7_75t_R _20702_ (.A(_05784_),
    .Y(_05839_));
 BUFx6f_ASAP7_75t_R _20703_ (.A(_05799_),
    .Y(_05840_));
 OA222x2_ASAP7_75t_R _20704_ (.A1(_01809_),
    .A2(_05839_),
    .B1(_05840_),
    .B2(_02004_),
    .C1(_05801_),
    .C2(_01960_),
    .Y(_05841_));
 AND4x1_ASAP7_75t_R _20705_ (.A(_05832_),
    .B(_05834_),
    .C(_05838_),
    .D(_05841_),
    .Y(_05842_));
 OAI21x1_ASAP7_75t_R _20706_ (.A1(_02189_),
    .A2(_05747_),
    .B(_05842_),
    .Y(_05843_));
 AO21x2_ASAP7_75t_R _20707_ (.A1(_05814_),
    .A2(_05828_),
    .B(_05843_),
    .Y(_05844_));
 BUFx12f_ASAP7_75t_R _20708_ (.A(_05806_),
    .Y(_05845_));
 BUFx6f_ASAP7_75t_R _20709_ (.A(_02227_),
    .Y(_05846_));
 AND2x2_ASAP7_75t_R _20710_ (.A(_14280_),
    .B(_18562_),
    .Y(_05847_));
 AO21x1_ASAP7_75t_R _20711_ (.A1(_05846_),
    .A2(_18564_),
    .B(_05847_),
    .Y(_05848_));
 NAND2x1_ASAP7_75t_R _20712_ (.A(_05845_),
    .B(_05848_),
    .Y(_05849_));
 OA21x2_ASAP7_75t_R _20713_ (.A1(_18562_),
    .A2(_05844_),
    .B(_05849_),
    .Y(_05850_));
 BUFx12f_ASAP7_75t_R _20714_ (.A(_05850_),
    .Y(_05851_));
 NOR3x1_ASAP7_75t_R _20715_ (.A(_05747_),
    .B(_05749_),
    .C(_05851_),
    .Y(_05852_));
 NOR2x1_ASAP7_75t_R _20716_ (.A(_05813_),
    .B(_05852_),
    .Y(_02341_));
 INVx2_ASAP7_75t_R _20717_ (.A(_05750_),
    .Y(_05853_));
 AND3x1_ASAP7_75t_R _20718_ (.A(_13448_),
    .B(_13542_),
    .C(_18568_),
    .Y(_05854_));
 AOI211x1_ASAP7_75t_R _20719_ (.A1(_13448_),
    .A2(_13543_),
    .B(_18568_),
    .C(_18573_),
    .Y(_05855_));
 OAI22x1_ASAP7_75t_R _20720_ (.A1(_13449_),
    .A2(_13543_),
    .B1(_14143_),
    .B2(_05044_),
    .Y(_05856_));
 OA31x2_ASAP7_75t_R _20721_ (.A1(_05854_),
    .A2(_05855_),
    .A3(_05856_),
    .B1(_05056_),
    .Y(_05857_));
 NAND2x1_ASAP7_75t_R _20722_ (.A(_18565_),
    .B(_05071_),
    .Y(_05858_));
 AOI211x1_ASAP7_75t_R _20723_ (.A1(_05028_),
    .A2(_05045_),
    .B(_05046_),
    .C(_05858_),
    .Y(_05859_));
 AO21x1_ASAP7_75t_R _20724_ (.A1(_05007_),
    .A2(_05008_),
    .B(_05067_),
    .Y(_05860_));
 AND3x1_ASAP7_75t_R _20725_ (.A(_18563_),
    .B(_05071_),
    .C(_05050_),
    .Y(_05861_));
 OR3x1_ASAP7_75t_R _20726_ (.A(_14143_),
    .B(_05860_),
    .C(_05861_),
    .Y(_05862_));
 AOI21x1_ASAP7_75t_R _20727_ (.A1(_05857_),
    .A2(_05859_),
    .B(_05862_),
    .Y(_05863_));
 AND3x1_ASAP7_75t_R _20728_ (.A(_05079_),
    .B(_05009_),
    .C(_05081_),
    .Y(_05864_));
 OR3x1_ASAP7_75t_R _20729_ (.A(_18573_),
    .B(_14143_),
    .C(_05775_),
    .Y(_05865_));
 AND2x2_ASAP7_75t_R _20730_ (.A(_13836_),
    .B(_05006_),
    .Y(_05866_));
 AND5x2_ASAP7_75t_R _20731_ (.A(_13769_),
    .B(_18583_),
    .C(_05127_),
    .D(_05131_),
    .E(_05866_),
    .Y(_05867_));
 NAND2x1_ASAP7_75t_R _20732_ (.A(_13448_),
    .B(_18563_),
    .Y(_05868_));
 AO21x1_ASAP7_75t_R _20733_ (.A1(_05142_),
    .A2(_05868_),
    .B(_14143_),
    .Y(_05869_));
 XNOR2x2_ASAP7_75t_R _20734_ (.A(_13448_),
    .B(_13612_),
    .Y(_05870_));
 AND4x1_ASAP7_75t_R _20735_ (.A(_05112_),
    .B(_05113_),
    .C(_05142_),
    .D(_05870_),
    .Y(_05871_));
 AO221x1_ASAP7_75t_R _20736_ (.A1(_05864_),
    .A2(_05865_),
    .B1(_05867_),
    .B2(_05869_),
    .C(_05871_),
    .Y(_05872_));
 OR2x2_ASAP7_75t_R _20737_ (.A(_13768_),
    .B(_05097_),
    .Y(_05873_));
 NAND2x1_ASAP7_75t_R _20738_ (.A(_13839_),
    .B(_05099_),
    .Y(_05874_));
 AND5x1_ASAP7_75t_R _20739_ (.A(_18578_),
    .B(_05006_),
    .C(_05007_),
    .D(_05008_),
    .E(_05874_),
    .Y(_05875_));
 AND2x2_ASAP7_75t_R _20740_ (.A(_13768_),
    .B(_05006_),
    .Y(_05876_));
 AND2x2_ASAP7_75t_R _20741_ (.A(_05044_),
    .B(_05115_),
    .Y(_05877_));
 AO32x1_ASAP7_75t_R _20742_ (.A1(_05876_),
    .A2(_05119_),
    .A3(_05877_),
    .B1(_05112_),
    .B2(_05113_),
    .Y(_05878_));
 AND2x2_ASAP7_75t_R _20743_ (.A(_05088_),
    .B(_05071_),
    .Y(_05879_));
 AO33x2_ASAP7_75t_R _20744_ (.A1(_05081_),
    .A2(_05873_),
    .A3(_05875_),
    .B1(_05758_),
    .B2(_05878_),
    .B3(_05879_),
    .Y(_05880_));
 OR4x1_ASAP7_75t_R _20745_ (.A(_18578_),
    .B(_14143_),
    .C(_05093_),
    .D(_05860_),
    .Y(_05881_));
 AOI21x1_ASAP7_75t_R _20746_ (.A1(_05087_),
    .A2(_05092_),
    .B(_05881_),
    .Y(_05882_));
 AND2x2_ASAP7_75t_R _20747_ (.A(_05076_),
    .B(_05106_),
    .Y(_05883_));
 OR5x2_ASAP7_75t_R _20748_ (.A(_13769_),
    .B(_18578_),
    .C(_14143_),
    .D(_05093_),
    .E(_05860_),
    .Y(_05884_));
 NOR3x1_ASAP7_75t_R _20749_ (.A(_05107_),
    .B(_05883_),
    .C(_05884_),
    .Y(_05885_));
 OR5x1_ASAP7_75t_R _20750_ (.A(_05863_),
    .B(_05872_),
    .C(_05880_),
    .D(_05882_),
    .E(_05885_),
    .Y(_05886_));
 AND4x1_ASAP7_75t_R _20751_ (.A(_13769_),
    .B(_18583_),
    .C(_05127_),
    .D(_05866_),
    .Y(_05887_));
 AND3x1_ASAP7_75t_R _20752_ (.A(_05004_),
    .B(_05009_),
    .C(_05025_),
    .Y(_05888_));
 AO221x1_ASAP7_75t_R _20753_ (.A1(_05126_),
    .A2(_05887_),
    .B1(_05867_),
    .B2(_05130_),
    .C(_05888_),
    .Y(_05889_));
 AND5x1_ASAP7_75t_R _20754_ (.A(_18568_),
    .B(_05701_),
    .C(_18608_),
    .D(_05079_),
    .E(_05081_),
    .Y(_05890_));
 AO21x1_ASAP7_75t_R _20755_ (.A1(_05072_),
    .A2(_05073_),
    .B(_05077_),
    .Y(_05891_));
 AND3x1_ASAP7_75t_R _20756_ (.A(_05112_),
    .B(_05138_),
    .C(_05875_),
    .Y(_05892_));
 OA21x2_ASAP7_75t_R _20757_ (.A1(_05137_),
    .A2(_05892_),
    .B(_04993_),
    .Y(_05893_));
 AO221x1_ASAP7_75t_R _20758_ (.A1(_04993_),
    .A2(_05889_),
    .B1(_05890_),
    .B2(_05891_),
    .C(_05893_),
    .Y(_05894_));
 AND5x1_ASAP7_75t_R _20759_ (.A(_02228_),
    .B(_05701_),
    .C(_05027_),
    .D(_05151_),
    .E(_05191_),
    .Y(_05895_));
 OA21x2_ASAP7_75t_R _20760_ (.A1(_05886_),
    .A2(_05894_),
    .B(_05895_),
    .Y(_05896_));
 BUFx12f_ASAP7_75t_R _20761_ (.A(_05896_),
    .Y(_05897_));
 OR2x2_ASAP7_75t_R _20762_ (.A(_05757_),
    .B(_05758_),
    .Y(_05898_));
 AOI21x1_ASAP7_75t_R _20763_ (.A1(_05879_),
    .A2(_05898_),
    .B(_05884_),
    .Y(_05899_));
 AO21x2_ASAP7_75t_R _20764_ (.A1(_05890_),
    .A2(_05756_),
    .B(_05899_),
    .Y(_05900_));
 OR3x2_ASAP7_75t_R _20765_ (.A(_05863_),
    .B(_05882_),
    .C(_05900_),
    .Y(_05901_));
 NAND3x2_ASAP7_75t_R _20766_ (.B(_05753_),
    .C(_05901_),
    .Y(_05902_),
    .A(_05897_));
 NAND2x1_ASAP7_75t_R _20767_ (.A(_05082_),
    .B(_05756_),
    .Y(_05903_));
 OR5x1_ASAP7_75t_R _20768_ (.A(_18578_),
    .B(_18610_),
    .C(_05093_),
    .D(_05792_),
    .E(_05067_),
    .Y(_05904_));
 AO21x1_ASAP7_75t_R _20769_ (.A1(_05759_),
    .A2(_05898_),
    .B(_05904_),
    .Y(_05905_));
 AND3x4_ASAP7_75t_R _20770_ (.A(_05095_),
    .B(_05903_),
    .C(_05905_),
    .Y(_05906_));
 BUFx6f_ASAP7_75t_R _20771_ (.A(_05906_),
    .Y(_05907_));
 OA21x2_ASAP7_75t_R _20772_ (.A1(_05078_),
    .A2(_05083_),
    .B(_05095_),
    .Y(_05908_));
 AND3x1_ASAP7_75t_R _20773_ (.A(_05009_),
    .B(_05081_),
    .C(_05101_),
    .Y(_05909_));
 AOI22x1_ASAP7_75t_R _20774_ (.A1(_05098_),
    .A2(_05909_),
    .B1(_05864_),
    .B2(_05105_),
    .Y(_05910_));
 AND5x2_ASAP7_75t_R _20775_ (.A(_18575_),
    .B(_05701_),
    .C(_05007_),
    .D(_05008_),
    .E(_05081_),
    .Y(_05911_));
 AND2x6_ASAP7_75t_R _20776_ (.A(_05044_),
    .B(_05911_),
    .Y(_05912_));
 AND3x1_ASAP7_75t_R _20777_ (.A(_05044_),
    .B(_05116_),
    .C(_05119_),
    .Y(_05913_));
 OAI21x1_ASAP7_75t_R _20778_ (.A1(_05912_),
    .A2(_05913_),
    .B(_05123_),
    .Y(_05914_));
 OR3x1_ASAP7_75t_R _20779_ (.A(_05107_),
    .B(_05883_),
    .C(_05904_),
    .Y(_05915_));
 AND3x4_ASAP7_75t_R _20780_ (.A(_05044_),
    .B(_05136_),
    .C(_05911_),
    .Y(_05916_));
 AND5x1_ASAP7_75t_R _20781_ (.A(_18575_),
    .B(_05009_),
    .C(_05081_),
    .D(_05101_),
    .E(_05138_),
    .Y(_05917_));
 OAI21x1_ASAP7_75t_R _20782_ (.A1(_05916_),
    .A2(_05917_),
    .B(_04993_),
    .Y(_05918_));
 OR5x1_ASAP7_75t_R _20783_ (.A(_18580_),
    .B(_18608_),
    .C(_05093_),
    .D(_05792_),
    .E(_05793_),
    .Y(_05919_));
 NAND2x1_ASAP7_75t_R _20784_ (.A(_18575_),
    .B(_18580_),
    .Y(_05920_));
 NAND2x1_ASAP7_75t_R _20785_ (.A(_18559_),
    .B(_05701_),
    .Y(_05921_));
 NAND2x1_ASAP7_75t_R _20786_ (.A(_18590_),
    .B(_05081_),
    .Y(_05922_));
 AO211x2_ASAP7_75t_R _20787_ (.A1(_14261_),
    .A2(_14271_),
    .B(_18585_),
    .C(_14144_),
    .Y(_05923_));
 OR4x1_ASAP7_75t_R _20788_ (.A(_05920_),
    .B(_05921_),
    .C(_05922_),
    .D(_05923_),
    .Y(_05924_));
 OR5x1_ASAP7_75t_R _20789_ (.A(_18559_),
    .B(_18590_),
    .C(_05793_),
    .D(_05920_),
    .E(_05923_),
    .Y(_05925_));
 AO32x1_ASAP7_75t_R _20790_ (.A1(_05919_),
    .A2(_05924_),
    .A3(_05925_),
    .B1(_05795_),
    .B2(_05702_),
    .Y(_05926_));
 AND5x1_ASAP7_75t_R _20791_ (.A(_05910_),
    .B(_05914_),
    .C(_05915_),
    .D(_05918_),
    .E(_05926_),
    .Y(_05927_));
 AND4x1_ASAP7_75t_R _20792_ (.A(_18583_),
    .B(_05701_),
    .C(_05007_),
    .D(_05008_),
    .Y(_05928_));
 AO33x2_ASAP7_75t_R _20793_ (.A1(_18565_),
    .A2(_05044_),
    .A3(_05911_),
    .B1(_05928_),
    .B2(_05073_),
    .B3(_05131_),
    .Y(_05929_));
 BUFx6f_ASAP7_75t_R _20794_ (.A(_13450_),
    .Y(_05930_));
 AND2x2_ASAP7_75t_R _20795_ (.A(_05930_),
    .B(_18563_),
    .Y(_05931_));
 AND4x1_ASAP7_75t_R _20796_ (.A(_18565_),
    .B(_05073_),
    .C(_05131_),
    .D(_05928_),
    .Y(_05932_));
 AO221x1_ASAP7_75t_R _20797_ (.A1(_13453_),
    .A2(_05929_),
    .B1(_05931_),
    .B2(_05912_),
    .C(_05932_),
    .Y(_05933_));
 AOI22x1_ASAP7_75t_R _20798_ (.A1(_05058_),
    .A2(_05069_),
    .B1(_05142_),
    .B2(_05933_),
    .Y(_05934_));
 OR2x2_ASAP7_75t_R _20799_ (.A(_04990_),
    .B(_05026_),
    .Y(_05935_));
 OR5x2_ASAP7_75t_R _20800_ (.A(_05150_),
    .B(_14144_),
    .C(_05935_),
    .D(_05119_),
    .E(_05159_),
    .Y(_05936_));
 AO31x2_ASAP7_75t_R _20801_ (.A1(_05908_),
    .A2(_05927_),
    .A3(_05934_),
    .B(_05936_),
    .Y(_05937_));
 AND2x4_ASAP7_75t_R _20802_ (.A(_05769_),
    .B(_05906_),
    .Y(_05938_));
 NOR2x2_ASAP7_75t_R _20803_ (.A(_05937_),
    .B(_05938_),
    .Y(_05939_));
 NAND2x2_ASAP7_75t_R _20804_ (.A(_05753_),
    .B(_05939_),
    .Y(_05940_));
 NOR2x2_ASAP7_75t_R _20805_ (.A(_05907_),
    .B(_05940_),
    .Y(_05941_));
 BUFx6f_ASAP7_75t_R _20806_ (.A(_05941_),
    .Y(_05942_));
 AO21x1_ASAP7_75t_R _20807_ (.A1(_05853_),
    .A2(_05902_),
    .B(_05942_),
    .Y(_05943_));
 AND3x4_ASAP7_75t_R _20808_ (.A(_05753_),
    .B(_05907_),
    .C(_05939_),
    .Y(_05944_));
 BUFx3_ASAP7_75t_R _20809_ (.A(_05944_),
    .Y(_05945_));
 AO32x1_ASAP7_75t_R _20810_ (.A1(_00747_),
    .A2(_05750_),
    .A3(_05940_),
    .B1(_05945_),
    .B2(_05811_),
    .Y(_05946_));
 AO21x1_ASAP7_75t_R _20811_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .A2(_05943_),
    .B(_05946_),
    .Y(_02342_));
 INVx1_ASAP7_75t_R _20812_ (.A(_02188_),
    .Y(_05947_));
 BUFx6f_ASAP7_75t_R _20813_ (.A(_05940_),
    .Y(_05948_));
 OR4x1_ASAP7_75t_R _20814_ (.A(_02134_),
    .B(_02145_),
    .C(_02156_),
    .D(_02167_),
    .Y(_05949_));
 OR3x2_ASAP7_75t_R _20815_ (.A(_05853_),
    .B(_02234_),
    .C(_05949_),
    .Y(_05950_));
 OR3x1_ASAP7_75t_R _20816_ (.A(_02127_),
    .B(_02128_),
    .C(_02129_),
    .Y(_05951_));
 BUFx6f_ASAP7_75t_R _20817_ (.A(_05951_),
    .Y(_05952_));
 OR3x1_ASAP7_75t_R _20818_ (.A(_02126_),
    .B(_05950_),
    .C(_05952_),
    .Y(_05953_));
 BUFx6f_ASAP7_75t_R _20819_ (.A(_05941_),
    .Y(_05954_));
 AO21x1_ASAP7_75t_R _20820_ (.A1(_05948_),
    .A2(_05953_),
    .B(_05954_),
    .Y(_05955_));
 NOR2x1_ASAP7_75t_R _20821_ (.A(_02126_),
    .B(_05952_),
    .Y(_05956_));
 INVx1_ASAP7_75t_R _20822_ (.A(_05950_),
    .Y(_05957_));
 AND2x6_ASAP7_75t_R _20823_ (.A(_05902_),
    .B(_05957_),
    .Y(_05958_));
 BUFx12f_ASAP7_75t_R _20824_ (.A(_05806_),
    .Y(_05959_));
 BUFx6f_ASAP7_75t_R _20825_ (.A(_02227_),
    .Y(_05960_));
 AND3x1_ASAP7_75t_R _20826_ (.A(_18074_),
    .B(_15228_),
    .C(_15230_),
    .Y(_05961_));
 AO21x1_ASAP7_75t_R _20827_ (.A1(_05960_),
    .A2(_18604_),
    .B(_05961_),
    .Y(_05962_));
 AND2x6_ASAP7_75t_R _20828_ (.A(_05702_),
    .B(_05752_),
    .Y(_05963_));
 BUFx12f_ASAP7_75t_R _20829_ (.A(_05744_),
    .Y(_05964_));
 BUFx12f_ASAP7_75t_R _20830_ (.A(_05798_),
    .Y(_05965_));
 BUFx6f_ASAP7_75t_R _20831_ (.A(_05965_),
    .Y(_05966_));
 OAI22x1_ASAP7_75t_R _20832_ (.A1(_02188_),
    .A2(_05964_),
    .B1(_05966_),
    .B2(_02125_),
    .Y(_05967_));
 INVx1_ASAP7_75t_R _20833_ (.A(_02090_),
    .Y(_05968_));
 INVx1_ASAP7_75t_R _20834_ (.A(_02153_),
    .Y(_05969_));
 AO32x2_ASAP7_75t_R _20835_ (.A1(_05968_),
    .A2(_18553_),
    .A3(_05816_),
    .B1(_05827_),
    .B2(_05969_),
    .Y(_05970_));
 BUFx6f_ASAP7_75t_R _20836_ (.A(_05763_),
    .Y(_05971_));
 AOI22x1_ASAP7_75t_R _20837_ (.A1(_05754_),
    .A2(_05967_),
    .B1(_05970_),
    .B2(_05971_),
    .Y(_05972_));
 OA222x2_ASAP7_75t_R _20838_ (.A1(_01905_),
    .A2(_05779_),
    .B1(_05800_),
    .B2(_02025_),
    .C1(_05831_),
    .C2(_02052_),
    .Y(_05973_));
 INVx1_ASAP7_75t_R _20839_ (.A(net84),
    .Y(_05974_));
 BUFx6f_ASAP7_75t_R _20840_ (.A(_05773_),
    .Y(_05975_));
 OA21x2_ASAP7_75t_R _20841_ (.A1(_01993_),
    .A2(_05781_),
    .B(_05745_),
    .Y(_05976_));
 OA22x2_ASAP7_75t_R _20842_ (.A1(_01830_),
    .A2(_05784_),
    .B1(_05789_),
    .B2(_01955_),
    .Y(_05977_));
 OA211x2_ASAP7_75t_R _20843_ (.A1(_05974_),
    .A2(_05975_),
    .B(_05976_),
    .C(_05977_),
    .Y(_05978_));
 OA211x2_ASAP7_75t_R _20844_ (.A1(_01405_),
    .A2(_05786_),
    .B(_05973_),
    .C(_05978_),
    .Y(_05979_));
 OA21x2_ASAP7_75t_R _20845_ (.A1(_05963_),
    .A2(_05972_),
    .B(_05979_),
    .Y(_05980_));
 AOI22x1_ASAP7_75t_R _20846_ (.A1(_05959_),
    .A2(_05962_),
    .B1(_05980_),
    .B2(_18604_),
    .Y(_05981_));
 AO32x1_ASAP7_75t_R _20847_ (.A1(_02188_),
    .A2(_05956_),
    .A3(_05958_),
    .B1(_05945_),
    .B2(_05981_),
    .Y(_05982_));
 AO21x1_ASAP7_75t_R _20848_ (.A1(_05947_),
    .A2(_05955_),
    .B(_05982_),
    .Y(_02343_));
 INVx1_ASAP7_75t_R _20849_ (.A(_02187_),
    .Y(_05983_));
 OR4x1_ASAP7_75t_R _20850_ (.A(_00747_),
    .B(_05853_),
    .C(_02178_),
    .D(_05949_),
    .Y(_05984_));
 OR4x1_ASAP7_75t_R _20851_ (.A(_02126_),
    .B(_02188_),
    .C(_05952_),
    .D(_05984_),
    .Y(_05985_));
 AO21x1_ASAP7_75t_R _20852_ (.A1(_05948_),
    .A2(_05985_),
    .B(_05954_),
    .Y(_05986_));
 BUFx6f_ASAP7_75t_R _20853_ (.A(_05940_),
    .Y(_05987_));
 INVx1_ASAP7_75t_R _20854_ (.A(_05985_),
    .Y(_05988_));
 BUFx6f_ASAP7_75t_R _20855_ (.A(_14280_),
    .Y(_05989_));
 AND3x1_ASAP7_75t_R _20856_ (.A(_05989_),
    .B(_14378_),
    .C(_14387_),
    .Y(_05990_));
 AO21x1_ASAP7_75t_R _20857_ (.A1(_05846_),
    .A2(_18609_),
    .B(_05990_),
    .Y(_05991_));
 BUFx12f_ASAP7_75t_R _20858_ (.A(_05767_),
    .Y(_05992_));
 INVx2_ASAP7_75t_R _20859_ (.A(_02124_),
    .Y(_05993_));
 BUFx3_ASAP7_75t_R _20860_ (.A(_13453_),
    .Y(_05994_));
 BUFx6f_ASAP7_75t_R _20861_ (.A(_05130_),
    .Y(_05995_));
 BUFx6f_ASAP7_75t_R _20862_ (.A(_05138_),
    .Y(_05996_));
 AO32x1_ASAP7_75t_R _20863_ (.A1(_05993_),
    .A2(_05994_),
    .A3(_05995_),
    .B1(_05996_),
    .B2(_05983_),
    .Y(_05997_));
 BUFx6f_ASAP7_75t_R _20864_ (.A(_02152_),
    .Y(_05998_));
 BUFx12f_ASAP7_75t_R _20865_ (.A(_05744_),
    .Y(_05999_));
 OAI22x1_ASAP7_75t_R _20866_ (.A1(_05998_),
    .A2(_05999_),
    .B1(_05965_),
    .B2(_02089_),
    .Y(_06000_));
 BUFx3_ASAP7_75t_R _20867_ (.A(_05762_),
    .Y(_06001_));
 AO32x1_ASAP7_75t_R _20868_ (.A1(_05821_),
    .A2(_05822_),
    .A3(_05997_),
    .B1(_06000_),
    .B2(_06001_),
    .Y(_06002_));
 NAND2x1_ASAP7_75t_R _20869_ (.A(_05992_),
    .B(_06002_),
    .Y(_06003_));
 BUFx6f_ASAP7_75t_R _20870_ (.A(_05839_),
    .Y(_06004_));
 BUFx6f_ASAP7_75t_R _20871_ (.A(_05840_),
    .Y(_06005_));
 NAND2x2_ASAP7_75t_R _20872_ (.A(_05123_),
    .B(_05114_),
    .Y(_06006_));
 BUFx6f_ASAP7_75t_R _20873_ (.A(_06006_),
    .Y(_06007_));
 OA222x2_ASAP7_75t_R _20874_ (.A1(_01829_),
    .A2(_06004_),
    .B1(_06005_),
    .B2(_02024_),
    .C1(_06007_),
    .C2(_01918_),
    .Y(_06008_));
 BUFx6f_ASAP7_75t_R _20875_ (.A(_05830_),
    .Y(_06009_));
 BUFx6f_ASAP7_75t_R _20876_ (.A(_06009_),
    .Y(_06010_));
 OR5x1_ASAP7_75t_R _20877_ (.A(_13449_),
    .B(_13543_),
    .C(_18565_),
    .D(_18568_),
    .E(_14144_),
    .Y(_06011_));
 OR3x1_ASAP7_75t_R _20878_ (.A(_18573_),
    .B(_18578_),
    .C(_18585_),
    .Y(_06012_));
 OR5x2_ASAP7_75t_R _20879_ (.A(_14144_),
    .B(_18608_),
    .C(_06011_),
    .D(_06012_),
    .E(_05922_),
    .Y(_06013_));
 BUFx6f_ASAP7_75t_R _20880_ (.A(_06013_),
    .Y(_06014_));
 BUFx6f_ASAP7_75t_R _20881_ (.A(_06014_),
    .Y(_06015_));
 OA222x2_ASAP7_75t_R _20882_ (.A1(_01954_),
    .A2(_05790_),
    .B1(_06010_),
    .B2(_02051_),
    .C1(_06015_),
    .C2(_05444_),
    .Y(_06016_));
 INVx1_ASAP7_75t_R _20883_ (.A(net85),
    .Y(_06017_));
 NAND2x2_ASAP7_75t_R _20884_ (.A(_05114_),
    .B(_05777_),
    .Y(_06018_));
 OA222x2_ASAP7_75t_R _20885_ (.A1(_06017_),
    .A2(_05773_),
    .B1(_05837_),
    .B2(_01992_),
    .C1(_06018_),
    .C2(_00331_),
    .Y(_06019_));
 NAND2x2_ASAP7_75t_R _20886_ (.A(_05134_),
    .B(_05777_),
    .Y(_06020_));
 OA22x2_ASAP7_75t_R _20887_ (.A1(_01904_),
    .A2(_05779_),
    .B1(_06020_),
    .B2(_02060_),
    .Y(_06021_));
 OA211x2_ASAP7_75t_R _20888_ (.A1(_00746_),
    .A2(_05786_),
    .B(_06019_),
    .C(_06021_),
    .Y(_06022_));
 AND5x2_ASAP7_75t_R _20889_ (.A(_05747_),
    .B(_06003_),
    .C(_06008_),
    .D(_06016_),
    .E(_06022_),
    .Y(_06023_));
 AOI22x1_ASAP7_75t_R _20890_ (.A1(_05845_),
    .A2(_05991_),
    .B1(_06023_),
    .B2(_18609_),
    .Y(_06024_));
 BUFx12f_ASAP7_75t_R _20891_ (.A(_06024_),
    .Y(_06025_));
 BUFx6f_ASAP7_75t_R _20892_ (.A(_05944_),
    .Y(_06026_));
 AO32x1_ASAP7_75t_R _20893_ (.A1(_02187_),
    .A2(_05987_),
    .A3(_05988_),
    .B1(_06025_),
    .B2(_06026_),
    .Y(_06027_));
 AO21x1_ASAP7_75t_R _20894_ (.A1(_05983_),
    .A2(_05986_),
    .B(_06027_),
    .Y(_02344_));
 INVx1_ASAP7_75t_R _20895_ (.A(_02186_),
    .Y(_06028_));
 OR3x2_ASAP7_75t_R _20896_ (.A(_02126_),
    .B(_02187_),
    .C(_02188_),
    .Y(_06029_));
 OR3x1_ASAP7_75t_R _20897_ (.A(_05950_),
    .B(_05952_),
    .C(_06029_),
    .Y(_06030_));
 AO21x1_ASAP7_75t_R _20898_ (.A1(_05948_),
    .A2(_06030_),
    .B(_05954_),
    .Y(_06031_));
 NOR2x1_ASAP7_75t_R _20899_ (.A(_05952_),
    .B(_06029_),
    .Y(_06032_));
 AND3x1_ASAP7_75t_R _20900_ (.A(_13269_),
    .B(_13293_),
    .C(_05989_),
    .Y(_06033_));
 AO21x1_ASAP7_75t_R _20901_ (.A1(_05846_),
    .A2(_18613_),
    .B(_06033_),
    .Y(_06034_));
 OAI22x1_ASAP7_75t_R _20902_ (.A1(_02186_),
    .A2(_05964_),
    .B1(_05966_),
    .B2(_02123_),
    .Y(_06035_));
 INVx1_ASAP7_75t_R _20903_ (.A(_02088_),
    .Y(_06036_));
 INVx2_ASAP7_75t_R _20904_ (.A(_02151_),
    .Y(_06037_));
 AO32x2_ASAP7_75t_R _20905_ (.A1(_06036_),
    .A2(_18553_),
    .A3(_05816_),
    .B1(_05827_),
    .B2(_06037_),
    .Y(_06038_));
 AOI22x1_ASAP7_75t_R _20906_ (.A1(_05754_),
    .A2(_06035_),
    .B1(_06038_),
    .B2(_05971_),
    .Y(_06039_));
 BUFx6f_ASAP7_75t_R _20907_ (.A(_05786_),
    .Y(_06040_));
 OA21x2_ASAP7_75t_R _20908_ (.A1(_00745_),
    .A2(_06040_),
    .B(_05140_),
    .Y(_06041_));
 OA22x2_ASAP7_75t_R _20909_ (.A1(_02023_),
    .A2(_06005_),
    .B1(_06018_),
    .B2(_00332_),
    .Y(_06042_));
 OA22x2_ASAP7_75t_R _20910_ (.A1(_01953_),
    .A2(_05791_),
    .B1(_06010_),
    .B2(_02050_),
    .Y(_06043_));
 INVx1_ASAP7_75t_R _20911_ (.A(net86),
    .Y(_06044_));
 BUFx6f_ASAP7_75t_R _20912_ (.A(_05781_),
    .Y(_06045_));
 OA222x2_ASAP7_75t_R _20913_ (.A1(_06044_),
    .A2(_05975_),
    .B1(_06045_),
    .B2(_01991_),
    .C1(_06020_),
    .C2(_02059_),
    .Y(_06046_));
 BUFx6f_ASAP7_75t_R _20914_ (.A(_05836_),
    .Y(_06047_));
 OA22x2_ASAP7_75t_R _20915_ (.A1(_01903_),
    .A2(_06047_),
    .B1(_06004_),
    .B2(_01828_),
    .Y(_06048_));
 AND4x1_ASAP7_75t_R _20916_ (.A(_06042_),
    .B(_06043_),
    .C(_06046_),
    .D(_06048_),
    .Y(_06049_));
 OA211x2_ASAP7_75t_R _20917_ (.A1(_05963_),
    .A2(_06039_),
    .B(_06041_),
    .C(_06049_),
    .Y(_06050_));
 AOI22x1_ASAP7_75t_R _20918_ (.A1(_05845_),
    .A2(_06034_),
    .B1(_06050_),
    .B2(_18613_),
    .Y(_06051_));
 BUFx12f_ASAP7_75t_R _20919_ (.A(_06051_),
    .Y(_06052_));
 AO32x1_ASAP7_75t_R _20920_ (.A1(_02186_),
    .A2(_05958_),
    .A3(_06032_),
    .B1(_06052_),
    .B2(_06026_),
    .Y(_06053_));
 AO21x1_ASAP7_75t_R _20921_ (.A1(_06028_),
    .A2(_06031_),
    .B(_06053_),
    .Y(_02345_));
 INVx1_ASAP7_75t_R _20922_ (.A(_02185_),
    .Y(_06054_));
 OR3x1_ASAP7_75t_R _20923_ (.A(_02186_),
    .B(_05952_),
    .C(_06029_),
    .Y(_06055_));
 OR2x2_ASAP7_75t_R _20924_ (.A(_05984_),
    .B(_06055_),
    .Y(_06056_));
 AO21x1_ASAP7_75t_R _20925_ (.A1(_05948_),
    .A2(_06056_),
    .B(_05954_),
    .Y(_06057_));
 BUFx12f_ASAP7_75t_R _20926_ (.A(_05806_),
    .Y(_06058_));
 BUFx6f_ASAP7_75t_R _20927_ (.A(_02227_),
    .Y(_06059_));
 BUFx6f_ASAP7_75t_R _20928_ (.A(_14280_),
    .Y(_06060_));
 AND3x1_ASAP7_75t_R _20929_ (.A(_06060_),
    .B(_15430_),
    .C(_15432_),
    .Y(_06061_));
 AO21x1_ASAP7_75t_R _20930_ (.A1(_06059_),
    .A2(_18618_),
    .B(_06061_),
    .Y(_06062_));
 BUFx6f_ASAP7_75t_R _20931_ (.A(_05058_),
    .Y(_06063_));
 BUFx3_ASAP7_75t_R _20932_ (.A(_05069_),
    .Y(_06064_));
 INVx2_ASAP7_75t_R _20933_ (.A(_02122_),
    .Y(_06065_));
 BUFx6f_ASAP7_75t_R _20934_ (.A(_05995_),
    .Y(_06066_));
 BUFx6f_ASAP7_75t_R _20935_ (.A(_05996_),
    .Y(_06067_));
 AO32x1_ASAP7_75t_R _20936_ (.A1(_06065_),
    .A2(_13454_),
    .A3(_06066_),
    .B1(_06067_),
    .B2(_06054_),
    .Y(_06068_));
 INVx1_ASAP7_75t_R _20937_ (.A(_02087_),
    .Y(_06069_));
 INVx2_ASAP7_75t_R _20938_ (.A(_02150_),
    .Y(_06070_));
 AO32x1_ASAP7_75t_R _20939_ (.A1(_06069_),
    .A2(_13454_),
    .A3(_05815_),
    .B1(_05826_),
    .B2(_06070_),
    .Y(_06071_));
 AO32x1_ASAP7_75t_R _20940_ (.A1(_06063_),
    .A2(_06064_),
    .A3(_06068_),
    .B1(_06071_),
    .B2(_05763_),
    .Y(_06072_));
 NAND2x1_ASAP7_75t_R _20941_ (.A(_05814_),
    .B(_06072_),
    .Y(_06073_));
 OA222x2_ASAP7_75t_R _20942_ (.A1(_01902_),
    .A2(_05836_),
    .B1(_06020_),
    .B2(_02058_),
    .C1(_05830_),
    .C2(_02049_),
    .Y(_06074_));
 OA21x2_ASAP7_75t_R _20943_ (.A1(_01827_),
    .A2(_05785_),
    .B(_06074_),
    .Y(_06075_));
 OA21x2_ASAP7_75t_R _20944_ (.A1(_01990_),
    .A2(_06045_),
    .B(_05746_),
    .Y(_06076_));
 AND2x6_ASAP7_75t_R _20945_ (.A(_05123_),
    .B(_05120_),
    .Y(_06077_));
 NAND2x1_ASAP7_75t_R _20946_ (.A(net87),
    .B(_06077_),
    .Y(_06078_));
 OA22x2_ASAP7_75t_R _20947_ (.A1(_02022_),
    .A2(_05800_),
    .B1(_05790_),
    .B2(_01952_),
    .Y(_06079_));
 AND4x1_ASAP7_75t_R _20948_ (.A(_06075_),
    .B(_06076_),
    .C(_06078_),
    .D(_06079_),
    .Y(_06080_));
 OA211x2_ASAP7_75t_R _20949_ (.A1(_01406_),
    .A2(_06040_),
    .B(_06073_),
    .C(_06080_),
    .Y(_06081_));
 AOI22x1_ASAP7_75t_R _20950_ (.A1(_06058_),
    .A2(_06062_),
    .B1(_06081_),
    .B2(_18618_),
    .Y(_06082_));
 AO21x2_ASAP7_75t_R _20951_ (.A1(_05753_),
    .A2(_05939_),
    .B(_05984_),
    .Y(_06083_));
 OR3x1_ASAP7_75t_R _20952_ (.A(_06054_),
    .B(_06055_),
    .C(_06083_),
    .Y(_06084_));
 INVx1_ASAP7_75t_R _20953_ (.A(_06084_),
    .Y(_06085_));
 AO21x1_ASAP7_75t_R _20954_ (.A1(_06026_),
    .A2(_06082_),
    .B(_06085_),
    .Y(_06086_));
 AO21x1_ASAP7_75t_R _20955_ (.A1(_06054_),
    .A2(_06057_),
    .B(_06086_),
    .Y(_02346_));
 INVx1_ASAP7_75t_R _20956_ (.A(_02184_),
    .Y(_06087_));
 OR4x1_ASAP7_75t_R _20957_ (.A(_02185_),
    .B(_02186_),
    .C(_05952_),
    .D(_06029_),
    .Y(_06088_));
 BUFx6f_ASAP7_75t_R _20958_ (.A(_06088_),
    .Y(_06089_));
 OR2x2_ASAP7_75t_R _20959_ (.A(_05950_),
    .B(_06089_),
    .Y(_06090_));
 AO21x1_ASAP7_75t_R _20960_ (.A1(_05948_),
    .A2(_06090_),
    .B(_05954_),
    .Y(_06091_));
 INVx2_ASAP7_75t_R _20961_ (.A(_06089_),
    .Y(_06092_));
 AND2x2_ASAP7_75t_R _20962_ (.A(_18074_),
    .B(_18625_),
    .Y(_06093_));
 AO21x1_ASAP7_75t_R _20963_ (.A1(_05960_),
    .A2(_18623_),
    .B(_06093_),
    .Y(_06094_));
 BUFx6f_ASAP7_75t_R _20964_ (.A(_05786_),
    .Y(_06095_));
 INVx1_ASAP7_75t_R _20965_ (.A(_02121_),
    .Y(_06096_));
 AO32x1_ASAP7_75t_R _20966_ (.A1(_06096_),
    .A2(_05994_),
    .A3(_05995_),
    .B1(_05996_),
    .B2(_06087_),
    .Y(_06097_));
 OAI22x1_ASAP7_75t_R _20967_ (.A1(_02149_),
    .A2(_05999_),
    .B1(_05798_),
    .B2(_02086_),
    .Y(_06098_));
 AO32x1_ASAP7_75t_R _20968_ (.A1(_05821_),
    .A2(_05822_),
    .A3(_06097_),
    .B1(_06098_),
    .B2(_05762_),
    .Y(_06099_));
 NAND2x1_ASAP7_75t_R _20969_ (.A(_05992_),
    .B(_06099_),
    .Y(_06100_));
 OA222x2_ASAP7_75t_R _20970_ (.A1(_01901_),
    .A2(_05836_),
    .B1(_05840_),
    .B2(_02021_),
    .C1(_06009_),
    .C2(_02048_),
    .Y(_06101_));
 OA21x2_ASAP7_75t_R _20971_ (.A1(_01989_),
    .A2(_05782_),
    .B(_05746_),
    .Y(_06102_));
 NAND2x1_ASAP7_75t_R _20972_ (.A(net88),
    .B(_06077_),
    .Y(_06103_));
 BUFx6f_ASAP7_75t_R _20973_ (.A(_05789_),
    .Y(_06104_));
 OA22x2_ASAP7_75t_R _20974_ (.A1(_01826_),
    .A2(_05785_),
    .B1(_06104_),
    .B2(_01951_),
    .Y(_06105_));
 AND4x1_ASAP7_75t_R _20975_ (.A(_06101_),
    .B(_06102_),
    .C(_06103_),
    .D(_06105_),
    .Y(_06106_));
 OA211x2_ASAP7_75t_R _20976_ (.A1(_01407_),
    .A2(_06095_),
    .B(_06100_),
    .C(_06106_),
    .Y(_06107_));
 AOI22x1_ASAP7_75t_R _20977_ (.A1(_05959_),
    .A2(_06094_),
    .B1(_06107_),
    .B2(_18623_),
    .Y(_06108_));
 AO32x1_ASAP7_75t_R _20978_ (.A1(_02184_),
    .A2(_05958_),
    .A3(_06092_),
    .B1(_06108_),
    .B2(_06026_),
    .Y(_06109_));
 AO21x1_ASAP7_75t_R _20979_ (.A1(_06087_),
    .A2(_06091_),
    .B(_06109_),
    .Y(_02347_));
 INVx1_ASAP7_75t_R _20980_ (.A(_02183_),
    .Y(_06110_));
 OR3x1_ASAP7_75t_R _20981_ (.A(_02184_),
    .B(_05984_),
    .C(_06089_),
    .Y(_06111_));
 AO21x1_ASAP7_75t_R _20982_ (.A1(_05948_),
    .A2(_06111_),
    .B(_05954_),
    .Y(_06112_));
 OR2x2_ASAP7_75t_R _20983_ (.A(_05984_),
    .B(_06089_),
    .Y(_06113_));
 NOR2x1_ASAP7_75t_R _20984_ (.A(_02184_),
    .B(_06113_),
    .Y(_06114_));
 AND2x2_ASAP7_75t_R _20985_ (.A(_06060_),
    .B(_18630_),
    .Y(_06115_));
 AO21x1_ASAP7_75t_R _20986_ (.A1(_06059_),
    .A2(_18628_),
    .B(_06115_),
    .Y(_06116_));
 OAI22x1_ASAP7_75t_R _20987_ (.A1(_02183_),
    .A2(_05964_),
    .B1(_05966_),
    .B2(_02120_),
    .Y(_06117_));
 INVx1_ASAP7_75t_R _20988_ (.A(_02085_),
    .Y(_06118_));
 BUFx6f_ASAP7_75t_R _20989_ (.A(_13453_),
    .Y(_06119_));
 INVx1_ASAP7_75t_R _20990_ (.A(_02148_),
    .Y(_06120_));
 AO32x1_ASAP7_75t_R _20991_ (.A1(_06118_),
    .A2(_06119_),
    .A3(_05816_),
    .B1(_05827_),
    .B2(_06120_),
    .Y(_06121_));
 AO32x1_ASAP7_75t_R _20992_ (.A1(_06063_),
    .A2(_06064_),
    .A3(_06117_),
    .B1(_06121_),
    .B2(_05971_),
    .Y(_06122_));
 NAND2x1_ASAP7_75t_R _20993_ (.A(_05814_),
    .B(_06122_),
    .Y(_06123_));
 OA222x2_ASAP7_75t_R _20994_ (.A1(_01900_),
    .A2(_06047_),
    .B1(_06020_),
    .B2(_02057_),
    .C1(_06010_),
    .C2(_02047_),
    .Y(_06124_));
 INVx1_ASAP7_75t_R _20995_ (.A(net89),
    .Y(_06125_));
 OA21x2_ASAP7_75t_R _20996_ (.A1(_01988_),
    .A2(_05782_),
    .B(_05746_),
    .Y(_06126_));
 OA22x2_ASAP7_75t_R _20997_ (.A1(_02020_),
    .A2(_05800_),
    .B1(_05790_),
    .B2(_01950_),
    .Y(_06127_));
 OA211x2_ASAP7_75t_R _20998_ (.A1(_06125_),
    .A2(_05975_),
    .B(_06126_),
    .C(_06127_),
    .Y(_06128_));
 OA211x2_ASAP7_75t_R _20999_ (.A1(_01825_),
    .A2(_06004_),
    .B(_06124_),
    .C(_06128_),
    .Y(_06129_));
 OA211x2_ASAP7_75t_R _21000_ (.A1(_01408_),
    .A2(_06040_),
    .B(_06123_),
    .C(_06129_),
    .Y(_06130_));
 AOI22x1_ASAP7_75t_R _21001_ (.A1(_06058_),
    .A2(_06116_),
    .B1(_06130_),
    .B2(_18628_),
    .Y(_06131_));
 AO32x1_ASAP7_75t_R _21002_ (.A1(_02183_),
    .A2(_05987_),
    .A3(_06114_),
    .B1(_06131_),
    .B2(_06026_),
    .Y(_06132_));
 AO21x1_ASAP7_75t_R _21003_ (.A1(_06110_),
    .A2(_06112_),
    .B(_06132_),
    .Y(_02348_));
 OR3x2_ASAP7_75t_R _21004_ (.A(_05882_),
    .B(_05900_),
    .C(_05902_),
    .Y(_06133_));
 BUFx6f_ASAP7_75t_R _21005_ (.A(_06133_),
    .Y(_06134_));
 NAND2x2_ASAP7_75t_R _21006_ (.A(_05958_),
    .B(_06092_),
    .Y(_06135_));
 OR3x1_ASAP7_75t_R _21007_ (.A(_02183_),
    .B(_02184_),
    .C(_06135_),
    .Y(_06136_));
 AND3x1_ASAP7_75t_R _21008_ (.A(_02182_),
    .B(_06134_),
    .C(_06136_),
    .Y(_06137_));
 AND2x2_ASAP7_75t_R _21009_ (.A(_05989_),
    .B(_18635_),
    .Y(_06138_));
 AO21x1_ASAP7_75t_R _21010_ (.A1(_05846_),
    .A2(_18633_),
    .B(_06138_),
    .Y(_06139_));
 BUFx6f_ASAP7_75t_R _21011_ (.A(_05745_),
    .Y(_06140_));
 OA222x2_ASAP7_75t_R _21012_ (.A1(_02019_),
    .A2(_05840_),
    .B1(_06104_),
    .B2(_01949_),
    .C1(_05430_),
    .C2(_06015_),
    .Y(_06141_));
 INVx1_ASAP7_75t_R _21013_ (.A(net90),
    .Y(_06142_));
 OA222x2_ASAP7_75t_R _21014_ (.A1(_06142_),
    .A2(_05774_),
    .B1(_05782_),
    .B2(_01987_),
    .C1(_06007_),
    .C2(_01924_),
    .Y(_06143_));
 OA222x2_ASAP7_75t_R _21015_ (.A1(_01899_),
    .A2(_05779_),
    .B1(_06009_),
    .B2(_02046_),
    .C1(_05839_),
    .C2(_01824_),
    .Y(_06144_));
 AND4x1_ASAP7_75t_R _21016_ (.A(_06140_),
    .B(_06141_),
    .C(_06143_),
    .D(_06144_),
    .Y(_06145_));
 OAI22x1_ASAP7_75t_R _21017_ (.A1(_02182_),
    .A2(_05999_),
    .B1(_05965_),
    .B2(_02119_),
    .Y(_06146_));
 INVx1_ASAP7_75t_R _21018_ (.A(_02084_),
    .Y(_06147_));
 INVx2_ASAP7_75t_R _21019_ (.A(_02147_),
    .Y(_06148_));
 AO32x1_ASAP7_75t_R _21020_ (.A1(_06147_),
    .A2(_13454_),
    .A3(_05815_),
    .B1(_05826_),
    .B2(_06148_),
    .Y(_06149_));
 AO32x1_ASAP7_75t_R _21021_ (.A1(_05821_),
    .A2(_05822_),
    .A3(_06146_),
    .B1(_06149_),
    .B2(_06001_),
    .Y(_06150_));
 NAND2x1_ASAP7_75t_R _21022_ (.A(_05992_),
    .B(_06150_),
    .Y(_06151_));
 OA211x2_ASAP7_75t_R _21023_ (.A1(_01409_),
    .A2(_06040_),
    .B(_06145_),
    .C(_06151_),
    .Y(_06152_));
 AOI22x1_ASAP7_75t_R _21024_ (.A1(_05845_),
    .A2(_06139_),
    .B1(_06152_),
    .B2(_18633_),
    .Y(_06153_));
 OR3x2_ASAP7_75t_R _21025_ (.A(_02182_),
    .B(_02183_),
    .C(_02184_),
    .Y(_06154_));
 OAI22x1_ASAP7_75t_R _21026_ (.A1(_06134_),
    .A2(_06153_),
    .B1(_06154_),
    .B2(_06135_),
    .Y(_06155_));
 NOR2x1_ASAP7_75t_R _21027_ (.A(_06137_),
    .B(_06155_),
    .Y(_02349_));
 INVx1_ASAP7_75t_R _21028_ (.A(_02181_),
    .Y(_06156_));
 OR3x1_ASAP7_75t_R _21029_ (.A(_05984_),
    .B(_06089_),
    .C(_06154_),
    .Y(_06157_));
 AO21x1_ASAP7_75t_R _21030_ (.A1(_05948_),
    .A2(_06157_),
    .B(_05954_),
    .Y(_06158_));
 BUFx6f_ASAP7_75t_R _21031_ (.A(_05940_),
    .Y(_06159_));
 INVx1_ASAP7_75t_R _21032_ (.A(_06157_),
    .Y(_06160_));
 AND3x1_ASAP7_75t_R _21033_ (.A(_05989_),
    .B(_15944_),
    .C(_15946_),
    .Y(_06161_));
 AO21x1_ASAP7_75t_R _21034_ (.A1(_05846_),
    .A2(_18638_),
    .B(_06161_),
    .Y(_06162_));
 INVx1_ASAP7_75t_R _21035_ (.A(_02118_),
    .Y(_06163_));
 AO32x2_ASAP7_75t_R _21036_ (.A1(_06163_),
    .A2(_13454_),
    .A3(_06066_),
    .B1(_06067_),
    .B2(_06156_),
    .Y(_06164_));
 INVx2_ASAP7_75t_R _21037_ (.A(_02083_),
    .Y(_06165_));
 INVx1_ASAP7_75t_R _21038_ (.A(_02146_),
    .Y(_06166_));
 AO32x1_ASAP7_75t_R _21039_ (.A1(_06165_),
    .A2(_06119_),
    .A3(_06066_),
    .B1(_06067_),
    .B2(_06166_),
    .Y(_06167_));
 AOI22x1_ASAP7_75t_R _21040_ (.A1(_05754_),
    .A2(_06164_),
    .B1(_06167_),
    .B2(_05763_),
    .Y(_06168_));
 OR2x2_ASAP7_75t_R _21041_ (.A(_01410_),
    .B(_05786_),
    .Y(_06169_));
 OA22x2_ASAP7_75t_R _21042_ (.A1(_02018_),
    .A2(_05799_),
    .B1(_06018_),
    .B2(_01832_),
    .Y(_06170_));
 OA22x2_ASAP7_75t_R _21043_ (.A1(_01823_),
    .A2(_05784_),
    .B1(_05830_),
    .B2(_02045_),
    .Y(_06171_));
 INVx1_ASAP7_75t_R _21044_ (.A(net91),
    .Y(_06172_));
 OA222x2_ASAP7_75t_R _21045_ (.A1(_06172_),
    .A2(_05773_),
    .B1(_05781_),
    .B2(_01986_),
    .C1(_06006_),
    .C2(_01915_),
    .Y(_06173_));
 OA21x2_ASAP7_75t_R _21046_ (.A1(_05429_),
    .A2(_06014_),
    .B(_05745_),
    .Y(_06174_));
 OA221x2_ASAP7_75t_R _21047_ (.A1(_01898_),
    .A2(_05778_),
    .B1(_05789_),
    .B2(_01948_),
    .C(_06174_),
    .Y(_06175_));
 AND5x2_ASAP7_75t_R _21048_ (.A(_06169_),
    .B(_06170_),
    .C(_06171_),
    .D(_06173_),
    .E(_06175_),
    .Y(_06176_));
 OA21x2_ASAP7_75t_R _21049_ (.A1(_05963_),
    .A2(_06168_),
    .B(_06176_),
    .Y(_06177_));
 AOI22x1_ASAP7_75t_R _21050_ (.A1(_05845_),
    .A2(_06162_),
    .B1(_06177_),
    .B2(_18638_),
    .Y(_06178_));
 BUFx12f_ASAP7_75t_R _21051_ (.A(_06178_),
    .Y(_06179_));
 AO32x1_ASAP7_75t_R _21052_ (.A1(_02181_),
    .A2(_06159_),
    .A3(_06160_),
    .B1(_06179_),
    .B2(_06026_),
    .Y(_06180_));
 AO21x1_ASAP7_75t_R _21053_ (.A1(_06156_),
    .A2(_06158_),
    .B(_06180_),
    .Y(_02350_));
 AND2x2_ASAP7_75t_R _21054_ (.A(_05989_),
    .B(_18645_),
    .Y(_06181_));
 AO21x1_ASAP7_75t_R _21055_ (.A1(_06059_),
    .A2(_18643_),
    .B(_06181_),
    .Y(_06182_));
 OA222x2_ASAP7_75t_R _21056_ (.A1(_02017_),
    .A2(_06005_),
    .B1(_05790_),
    .B2(_01947_),
    .C1(_05427_),
    .C2(_06015_),
    .Y(_06183_));
 INVx1_ASAP7_75t_R _21057_ (.A(net92),
    .Y(_06184_));
 OA222x2_ASAP7_75t_R _21058_ (.A1(_06184_),
    .A2(_05975_),
    .B1(_06045_),
    .B2(_01985_),
    .C1(_06007_),
    .C2(_01914_),
    .Y(_06185_));
 OA222x2_ASAP7_75t_R _21059_ (.A1(_01897_),
    .A2(_06047_),
    .B1(_05831_),
    .B2(_02044_),
    .C1(_06004_),
    .C2(_01822_),
    .Y(_06186_));
 AND4x1_ASAP7_75t_R _21060_ (.A(_05747_),
    .B(_06183_),
    .C(_06185_),
    .D(_06186_),
    .Y(_06187_));
 BUFx3_ASAP7_75t_R _21061_ (.A(_02117_),
    .Y(_06188_));
 OAI22x1_ASAP7_75t_R _21062_ (.A1(_02180_),
    .A2(_05964_),
    .B1(_05966_),
    .B2(_06188_),
    .Y(_06189_));
 INVx1_ASAP7_75t_R _21063_ (.A(_02081_),
    .Y(_06190_));
 INVx1_ASAP7_75t_R _21064_ (.A(_02144_),
    .Y(_06191_));
 AO32x1_ASAP7_75t_R _21065_ (.A1(_06190_),
    .A2(_06119_),
    .A3(_06066_),
    .B1(_06067_),
    .B2(_06191_),
    .Y(_06192_));
 AO32x1_ASAP7_75t_R _21066_ (.A1(_06063_),
    .A2(_06064_),
    .A3(_06189_),
    .B1(_06192_),
    .B2(_05763_),
    .Y(_06193_));
 NAND2x1_ASAP7_75t_R _21067_ (.A(_05814_),
    .B(_06193_),
    .Y(_06194_));
 OA211x2_ASAP7_75t_R _21068_ (.A1(_01411_),
    .A2(_06040_),
    .B(_06187_),
    .C(_06194_),
    .Y(_06195_));
 AOI22x1_ASAP7_75t_R _21069_ (.A1(_06058_),
    .A2(_06182_),
    .B1(_06195_),
    .B2(_18643_),
    .Y(_06196_));
 BUFx12f_ASAP7_75t_R _21070_ (.A(_06196_),
    .Y(_06197_));
 OR3x1_ASAP7_75t_R _21071_ (.A(_02181_),
    .B(_06135_),
    .C(_06154_),
    .Y(_06198_));
 OR2x2_ASAP7_75t_R _21072_ (.A(_02180_),
    .B(_06198_),
    .Y(_06199_));
 NAND3x1_ASAP7_75t_R _21073_ (.A(_02180_),
    .B(_06134_),
    .C(_06198_),
    .Y(_06200_));
 OA211x2_ASAP7_75t_R _21074_ (.A1(_06134_),
    .A2(_06197_),
    .B(_06199_),
    .C(_06200_),
    .Y(_02351_));
 INVx1_ASAP7_75t_R _21075_ (.A(_02179_),
    .Y(_06201_));
 OR3x1_ASAP7_75t_R _21076_ (.A(_02180_),
    .B(_02181_),
    .C(_06157_),
    .Y(_06202_));
 AO21x1_ASAP7_75t_R _21077_ (.A1(_05948_),
    .A2(_06202_),
    .B(_05954_),
    .Y(_06203_));
 INVx1_ASAP7_75t_R _21078_ (.A(_06202_),
    .Y(_06204_));
 AND3x1_ASAP7_75t_R _21079_ (.A(_18074_),
    .B(_16191_),
    .C(_16194_),
    .Y(_06205_));
 AO21x1_ASAP7_75t_R _21080_ (.A1(_05960_),
    .A2(_18648_),
    .B(_06205_),
    .Y(_06206_));
 OA222x2_ASAP7_75t_R _21081_ (.A1(_02016_),
    .A2(_05840_),
    .B1(_06104_),
    .B2(_01946_),
    .C1(_05426_),
    .C2(_06015_),
    .Y(_06207_));
 INVx1_ASAP7_75t_R _21082_ (.A(net93),
    .Y(_06208_));
 OA222x2_ASAP7_75t_R _21083_ (.A1(_06208_),
    .A2(_05774_),
    .B1(_05782_),
    .B2(_01984_),
    .C1(_06007_),
    .C2(_01913_),
    .Y(_06209_));
 OA222x2_ASAP7_75t_R _21084_ (.A1(_01896_),
    .A2(_05779_),
    .B1(_06009_),
    .B2(_02043_),
    .C1(_05839_),
    .C2(_01821_),
    .Y(_06210_));
 AND4x1_ASAP7_75t_R _21085_ (.A(_06140_),
    .B(_06207_),
    .C(_06209_),
    .D(_06210_),
    .Y(_06211_));
 OAI22x1_ASAP7_75t_R _21086_ (.A1(_02179_),
    .A2(_05999_),
    .B1(_05965_),
    .B2(_02116_),
    .Y(_06212_));
 INVx2_ASAP7_75t_R _21087_ (.A(_02080_),
    .Y(_06213_));
 INVx1_ASAP7_75t_R _21088_ (.A(_02143_),
    .Y(_06214_));
 AO32x1_ASAP7_75t_R _21089_ (.A1(_06213_),
    .A2(_13454_),
    .A3(_05815_),
    .B1(_05826_),
    .B2(_06214_),
    .Y(_06215_));
 AO32x1_ASAP7_75t_R _21090_ (.A1(_06063_),
    .A2(_06064_),
    .A3(_06212_),
    .B1(_06215_),
    .B2(_06001_),
    .Y(_06216_));
 NAND2x1_ASAP7_75t_R _21091_ (.A(_05992_),
    .B(_06216_),
    .Y(_06217_));
 OA211x2_ASAP7_75t_R _21092_ (.A1(_01412_),
    .A2(_06040_),
    .B(_06211_),
    .C(_06217_),
    .Y(_06218_));
 AOI22x1_ASAP7_75t_R _21093_ (.A1(_05959_),
    .A2(_06206_),
    .B1(_06218_),
    .B2(_18648_),
    .Y(_06219_));
 AO32x1_ASAP7_75t_R _21094_ (.A1(_02179_),
    .A2(_06159_),
    .A3(_06204_),
    .B1(_06219_),
    .B2(_06026_),
    .Y(_06220_));
 AO21x1_ASAP7_75t_R _21095_ (.A1(_06201_),
    .A2(_06203_),
    .B(_06220_),
    .Y(_02352_));
 INVx1_ASAP7_75t_R _21096_ (.A(net94),
    .Y(_06221_));
 OA222x2_ASAP7_75t_R _21097_ (.A1(_06221_),
    .A2(_05975_),
    .B1(_06047_),
    .B2(_01895_),
    .C1(_06045_),
    .C2(_01983_),
    .Y(_06222_));
 OA22x2_ASAP7_75t_R _21098_ (.A1(_01820_),
    .A2(_06004_),
    .B1(_05791_),
    .B2(_01945_),
    .Y(_06223_));
 OA22x2_ASAP7_75t_R _21099_ (.A1(_02015_),
    .A2(_06005_),
    .B1(_06020_),
    .B2(_02056_),
    .Y(_06224_));
 OA22x2_ASAP7_75t_R _21100_ (.A1(_01961_),
    .A2(_05801_),
    .B1(_06010_),
    .B2(_00749_),
    .Y(_06225_));
 AO32x1_ASAP7_75t_R _21101_ (.A1(\cs_registers_i.mhpmcounter[1857] ),
    .A2(_05994_),
    .A3(_05815_),
    .B1(_05826_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .Y(_06226_));
 BUFx6f_ASAP7_75t_R _21102_ (.A(_02163_),
    .Y(_06227_));
 OAI22x1_ASAP7_75t_R _21103_ (.A1(_06227_),
    .A2(_05999_),
    .B1(_05965_),
    .B2(_02100_),
    .Y(_06228_));
 AO32x1_ASAP7_75t_R _21104_ (.A1(_05821_),
    .A2(_05822_),
    .A3(_06226_),
    .B1(_06228_),
    .B2(_06001_),
    .Y(_06229_));
 NAND2x1_ASAP7_75t_R _21105_ (.A(_05992_),
    .B(_06229_),
    .Y(_06230_));
 AND5x2_ASAP7_75t_R _21106_ (.A(_06222_),
    .B(_06223_),
    .C(_06224_),
    .D(_06225_),
    .E(_06230_),
    .Y(_06231_));
 AND2x2_ASAP7_75t_R _21107_ (.A(_14280_),
    .B(_18558_),
    .Y(_06232_));
 AO21x1_ASAP7_75t_R _21108_ (.A1(_02227_),
    .A2(_18560_),
    .B(_06232_),
    .Y(_06233_));
 AND2x2_ASAP7_75t_R _21109_ (.A(_05806_),
    .B(_06233_),
    .Y(_06234_));
 AOI21x1_ASAP7_75t_R _21110_ (.A1(_18560_),
    .A2(_06231_),
    .B(_06234_),
    .Y(_06235_));
 INVx1_ASAP7_75t_R _21111_ (.A(_02235_),
    .Y(_06236_));
 AND3x1_ASAP7_75t_R _21112_ (.A(_05750_),
    .B(_06236_),
    .C(_05902_),
    .Y(_06237_));
 AO221x1_ASAP7_75t_R _21113_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .A2(_05943_),
    .B1(_06026_),
    .B2(_06235_),
    .C(_06237_),
    .Y(_02353_));
 AND3x1_ASAP7_75t_R _21114_ (.A(_18074_),
    .B(_16326_),
    .C(_16328_),
    .Y(_06238_));
 AO21x1_ASAP7_75t_R _21115_ (.A1(_05960_),
    .A2(_18653_),
    .B(_06238_),
    .Y(_06239_));
 OAI22x1_ASAP7_75t_R _21116_ (.A1(_02177_),
    .A2(_05964_),
    .B1(_05966_),
    .B2(_02114_),
    .Y(_06240_));
 INVx1_ASAP7_75t_R _21117_ (.A(_02079_),
    .Y(_06241_));
 INVx2_ASAP7_75t_R _21118_ (.A(_02142_),
    .Y(_06242_));
 AO32x2_ASAP7_75t_R _21119_ (.A1(_06241_),
    .A2(_18553_),
    .A3(_05816_),
    .B1(_05827_),
    .B2(_06242_),
    .Y(_06243_));
 AOI22x1_ASAP7_75t_R _21120_ (.A1(_05754_),
    .A2(_06240_),
    .B1(_06243_),
    .B2(_05971_),
    .Y(_06244_));
 OA222x2_ASAP7_75t_R _21121_ (.A1(_01894_),
    .A2(_06047_),
    .B1(_06010_),
    .B2(_02042_),
    .C1(_06015_),
    .C2(_05483_),
    .Y(_06245_));
 OA21x2_ASAP7_75t_R _21122_ (.A1(_01944_),
    .A2(_05791_),
    .B(_06245_),
    .Y(_06246_));
 INVx1_ASAP7_75t_R _21123_ (.A(_01413_),
    .Y(_06247_));
 AO32x1_ASAP7_75t_R _21124_ (.A1(_06247_),
    .A2(_05121_),
    .A3(_05136_),
    .B1(_05123_),
    .B2(_05421_),
    .Y(_06248_));
 AOI22x1_ASAP7_75t_R _21125_ (.A1(net95),
    .A2(_06077_),
    .B1(_06248_),
    .B2(_05114_),
    .Y(_06249_));
 OA21x2_ASAP7_75t_R _21126_ (.A1(_01982_),
    .A2(_06045_),
    .B(_06249_),
    .Y(_06250_));
 OA21x2_ASAP7_75t_R _21127_ (.A1(_02014_),
    .A2(_06005_),
    .B(_05140_),
    .Y(_06251_));
 OA211x2_ASAP7_75t_R _21128_ (.A1(_01819_),
    .A2(_06004_),
    .B(_06250_),
    .C(_06251_),
    .Y(_06252_));
 OA211x2_ASAP7_75t_R _21129_ (.A1(_05963_),
    .A2(_06244_),
    .B(_06246_),
    .C(_06252_),
    .Y(_06253_));
 AOI22x1_ASAP7_75t_R _21130_ (.A1(_05959_),
    .A2(_06239_),
    .B1(_06253_),
    .B2(_18653_),
    .Y(_06254_));
 BUFx12f_ASAP7_75t_R _21131_ (.A(_06254_),
    .Y(_06255_));
 OR5x1_ASAP7_75t_R _21132_ (.A(_02180_),
    .B(_02181_),
    .C(_02182_),
    .D(_02183_),
    .E(_02184_),
    .Y(_06256_));
 OR2x2_ASAP7_75t_R _21133_ (.A(_02179_),
    .B(_06256_),
    .Y(_06257_));
 OR3x1_ASAP7_75t_R _21134_ (.A(_02177_),
    .B(_06135_),
    .C(_06257_),
    .Y(_06258_));
 AND2x2_ASAP7_75t_R _21135_ (.A(_02177_),
    .B(_06133_),
    .Y(_06259_));
 OAI21x1_ASAP7_75t_R _21136_ (.A1(_06135_),
    .A2(_06257_),
    .B(_06259_),
    .Y(_06260_));
 OA211x2_ASAP7_75t_R _21137_ (.A1(_06134_),
    .A2(_06255_),
    .B(_06258_),
    .C(_06260_),
    .Y(_02354_));
 AND3x1_ASAP7_75t_R _21138_ (.A(_05989_),
    .B(_16449_),
    .C(_16451_),
    .Y(_06261_));
 AO21x1_ASAP7_75t_R _21139_ (.A1(_05846_),
    .A2(_18658_),
    .B(_06261_),
    .Y(_06262_));
 OA22x2_ASAP7_75t_R _21140_ (.A1(_02013_),
    .A2(_05800_),
    .B1(_06018_),
    .B2(_01833_),
    .Y(_06263_));
 OA22x2_ASAP7_75t_R _21141_ (.A1(_01818_),
    .A2(_05785_),
    .B1(_05831_),
    .B2(_02041_),
    .Y(_06264_));
 INVx1_ASAP7_75t_R _21142_ (.A(net96),
    .Y(_06265_));
 OA222x2_ASAP7_75t_R _21143_ (.A1(_06265_),
    .A2(_05774_),
    .B1(_05782_),
    .B2(_01981_),
    .C1(_06007_),
    .C2(_01911_),
    .Y(_06266_));
 INVx1_ASAP7_75t_R _21144_ (.A(net161),
    .Y(_06267_));
 OA22x2_ASAP7_75t_R _21145_ (.A1(_01893_),
    .A2(_05778_),
    .B1(_05789_),
    .B2(_01943_),
    .Y(_06268_));
 OA211x2_ASAP7_75t_R _21146_ (.A1(_06267_),
    .A2(_06015_),
    .B(_06268_),
    .C(_05746_),
    .Y(_06269_));
 AND4x1_ASAP7_75t_R _21147_ (.A(_06263_),
    .B(_06264_),
    .C(_06266_),
    .D(_06269_),
    .Y(_06270_));
 OAI22x1_ASAP7_75t_R _21148_ (.A1(_02176_),
    .A2(_05964_),
    .B1(_05965_),
    .B2(_02113_),
    .Y(_06271_));
 OAI22x1_ASAP7_75t_R _21149_ (.A1(_02141_),
    .A2(_05999_),
    .B1(_05965_),
    .B2(_02078_),
    .Y(_06272_));
 AO32x1_ASAP7_75t_R _21150_ (.A1(_06063_),
    .A2(_06064_),
    .A3(_06271_),
    .B1(_06272_),
    .B2(_06001_),
    .Y(_06273_));
 NAND2x1_ASAP7_75t_R _21151_ (.A(_05814_),
    .B(_06273_),
    .Y(_06274_));
 OA211x2_ASAP7_75t_R _21152_ (.A1(_01414_),
    .A2(_06040_),
    .B(_06270_),
    .C(_06274_),
    .Y(_06275_));
 AOI22x1_ASAP7_75t_R _21153_ (.A1(_05845_),
    .A2(_06262_),
    .B1(_06275_),
    .B2(_18658_),
    .Y(_06276_));
 BUFx12f_ASAP7_75t_R _21154_ (.A(_06276_),
    .Y(_06277_));
 INVx1_ASAP7_75t_R _21155_ (.A(_05940_),
    .Y(_06278_));
 OR3x1_ASAP7_75t_R _21156_ (.A(_02177_),
    .B(_02179_),
    .C(_06256_),
    .Y(_06279_));
 OR4x1_ASAP7_75t_R _21157_ (.A(_02176_),
    .B(_06278_),
    .C(_06113_),
    .D(_06279_),
    .Y(_06280_));
 OR3x1_ASAP7_75t_R _21158_ (.A(_06083_),
    .B(_06089_),
    .C(_06279_),
    .Y(_06281_));
 NAND3x1_ASAP7_75t_R _21159_ (.A(_02176_),
    .B(_06134_),
    .C(_06281_),
    .Y(_06282_));
 OA211x2_ASAP7_75t_R _21160_ (.A1(_06134_),
    .A2(_06277_),
    .B(_06280_),
    .C(_06282_),
    .Y(_02355_));
 AND2x2_ASAP7_75t_R _21161_ (.A(_06060_),
    .B(_18665_),
    .Y(_06283_));
 AO21x1_ASAP7_75t_R _21162_ (.A1(_06059_),
    .A2(_18663_),
    .B(_06283_),
    .Y(_06284_));
 OA222x2_ASAP7_75t_R _21163_ (.A1(_02012_),
    .A2(_05840_),
    .B1(_06104_),
    .B2(_01942_),
    .C1(_05424_),
    .C2(_06014_),
    .Y(_06285_));
 INVx1_ASAP7_75t_R _21164_ (.A(net97),
    .Y(_06286_));
 OA222x2_ASAP7_75t_R _21165_ (.A1(_06286_),
    .A2(_05774_),
    .B1(_05837_),
    .B2(_01980_),
    .C1(_06006_),
    .C2(_01910_),
    .Y(_06287_));
 OA222x2_ASAP7_75t_R _21166_ (.A1(_01892_),
    .A2(_05836_),
    .B1(_06009_),
    .B2(_02040_),
    .C1(_05839_),
    .C2(_01817_),
    .Y(_06288_));
 AND4x1_ASAP7_75t_R _21167_ (.A(_06140_),
    .B(_06285_),
    .C(_06287_),
    .D(_06288_),
    .Y(_06289_));
 OAI22x1_ASAP7_75t_R _21168_ (.A1(_02175_),
    .A2(_05999_),
    .B1(_05965_),
    .B2(_02112_),
    .Y(_06290_));
 INVx1_ASAP7_75t_R _21169_ (.A(_02077_),
    .Y(_06291_));
 INVx1_ASAP7_75t_R _21170_ (.A(_02140_),
    .Y(_06292_));
 AO32x1_ASAP7_75t_R _21171_ (.A1(_06291_),
    .A2(_05994_),
    .A3(_05995_),
    .B1(_05996_),
    .B2(_06292_),
    .Y(_06293_));
 AO32x1_ASAP7_75t_R _21172_ (.A1(_05821_),
    .A2(_05822_),
    .A3(_06290_),
    .B1(_06293_),
    .B2(_06001_),
    .Y(_06294_));
 NAND2x1_ASAP7_75t_R _21173_ (.A(_05992_),
    .B(_06294_),
    .Y(_06295_));
 OA211x2_ASAP7_75t_R _21174_ (.A1(_01415_),
    .A2(_06095_),
    .B(_06289_),
    .C(_06295_),
    .Y(_06296_));
 AOI22x1_ASAP7_75t_R _21175_ (.A1(_06058_),
    .A2(_06284_),
    .B1(_06296_),
    .B2(_18663_),
    .Y(_06297_));
 BUFx12f_ASAP7_75t_R _21176_ (.A(_06297_),
    .Y(_06298_));
 NAND2x1_ASAP7_75t_R _21177_ (.A(_05902_),
    .B(_05957_),
    .Y(_06299_));
 OR4x1_ASAP7_75t_R _21178_ (.A(_02176_),
    .B(_02177_),
    .C(_02179_),
    .D(_06256_),
    .Y(_06300_));
 OR3x1_ASAP7_75t_R _21179_ (.A(_06299_),
    .B(_06089_),
    .C(_06300_),
    .Y(_06301_));
 OR2x2_ASAP7_75t_R _21180_ (.A(_02175_),
    .B(_06301_),
    .Y(_06302_));
 NAND3x1_ASAP7_75t_R _21181_ (.A(_02175_),
    .B(_06133_),
    .C(_06301_),
    .Y(_06303_));
 OA211x2_ASAP7_75t_R _21182_ (.A1(_06134_),
    .A2(_06298_),
    .B(_06302_),
    .C(_06303_),
    .Y(_02356_));
 INVx1_ASAP7_75t_R _21183_ (.A(_02174_),
    .Y(_06304_));
 OR3x1_ASAP7_75t_R _21184_ (.A(_02175_),
    .B(_06089_),
    .C(_06300_),
    .Y(_06305_));
 OR2x2_ASAP7_75t_R _21185_ (.A(_05984_),
    .B(_06305_),
    .Y(_06306_));
 AO21x1_ASAP7_75t_R _21186_ (.A1(_05987_),
    .A2(_06306_),
    .B(_05954_),
    .Y(_06307_));
 INVx1_ASAP7_75t_R _21187_ (.A(_06306_),
    .Y(_06308_));
 AND3x1_ASAP7_75t_R _21188_ (.A(_06060_),
    .B(_16697_),
    .C(_16700_),
    .Y(_06309_));
 AO21x1_ASAP7_75t_R _21189_ (.A1(_06059_),
    .A2(_18668_),
    .B(_06309_),
    .Y(_06310_));
 OA222x2_ASAP7_75t_R _21190_ (.A1(_02011_),
    .A2(_05840_),
    .B1(_06104_),
    .B2(_01941_),
    .C1(_05423_),
    .C2(_06014_),
    .Y(_06311_));
 INVx1_ASAP7_75t_R _21191_ (.A(net98),
    .Y(_06312_));
 OA222x2_ASAP7_75t_R _21192_ (.A1(_06312_),
    .A2(_05773_),
    .B1(_05837_),
    .B2(_01979_),
    .C1(_06006_),
    .C2(_01909_),
    .Y(_06313_));
 OA222x2_ASAP7_75t_R _21193_ (.A1(_01891_),
    .A2(_05836_),
    .B1(_06009_),
    .B2(_02039_),
    .C1(_05839_),
    .C2(_01816_),
    .Y(_06314_));
 AND4x1_ASAP7_75t_R _21194_ (.A(_06140_),
    .B(_06311_),
    .C(_06313_),
    .D(_06314_),
    .Y(_06315_));
 INVx1_ASAP7_75t_R _21195_ (.A(_02111_),
    .Y(_06316_));
 AO32x1_ASAP7_75t_R _21196_ (.A1(_06316_),
    .A2(_05994_),
    .A3(_05995_),
    .B1(_05996_),
    .B2(_06304_),
    .Y(_06317_));
 BUFx6f_ASAP7_75t_R _21197_ (.A(_02139_),
    .Y(_06318_));
 OAI22x1_ASAP7_75t_R _21198_ (.A1(_06318_),
    .A2(_05999_),
    .B1(_05798_),
    .B2(_02076_),
    .Y(_06319_));
 AO32x1_ASAP7_75t_R _21199_ (.A1(_05821_),
    .A2(_05822_),
    .A3(_06317_),
    .B1(_06319_),
    .B2(_05762_),
    .Y(_06320_));
 NAND2x1_ASAP7_75t_R _21200_ (.A(_05992_),
    .B(_06320_),
    .Y(_06321_));
 OA211x2_ASAP7_75t_R _21201_ (.A1(_00007_),
    .A2(_06095_),
    .B(_06315_),
    .C(_06321_),
    .Y(_06322_));
 AOI22x1_ASAP7_75t_R _21202_ (.A1(_06058_),
    .A2(_06310_),
    .B1(_06322_),
    .B2(_18668_),
    .Y(_06323_));
 AO32x1_ASAP7_75t_R _21203_ (.A1(_02174_),
    .A2(_06159_),
    .A3(_06308_),
    .B1(_06323_),
    .B2(_06026_),
    .Y(_06324_));
 AO21x1_ASAP7_75t_R _21204_ (.A1(_06304_),
    .A2(_06307_),
    .B(_06324_),
    .Y(_02357_));
 AND2x4_ASAP7_75t_R _21205_ (.A(_05148_),
    .B(_05748_),
    .Y(_06325_));
 OA211x2_ASAP7_75t_R _21206_ (.A1(_05754_),
    .A2(_05971_),
    .B(_05753_),
    .C(_06325_),
    .Y(_06326_));
 AND2x4_ASAP7_75t_R _21207_ (.A(_05770_),
    .B(_06326_),
    .Y(_06327_));
 AND3x1_ASAP7_75t_R _21208_ (.A(_05989_),
    .B(_16820_),
    .C(_16822_),
    .Y(_06328_));
 AO21x1_ASAP7_75t_R _21209_ (.A1(_05846_),
    .A2(_18673_),
    .B(_06328_),
    .Y(_06329_));
 INVx1_ASAP7_75t_R _21210_ (.A(net164),
    .Y(_06330_));
 OA222x2_ASAP7_75t_R _21211_ (.A1(_02010_),
    .A2(_05840_),
    .B1(_06104_),
    .B2(_01940_),
    .C1(_06330_),
    .C2(_06014_),
    .Y(_06331_));
 INVx1_ASAP7_75t_R _21212_ (.A(net99),
    .Y(_06332_));
 OA222x2_ASAP7_75t_R _21213_ (.A1(_06332_),
    .A2(_05773_),
    .B1(_05837_),
    .B2(_01978_),
    .C1(_06006_),
    .C2(_01908_),
    .Y(_06333_));
 OA222x2_ASAP7_75t_R _21214_ (.A1(_01890_),
    .A2(_05836_),
    .B1(_06009_),
    .B2(_02038_),
    .C1(_05839_),
    .C2(_01815_),
    .Y(_06334_));
 AND4x1_ASAP7_75t_R _21215_ (.A(_06140_),
    .B(_06331_),
    .C(_06333_),
    .D(_06334_),
    .Y(_06335_));
 OAI22x1_ASAP7_75t_R _21216_ (.A1(_02173_),
    .A2(_05999_),
    .B1(_05798_),
    .B2(_02110_),
    .Y(_06336_));
 INVx1_ASAP7_75t_R _21217_ (.A(_02075_),
    .Y(_06337_));
 INVx2_ASAP7_75t_R _21218_ (.A(_02138_),
    .Y(_06338_));
 AO32x1_ASAP7_75t_R _21219_ (.A1(_06337_),
    .A2(_05994_),
    .A3(_05995_),
    .B1(_05996_),
    .B2(_06338_),
    .Y(_06339_));
 AO32x1_ASAP7_75t_R _21220_ (.A1(_05821_),
    .A2(_05822_),
    .A3(_06336_),
    .B1(_06339_),
    .B2(_05762_),
    .Y(_06340_));
 NAND2x1_ASAP7_75t_R _21221_ (.A(_05992_),
    .B(_06340_),
    .Y(_06341_));
 OA211x2_ASAP7_75t_R _21222_ (.A1(_00008_),
    .A2(_06095_),
    .B(_06335_),
    .C(_06341_),
    .Y(_06342_));
 AOI22x1_ASAP7_75t_R _21223_ (.A1(_06058_),
    .A2(_06329_),
    .B1(_06342_),
    .B2(_18673_),
    .Y(_06343_));
 INVx4_ASAP7_75t_R _21224_ (.A(_06343_),
    .Y(_06344_));
 OR3x1_ASAP7_75t_R _21225_ (.A(_02174_),
    .B(_06299_),
    .C(_06305_),
    .Y(_06345_));
 NOR2x1_ASAP7_75t_R _21226_ (.A(_02173_),
    .B(_06345_),
    .Y(_06346_));
 AND3x1_ASAP7_75t_R _21227_ (.A(_02173_),
    .B(_06134_),
    .C(_06345_),
    .Y(_06347_));
 AOI211x1_ASAP7_75t_R _21228_ (.A1(_06327_),
    .A2(_06344_),
    .B(_06346_),
    .C(_06347_),
    .Y(_02358_));
 INVx1_ASAP7_75t_R _21229_ (.A(_02172_),
    .Y(_06348_));
 OR3x2_ASAP7_75t_R _21230_ (.A(_02173_),
    .B(_02174_),
    .C(_06306_),
    .Y(_06349_));
 AO21x1_ASAP7_75t_R _21231_ (.A1(_05987_),
    .A2(_06349_),
    .B(_05954_),
    .Y(_06350_));
 INVx1_ASAP7_75t_R _21232_ (.A(_06349_),
    .Y(_06351_));
 AND2x2_ASAP7_75t_R _21233_ (.A(_06060_),
    .B(_18680_),
    .Y(_06352_));
 AO21x1_ASAP7_75t_R _21234_ (.A1(_06059_),
    .A2(_18678_),
    .B(_06352_),
    .Y(_06353_));
 INVx1_ASAP7_75t_R _21235_ (.A(net165),
    .Y(_06354_));
 OA222x2_ASAP7_75t_R _21236_ (.A1(_02009_),
    .A2(_05840_),
    .B1(_06104_),
    .B2(_01939_),
    .C1(_06354_),
    .C2(_06014_),
    .Y(_06355_));
 INVx1_ASAP7_75t_R _21237_ (.A(net100),
    .Y(_06356_));
 OA222x2_ASAP7_75t_R _21238_ (.A1(_06356_),
    .A2(_05774_),
    .B1(_05837_),
    .B2(_01977_),
    .C1(_06007_),
    .C2(_01907_),
    .Y(_06357_));
 OA222x2_ASAP7_75t_R _21239_ (.A1(_01889_),
    .A2(_05836_),
    .B1(_06009_),
    .B2(_02037_),
    .C1(_05839_),
    .C2(_01814_),
    .Y(_06358_));
 AND4x1_ASAP7_75t_R _21240_ (.A(_06140_),
    .B(_06355_),
    .C(_06357_),
    .D(_06358_),
    .Y(_06359_));
 INVx2_ASAP7_75t_R _21241_ (.A(_02109_),
    .Y(_06360_));
 AO32x1_ASAP7_75t_R _21242_ (.A1(_06360_),
    .A2(_05994_),
    .A3(_05815_),
    .B1(_05826_),
    .B2(_06348_),
    .Y(_06361_));
 OAI22x1_ASAP7_75t_R _21243_ (.A1(_02137_),
    .A2(_05999_),
    .B1(_05965_),
    .B2(_02074_),
    .Y(_06362_));
 AO32x1_ASAP7_75t_R _21244_ (.A1(_05821_),
    .A2(_05822_),
    .A3(_06361_),
    .B1(_06362_),
    .B2(_06001_),
    .Y(_06363_));
 NAND2x1_ASAP7_75t_R _21245_ (.A(_05992_),
    .B(_06363_),
    .Y(_06364_));
 OA211x2_ASAP7_75t_R _21246_ (.A1(_00009_),
    .A2(_06095_),
    .B(_06359_),
    .C(_06364_),
    .Y(_06365_));
 AOI22x1_ASAP7_75t_R _21247_ (.A1(_06058_),
    .A2(_06353_),
    .B1(_06365_),
    .B2(_18678_),
    .Y(_06366_));
 AO32x1_ASAP7_75t_R _21248_ (.A1(_02172_),
    .A2(_06159_),
    .A3(_06351_),
    .B1(_06366_),
    .B2(_05945_),
    .Y(_06367_));
 AO21x1_ASAP7_75t_R _21249_ (.A1(_06348_),
    .A2(_06350_),
    .B(_06367_),
    .Y(_02359_));
 INVx2_ASAP7_75t_R _21250_ (.A(_02171_),
    .Y(_06368_));
 OR2x6_ASAP7_75t_R _21251_ (.A(_05853_),
    .B(_02234_),
    .Y(_06369_));
 OR5x1_ASAP7_75t_R _21252_ (.A(_02172_),
    .B(_02173_),
    .C(_02174_),
    .D(_02175_),
    .E(_05949_),
    .Y(_06370_));
 OR4x1_ASAP7_75t_R _21253_ (.A(_06369_),
    .B(_06089_),
    .C(_06300_),
    .D(_06370_),
    .Y(_06371_));
 AO21x1_ASAP7_75t_R _21254_ (.A1(_05987_),
    .A2(_06371_),
    .B(_05942_),
    .Y(_06372_));
 INVx1_ASAP7_75t_R _21255_ (.A(_06371_),
    .Y(_06373_));
 AND2x2_ASAP7_75t_R _21256_ (.A(_05989_),
    .B(_18685_),
    .Y(_06374_));
 AO21x1_ASAP7_75t_R _21257_ (.A1(_06059_),
    .A2(_18683_),
    .B(_06374_),
    .Y(_06375_));
 INVx2_ASAP7_75t_R _21258_ (.A(_02108_),
    .Y(_06376_));
 AO32x1_ASAP7_75t_R _21259_ (.A1(_06376_),
    .A2(_13454_),
    .A3(_05815_),
    .B1(_05826_),
    .B2(_06368_),
    .Y(_06377_));
 INVx1_ASAP7_75t_R _21260_ (.A(_02073_),
    .Y(_06378_));
 INVx1_ASAP7_75t_R _21261_ (.A(_02136_),
    .Y(_06379_));
 AO32x1_ASAP7_75t_R _21262_ (.A1(_06378_),
    .A2(_05994_),
    .A3(_05995_),
    .B1(_05996_),
    .B2(_06379_),
    .Y(_06380_));
 AO32x1_ASAP7_75t_R _21263_ (.A1(_05821_),
    .A2(_05822_),
    .A3(_06377_),
    .B1(_06380_),
    .B2(_06001_),
    .Y(_06381_));
 NAND2x1_ASAP7_75t_R _21264_ (.A(_05992_),
    .B(_06381_),
    .Y(_06382_));
 INVx1_ASAP7_75t_R _21265_ (.A(net152),
    .Y(_06383_));
 OA222x2_ASAP7_75t_R _21266_ (.A1(_02008_),
    .A2(_05840_),
    .B1(_06104_),
    .B2(_01938_),
    .C1(_06383_),
    .C2(_06014_),
    .Y(_06384_));
 INVx1_ASAP7_75t_R _21267_ (.A(net101),
    .Y(_06385_));
 OA222x2_ASAP7_75t_R _21268_ (.A1(_06385_),
    .A2(_05773_),
    .B1(_05837_),
    .B2(_01976_),
    .C1(_06006_),
    .C2(_01923_),
    .Y(_06386_));
 OA222x2_ASAP7_75t_R _21269_ (.A1(_01888_),
    .A2(_05836_),
    .B1(_06009_),
    .B2(_02036_),
    .C1(_05839_),
    .C2(_01813_),
    .Y(_06387_));
 AND4x1_ASAP7_75t_R _21270_ (.A(_06140_),
    .B(_06384_),
    .C(_06386_),
    .D(_06387_),
    .Y(_06388_));
 OA211x2_ASAP7_75t_R _21271_ (.A1(_00010_),
    .A2(_06095_),
    .B(_06382_),
    .C(_06388_),
    .Y(_06389_));
 AOI22x1_ASAP7_75t_R _21272_ (.A1(_06058_),
    .A2(_06375_),
    .B1(_06389_),
    .B2(_18683_),
    .Y(_06390_));
 BUFx12f_ASAP7_75t_R _21273_ (.A(_06390_),
    .Y(_06391_));
 AO32x1_ASAP7_75t_R _21274_ (.A1(_02171_),
    .A2(_06159_),
    .A3(_06373_),
    .B1(_06391_),
    .B2(_05945_),
    .Y(_06392_));
 AO21x1_ASAP7_75t_R _21275_ (.A1(_06368_),
    .A2(_06372_),
    .B(_06392_),
    .Y(_02360_));
 INVx1_ASAP7_75t_R _21276_ (.A(_02170_),
    .Y(_06393_));
 OR3x1_ASAP7_75t_R _21277_ (.A(_02171_),
    .B(_02172_),
    .C(_06349_),
    .Y(_06394_));
 AO21x1_ASAP7_75t_R _21278_ (.A1(_05987_),
    .A2(_06394_),
    .B(_05942_),
    .Y(_06395_));
 AND3x1_ASAP7_75t_R _21279_ (.A(_06348_),
    .B(_05940_),
    .C(_06351_),
    .Y(_06396_));
 AND3x1_ASAP7_75t_R _21280_ (.A(_06060_),
    .B(_04418_),
    .C(_04421_),
    .Y(_06397_));
 AO21x1_ASAP7_75t_R _21281_ (.A1(_06059_),
    .A2(_18688_),
    .B(_06397_),
    .Y(_06398_));
 INVx1_ASAP7_75t_R _21282_ (.A(net153),
    .Y(_06399_));
 OA222x2_ASAP7_75t_R _21283_ (.A1(_02007_),
    .A2(_05799_),
    .B1(_05789_),
    .B2(_01937_),
    .C1(_06399_),
    .C2(_06014_),
    .Y(_06400_));
 INVx1_ASAP7_75t_R _21284_ (.A(net102),
    .Y(_06401_));
 OA222x2_ASAP7_75t_R _21285_ (.A1(_06401_),
    .A2(_05773_),
    .B1(_05837_),
    .B2(_01975_),
    .C1(_06006_),
    .C2(_01922_),
    .Y(_06402_));
 OA222x2_ASAP7_75t_R _21286_ (.A1(_01887_),
    .A2(_05778_),
    .B1(_05830_),
    .B2(_02035_),
    .C1(_05784_),
    .C2(_01812_),
    .Y(_06403_));
 AND4x1_ASAP7_75t_R _21287_ (.A(_06140_),
    .B(_06400_),
    .C(_06402_),
    .D(_06403_),
    .Y(_06404_));
 INVx2_ASAP7_75t_R _21288_ (.A(_02107_),
    .Y(_06405_));
 AO32x1_ASAP7_75t_R _21289_ (.A1(_06405_),
    .A2(_13453_),
    .A3(_05995_),
    .B1(_05996_),
    .B2(_06393_),
    .Y(_06406_));
 OAI22x1_ASAP7_75t_R _21290_ (.A1(_02135_),
    .A2(_05744_),
    .B1(_05798_),
    .B2(_02072_),
    .Y(_06407_));
 AO32x2_ASAP7_75t_R _21291_ (.A1(_05058_),
    .A2(_05069_),
    .A3(_06406_),
    .B1(_06407_),
    .B2(_05762_),
    .Y(_06408_));
 NAND2x1_ASAP7_75t_R _21292_ (.A(_05767_),
    .B(_06408_),
    .Y(_06409_));
 OA211x2_ASAP7_75t_R _21293_ (.A1(_00011_),
    .A2(_06095_),
    .B(_06404_),
    .C(_06409_),
    .Y(_06410_));
 AOI22x1_ASAP7_75t_R _21294_ (.A1(_06058_),
    .A2(_06398_),
    .B1(_06410_),
    .B2(_18688_),
    .Y(_06411_));
 AO32x1_ASAP7_75t_R _21295_ (.A1(_02170_),
    .A2(_06368_),
    .A3(_06396_),
    .B1(_06411_),
    .B2(_05945_),
    .Y(_06412_));
 AO21x1_ASAP7_75t_R _21296_ (.A1(_06393_),
    .A2(_06395_),
    .B(_06412_),
    .Y(_02361_));
 INVx1_ASAP7_75t_R _21297_ (.A(_02169_),
    .Y(_06413_));
 OR3x1_ASAP7_75t_R _21298_ (.A(_02170_),
    .B(_02171_),
    .C(_06371_),
    .Y(_06414_));
 AO21x1_ASAP7_75t_R _21299_ (.A1(_05987_),
    .A2(_06414_),
    .B(_05942_),
    .Y(_06415_));
 AND2x2_ASAP7_75t_R _21300_ (.A(_06060_),
    .B(_18695_),
    .Y(_06416_));
 AO21x1_ASAP7_75t_R _21301_ (.A1(_05960_),
    .A2(_18693_),
    .B(_06416_),
    .Y(_06417_));
 INVx1_ASAP7_75t_R _21302_ (.A(net154),
    .Y(_06418_));
 OA222x2_ASAP7_75t_R _21303_ (.A1(_02006_),
    .A2(_05799_),
    .B1(_05789_),
    .B2(_01936_),
    .C1(_06418_),
    .C2(_06014_),
    .Y(_06419_));
 INVx1_ASAP7_75t_R _21304_ (.A(net103),
    .Y(_06420_));
 OA222x2_ASAP7_75t_R _21305_ (.A1(_06420_),
    .A2(_05773_),
    .B1(_05837_),
    .B2(_01974_),
    .C1(_06006_),
    .C2(_01921_),
    .Y(_06421_));
 OA222x2_ASAP7_75t_R _21306_ (.A1(_01886_),
    .A2(_05836_),
    .B1(_06009_),
    .B2(_02034_),
    .C1(_05784_),
    .C2(_01811_),
    .Y(_06422_));
 AND4x1_ASAP7_75t_R _21307_ (.A(_06140_),
    .B(_06419_),
    .C(_06421_),
    .D(_06422_),
    .Y(_06423_));
 INVx2_ASAP7_75t_R _21308_ (.A(_02106_),
    .Y(_06424_));
 AO32x1_ASAP7_75t_R _21309_ (.A1(_06424_),
    .A2(_05994_),
    .A3(_05995_),
    .B1(_05996_),
    .B2(_06413_),
    .Y(_06425_));
 INVx1_ASAP7_75t_R _21310_ (.A(_02070_),
    .Y(_06426_));
 INVx2_ASAP7_75t_R _21311_ (.A(_02133_),
    .Y(_06427_));
 AO32x1_ASAP7_75t_R _21312_ (.A1(_06426_),
    .A2(_05994_),
    .A3(_05995_),
    .B1(_05996_),
    .B2(_06427_),
    .Y(_06428_));
 AO32x2_ASAP7_75t_R _21313_ (.A1(_05058_),
    .A2(_05069_),
    .A3(_06425_),
    .B1(_06428_),
    .B2(_05762_),
    .Y(_06429_));
 NAND2x1_ASAP7_75t_R _21314_ (.A(_05767_),
    .B(_06429_),
    .Y(_06430_));
 OA211x2_ASAP7_75t_R _21315_ (.A1(_00012_),
    .A2(_06095_),
    .B(_06423_),
    .C(_06430_),
    .Y(_06431_));
 AOI22x1_ASAP7_75t_R _21316_ (.A1(_05959_),
    .A2(_06417_),
    .B1(_06431_),
    .B2(_18693_),
    .Y(_06432_));
 AND5x1_ASAP7_75t_R _21317_ (.A(_02169_),
    .B(_06393_),
    .C(_06368_),
    .D(_05940_),
    .E(_06373_),
    .Y(_06433_));
 AO21x1_ASAP7_75t_R _21318_ (.A1(_06026_),
    .A2(_06432_),
    .B(_06433_),
    .Y(_06434_));
 AO21x1_ASAP7_75t_R _21319_ (.A1(_06413_),
    .A2(_06415_),
    .B(_06434_),
    .Y(_02362_));
 INVx1_ASAP7_75t_R _21320_ (.A(_02168_),
    .Y(_06435_));
 OR3x2_ASAP7_75t_R _21321_ (.A(_02169_),
    .B(_02170_),
    .C(_02171_),
    .Y(_06436_));
 OR3x1_ASAP7_75t_R _21322_ (.A(_02172_),
    .B(_06349_),
    .C(_06436_),
    .Y(_06437_));
 AO21x1_ASAP7_75t_R _21323_ (.A1(_05987_),
    .A2(_06437_),
    .B(_05942_),
    .Y(_06438_));
 INVx1_ASAP7_75t_R _21324_ (.A(_06436_),
    .Y(_06439_));
 AND3x1_ASAP7_75t_R _21325_ (.A(_06060_),
    .B(_04666_),
    .C(_04669_),
    .Y(_06440_));
 AO21x1_ASAP7_75t_R _21326_ (.A1(_05960_),
    .A2(_18698_),
    .B(_06440_),
    .Y(_06441_));
 INVx1_ASAP7_75t_R _21327_ (.A(net155),
    .Y(_06442_));
 OA222x2_ASAP7_75t_R _21328_ (.A1(_02005_),
    .A2(_05800_),
    .B1(_05790_),
    .B2(_01935_),
    .C1(_06442_),
    .C2(_06015_),
    .Y(_06443_));
 INVx1_ASAP7_75t_R _21329_ (.A(net104),
    .Y(_06444_));
 OA222x2_ASAP7_75t_R _21330_ (.A1(_06444_),
    .A2(_05774_),
    .B1(_05782_),
    .B2(_01973_),
    .C1(_06007_),
    .C2(_01920_),
    .Y(_06445_));
 OA222x2_ASAP7_75t_R _21331_ (.A1(_01885_),
    .A2(_05779_),
    .B1(_05831_),
    .B2(_02033_),
    .C1(_05785_),
    .C2(_01810_),
    .Y(_06446_));
 AND4x1_ASAP7_75t_R _21332_ (.A(_05747_),
    .B(_06443_),
    .C(_06445_),
    .D(_06446_),
    .Y(_06447_));
 INVx2_ASAP7_75t_R _21333_ (.A(_02105_),
    .Y(_06448_));
 AO32x1_ASAP7_75t_R _21334_ (.A1(_06448_),
    .A2(_13454_),
    .A3(_05815_),
    .B1(_05826_),
    .B2(_06435_),
    .Y(_06449_));
 OAI22x1_ASAP7_75t_R _21335_ (.A1(_02132_),
    .A2(_05964_),
    .B1(_05965_),
    .B2(_02069_),
    .Y(_06450_));
 AO32x2_ASAP7_75t_R _21336_ (.A1(_06063_),
    .A2(_06064_),
    .A3(_06449_),
    .B1(_06450_),
    .B2(_06001_),
    .Y(_06451_));
 NAND2x1_ASAP7_75t_R _21337_ (.A(_05814_),
    .B(_06451_),
    .Y(_06452_));
 OA211x2_ASAP7_75t_R _21338_ (.A1(_00013_),
    .A2(_06040_),
    .B(_06447_),
    .C(_06452_),
    .Y(_06453_));
 AOI22x1_ASAP7_75t_R _21339_ (.A1(_05959_),
    .A2(_06441_),
    .B1(_06453_),
    .B2(_18698_),
    .Y(_06454_));
 AO32x1_ASAP7_75t_R _21340_ (.A1(_02168_),
    .A2(_06396_),
    .A3(_06439_),
    .B1(_06454_),
    .B2(_05945_),
    .Y(_06455_));
 AO21x1_ASAP7_75t_R _21341_ (.A1(_06435_),
    .A2(_06438_),
    .B(_06455_),
    .Y(_02363_));
 AO21x1_ASAP7_75t_R _21342_ (.A1(_05902_),
    .A2(_06369_),
    .B(_05941_),
    .Y(_06456_));
 OAI21x1_ASAP7_75t_R _21343_ (.A1(_06326_),
    .A2(_06369_),
    .B(_02167_),
    .Y(_06457_));
 OA21x2_ASAP7_75t_R _21344_ (.A1(_02167_),
    .A2(_06456_),
    .B(_06457_),
    .Y(_06458_));
 AO21x1_ASAP7_75t_R _21345_ (.A1(_05851_),
    .A2(_06327_),
    .B(_06458_),
    .Y(_02364_));
 INVx1_ASAP7_75t_R _21346_ (.A(_02166_),
    .Y(_06459_));
 OR3x1_ASAP7_75t_R _21347_ (.A(_02168_),
    .B(_06371_),
    .C(_06436_),
    .Y(_06460_));
 AO21x1_ASAP7_75t_R _21348_ (.A1(_05987_),
    .A2(_06460_),
    .B(_05942_),
    .Y(_06461_));
 INVx1_ASAP7_75t_R _21349_ (.A(_06460_),
    .Y(_06462_));
 AND3x1_ASAP7_75t_R _21350_ (.A(_06060_),
    .B(_04788_),
    .C(_04790_),
    .Y(_06463_));
 AO21x1_ASAP7_75t_R _21351_ (.A1(_06059_),
    .A2(_18703_),
    .B(_06463_),
    .Y(_06464_));
 INVx1_ASAP7_75t_R _21352_ (.A(_02103_),
    .Y(_06465_));
 AO32x1_ASAP7_75t_R _21353_ (.A1(_06465_),
    .A2(_06119_),
    .A3(_06066_),
    .B1(_06067_),
    .B2(_06459_),
    .Y(_06466_));
 INVx1_ASAP7_75t_R _21354_ (.A(_02068_),
    .Y(_06467_));
 INVx1_ASAP7_75t_R _21355_ (.A(_02131_),
    .Y(_06468_));
 AO32x1_ASAP7_75t_R _21356_ (.A1(_06467_),
    .A2(_06119_),
    .A3(_06066_),
    .B1(_06067_),
    .B2(_06468_),
    .Y(_06469_));
 AO32x2_ASAP7_75t_R _21357_ (.A1(_06063_),
    .A2(_06064_),
    .A3(_06466_),
    .B1(_06469_),
    .B2(_05763_),
    .Y(_06470_));
 NAND2x1_ASAP7_75t_R _21358_ (.A(_05814_),
    .B(_06470_),
    .Y(_06471_));
 OA22x2_ASAP7_75t_R _21359_ (.A1(_01808_),
    .A2(_06004_),
    .B1(_06010_),
    .B2(_02031_),
    .Y(_06472_));
 OA222x2_ASAP7_75t_R _21360_ (.A1(_01883_),
    .A2(_06047_),
    .B1(_06007_),
    .B2(_01919_),
    .C1(_06015_),
    .C2(_05418_),
    .Y(_06473_));
 OA22x2_ASAP7_75t_R _21361_ (.A1(_02003_),
    .A2(_06005_),
    .B1(_05791_),
    .B2(_01933_),
    .Y(_06474_));
 NAND2x1_ASAP7_75t_R _21362_ (.A(net106),
    .B(_06077_),
    .Y(_06475_));
 OA211x2_ASAP7_75t_R _21363_ (.A1(_01971_),
    .A2(_06045_),
    .B(_06475_),
    .C(_05140_),
    .Y(_06476_));
 OA211x2_ASAP7_75t_R _21364_ (.A1(_00014_),
    .A2(_06095_),
    .B(_06020_),
    .C(_06476_),
    .Y(_06477_));
 AND5x2_ASAP7_75t_R _21365_ (.A(_06471_),
    .B(_06472_),
    .C(_06473_),
    .D(_06474_),
    .E(_06477_),
    .Y(_06478_));
 AOI22x1_ASAP7_75t_R _21366_ (.A1(_05845_),
    .A2(_06464_),
    .B1(_06478_),
    .B2(_18703_),
    .Y(_06479_));
 BUFx12f_ASAP7_75t_R _21367_ (.A(_06479_),
    .Y(_06480_));
 AO32x1_ASAP7_75t_R _21368_ (.A1(_02166_),
    .A2(_06159_),
    .A3(_06462_),
    .B1(_06480_),
    .B2(_05945_),
    .Y(_06481_));
 AO21x1_ASAP7_75t_R _21369_ (.A1(_06459_),
    .A2(_06461_),
    .B(_06481_),
    .Y(_02365_));
 INVx1_ASAP7_75t_R _21370_ (.A(_02165_),
    .Y(_06482_));
 OR3x1_ASAP7_75t_R _21371_ (.A(_02166_),
    .B(_02168_),
    .C(_06436_),
    .Y(_06483_));
 OR3x1_ASAP7_75t_R _21372_ (.A(_02172_),
    .B(_06349_),
    .C(_06483_),
    .Y(_06484_));
 AO21x1_ASAP7_75t_R _21373_ (.A1(_05987_),
    .A2(_06484_),
    .B(_05942_),
    .Y(_06485_));
 INVx1_ASAP7_75t_R _21374_ (.A(_06483_),
    .Y(_06486_));
 AND2x2_ASAP7_75t_R _21375_ (.A(_05989_),
    .B(_18072_),
    .Y(_06487_));
 AO21x1_ASAP7_75t_R _21376_ (.A1(_05846_),
    .A2(_18070_),
    .B(_06487_),
    .Y(_06488_));
 INVx1_ASAP7_75t_R _21377_ (.A(_02102_),
    .Y(_06489_));
 AO32x1_ASAP7_75t_R _21378_ (.A1(_06489_),
    .A2(_13454_),
    .A3(_05815_),
    .B1(_05826_),
    .B2(_06482_),
    .Y(_06490_));
 INVx1_ASAP7_75t_R _21379_ (.A(_02067_),
    .Y(_06491_));
 INVx1_ASAP7_75t_R _21380_ (.A(_02130_),
    .Y(_06492_));
 AO32x1_ASAP7_75t_R _21381_ (.A1(_06491_),
    .A2(_13454_),
    .A3(_05815_),
    .B1(_05826_),
    .B2(_06492_),
    .Y(_06493_));
 AO32x2_ASAP7_75t_R _21382_ (.A1(_06063_),
    .A2(_06064_),
    .A3(_06490_),
    .B1(_06493_),
    .B2(_06001_),
    .Y(_06494_));
 NAND2x1_ASAP7_75t_R _21383_ (.A(_05814_),
    .B(_06494_),
    .Y(_06495_));
 OA22x2_ASAP7_75t_R _21384_ (.A1(_01807_),
    .A2(_05785_),
    .B1(_05831_),
    .B2(_02030_),
    .Y(_06496_));
 OA22x2_ASAP7_75t_R _21385_ (.A1(_02002_),
    .A2(_05800_),
    .B1(_05801_),
    .B2(_01957_),
    .Y(_06497_));
 OA21x2_ASAP7_75t_R _21386_ (.A1(_01970_),
    .A2(_05782_),
    .B(_05746_),
    .Y(_06498_));
 NAND2x1_ASAP7_75t_R _21387_ (.A(net107),
    .B(_06077_),
    .Y(_06499_));
 OA22x2_ASAP7_75t_R _21388_ (.A1(_01882_),
    .A2(_05779_),
    .B1(_06104_),
    .B2(_01932_),
    .Y(_06500_));
 AND5x1_ASAP7_75t_R _21389_ (.A(_06496_),
    .B(_06497_),
    .C(_06498_),
    .D(_06499_),
    .E(_06500_),
    .Y(_06501_));
 OA211x2_ASAP7_75t_R _21390_ (.A1(_00015_),
    .A2(_06040_),
    .B(_06495_),
    .C(_06501_),
    .Y(_06502_));
 AOI22x1_ASAP7_75t_R _21391_ (.A1(_05845_),
    .A2(_06488_),
    .B1(_06502_),
    .B2(_18070_),
    .Y(_06503_));
 BUFx12f_ASAP7_75t_R _21392_ (.A(_06503_),
    .Y(_06504_));
 AO32x1_ASAP7_75t_R _21393_ (.A1(_02165_),
    .A2(_06396_),
    .A3(_06486_),
    .B1(_06504_),
    .B2(_05945_),
    .Y(_06505_));
 AO21x1_ASAP7_75t_R _21394_ (.A1(_06482_),
    .A2(_06485_),
    .B(_06505_),
    .Y(_02366_));
 BUFx6f_ASAP7_75t_R _21395_ (.A(_06159_),
    .Y(_06506_));
 NOR2x2_ASAP7_75t_R _21396_ (.A(_05906_),
    .B(_05937_),
    .Y(_06507_));
 AND2x6_ASAP7_75t_R _21397_ (.A(_05753_),
    .B(_06507_),
    .Y(_06508_));
 NOR2x2_ASAP7_75t_R _21398_ (.A(_05750_),
    .B(_06508_),
    .Y(_06509_));
 OR5x2_ASAP7_75t_R _21399_ (.A(_02165_),
    .B(_06089_),
    .C(_06300_),
    .D(_06370_),
    .E(_06483_),
    .Y(_06510_));
 OR3x1_ASAP7_75t_R _21400_ (.A(_05764_),
    .B(_02234_),
    .C(_06510_),
    .Y(_06511_));
 OAI21x1_ASAP7_75t_R _21401_ (.A1(_02234_),
    .A2(_06510_),
    .B(_05764_),
    .Y(_06512_));
 OAI21x1_ASAP7_75t_R _21402_ (.A1(_06509_),
    .A2(_06511_),
    .B(_06512_),
    .Y(_06513_));
 BUFx6f_ASAP7_75t_R _21403_ (.A(_06508_),
    .Y(_06514_));
 AO21x1_ASAP7_75t_R _21404_ (.A1(_05750_),
    .A2(_05902_),
    .B(_06508_),
    .Y(_06515_));
 BUFx6f_ASAP7_75t_R _21405_ (.A(_06515_),
    .Y(_06516_));
 BUFx12f_ASAP7_75t_R _21406_ (.A(_06516_),
    .Y(_06517_));
 NOR2x1_ASAP7_75t_R _21407_ (.A(_02164_),
    .B(_06517_),
    .Y(_06518_));
 AO21x1_ASAP7_75t_R _21408_ (.A1(_05811_),
    .A2(_06514_),
    .B(_06518_),
    .Y(_06519_));
 AO21x1_ASAP7_75t_R _21409_ (.A1(_06506_),
    .A2(_06513_),
    .B(_06519_),
    .Y(_02367_));
 INVx1_ASAP7_75t_R _21410_ (.A(_06227_),
    .Y(_06520_));
 OR3x1_ASAP7_75t_R _21411_ (.A(_00747_),
    .B(_02164_),
    .C(_02178_),
    .Y(_06521_));
 NOR2x1_ASAP7_75t_R _21412_ (.A(_06510_),
    .B(_06521_),
    .Y(_06522_));
 INVx1_ASAP7_75t_R _21413_ (.A(_06522_),
    .Y(_06523_));
 AO21x2_ASAP7_75t_R _21414_ (.A1(_05753_),
    .A2(_06507_),
    .B(_05750_),
    .Y(_06524_));
 BUFx6f_ASAP7_75t_R _21415_ (.A(_06524_),
    .Y(_06525_));
 AND3x1_ASAP7_75t_R _21416_ (.A(_06227_),
    .B(_06525_),
    .C(_06522_),
    .Y(_06526_));
 AO21x1_ASAP7_75t_R _21417_ (.A1(_06520_),
    .A2(_06523_),
    .B(_06526_),
    .Y(_06527_));
 NOR2x1_ASAP7_75t_R _21418_ (.A(_06227_),
    .B(_06517_),
    .Y(_06528_));
 AO21x1_ASAP7_75t_R _21419_ (.A1(_06235_),
    .A2(_06514_),
    .B(_06528_),
    .Y(_06529_));
 AO21x1_ASAP7_75t_R _21420_ (.A1(_06506_),
    .A2(_06527_),
    .B(_06529_),
    .Y(_02368_));
 OR4x1_ASAP7_75t_R _21421_ (.A(_06227_),
    .B(_02164_),
    .C(_02234_),
    .D(_06510_),
    .Y(_06530_));
 OAI21x1_ASAP7_75t_R _21422_ (.A1(_06509_),
    .A2(_06530_),
    .B(_05823_),
    .Y(_06531_));
 OA21x2_ASAP7_75t_R _21423_ (.A1(_05823_),
    .A2(_06530_),
    .B(_06531_),
    .Y(_06532_));
 NOR2x1_ASAP7_75t_R _21424_ (.A(_05823_),
    .B(_06517_),
    .Y(_06533_));
 AO21x1_ASAP7_75t_R _21425_ (.A1(_05851_),
    .A2(_06514_),
    .B(_06533_),
    .Y(_06534_));
 AO21x1_ASAP7_75t_R _21426_ (.A1(_06506_),
    .A2(_06532_),
    .B(_06534_),
    .Y(_02369_));
 INVx1_ASAP7_75t_R _21427_ (.A(_02161_),
    .Y(_06535_));
 OR3x1_ASAP7_75t_R _21428_ (.A(_05823_),
    .B(_06227_),
    .C(_06523_),
    .Y(_06536_));
 INVx1_ASAP7_75t_R _21429_ (.A(_06536_),
    .Y(_06537_));
 AND3x1_ASAP7_75t_R _21430_ (.A(_02161_),
    .B(_06525_),
    .C(_06537_),
    .Y(_06538_));
 AO21x1_ASAP7_75t_R _21431_ (.A1(_06535_),
    .A2(_06536_),
    .B(_06538_),
    .Y(_06539_));
 AND2x2_ASAP7_75t_R _21432_ (.A(_05989_),
    .B(_18567_),
    .Y(_06540_));
 AO21x1_ASAP7_75t_R _21433_ (.A1(_05846_),
    .A2(_18569_),
    .B(_06540_),
    .Y(_06541_));
 OAI22x1_ASAP7_75t_R _21434_ (.A1(_02156_),
    .A2(_05964_),
    .B1(_05966_),
    .B2(_02093_),
    .Y(_06542_));
 INVx1_ASAP7_75t_R _21435_ (.A(_02098_),
    .Y(_06543_));
 AO32x1_ASAP7_75t_R _21436_ (.A1(_06543_),
    .A2(_18553_),
    .A3(_05816_),
    .B1(_05827_),
    .B2(_06535_),
    .Y(_06544_));
 AOI22x1_ASAP7_75t_R _21437_ (.A1(_05754_),
    .A2(_06542_),
    .B1(_06544_),
    .B2(_05971_),
    .Y(_06545_));
 OA222x2_ASAP7_75t_R _21438_ (.A1(_02001_),
    .A2(_05800_),
    .B1(_05801_),
    .B2(_01959_),
    .C1(_00759_),
    .C2(_06018_),
    .Y(_06546_));
 OA22x2_ASAP7_75t_R _21439_ (.A1(_01881_),
    .A2(_06047_),
    .B1(_05790_),
    .B2(_01931_),
    .Y(_06547_));
 OA21x2_ASAP7_75t_R _21440_ (.A1(_01806_),
    .A2(_05785_),
    .B(_05746_),
    .Y(_06548_));
 AND3x1_ASAP7_75t_R _21441_ (.A(_06546_),
    .B(_06547_),
    .C(_06548_),
    .Y(_06549_));
 INVx1_ASAP7_75t_R _21442_ (.A(net108),
    .Y(_06550_));
 OA222x2_ASAP7_75t_R _21443_ (.A1(_06550_),
    .A2(_05774_),
    .B1(_05782_),
    .B2(_01969_),
    .C1(_05831_),
    .C2(_01399_),
    .Y(_06551_));
 OR2x2_ASAP7_75t_R _21444_ (.A(_05443_),
    .B(_06015_),
    .Y(_06552_));
 OA211x2_ASAP7_75t_R _21445_ (.A1(_01916_),
    .A2(_06007_),
    .B(_06551_),
    .C(_06552_),
    .Y(_06553_));
 OA211x2_ASAP7_75t_R _21446_ (.A1(_05963_),
    .A2(_06545_),
    .B(_06549_),
    .C(_06553_),
    .Y(_06554_));
 AOI22x1_ASAP7_75t_R _21447_ (.A1(_05845_),
    .A2(_06541_),
    .B1(_06554_),
    .B2(_18569_),
    .Y(_06555_));
 BUFx12f_ASAP7_75t_R _21448_ (.A(_06555_),
    .Y(_06556_));
 NOR2x1_ASAP7_75t_R _21449_ (.A(_02161_),
    .B(_06517_),
    .Y(_06557_));
 AO21x1_ASAP7_75t_R _21450_ (.A1(_06514_),
    .A2(_06556_),
    .B(_06557_),
    .Y(_06558_));
 AO21x1_ASAP7_75t_R _21451_ (.A1(_06506_),
    .A2(_06539_),
    .B(_06558_),
    .Y(_02370_));
 OR3x1_ASAP7_75t_R _21452_ (.A(_02161_),
    .B(_05823_),
    .C(_06530_),
    .Y(_06559_));
 INVx1_ASAP7_75t_R _21453_ (.A(_06559_),
    .Y(_06560_));
 INVx1_ASAP7_75t_R _21454_ (.A(_02160_),
    .Y(_06561_));
 OR5x1_ASAP7_75t_R _21455_ (.A(_06561_),
    .B(_02161_),
    .C(_05823_),
    .D(_06509_),
    .E(_06530_),
    .Y(_06562_));
 OAI21x1_ASAP7_75t_R _21456_ (.A1(_02160_),
    .A2(_06560_),
    .B(_06562_),
    .Y(_06563_));
 AND2x2_ASAP7_75t_R _21457_ (.A(_18074_),
    .B(_18572_),
    .Y(_06564_));
 AO21x1_ASAP7_75t_R _21458_ (.A1(_05960_),
    .A2(_18574_),
    .B(_06564_),
    .Y(_06565_));
 INVx1_ASAP7_75t_R _21459_ (.A(net109),
    .Y(_06566_));
 OA21x2_ASAP7_75t_R _21460_ (.A1(_01968_),
    .A2(_06045_),
    .B(_06140_),
    .Y(_06567_));
 OA22x2_ASAP7_75t_R _21461_ (.A1(_02000_),
    .A2(_06005_),
    .B1(_06010_),
    .B2(_01400_),
    .Y(_06568_));
 OA211x2_ASAP7_75t_R _21462_ (.A1(_06566_),
    .A2(_05975_),
    .B(_06567_),
    .C(_06568_),
    .Y(_06569_));
 OA22x2_ASAP7_75t_R _21463_ (.A1(_01880_),
    .A2(_06047_),
    .B1(_05791_),
    .B2(_01930_),
    .Y(_06570_));
 OA22x2_ASAP7_75t_R _21464_ (.A1(_01805_),
    .A2(_06004_),
    .B1(_05801_),
    .B2(_01958_),
    .Y(_06571_));
 INVx2_ASAP7_75t_R _21465_ (.A(_02082_),
    .Y(_06572_));
 INVx1_ASAP7_75t_R _21466_ (.A(_02145_),
    .Y(_06573_));
 AO32x1_ASAP7_75t_R _21467_ (.A1(_06572_),
    .A2(_06119_),
    .A3(_06066_),
    .B1(_06067_),
    .B2(_06573_),
    .Y(_06574_));
 INVx2_ASAP7_75t_R _21468_ (.A(_02097_),
    .Y(_06575_));
 AO32x1_ASAP7_75t_R _21469_ (.A1(_06575_),
    .A2(_06119_),
    .A3(_06066_),
    .B1(_06067_),
    .B2(_06561_),
    .Y(_06576_));
 AO32x1_ASAP7_75t_R _21470_ (.A1(_06063_),
    .A2(_06064_),
    .A3(_06574_),
    .B1(_06576_),
    .B2(_05763_),
    .Y(_06577_));
 NAND2x1_ASAP7_75t_R _21471_ (.A(_05814_),
    .B(_06577_),
    .Y(_06578_));
 AND4x1_ASAP7_75t_R _21472_ (.A(_06569_),
    .B(_06570_),
    .C(_06571_),
    .D(_06578_),
    .Y(_06579_));
 AOI22x1_ASAP7_75t_R _21473_ (.A1(_05959_),
    .A2(_06565_),
    .B1(_06579_),
    .B2(_18574_),
    .Y(_06580_));
 NOR2x1_ASAP7_75t_R _21474_ (.A(_02160_),
    .B(_06517_),
    .Y(_06581_));
 AO21x1_ASAP7_75t_R _21475_ (.A1(_06514_),
    .A2(_06580_),
    .B(_06581_),
    .Y(_06582_));
 AO21x1_ASAP7_75t_R _21476_ (.A1(_06506_),
    .A2(_06563_),
    .B(_06582_),
    .Y(_02371_));
 INVx1_ASAP7_75t_R _21477_ (.A(_02159_),
    .Y(_06583_));
 OR3x1_ASAP7_75t_R _21478_ (.A(_02160_),
    .B(_02161_),
    .C(_06536_),
    .Y(_06584_));
 BUFx6f_ASAP7_75t_R _21479_ (.A(_06524_),
    .Y(_06585_));
 AND5x1_ASAP7_75t_R _21480_ (.A(_02159_),
    .B(_06561_),
    .C(_06535_),
    .D(_06585_),
    .E(_06537_),
    .Y(_06586_));
 AO21x1_ASAP7_75t_R _21481_ (.A1(_06583_),
    .A2(_06584_),
    .B(_06586_),
    .Y(_06587_));
 AND3x1_ASAP7_75t_R _21482_ (.A(_18074_),
    .B(_14899_),
    .C(_14902_),
    .Y(_06588_));
 AO21x1_ASAP7_75t_R _21483_ (.A1(_05960_),
    .A2(_18579_),
    .B(_06588_),
    .Y(_06589_));
 OAI22x1_ASAP7_75t_R _21484_ (.A1(_02134_),
    .A2(_05964_),
    .B1(_05966_),
    .B2(_02071_),
    .Y(_06590_));
 INVx1_ASAP7_75t_R _21485_ (.A(_02096_),
    .Y(_06591_));
 AO32x2_ASAP7_75t_R _21486_ (.A1(_06591_),
    .A2(_18553_),
    .A3(_05816_),
    .B1(_05827_),
    .B2(_06583_),
    .Y(_06592_));
 AOI22x1_ASAP7_75t_R _21487_ (.A1(_05754_),
    .A2(_06590_),
    .B1(_06592_),
    .B2(_05971_),
    .Y(_06593_));
 OA22x2_ASAP7_75t_R _21488_ (.A1(_01999_),
    .A2(_06005_),
    .B1(_06010_),
    .B2(_01401_),
    .Y(_06594_));
 INVx1_ASAP7_75t_R _21489_ (.A(net110),
    .Y(_06595_));
 OA21x2_ASAP7_75t_R _21490_ (.A1(_01967_),
    .A2(_06045_),
    .B(_05746_),
    .Y(_06596_));
 OA222x2_ASAP7_75t_R _21491_ (.A1(_01879_),
    .A2(_05779_),
    .B1(_05790_),
    .B2(_01929_),
    .C1(_05785_),
    .C2(_01804_),
    .Y(_06597_));
 OA211x2_ASAP7_75t_R _21492_ (.A1(_06595_),
    .A2(_05975_),
    .B(_06596_),
    .C(_06597_),
    .Y(_06598_));
 OA211x2_ASAP7_75t_R _21493_ (.A1(_05963_),
    .A2(_06593_),
    .B(_06594_),
    .C(_06598_),
    .Y(_06599_));
 AOI22x1_ASAP7_75t_R _21494_ (.A1(_05959_),
    .A2(_06589_),
    .B1(_06599_),
    .B2(_18579_),
    .Y(_06600_));
 NOR2x1_ASAP7_75t_R _21495_ (.A(_02159_),
    .B(_06517_),
    .Y(_06601_));
 AO21x1_ASAP7_75t_R _21496_ (.A1(_06514_),
    .A2(_06600_),
    .B(_06601_),
    .Y(_06602_));
 AO21x1_ASAP7_75t_R _21497_ (.A1(_06506_),
    .A2(_06587_),
    .B(_06602_),
    .Y(_02372_));
 INVx1_ASAP7_75t_R _21498_ (.A(_02158_),
    .Y(_06603_));
 OR4x1_ASAP7_75t_R _21499_ (.A(_02159_),
    .B(_02160_),
    .C(_02161_),
    .D(_05823_),
    .Y(_06604_));
 OR2x2_ASAP7_75t_R _21500_ (.A(_06530_),
    .B(_06604_),
    .Y(_06605_));
 NOR2x1_ASAP7_75t_R _21501_ (.A(_06530_),
    .B(_06604_),
    .Y(_06606_));
 AND3x1_ASAP7_75t_R _21502_ (.A(_02158_),
    .B(_06525_),
    .C(_06606_),
    .Y(_06607_));
 AO21x1_ASAP7_75t_R _21503_ (.A1(_06603_),
    .A2(_06605_),
    .B(_06607_),
    .Y(_06608_));
 AND3x1_ASAP7_75t_R _21504_ (.A(_18074_),
    .B(_14965_),
    .C(_14970_),
    .Y(_06609_));
 AO21x1_ASAP7_75t_R _21505_ (.A1(_05960_),
    .A2(_18584_),
    .B(_06609_),
    .Y(_06610_));
 INVx1_ASAP7_75t_R _21506_ (.A(_02066_),
    .Y(_06611_));
 INVx1_ASAP7_75t_R _21507_ (.A(_02129_),
    .Y(_06612_));
 AO32x1_ASAP7_75t_R _21508_ (.A1(_06611_),
    .A2(_06119_),
    .A3(_06066_),
    .B1(_06067_),
    .B2(_06612_),
    .Y(_06613_));
 INVx1_ASAP7_75t_R _21509_ (.A(_02095_),
    .Y(_06614_));
 AO32x2_ASAP7_75t_R _21510_ (.A1(_06614_),
    .A2(_06119_),
    .A3(_05816_),
    .B1(_05827_),
    .B2(_06603_),
    .Y(_06615_));
 AOI22x1_ASAP7_75t_R _21511_ (.A1(_05754_),
    .A2(_06613_),
    .B1(_06615_),
    .B2(_05971_),
    .Y(_06616_));
 OA222x2_ASAP7_75t_R _21512_ (.A1(_01928_),
    .A2(_05790_),
    .B1(_06020_),
    .B2(_02055_),
    .C1(_05831_),
    .C2(_01402_),
    .Y(_06617_));
 OA21x2_ASAP7_75t_R _21513_ (.A1(_01998_),
    .A2(_06005_),
    .B(_06617_),
    .Y(_06618_));
 INVx1_ASAP7_75t_R _21514_ (.A(net111),
    .Y(_06619_));
 OA21x2_ASAP7_75t_R _21515_ (.A1(_01966_),
    .A2(_05782_),
    .B(_05746_),
    .Y(_06620_));
 OA22x2_ASAP7_75t_R _21516_ (.A1(_01878_),
    .A2(_05779_),
    .B1(_05785_),
    .B2(_01803_),
    .Y(_06621_));
 OA211x2_ASAP7_75t_R _21517_ (.A1(_06619_),
    .A2(_05975_),
    .B(_06620_),
    .C(_06621_),
    .Y(_06622_));
 OA211x2_ASAP7_75t_R _21518_ (.A1(_05963_),
    .A2(_06616_),
    .B(_06618_),
    .C(_06622_),
    .Y(_06623_));
 AOI22x1_ASAP7_75t_R _21519_ (.A1(_05959_),
    .A2(_06610_),
    .B1(_06623_),
    .B2(_18584_),
    .Y(_06624_));
 NOR2x1_ASAP7_75t_R _21520_ (.A(_02158_),
    .B(_06517_),
    .Y(_06625_));
 AO21x1_ASAP7_75t_R _21521_ (.A1(_06514_),
    .A2(_06624_),
    .B(_06625_),
    .Y(_06626_));
 AO21x1_ASAP7_75t_R _21522_ (.A1(_06506_),
    .A2(_06608_),
    .B(_06626_),
    .Y(_02373_));
 OR3x1_ASAP7_75t_R _21523_ (.A(_02158_),
    .B(_02159_),
    .C(_06584_),
    .Y(_06627_));
 INVx1_ASAP7_75t_R _21524_ (.A(_06627_),
    .Y(_06628_));
 INVx1_ASAP7_75t_R _21525_ (.A(_02157_),
    .Y(_06629_));
 OR3x1_ASAP7_75t_R _21526_ (.A(_06629_),
    .B(_06509_),
    .C(_06627_),
    .Y(_06630_));
 OAI21x1_ASAP7_75t_R _21527_ (.A1(_02157_),
    .A2(_06628_),
    .B(_06630_),
    .Y(_06631_));
 AND3x1_ASAP7_75t_R _21528_ (.A(_14280_),
    .B(_15024_),
    .C(_15026_),
    .Y(_06632_));
 AO21x1_ASAP7_75t_R _21529_ (.A1(_05846_),
    .A2(_18589_),
    .B(_06632_),
    .Y(_06633_));
 INVx1_ASAP7_75t_R _21530_ (.A(_02065_),
    .Y(_06634_));
 INVx1_ASAP7_75t_R _21531_ (.A(_02128_),
    .Y(_06635_));
 AO32x1_ASAP7_75t_R _21532_ (.A1(_06634_),
    .A2(_18553_),
    .A3(_05816_),
    .B1(_05827_),
    .B2(_06635_),
    .Y(_06636_));
 INVx1_ASAP7_75t_R _21533_ (.A(_02094_),
    .Y(_06637_));
 AO32x1_ASAP7_75t_R _21534_ (.A1(_06637_),
    .A2(_18553_),
    .A3(_05816_),
    .B1(_05827_),
    .B2(_06629_),
    .Y(_06638_));
 AOI22x1_ASAP7_75t_R _21535_ (.A1(_05754_),
    .A2(_06636_),
    .B1(_06638_),
    .B2(_05971_),
    .Y(_06639_));
 OA22x2_ASAP7_75t_R _21536_ (.A1(_02054_),
    .A2(_06020_),
    .B1(_06007_),
    .B2(_01917_),
    .Y(_06640_));
 OA211x2_ASAP7_75t_R _21537_ (.A1(_01927_),
    .A2(_05791_),
    .B(_06640_),
    .C(_05747_),
    .Y(_06641_));
 OA222x2_ASAP7_75t_R _21538_ (.A1(_01802_),
    .A2(_05785_),
    .B1(_05800_),
    .B2(_01997_),
    .C1(_05831_),
    .C2(_02029_),
    .Y(_06642_));
 INVx1_ASAP7_75t_R _21539_ (.A(net112),
    .Y(_06643_));
 INVx1_ASAP7_75t_R _21540_ (.A(net168),
    .Y(_06644_));
 OA222x2_ASAP7_75t_R _21541_ (.A1(_06643_),
    .A2(_05774_),
    .B1(_06045_),
    .B2(_01965_),
    .C1(_06015_),
    .C2(_06644_),
    .Y(_06645_));
 OA22x2_ASAP7_75t_R _21542_ (.A1(_01877_),
    .A2(_05779_),
    .B1(_06018_),
    .B2(_00333_),
    .Y(_06646_));
 AND3x1_ASAP7_75t_R _21543_ (.A(_06642_),
    .B(_06645_),
    .C(_06646_),
    .Y(_06647_));
 OA211x2_ASAP7_75t_R _21544_ (.A1(_05963_),
    .A2(_06639_),
    .B(_06641_),
    .C(_06647_),
    .Y(_06648_));
 AOI22x1_ASAP7_75t_R _21545_ (.A1(_05845_),
    .A2(_06633_),
    .B1(_06648_),
    .B2(_18589_),
    .Y(_06649_));
 BUFx12f_ASAP7_75t_R _21546_ (.A(_06649_),
    .Y(_06650_));
 NOR2x1_ASAP7_75t_R _21547_ (.A(_02157_),
    .B(_06517_),
    .Y(_06651_));
 AO21x1_ASAP7_75t_R _21548_ (.A1(_06514_),
    .A2(_06650_),
    .B(_06651_),
    .Y(_06652_));
 AO21x1_ASAP7_75t_R _21549_ (.A1(_06506_),
    .A2(_06631_),
    .B(_06652_),
    .Y(_02374_));
 INVx1_ASAP7_75t_R _21550_ (.A(_02156_),
    .Y(_06653_));
 OR4x1_ASAP7_75t_R _21551_ (.A(_00747_),
    .B(_05853_),
    .C(_02167_),
    .D(_02178_),
    .Y(_06654_));
 AO21x1_ASAP7_75t_R _21552_ (.A1(_05902_),
    .A2(_06654_),
    .B(_05942_),
    .Y(_06655_));
 INVx1_ASAP7_75t_R _21553_ (.A(_06654_),
    .Y(_06656_));
 AO32x1_ASAP7_75t_R _21554_ (.A1(_02156_),
    .A2(_06159_),
    .A3(_06656_),
    .B1(_06556_),
    .B2(_05945_),
    .Y(_06657_));
 AO21x1_ASAP7_75t_R _21555_ (.A1(_06653_),
    .A2(_06655_),
    .B(_06657_),
    .Y(_02375_));
 INVx1_ASAP7_75t_R _21556_ (.A(_02155_),
    .Y(_06658_));
 OR3x1_ASAP7_75t_R _21557_ (.A(_02157_),
    .B(_02158_),
    .C(_06605_),
    .Y(_06659_));
 AND5x1_ASAP7_75t_R _21558_ (.A(_02155_),
    .B(_06629_),
    .C(_06603_),
    .D(_06585_),
    .E(_06606_),
    .Y(_06660_));
 AO21x1_ASAP7_75t_R _21559_ (.A1(_06658_),
    .A2(_06659_),
    .B(_06660_),
    .Y(_06661_));
 AND2x2_ASAP7_75t_R _21560_ (.A(_18074_),
    .B(_18592_),
    .Y(_06662_));
 AO21x1_ASAP7_75t_R _21561_ (.A1(_05960_),
    .A2(_18594_),
    .B(_06662_),
    .Y(_06663_));
 INVx1_ASAP7_75t_R _21562_ (.A(net113),
    .Y(_06664_));
 OA222x2_ASAP7_75t_R _21563_ (.A1(_06664_),
    .A2(_05975_),
    .B1(_06047_),
    .B2(_01876_),
    .C1(_06045_),
    .C2(_01964_),
    .Y(_06665_));
 OA22x2_ASAP7_75t_R _21564_ (.A1(_01926_),
    .A2(_05791_),
    .B1(_06010_),
    .B2(_02028_),
    .Y(_06666_));
 OA222x2_ASAP7_75t_R _21565_ (.A1(_01801_),
    .A2(_06004_),
    .B1(_06005_),
    .B2(_01996_),
    .C1(_06020_),
    .C2(_02053_),
    .Y(_06667_));
 OA211x2_ASAP7_75t_R _21566_ (.A1(_01403_),
    .A2(_06040_),
    .B(_06667_),
    .C(_05140_),
    .Y(_06668_));
 OAI22x1_ASAP7_75t_R _21567_ (.A1(_02127_),
    .A2(_05964_),
    .B1(_05966_),
    .B2(_02064_),
    .Y(_06669_));
 INVx1_ASAP7_75t_R _21568_ (.A(_02092_),
    .Y(_06670_));
 AO32x1_ASAP7_75t_R _21569_ (.A1(_06670_),
    .A2(_06119_),
    .A3(_06066_),
    .B1(_06067_),
    .B2(_06658_),
    .Y(_06671_));
 AO32x2_ASAP7_75t_R _21570_ (.A1(_06063_),
    .A2(_06064_),
    .A3(_06669_),
    .B1(_06671_),
    .B2(_05763_),
    .Y(_06672_));
 NAND2x1_ASAP7_75t_R _21571_ (.A(_05814_),
    .B(_06672_),
    .Y(_06673_));
 AND4x1_ASAP7_75t_R _21572_ (.A(_06665_),
    .B(_06666_),
    .C(_06668_),
    .D(_06673_),
    .Y(_06674_));
 AOI22x1_ASAP7_75t_R _21573_ (.A1(_05959_),
    .A2(_06663_),
    .B1(_06674_),
    .B2(_18594_),
    .Y(_06675_));
 NOR2x1_ASAP7_75t_R _21574_ (.A(_02155_),
    .B(_06517_),
    .Y(_06676_));
 AO21x1_ASAP7_75t_R _21575_ (.A1(_06514_),
    .A2(_06675_),
    .B(_06676_),
    .Y(_06677_));
 AO21x1_ASAP7_75t_R _21576_ (.A1(_06506_),
    .A2(_06661_),
    .B(_06677_),
    .Y(_02376_));
 OR4x1_ASAP7_75t_R _21577_ (.A(_02155_),
    .B(_02157_),
    .C(_02158_),
    .D(_06604_),
    .Y(_06678_));
 INVx1_ASAP7_75t_R _21578_ (.A(_06678_),
    .Y(_06679_));
 AND3x1_ASAP7_75t_R _21579_ (.A(_06520_),
    .B(_06522_),
    .C(_06679_),
    .Y(_06680_));
 AND2x2_ASAP7_75t_R _21580_ (.A(_02154_),
    .B(_06680_),
    .Y(_06681_));
 NOR2x1_ASAP7_75t_R _21581_ (.A(_02154_),
    .B(_06680_),
    .Y(_06682_));
 AO21x1_ASAP7_75t_R _21582_ (.A1(_06525_),
    .A2(_06681_),
    .B(_06682_),
    .Y(_06683_));
 AND3x1_ASAP7_75t_R _21583_ (.A(_06060_),
    .B(_15157_),
    .C(_15160_),
    .Y(_06684_));
 AO21x1_ASAP7_75t_R _21584_ (.A1(_06059_),
    .A2(_18599_),
    .B(_06684_),
    .Y(_06685_));
 OA21x2_ASAP7_75t_R _21585_ (.A1(_18555_),
    .A2(_05752_),
    .B(_05702_),
    .Y(_06686_));
 AND3x1_ASAP7_75t_R _21586_ (.A(_02063_),
    .B(_18559_),
    .C(_05702_),
    .Y(_06687_));
 AO21x1_ASAP7_75t_R _21587_ (.A1(_02126_),
    .A2(_05921_),
    .B(_06687_),
    .Y(_06688_));
 AND3x1_ASAP7_75t_R _21588_ (.A(_02091_),
    .B(_18559_),
    .C(_05702_),
    .Y(_06689_));
 AO21x1_ASAP7_75t_R _21589_ (.A1(_02154_),
    .A2(_05921_),
    .B(_06689_),
    .Y(_06690_));
 OA22x2_ASAP7_75t_R _21590_ (.A1(_05769_),
    .A2(_06688_),
    .B1(_06690_),
    .B2(_05770_),
    .Y(_06691_));
 OA222x2_ASAP7_75t_R _21591_ (.A1(_01875_),
    .A2(_06047_),
    .B1(_05800_),
    .B2(_01995_),
    .C1(_05831_),
    .C2(_02027_),
    .Y(_06692_));
 INVx1_ASAP7_75t_R _21592_ (.A(net114),
    .Y(_06693_));
 OA21x2_ASAP7_75t_R _21593_ (.A1(_01963_),
    .A2(_05837_),
    .B(_05746_),
    .Y(_06694_));
 OA22x2_ASAP7_75t_R _21594_ (.A1(_01800_),
    .A2(_05839_),
    .B1(_06104_),
    .B2(_01925_),
    .Y(_06695_));
 OA211x2_ASAP7_75t_R _21595_ (.A1(_06693_),
    .A2(_05975_),
    .B(_06694_),
    .C(_06695_),
    .Y(_06696_));
 OA211x2_ASAP7_75t_R _21596_ (.A1(_01404_),
    .A2(_06095_),
    .B(_06692_),
    .C(_06696_),
    .Y(_06697_));
 OA21x2_ASAP7_75t_R _21597_ (.A1(_06686_),
    .A2(_06691_),
    .B(_06697_),
    .Y(_06698_));
 AOI22x1_ASAP7_75t_R _21598_ (.A1(_06058_),
    .A2(_06685_),
    .B1(_06698_),
    .B2(_18599_),
    .Y(_06699_));
 NOR2x1_ASAP7_75t_R _21599_ (.A(_02154_),
    .B(_06517_),
    .Y(_06700_));
 AO21x1_ASAP7_75t_R _21600_ (.A1(_06514_),
    .A2(_06699_),
    .B(_06700_),
    .Y(_06701_));
 AO21x1_ASAP7_75t_R _21601_ (.A1(_06506_),
    .A2(_06683_),
    .B(_06701_),
    .Y(_02377_));
 BUFx6f_ASAP7_75t_R _21602_ (.A(_06159_),
    .Y(_06702_));
 OR3x2_ASAP7_75t_R _21603_ (.A(_02154_),
    .B(_06530_),
    .C(_06678_),
    .Y(_06703_));
 INVx1_ASAP7_75t_R _21604_ (.A(_06703_),
    .Y(_06704_));
 AND3x1_ASAP7_75t_R _21605_ (.A(_02153_),
    .B(_06525_),
    .C(_06704_),
    .Y(_06705_));
 AO21x1_ASAP7_75t_R _21606_ (.A1(_05969_),
    .A2(_06703_),
    .B(_06705_),
    .Y(_06706_));
 BUFx6f_ASAP7_75t_R _21607_ (.A(_06508_),
    .Y(_06707_));
 BUFx12f_ASAP7_75t_R _21608_ (.A(_06516_),
    .Y(_06708_));
 NOR2x1_ASAP7_75t_R _21609_ (.A(_02153_),
    .B(_06708_),
    .Y(_06709_));
 AO21x1_ASAP7_75t_R _21610_ (.A1(_05981_),
    .A2(_06707_),
    .B(_06709_),
    .Y(_06710_));
 AO21x1_ASAP7_75t_R _21611_ (.A1(_06702_),
    .A2(_06706_),
    .B(_06710_),
    .Y(_02378_));
 INVx1_ASAP7_75t_R _21612_ (.A(_05998_),
    .Y(_06711_));
 OR5x2_ASAP7_75t_R _21613_ (.A(_02153_),
    .B(_02154_),
    .C(_06227_),
    .D(_06523_),
    .E(_06678_),
    .Y(_06712_));
 INVx1_ASAP7_75t_R _21614_ (.A(_06712_),
    .Y(_06713_));
 AND3x1_ASAP7_75t_R _21615_ (.A(_05998_),
    .B(_06525_),
    .C(_06713_),
    .Y(_06714_));
 AO21x1_ASAP7_75t_R _21616_ (.A1(_06711_),
    .A2(_06712_),
    .B(_06714_),
    .Y(_06715_));
 NOR2x1_ASAP7_75t_R _21617_ (.A(_05998_),
    .B(_06708_),
    .Y(_06716_));
 AO21x1_ASAP7_75t_R _21618_ (.A1(_06025_),
    .A2(_06707_),
    .B(_06716_),
    .Y(_06717_));
 AO21x1_ASAP7_75t_R _21619_ (.A1(_06702_),
    .A2(_06715_),
    .B(_06717_),
    .Y(_02379_));
 OR3x1_ASAP7_75t_R _21620_ (.A(_05998_),
    .B(_02153_),
    .C(_06703_),
    .Y(_06718_));
 INVx1_ASAP7_75t_R _21621_ (.A(_06718_),
    .Y(_06719_));
 AND3x1_ASAP7_75t_R _21622_ (.A(_02151_),
    .B(_06525_),
    .C(_06719_),
    .Y(_06720_));
 AO21x1_ASAP7_75t_R _21623_ (.A1(_06037_),
    .A2(_06718_),
    .B(_06720_),
    .Y(_06721_));
 NOR2x1_ASAP7_75t_R _21624_ (.A(_02151_),
    .B(_06708_),
    .Y(_06722_));
 AO21x1_ASAP7_75t_R _21625_ (.A1(_06052_),
    .A2(_06707_),
    .B(_06722_),
    .Y(_06723_));
 AO21x1_ASAP7_75t_R _21626_ (.A1(_06702_),
    .A2(_06721_),
    .B(_06723_),
    .Y(_02380_));
 OR3x1_ASAP7_75t_R _21627_ (.A(_02151_),
    .B(_05998_),
    .C(_06712_),
    .Y(_06724_));
 AND5x1_ASAP7_75t_R _21628_ (.A(_02150_),
    .B(_06037_),
    .C(_06711_),
    .D(_06585_),
    .E(_06713_),
    .Y(_06725_));
 AO21x1_ASAP7_75t_R _21629_ (.A1(_06070_),
    .A2(_06724_),
    .B(_06725_),
    .Y(_06726_));
 NOR2x1_ASAP7_75t_R _21630_ (.A(_02150_),
    .B(_06708_),
    .Y(_06727_));
 AO21x1_ASAP7_75t_R _21631_ (.A1(_06082_),
    .A2(_06707_),
    .B(_06727_),
    .Y(_06728_));
 AO21x1_ASAP7_75t_R _21632_ (.A1(_06702_),
    .A2(_06726_),
    .B(_06728_),
    .Y(_02381_));
 INVx1_ASAP7_75t_R _21633_ (.A(_02149_),
    .Y(_06729_));
 OR5x1_ASAP7_75t_R _21634_ (.A(_02150_),
    .B(_02151_),
    .C(_05998_),
    .D(_02153_),
    .E(_06703_),
    .Y(_06730_));
 AND5x1_ASAP7_75t_R _21635_ (.A(_02149_),
    .B(_06070_),
    .C(_06037_),
    .D(_06585_),
    .E(_06719_),
    .Y(_06731_));
 AO21x1_ASAP7_75t_R _21636_ (.A1(_06729_),
    .A2(_06730_),
    .B(_06731_),
    .Y(_06732_));
 NOR2x1_ASAP7_75t_R _21637_ (.A(_02149_),
    .B(_06708_),
    .Y(_06733_));
 AO21x1_ASAP7_75t_R _21638_ (.A1(_06108_),
    .A2(_06707_),
    .B(_06733_),
    .Y(_06734_));
 AO21x1_ASAP7_75t_R _21639_ (.A1(_06702_),
    .A2(_06732_),
    .B(_06734_),
    .Y(_02382_));
 OR3x1_ASAP7_75t_R _21640_ (.A(_02149_),
    .B(_02150_),
    .C(_06724_),
    .Y(_06735_));
 INVx1_ASAP7_75t_R _21641_ (.A(_06735_),
    .Y(_06736_));
 AND3x1_ASAP7_75t_R _21642_ (.A(_02148_),
    .B(_06525_),
    .C(_06736_),
    .Y(_06737_));
 AO21x1_ASAP7_75t_R _21643_ (.A1(_06120_),
    .A2(_06735_),
    .B(_06737_),
    .Y(_06738_));
 NOR2x1_ASAP7_75t_R _21644_ (.A(_02148_),
    .B(_06708_),
    .Y(_06739_));
 AO21x1_ASAP7_75t_R _21645_ (.A1(_06131_),
    .A2(_06707_),
    .B(_06739_),
    .Y(_06740_));
 AO21x1_ASAP7_75t_R _21646_ (.A1(_06702_),
    .A2(_06738_),
    .B(_06740_),
    .Y(_02383_));
 OR3x1_ASAP7_75t_R _21647_ (.A(_02148_),
    .B(_02149_),
    .C(_06730_),
    .Y(_06741_));
 INVx1_ASAP7_75t_R _21648_ (.A(_06741_),
    .Y(_06742_));
 AND3x1_ASAP7_75t_R _21649_ (.A(_02147_),
    .B(_06525_),
    .C(_06742_),
    .Y(_06743_));
 AO21x1_ASAP7_75t_R _21650_ (.A1(_06148_),
    .A2(_06741_),
    .B(_06743_),
    .Y(_06744_));
 NOR2x1_ASAP7_75t_R _21651_ (.A(_02147_),
    .B(_06708_),
    .Y(_06745_));
 AO21x1_ASAP7_75t_R _21652_ (.A1(_06153_),
    .A2(_06707_),
    .B(_06745_),
    .Y(_06746_));
 AO21x1_ASAP7_75t_R _21653_ (.A1(_06702_),
    .A2(_06744_),
    .B(_06746_),
    .Y(_02384_));
 OR3x1_ASAP7_75t_R _21654_ (.A(_02147_),
    .B(_02148_),
    .C(_06735_),
    .Y(_06747_));
 AND5x1_ASAP7_75t_R _21655_ (.A(_02146_),
    .B(_06148_),
    .C(_06120_),
    .D(_06585_),
    .E(_06736_),
    .Y(_06748_));
 AO21x1_ASAP7_75t_R _21656_ (.A1(_06166_),
    .A2(_06747_),
    .B(_06748_),
    .Y(_06749_));
 NOR2x1_ASAP7_75t_R _21657_ (.A(_02146_),
    .B(_06708_),
    .Y(_06750_));
 AO21x1_ASAP7_75t_R _21658_ (.A1(_06179_),
    .A2(_06707_),
    .B(_06750_),
    .Y(_06751_));
 AO21x1_ASAP7_75t_R _21659_ (.A1(_06702_),
    .A2(_06749_),
    .B(_06751_),
    .Y(_02385_));
 OR3x1_ASAP7_75t_R _21660_ (.A(_02156_),
    .B(_02167_),
    .C(_06369_),
    .Y(_06752_));
 AO21x1_ASAP7_75t_R _21661_ (.A1(_05902_),
    .A2(_06752_),
    .B(_05942_),
    .Y(_06753_));
 INVx1_ASAP7_75t_R _21662_ (.A(_06752_),
    .Y(_06754_));
 AO32x1_ASAP7_75t_R _21663_ (.A1(_02145_),
    .A2(_06159_),
    .A3(_06754_),
    .B1(_06580_),
    .B2(_05945_),
    .Y(_06755_));
 AO21x1_ASAP7_75t_R _21664_ (.A1(_06573_),
    .A2(_06753_),
    .B(_06755_),
    .Y(_02386_));
 OR3x1_ASAP7_75t_R _21665_ (.A(_02146_),
    .B(_02147_),
    .C(_06741_),
    .Y(_06756_));
 AND5x1_ASAP7_75t_R _21666_ (.A(_02144_),
    .B(_06166_),
    .C(_06148_),
    .D(_06524_),
    .E(_06742_),
    .Y(_06757_));
 AO21x1_ASAP7_75t_R _21667_ (.A1(_06191_),
    .A2(_06756_),
    .B(_06757_),
    .Y(_06758_));
 NOR2x1_ASAP7_75t_R _21668_ (.A(_02144_),
    .B(_06708_),
    .Y(_06759_));
 AO21x1_ASAP7_75t_R _21669_ (.A1(_06197_),
    .A2(_06707_),
    .B(_06759_),
    .Y(_06760_));
 AO21x1_ASAP7_75t_R _21670_ (.A1(_06702_),
    .A2(_06758_),
    .B(_06760_),
    .Y(_02387_));
 OR3x1_ASAP7_75t_R _21671_ (.A(_02144_),
    .B(_02146_),
    .C(_06747_),
    .Y(_06761_));
 INVx1_ASAP7_75t_R _21672_ (.A(_06761_),
    .Y(_06762_));
 AND3x1_ASAP7_75t_R _21673_ (.A(_02143_),
    .B(_06525_),
    .C(_06762_),
    .Y(_06763_));
 AO21x1_ASAP7_75t_R _21674_ (.A1(_06214_),
    .A2(_06761_),
    .B(_06763_),
    .Y(_06764_));
 NOR2x1_ASAP7_75t_R _21675_ (.A(_02143_),
    .B(_06708_),
    .Y(_06765_));
 AO21x1_ASAP7_75t_R _21676_ (.A1(_06219_),
    .A2(_06707_),
    .B(_06765_),
    .Y(_06766_));
 AO21x1_ASAP7_75t_R _21677_ (.A1(_06702_),
    .A2(_06764_),
    .B(_06766_),
    .Y(_02388_));
 BUFx6f_ASAP7_75t_R _21678_ (.A(_05940_),
    .Y(_06767_));
 OR3x1_ASAP7_75t_R _21679_ (.A(_02143_),
    .B(_02144_),
    .C(_06756_),
    .Y(_06768_));
 INVx1_ASAP7_75t_R _21680_ (.A(_06768_),
    .Y(_06769_));
 AND3x1_ASAP7_75t_R _21681_ (.A(_02142_),
    .B(_06585_),
    .C(_06769_),
    .Y(_06770_));
 AO21x1_ASAP7_75t_R _21682_ (.A1(_06242_),
    .A2(_06768_),
    .B(_06770_),
    .Y(_06771_));
 BUFx6f_ASAP7_75t_R _21683_ (.A(_06508_),
    .Y(_06772_));
 BUFx12f_ASAP7_75t_R _21684_ (.A(_06516_),
    .Y(_06773_));
 NOR2x1_ASAP7_75t_R _21685_ (.A(_02142_),
    .B(_06773_),
    .Y(_06774_));
 AO21x1_ASAP7_75t_R _21686_ (.A1(_06255_),
    .A2(_06772_),
    .B(_06774_),
    .Y(_06775_));
 AO21x1_ASAP7_75t_R _21687_ (.A1(_06767_),
    .A2(_06771_),
    .B(_06775_),
    .Y(_02389_));
 INVx1_ASAP7_75t_R _21688_ (.A(_02141_),
    .Y(_06776_));
 OR3x1_ASAP7_75t_R _21689_ (.A(_02142_),
    .B(_02143_),
    .C(_06761_),
    .Y(_06777_));
 AND5x1_ASAP7_75t_R _21690_ (.A(_02141_),
    .B(_06242_),
    .C(_06214_),
    .D(_06524_),
    .E(_06762_),
    .Y(_06778_));
 AO21x1_ASAP7_75t_R _21691_ (.A1(_06776_),
    .A2(_06777_),
    .B(_06778_),
    .Y(_06779_));
 NOR2x1_ASAP7_75t_R _21692_ (.A(_02141_),
    .B(_06773_),
    .Y(_06780_));
 AO21x1_ASAP7_75t_R _21693_ (.A1(_06277_),
    .A2(_06772_),
    .B(_06780_),
    .Y(_06781_));
 AO21x1_ASAP7_75t_R _21694_ (.A1(_06767_),
    .A2(_06779_),
    .B(_06781_),
    .Y(_02390_));
 OR3x1_ASAP7_75t_R _21695_ (.A(_02141_),
    .B(_02142_),
    .C(_06768_),
    .Y(_06782_));
 AND5x1_ASAP7_75t_R _21696_ (.A(_02140_),
    .B(_06776_),
    .C(_06242_),
    .D(_06524_),
    .E(_06769_),
    .Y(_06783_));
 AO21x1_ASAP7_75t_R _21697_ (.A1(_06292_),
    .A2(_06782_),
    .B(_06783_),
    .Y(_06784_));
 NOR2x1_ASAP7_75t_R _21698_ (.A(_02140_),
    .B(_06773_),
    .Y(_06785_));
 AO21x1_ASAP7_75t_R _21699_ (.A1(_06298_),
    .A2(_06772_),
    .B(_06785_),
    .Y(_06786_));
 AO21x1_ASAP7_75t_R _21700_ (.A1(_06767_),
    .A2(_06784_),
    .B(_06786_),
    .Y(_02391_));
 INVx1_ASAP7_75t_R _21701_ (.A(_06318_),
    .Y(_06787_));
 OR3x2_ASAP7_75t_R _21702_ (.A(_02140_),
    .B(_02141_),
    .C(_06777_),
    .Y(_06788_));
 INVx1_ASAP7_75t_R _21703_ (.A(_06788_),
    .Y(_06789_));
 AND3x1_ASAP7_75t_R _21704_ (.A(_06318_),
    .B(_06585_),
    .C(_06789_),
    .Y(_06790_));
 AO21x1_ASAP7_75t_R _21705_ (.A1(_06787_),
    .A2(_06788_),
    .B(_06790_),
    .Y(_06791_));
 NOR2x1_ASAP7_75t_R _21706_ (.A(_06318_),
    .B(_06773_),
    .Y(_06792_));
 AO21x1_ASAP7_75t_R _21707_ (.A1(_06323_),
    .A2(_06772_),
    .B(_06792_),
    .Y(_06793_));
 AO21x1_ASAP7_75t_R _21708_ (.A1(_06767_),
    .A2(_06791_),
    .B(_06793_),
    .Y(_02392_));
 OR3x1_ASAP7_75t_R _21709_ (.A(_06318_),
    .B(_02140_),
    .C(_06782_),
    .Y(_06794_));
 INVx1_ASAP7_75t_R _21710_ (.A(_06794_),
    .Y(_06795_));
 AND3x1_ASAP7_75t_R _21711_ (.A(_02138_),
    .B(_06585_),
    .C(_06795_),
    .Y(_06796_));
 AO21x1_ASAP7_75t_R _21712_ (.A1(_06338_),
    .A2(_06794_),
    .B(_06796_),
    .Y(_06797_));
 NOR2x1_ASAP7_75t_R _21713_ (.A(_02138_),
    .B(_06773_),
    .Y(_06798_));
 AO21x1_ASAP7_75t_R _21714_ (.A1(_06343_),
    .A2(_06772_),
    .B(_06798_),
    .Y(_06799_));
 AO21x1_ASAP7_75t_R _21715_ (.A1(_06767_),
    .A2(_06797_),
    .B(_06799_),
    .Y(_02393_));
 INVx1_ASAP7_75t_R _21716_ (.A(_02137_),
    .Y(_06800_));
 OR3x1_ASAP7_75t_R _21717_ (.A(_02138_),
    .B(_06318_),
    .C(_06788_),
    .Y(_06801_));
 AND5x1_ASAP7_75t_R _21718_ (.A(_02137_),
    .B(_06338_),
    .C(_06787_),
    .D(_06524_),
    .E(_06789_),
    .Y(_06802_));
 AO21x1_ASAP7_75t_R _21719_ (.A1(_06800_),
    .A2(_06801_),
    .B(_06802_),
    .Y(_06803_));
 NOR2x1_ASAP7_75t_R _21720_ (.A(_02137_),
    .B(_06773_),
    .Y(_06804_));
 AO21x1_ASAP7_75t_R _21721_ (.A1(_06366_),
    .A2(_06772_),
    .B(_06804_),
    .Y(_06805_));
 AO21x1_ASAP7_75t_R _21722_ (.A1(_06767_),
    .A2(_06803_),
    .B(_06805_),
    .Y(_02394_));
 OR3x1_ASAP7_75t_R _21723_ (.A(_02137_),
    .B(_02138_),
    .C(_06794_),
    .Y(_06806_));
 AND5x1_ASAP7_75t_R _21724_ (.A(_02136_),
    .B(_06800_),
    .C(_06338_),
    .D(_06524_),
    .E(_06795_),
    .Y(_06807_));
 AO21x1_ASAP7_75t_R _21725_ (.A1(_06379_),
    .A2(_06806_),
    .B(_06807_),
    .Y(_06808_));
 NOR2x1_ASAP7_75t_R _21726_ (.A(_02136_),
    .B(_06773_),
    .Y(_06809_));
 AO21x1_ASAP7_75t_R _21727_ (.A1(_06391_),
    .A2(_06772_),
    .B(_06809_),
    .Y(_06810_));
 AO21x1_ASAP7_75t_R _21728_ (.A1(_06767_),
    .A2(_06808_),
    .B(_06810_),
    .Y(_02395_));
 INVx1_ASAP7_75t_R _21729_ (.A(_02135_),
    .Y(_06811_));
 OR5x2_ASAP7_75t_R _21730_ (.A(_02136_),
    .B(_02137_),
    .C(_02138_),
    .D(_06318_),
    .E(_06788_),
    .Y(_06812_));
 INVx1_ASAP7_75t_R _21731_ (.A(_06812_),
    .Y(_06813_));
 AND3x1_ASAP7_75t_R _21732_ (.A(_02135_),
    .B(_06585_),
    .C(_06813_),
    .Y(_06814_));
 AO21x1_ASAP7_75t_R _21733_ (.A1(_06811_),
    .A2(_06812_),
    .B(_06814_),
    .Y(_06815_));
 NOR2x1_ASAP7_75t_R _21734_ (.A(_02135_),
    .B(_06773_),
    .Y(_06816_));
 AO21x1_ASAP7_75t_R _21735_ (.A1(_06411_),
    .A2(_06772_),
    .B(_06816_),
    .Y(_06817_));
 AO21x1_ASAP7_75t_R _21736_ (.A1(_06767_),
    .A2(_06815_),
    .B(_06817_),
    .Y(_02396_));
 OR3x1_ASAP7_75t_R _21737_ (.A(_02145_),
    .B(_02156_),
    .C(_06654_),
    .Y(_06818_));
 AO21x1_ASAP7_75t_R _21738_ (.A1(_05940_),
    .A2(_06818_),
    .B(_05941_),
    .Y(_06819_));
 NAND2x1_ASAP7_75t_R _21739_ (.A(_02134_),
    .B(_06819_),
    .Y(_06820_));
 OA211x2_ASAP7_75t_R _21740_ (.A1(_06134_),
    .A2(_06600_),
    .B(_06820_),
    .C(_06083_),
    .Y(_02397_));
 OR3x1_ASAP7_75t_R _21741_ (.A(_02135_),
    .B(_02136_),
    .C(_06806_),
    .Y(_06821_));
 INVx1_ASAP7_75t_R _21742_ (.A(_06821_),
    .Y(_06822_));
 AND3x1_ASAP7_75t_R _21743_ (.A(_02133_),
    .B(_06585_),
    .C(_06822_),
    .Y(_06823_));
 AO21x1_ASAP7_75t_R _21744_ (.A1(_06427_),
    .A2(_06821_),
    .B(_06823_),
    .Y(_06824_));
 NOR2x1_ASAP7_75t_R _21745_ (.A(_02133_),
    .B(_06773_),
    .Y(_06825_));
 AO21x1_ASAP7_75t_R _21746_ (.A1(_06432_),
    .A2(_06772_),
    .B(_06825_),
    .Y(_06826_));
 AO21x1_ASAP7_75t_R _21747_ (.A1(_06767_),
    .A2(_06824_),
    .B(_06826_),
    .Y(_02398_));
 INVx1_ASAP7_75t_R _21748_ (.A(_02132_),
    .Y(_06827_));
 OR3x1_ASAP7_75t_R _21749_ (.A(_02133_),
    .B(_02135_),
    .C(_06812_),
    .Y(_06828_));
 AND5x1_ASAP7_75t_R _21750_ (.A(_02132_),
    .B(_06427_),
    .C(_06811_),
    .D(_06524_),
    .E(_06813_),
    .Y(_06829_));
 AO21x1_ASAP7_75t_R _21751_ (.A1(_06827_),
    .A2(_06828_),
    .B(_06829_),
    .Y(_06830_));
 NOR2x1_ASAP7_75t_R _21752_ (.A(_02132_),
    .B(_06773_),
    .Y(_06831_));
 AO21x1_ASAP7_75t_R _21753_ (.A1(_06454_),
    .A2(_06772_),
    .B(_06831_),
    .Y(_06832_));
 AO21x1_ASAP7_75t_R _21754_ (.A1(_06767_),
    .A2(_06830_),
    .B(_06832_),
    .Y(_02399_));
 AND3x1_ASAP7_75t_R _21755_ (.A(_06827_),
    .B(_06427_),
    .C(_06822_),
    .Y(_06833_));
 OR5x1_ASAP7_75t_R _21756_ (.A(_06468_),
    .B(_02132_),
    .C(_02133_),
    .D(_06509_),
    .E(_06821_),
    .Y(_06834_));
 OAI21x1_ASAP7_75t_R _21757_ (.A1(_02131_),
    .A2(_06833_),
    .B(_06834_),
    .Y(_06835_));
 NOR2x1_ASAP7_75t_R _21758_ (.A(_02131_),
    .B(_06516_),
    .Y(_06836_));
 AO21x1_ASAP7_75t_R _21759_ (.A1(_06480_),
    .A2(_06508_),
    .B(_06836_),
    .Y(_06837_));
 AO21x1_ASAP7_75t_R _21760_ (.A1(_05948_),
    .A2(_06835_),
    .B(_06837_),
    .Y(_02400_));
 AND5x1_ASAP7_75t_R _21761_ (.A(_06468_),
    .B(_06827_),
    .C(_06427_),
    .D(_06811_),
    .E(_06813_),
    .Y(_06838_));
 OR5x1_ASAP7_75t_R _21762_ (.A(_06492_),
    .B(_02131_),
    .C(_02132_),
    .D(_06509_),
    .E(_06828_),
    .Y(_06839_));
 OAI21x1_ASAP7_75t_R _21763_ (.A1(_02130_),
    .A2(_06838_),
    .B(_06839_),
    .Y(_06840_));
 NOR2x1_ASAP7_75t_R _21764_ (.A(_02130_),
    .B(_06516_),
    .Y(_06841_));
 AO21x1_ASAP7_75t_R _21765_ (.A1(_06504_),
    .A2(_06508_),
    .B(_06841_),
    .Y(_06842_));
 AO21x1_ASAP7_75t_R _21766_ (.A1(_05948_),
    .A2(_06840_),
    .B(_06842_),
    .Y(_02401_));
 AO21x1_ASAP7_75t_R _21767_ (.A1(_05902_),
    .A2(_05950_),
    .B(_05942_),
    .Y(_06843_));
 AO32x1_ASAP7_75t_R _21768_ (.A1(_05907_),
    .A2(_06278_),
    .A3(_06624_),
    .B1(_05958_),
    .B2(_02129_),
    .Y(_06844_));
 AO21x1_ASAP7_75t_R _21769_ (.A1(_06612_),
    .A2(_06843_),
    .B(_06844_),
    .Y(_02402_));
 OA211x2_ASAP7_75t_R _21770_ (.A1(_02129_),
    .A2(_06083_),
    .B(_06133_),
    .C(_06635_),
    .Y(_06845_));
 INVx1_ASAP7_75t_R _21771_ (.A(_06083_),
    .Y(_06846_));
 AO32x1_ASAP7_75t_R _21772_ (.A1(_02128_),
    .A2(_06612_),
    .A3(_06846_),
    .B1(_06650_),
    .B2(_05944_),
    .Y(_06847_));
 OR2x2_ASAP7_75t_R _21773_ (.A(_06845_),
    .B(_06847_),
    .Y(_02403_));
 OR3x1_ASAP7_75t_R _21774_ (.A(_02128_),
    .B(_02129_),
    .C(_06299_),
    .Y(_06848_));
 NOR2x1_ASAP7_75t_R _21775_ (.A(_02127_),
    .B(_06327_),
    .Y(_06849_));
 INVx1_ASAP7_75t_R _21776_ (.A(_06848_),
    .Y(_06850_));
 AO32x1_ASAP7_75t_R _21777_ (.A1(_05907_),
    .A2(_06278_),
    .A3(_06675_),
    .B1(_06850_),
    .B2(_02127_),
    .Y(_06851_));
 AO21x1_ASAP7_75t_R _21778_ (.A1(_06848_),
    .A2(_06849_),
    .B(_06851_),
    .Y(_02404_));
 NOR2x1_ASAP7_75t_R _21779_ (.A(_05952_),
    .B(_06083_),
    .Y(_06852_));
 INVx1_ASAP7_75t_R _21780_ (.A(_02126_),
    .Y(_06853_));
 OA211x2_ASAP7_75t_R _21781_ (.A1(_05952_),
    .A2(_06083_),
    .B(_06853_),
    .C(_06133_),
    .Y(_06854_));
 AO221x1_ASAP7_75t_R _21782_ (.A1(_06327_),
    .A2(_06699_),
    .B1(_06852_),
    .B2(_02126_),
    .C(_06854_),
    .Y(_02405_));
 NAND2x1_ASAP7_75t_R _21783_ (.A(_14588_),
    .B(_14544_),
    .Y(_06855_));
 OR3x1_ASAP7_75t_R _21784_ (.A(_02222_),
    .B(_14603_),
    .C(_06855_),
    .Y(_06856_));
 AO21x2_ASAP7_75t_R _21785_ (.A1(_05229_),
    .A2(_05230_),
    .B(_06856_),
    .Y(_06857_));
 AND2x4_ASAP7_75t_R _21786_ (.A(net1975),
    .B(_01389_),
    .Y(_06858_));
 AND3x1_ASAP7_75t_R _21787_ (.A(_14580_),
    .B(_14587_),
    .C(_14598_),
    .Y(_06859_));
 BUFx6f_ASAP7_75t_R _21788_ (.A(_06859_),
    .Y(_06860_));
 OAI22x1_ASAP7_75t_R _21789_ (.A1(net1974),
    .A2(_14603_),
    .B1(_06858_),
    .B2(_06860_),
    .Y(_06861_));
 NAND2x1_ASAP7_75t_R _21790_ (.A(_06860_),
    .B(_14605_),
    .Y(_06862_));
 AO21x1_ASAP7_75t_R _21791_ (.A1(net1975),
    .A2(_06862_),
    .B(net1974),
    .Y(_06863_));
 OR2x2_ASAP7_75t_R _21792_ (.A(net1975),
    .B(_14604_),
    .Y(_06864_));
 AND4x1_ASAP7_75t_R _21793_ (.A(_14566_),
    .B(_14580_),
    .C(_14587_),
    .D(_14590_),
    .Y(_06865_));
 AO21x1_ASAP7_75t_R _21794_ (.A1(_06863_),
    .A2(_06864_),
    .B(_06865_),
    .Y(_06866_));
 XNOR2x2_ASAP7_75t_R _21795_ (.A(_18072_),
    .B(_06866_),
    .Y(_06867_));
 NOR2x1_ASAP7_75t_R _21796_ (.A(_01390_),
    .B(_06867_),
    .Y(_06868_));
 AO221x1_ASAP7_75t_R _21797_ (.A1(_01390_),
    .A2(\alu_adder_result_ex[31] ),
    .B1(_06861_),
    .B2(_14605_),
    .C(_06868_),
    .Y(_06869_));
 INVx1_ASAP7_75t_R _21798_ (.A(_01390_),
    .Y(_06870_));
 NOR3x1_ASAP7_75t_R _21799_ (.A(_14576_),
    .B(_14609_),
    .C(_14617_),
    .Y(_06871_));
 OR5x1_ASAP7_75t_R _21800_ (.A(_02221_),
    .B(_14576_),
    .C(_14609_),
    .D(_14614_),
    .E(_14615_),
    .Y(_06872_));
 OA21x2_ASAP7_75t_R _21801_ (.A1(_02222_),
    .A2(_06860_),
    .B(_06872_),
    .Y(_06873_));
 OA22x2_ASAP7_75t_R _21802_ (.A1(_06871_),
    .A2(_06858_),
    .B1(_06873_),
    .B2(_06855_),
    .Y(_06874_));
 OR3x1_ASAP7_75t_R _21803_ (.A(_14603_),
    .B(_06855_),
    .C(_06858_),
    .Y(_06875_));
 NAND2x1_ASAP7_75t_R _21804_ (.A(_06874_),
    .B(_06875_),
    .Y(_06876_));
 OR2x2_ASAP7_75t_R _21805_ (.A(_06870_),
    .B(_06876_),
    .Y(_06877_));
 OR3x1_ASAP7_75t_R _21806_ (.A(_01390_),
    .B(_06867_),
    .C(_06876_),
    .Y(_06878_));
 OA21x2_ASAP7_75t_R _21807_ (.A1(net1952),
    .A2(_06877_),
    .B(_06878_),
    .Y(_06879_));
 NOR2x1_ASAP7_75t_R _21808_ (.A(_02222_),
    .B(_14603_),
    .Y(_06880_));
 AND2x4_ASAP7_75t_R _21809_ (.A(_14605_),
    .B(_06880_),
    .Y(_06881_));
 AOI22x1_ASAP7_75t_R _21810_ (.A1(_06869_),
    .A2(_06879_),
    .B1(_06881_),
    .B2(_05232_),
    .Y(_06882_));
 NAND2x2_ASAP7_75t_R _21811_ (.A(_13235_),
    .B(_05192_),
    .Y(_06883_));
 OR2x6_ASAP7_75t_R _21812_ (.A(_14592_),
    .B(_06883_),
    .Y(_06884_));
 AOI21x1_ASAP7_75t_R _21813_ (.A1(_06857_),
    .A2(_06882_),
    .B(_06884_),
    .Y(_06885_));
 AOI211x1_ASAP7_75t_R _21814_ (.A1(_14605_),
    .A2(_06861_),
    .B(_06876_),
    .C(_06881_),
    .Y(_06886_));
 AND5x1_ASAP7_75t_R _21815_ (.A(_04246_),
    .B(_04729_),
    .C(net1952),
    .D(_04983_),
    .E(_06886_),
    .Y(_06887_));
 NAND3x1_ASAP7_75t_R _21816_ (.A(_05229_),
    .B(_05230_),
    .C(_06887_),
    .Y(_06888_));
 NAND2x1_ASAP7_75t_R _21817_ (.A(_05730_),
    .B(_04987_),
    .Y(_06889_));
 OA211x2_ASAP7_75t_R _21818_ (.A1(_02194_),
    .A2(_14119_),
    .B(_02199_),
    .C(_01397_),
    .Y(_06890_));
 NAND2x1_ASAP7_75t_R _21819_ (.A(_14623_),
    .B(_06890_),
    .Y(_06891_));
 OAI21x1_ASAP7_75t_R _21820_ (.A1(_05181_),
    .A2(_06889_),
    .B(_06891_),
    .Y(_06892_));
 AO21x1_ASAP7_75t_R _21821_ (.A1(_14623_),
    .A2(_06890_),
    .B(_13294_),
    .Y(_06893_));
 OR3x1_ASAP7_75t_R _21822_ (.A(_13235_),
    .B(_14543_),
    .C(_14623_),
    .Y(_06894_));
 AO21x1_ASAP7_75t_R _21823_ (.A1(_06893_),
    .A2(_06894_),
    .B(_05395_),
    .Y(_06895_));
 AO32x1_ASAP7_75t_R _21824_ (.A1(_13234_),
    .A2(_05730_),
    .A3(_04987_),
    .B1(_05192_),
    .B2(_06895_),
    .Y(_06896_));
 OA21x2_ASAP7_75t_R _21825_ (.A1(_13235_),
    .A2(_06892_),
    .B(_06896_),
    .Y(_06897_));
 INVx1_ASAP7_75t_R _21826_ (.A(_06897_),
    .Y(_06898_));
 OAI21x1_ASAP7_75t_R _21827_ (.A1(_06888_),
    .A2(_06884_),
    .B(_06898_),
    .Y(_06899_));
 NOR3x1_ASAP7_75t_R _21828_ (.A(_05102_),
    .B(_05111_),
    .C(_05124_),
    .Y(_06900_));
 OA21x2_ASAP7_75t_R _21829_ (.A1(_05104_),
    .A2(_05135_),
    .B(_05140_),
    .Y(_06901_));
 NAND2x1_ASAP7_75t_R _21830_ (.A(_05142_),
    .B(_05146_),
    .Y(_06902_));
 AND5x2_ASAP7_75t_R _21831_ (.A(_05769_),
    .B(_05908_),
    .C(_06900_),
    .D(_06901_),
    .E(_06902_),
    .Y(_06903_));
 OA21x2_ASAP7_75t_R _21832_ (.A1(_05935_),
    .A2(_06903_),
    .B(_14120_),
    .Y(_06904_));
 NAND2x2_ASAP7_75t_R _21833_ (.A(_04987_),
    .B(_05191_),
    .Y(_06905_));
 AND3x4_ASAP7_75t_R _21834_ (.A(_05897_),
    .B(_05768_),
    .C(_05901_),
    .Y(_06906_));
 INVx1_ASAP7_75t_R _21835_ (.A(_02189_),
    .Y(_06907_));
 INVx1_ASAP7_75t_R _21836_ (.A(_05184_),
    .Y(_06908_));
 OR3x1_ASAP7_75t_R _21837_ (.A(_05152_),
    .B(_06907_),
    .C(_06908_),
    .Y(_06909_));
 AND3x1_ASAP7_75t_R _21838_ (.A(_13228_),
    .B(_13265_),
    .C(_14103_),
    .Y(_06910_));
 OR2x2_ASAP7_75t_R _21839_ (.A(_06909_),
    .B(_06910_),
    .Y(_06911_));
 AND3x1_ASAP7_75t_R _21840_ (.A(_02228_),
    .B(_14120_),
    .C(_05119_),
    .Y(_06912_));
 OR5x2_ASAP7_75t_R _21841_ (.A(_06904_),
    .B(_06905_),
    .C(_06906_),
    .D(_06911_),
    .E(_06912_),
    .Y(_06913_));
 OR3x2_ASAP7_75t_R _21842_ (.A(_06885_),
    .B(_06899_),
    .C(_06913_),
    .Y(_06914_));
 BUFx6f_ASAP7_75t_R _21843_ (.A(_06914_),
    .Y(_06915_));
 AND2x6_ASAP7_75t_R _21844_ (.A(_05768_),
    .B(_05939_),
    .Y(_06916_));
 NAND2x1_ASAP7_75t_R _21845_ (.A(_05907_),
    .B(_06916_),
    .Y(_06917_));
 AND2x2_ASAP7_75t_R _21846_ (.A(_06915_),
    .B(_06917_),
    .Y(_06918_));
 NOR3x1_ASAP7_75t_R _21847_ (.A(_06885_),
    .B(_06899_),
    .C(_06913_),
    .Y(_06919_));
 BUFx6f_ASAP7_75t_R _21848_ (.A(_06919_),
    .Y(_06920_));
 BUFx6f_ASAP7_75t_R _21849_ (.A(_06920_),
    .Y(_06921_));
 AO32x1_ASAP7_75t_R _21850_ (.A1(_05907_),
    .A2(_05811_),
    .A3(_06916_),
    .B1(_06921_),
    .B2(_00748_),
    .Y(_06922_));
 AO21x1_ASAP7_75t_R _21851_ (.A1(\cs_registers_i.mhpmcounter[1856] ),
    .A2(_06918_),
    .B(_06922_),
    .Y(_02406_));
 INVx2_ASAP7_75t_R _21852_ (.A(_05981_),
    .Y(_06923_));
 BUFx12f_ASAP7_75t_R _21853_ (.A(_06917_),
    .Y(_06924_));
 BUFx12f_ASAP7_75t_R _21854_ (.A(_06924_),
    .Y(_06925_));
 OR4x1_ASAP7_75t_R _21855_ (.A(_02063_),
    .B(_02064_),
    .C(_02065_),
    .D(_02066_),
    .Y(_06926_));
 OR4x1_ASAP7_75t_R _21856_ (.A(_02071_),
    .B(_02082_),
    .C(_02093_),
    .D(_02104_),
    .Y(_06927_));
 OR5x2_ASAP7_75t_R _21857_ (.A(_02232_),
    .B(_06885_),
    .C(_06899_),
    .D(_06913_),
    .E(_06927_),
    .Y(_06928_));
 OA21x2_ASAP7_75t_R _21858_ (.A1(_06926_),
    .A2(_06928_),
    .B(_02125_),
    .Y(_06929_));
 NOR2x1_ASAP7_75t_R _21859_ (.A(_05907_),
    .B(_06920_),
    .Y(_06930_));
 BUFx6f_ASAP7_75t_R _21860_ (.A(_06930_),
    .Y(_06931_));
 NAND2x1_ASAP7_75t_R _21861_ (.A(_05766_),
    .B(_05767_),
    .Y(_06932_));
 OR3x2_ASAP7_75t_R _21862_ (.A(_06932_),
    .B(_05937_),
    .C(_05938_),
    .Y(_06933_));
 BUFx6f_ASAP7_75t_R _21863_ (.A(_06933_),
    .Y(_06934_));
 OA21x2_ASAP7_75t_R _21864_ (.A1(_06926_),
    .A2(_06928_),
    .B(_06934_),
    .Y(_06935_));
 NOR3x1_ASAP7_75t_R _21865_ (.A(_02125_),
    .B(_06931_),
    .C(_06935_),
    .Y(_06936_));
 OAI22x1_ASAP7_75t_R _21866_ (.A1(_06923_),
    .A2(_06925_),
    .B1(_06929_),
    .B2(_06936_),
    .Y(_02407_));
 INVx4_ASAP7_75t_R _21867_ (.A(_06024_),
    .Y(_06937_));
 BUFx6f_ASAP7_75t_R _21868_ (.A(_06919_),
    .Y(_06938_));
 INVx2_ASAP7_75t_R _21869_ (.A(_02071_),
    .Y(_06939_));
 NOR2x1_ASAP7_75t_R _21870_ (.A(_02093_),
    .B(_02104_),
    .Y(_06940_));
 AND3x4_ASAP7_75t_R _21871_ (.A(_06939_),
    .B(_06572_),
    .C(_06940_),
    .Y(_06941_));
 OR5x2_ASAP7_75t_R _21872_ (.A(_02063_),
    .B(_02064_),
    .C(_02065_),
    .D(_02066_),
    .E(_02125_),
    .Y(_06942_));
 INVx1_ASAP7_75t_R _21873_ (.A(_06942_),
    .Y(_06943_));
 NOR2x2_ASAP7_75t_R _21874_ (.A(_00748_),
    .B(_02115_),
    .Y(_06944_));
 AND4x1_ASAP7_75t_R _21875_ (.A(_06938_),
    .B(_06941_),
    .C(_06943_),
    .D(_06944_),
    .Y(_06945_));
 NOR2x1_ASAP7_75t_R _21876_ (.A(_05993_),
    .B(_06945_),
    .Y(_06946_));
 BUFx6f_ASAP7_75t_R _21877_ (.A(_06916_),
    .Y(_06947_));
 OR2x6_ASAP7_75t_R _21878_ (.A(_05907_),
    .B(_06920_),
    .Y(_06948_));
 BUFx6f_ASAP7_75t_R _21879_ (.A(_06948_),
    .Y(_06949_));
 OA211x2_ASAP7_75t_R _21880_ (.A1(_06947_),
    .A2(_06945_),
    .B(_06949_),
    .C(_05993_),
    .Y(_06950_));
 OAI22x1_ASAP7_75t_R _21881_ (.A1(_06937_),
    .A2(_06925_),
    .B1(_06946_),
    .B2(_06950_),
    .Y(_02408_));
 AND3x4_ASAP7_75t_R _21882_ (.A(_05768_),
    .B(_05907_),
    .C(_05939_),
    .Y(_06951_));
 OR2x2_ASAP7_75t_R _21883_ (.A(_02124_),
    .B(_06942_),
    .Y(_06952_));
 OAI21x1_ASAP7_75t_R _21884_ (.A1(_06928_),
    .A2(_06952_),
    .B(_02123_),
    .Y(_06953_));
 OA21x2_ASAP7_75t_R _21885_ (.A1(_06928_),
    .A2(_06952_),
    .B(_06933_),
    .Y(_06954_));
 OR3x1_ASAP7_75t_R _21886_ (.A(_02123_),
    .B(_06930_),
    .C(_06954_),
    .Y(_06955_));
 AO22x1_ASAP7_75t_R _21887_ (.A1(_06052_),
    .A2(_06951_),
    .B1(_06953_),
    .B2(_06955_),
    .Y(_02409_));
 BUFx6f_ASAP7_75t_R _21888_ (.A(_06933_),
    .Y(_06956_));
 OR2x2_ASAP7_75t_R _21889_ (.A(_00748_),
    .B(_02115_),
    .Y(_06957_));
 OR5x2_ASAP7_75t_R _21890_ (.A(_02123_),
    .B(_02124_),
    .C(_06927_),
    .D(_06942_),
    .E(_06957_),
    .Y(_06958_));
 OR2x2_ASAP7_75t_R _21891_ (.A(_06914_),
    .B(_06958_),
    .Y(_06959_));
 AO21x1_ASAP7_75t_R _21892_ (.A1(_06956_),
    .A2(_06959_),
    .B(_06931_),
    .Y(_06960_));
 INVx3_ASAP7_75t_R _21893_ (.A(_06082_),
    .Y(_06961_));
 OAI22x1_ASAP7_75t_R _21894_ (.A1(_06961_),
    .A2(_06924_),
    .B1(_06959_),
    .B2(_06065_),
    .Y(_06962_));
 AO21x1_ASAP7_75t_R _21895_ (.A1(_06065_),
    .A2(_06960_),
    .B(_06962_),
    .Y(_02410_));
 OR4x1_ASAP7_75t_R _21896_ (.A(_02123_),
    .B(_02124_),
    .C(_06927_),
    .D(_06942_),
    .Y(_06963_));
 OR2x6_ASAP7_75t_R _21897_ (.A(_02232_),
    .B(_06963_),
    .Y(_06964_));
 OR3x1_ASAP7_75t_R _21898_ (.A(_02122_),
    .B(_06914_),
    .C(_06964_),
    .Y(_06965_));
 AO21x1_ASAP7_75t_R _21899_ (.A1(_06934_),
    .A2(_06965_),
    .B(_06931_),
    .Y(_06966_));
 NOR2x1_ASAP7_75t_R _21900_ (.A(_06096_),
    .B(_06965_),
    .Y(_06967_));
 AO221x1_ASAP7_75t_R _21901_ (.A1(_06108_),
    .A2(_06951_),
    .B1(_06966_),
    .B2(_06096_),
    .C(_06967_),
    .Y(_02411_));
 INVx3_ASAP7_75t_R _21902_ (.A(_06131_),
    .Y(_06968_));
 OR4x1_ASAP7_75t_R _21903_ (.A(_02121_),
    .B(_02122_),
    .C(_06914_),
    .D(_06958_),
    .Y(_06969_));
 AND2x2_ASAP7_75t_R _21904_ (.A(_02120_),
    .B(_06969_),
    .Y(_06970_));
 BUFx6f_ASAP7_75t_R _21905_ (.A(_06934_),
    .Y(_06971_));
 AOI211x1_ASAP7_75t_R _21906_ (.A1(_06971_),
    .A2(_06969_),
    .B(_06931_),
    .C(_02120_),
    .Y(_06972_));
 OAI22x1_ASAP7_75t_R _21907_ (.A1(_06968_),
    .A2(_06925_),
    .B1(_06970_),
    .B2(_06972_),
    .Y(_02412_));
 INVx3_ASAP7_75t_R _21908_ (.A(_06153_),
    .Y(_06973_));
 OR3x1_ASAP7_75t_R _21909_ (.A(_02120_),
    .B(_02121_),
    .C(_02122_),
    .Y(_06974_));
 OR3x1_ASAP7_75t_R _21910_ (.A(_06915_),
    .B(_06964_),
    .C(_06974_),
    .Y(_06975_));
 AND2x2_ASAP7_75t_R _21911_ (.A(_02119_),
    .B(_06975_),
    .Y(_06976_));
 AOI211x1_ASAP7_75t_R _21912_ (.A1(_06971_),
    .A2(_06975_),
    .B(_06931_),
    .C(_02119_),
    .Y(_06977_));
 OAI22x1_ASAP7_75t_R _21913_ (.A1(_06973_),
    .A2(_06925_),
    .B1(_06976_),
    .B2(_06977_),
    .Y(_02413_));
 INVx3_ASAP7_75t_R _21914_ (.A(_06178_),
    .Y(_06978_));
 BUFx6f_ASAP7_75t_R _21915_ (.A(_06920_),
    .Y(_06979_));
 OR3x1_ASAP7_75t_R _21916_ (.A(_02119_),
    .B(_06963_),
    .C(_06974_),
    .Y(_06980_));
 INVx1_ASAP7_75t_R _21917_ (.A(_06980_),
    .Y(_06981_));
 AND3x1_ASAP7_75t_R _21918_ (.A(_06979_),
    .B(_06944_),
    .C(_06981_),
    .Y(_06982_));
 NOR2x1_ASAP7_75t_R _21919_ (.A(_06163_),
    .B(_06982_),
    .Y(_06983_));
 OA211x2_ASAP7_75t_R _21920_ (.A1(_06947_),
    .A2(_06982_),
    .B(_06949_),
    .C(_06163_),
    .Y(_06984_));
 OAI22x1_ASAP7_75t_R _21921_ (.A1(_06978_),
    .A2(_06925_),
    .B1(_06983_),
    .B2(_06984_),
    .Y(_02414_));
 NOR2x1_ASAP7_75t_R _21922_ (.A(_05882_),
    .B(_05900_),
    .Y(_06985_));
 AND2x4_ASAP7_75t_R _21923_ (.A(_06985_),
    .B(_06906_),
    .Y(_06986_));
 BUFx6f_ASAP7_75t_R _21924_ (.A(_06938_),
    .Y(_06987_));
 NOR2x1_ASAP7_75t_R _21925_ (.A(_06985_),
    .B(_06987_),
    .Y(_06988_));
 INVx1_ASAP7_75t_R _21926_ (.A(_06188_),
    .Y(_06989_));
 OR5x2_ASAP7_75t_R _21927_ (.A(_02118_),
    .B(_02119_),
    .C(_02120_),
    .D(_02121_),
    .E(_02122_),
    .Y(_06990_));
 NOR2x1_ASAP7_75t_R _21928_ (.A(_06964_),
    .B(_06990_),
    .Y(_06991_));
 AOI211x1_ASAP7_75t_R _21929_ (.A1(_06938_),
    .A2(_06991_),
    .B(_06188_),
    .C(_06906_),
    .Y(_06992_));
 AND3x1_ASAP7_75t_R _21930_ (.A(_06188_),
    .B(_06938_),
    .C(_06991_),
    .Y(_06993_));
 OR2x2_ASAP7_75t_R _21931_ (.A(_06992_),
    .B(_06993_),
    .Y(_06994_));
 AO221x1_ASAP7_75t_R _21932_ (.A1(_06197_),
    .A2(_06986_),
    .B1(_06988_),
    .B2(_06989_),
    .C(_06994_),
    .Y(_02415_));
 INVx4_ASAP7_75t_R _21933_ (.A(_06219_),
    .Y(_06995_));
 OR4x1_ASAP7_75t_R _21934_ (.A(_06188_),
    .B(_06915_),
    .C(_06958_),
    .D(_06990_),
    .Y(_06996_));
 AND2x2_ASAP7_75t_R _21935_ (.A(_02116_),
    .B(_06996_),
    .Y(_06997_));
 AOI211x1_ASAP7_75t_R _21936_ (.A1(_06971_),
    .A2(_06996_),
    .B(_06931_),
    .C(_02116_),
    .Y(_06998_));
 OAI22x1_ASAP7_75t_R _21937_ (.A1(_06995_),
    .A2(_06925_),
    .B1(_06997_),
    .B2(_06998_),
    .Y(_02416_));
 NAND2x1_ASAP7_75t_R _21938_ (.A(_06235_),
    .B(_06951_),
    .Y(_06999_));
 OA211x2_ASAP7_75t_R _21939_ (.A1(_02115_),
    .A2(_06951_),
    .B(_06999_),
    .C(_06915_),
    .Y(_07000_));
 AOI21x1_ASAP7_75t_R _21940_ (.A1(_02233_),
    .A2(_06987_),
    .B(_07000_),
    .Y(_02417_));
 INVx1_ASAP7_75t_R _21941_ (.A(_06255_),
    .Y(_07001_));
 OR3x1_ASAP7_75t_R _21942_ (.A(_02116_),
    .B(_06188_),
    .C(_06990_),
    .Y(_07002_));
 OR3x1_ASAP7_75t_R _21943_ (.A(_06915_),
    .B(_06964_),
    .C(_07002_),
    .Y(_07003_));
 AND2x2_ASAP7_75t_R _21944_ (.A(_02114_),
    .B(_07003_),
    .Y(_07004_));
 AOI211x1_ASAP7_75t_R _21945_ (.A1(_06971_),
    .A2(_07003_),
    .B(_06931_),
    .C(_02114_),
    .Y(_07005_));
 OAI22x1_ASAP7_75t_R _21946_ (.A1(_07001_),
    .A2(_06925_),
    .B1(_07004_),
    .B2(_07005_),
    .Y(_02418_));
 INVx3_ASAP7_75t_R _21947_ (.A(_06276_),
    .Y(_07006_));
 OR4x1_ASAP7_75t_R _21948_ (.A(_02114_),
    .B(_06915_),
    .C(_06958_),
    .D(_07002_),
    .Y(_07007_));
 AND2x2_ASAP7_75t_R _21949_ (.A(_02113_),
    .B(_07007_),
    .Y(_07008_));
 AOI211x1_ASAP7_75t_R _21950_ (.A1(_06971_),
    .A2(_07007_),
    .B(_06931_),
    .C(_02113_),
    .Y(_07009_));
 OAI22x1_ASAP7_75t_R _21951_ (.A1(_07006_),
    .A2(_06925_),
    .B1(_07008_),
    .B2(_07009_),
    .Y(_02419_));
 INVx1_ASAP7_75t_R _21952_ (.A(_02112_),
    .Y(_07010_));
 OR5x2_ASAP7_75t_R _21953_ (.A(_02113_),
    .B(_02114_),
    .C(_02116_),
    .D(_06188_),
    .E(_06990_),
    .Y(_07011_));
 NOR2x1_ASAP7_75t_R _21954_ (.A(_06964_),
    .B(_07011_),
    .Y(_07012_));
 AND2x4_ASAP7_75t_R _21955_ (.A(_06921_),
    .B(_07012_),
    .Y(_07013_));
 OAI21x1_ASAP7_75t_R _21956_ (.A1(_06947_),
    .A2(_07013_),
    .B(_06949_),
    .Y(_07014_));
 AO32x1_ASAP7_75t_R _21957_ (.A1(_02112_),
    .A2(_06987_),
    .A3(_07012_),
    .B1(_06951_),
    .B2(_06298_),
    .Y(_07015_));
 AO21x1_ASAP7_75t_R _21958_ (.A1(_07010_),
    .A2(_07014_),
    .B(_07015_),
    .Y(_02420_));
 INVx3_ASAP7_75t_R _21959_ (.A(_06323_),
    .Y(_07016_));
 NOR2x1_ASAP7_75t_R _21960_ (.A(_06958_),
    .B(_07011_),
    .Y(_07017_));
 AND3x1_ASAP7_75t_R _21961_ (.A(_07010_),
    .B(_06979_),
    .C(_07017_),
    .Y(_07018_));
 NOR2x1_ASAP7_75t_R _21962_ (.A(_06316_),
    .B(_07018_),
    .Y(_07019_));
 OA211x2_ASAP7_75t_R _21963_ (.A1(_06947_),
    .A2(_07018_),
    .B(_06949_),
    .C(_06316_),
    .Y(_07020_));
 OAI22x1_ASAP7_75t_R _21964_ (.A1(_07016_),
    .A2(_06925_),
    .B1(_07019_),
    .B2(_07020_),
    .Y(_02421_));
 INVx1_ASAP7_75t_R _21965_ (.A(_02110_),
    .Y(_07021_));
 NOR2x1_ASAP7_75t_R _21966_ (.A(_02111_),
    .B(_02112_),
    .Y(_07022_));
 AND3x1_ASAP7_75t_R _21967_ (.A(_06979_),
    .B(_07012_),
    .C(_07022_),
    .Y(_07023_));
 NOR2x1_ASAP7_75t_R _21968_ (.A(_07021_),
    .B(_07023_),
    .Y(_07024_));
 OA211x2_ASAP7_75t_R _21969_ (.A1(_06947_),
    .A2(_07023_),
    .B(_06949_),
    .C(_07021_),
    .Y(_07025_));
 OAI22x1_ASAP7_75t_R _21970_ (.A1(_06344_),
    .A2(_06925_),
    .B1(_07024_),
    .B2(_07025_),
    .Y(_02422_));
 INVx3_ASAP7_75t_R _21971_ (.A(_06366_),
    .Y(_07026_));
 AND4x1_ASAP7_75t_R _21972_ (.A(_07021_),
    .B(_06938_),
    .C(_07017_),
    .D(_07022_),
    .Y(_07027_));
 NOR2x1_ASAP7_75t_R _21973_ (.A(_06360_),
    .B(_07027_),
    .Y(_07028_));
 OA211x2_ASAP7_75t_R _21974_ (.A1(_06947_),
    .A2(_07027_),
    .B(_06949_),
    .C(_06360_),
    .Y(_07029_));
 OAI22x1_ASAP7_75t_R _21975_ (.A1(_07026_),
    .A2(_06924_),
    .B1(_07028_),
    .B2(_07029_),
    .Y(_02423_));
 OR2x2_ASAP7_75t_R _21976_ (.A(_05937_),
    .B(_05938_),
    .Y(_07030_));
 OR3x2_ASAP7_75t_R _21977_ (.A(_02232_),
    .B(_06963_),
    .C(_07011_),
    .Y(_07031_));
 OR4x1_ASAP7_75t_R _21978_ (.A(_02109_),
    .B(_02110_),
    .C(_02111_),
    .D(_02112_),
    .Y(_07032_));
 OA33x2_ASAP7_75t_R _21979_ (.A1(_05966_),
    .A2(_05963_),
    .A3(_07030_),
    .B1(_06914_),
    .B2(_07031_),
    .B3(_07032_),
    .Y(_07033_));
 INVx1_ASAP7_75t_R _21980_ (.A(_07032_),
    .Y(_07034_));
 AND4x1_ASAP7_75t_R _21981_ (.A(_02108_),
    .B(_06938_),
    .C(_07012_),
    .D(_07034_),
    .Y(_07035_));
 AO21x1_ASAP7_75t_R _21982_ (.A1(_06376_),
    .A2(_07033_),
    .B(_07035_),
    .Y(_07036_));
 AO221x1_ASAP7_75t_R _21983_ (.A1(_06391_),
    .A2(_06986_),
    .B1(_06988_),
    .B2(_06376_),
    .C(_07036_),
    .Y(_02424_));
 INVx2_ASAP7_75t_R _21984_ (.A(_06411_),
    .Y(_07037_));
 AND4x1_ASAP7_75t_R _21985_ (.A(_06376_),
    .B(_06938_),
    .C(_07017_),
    .D(_07034_),
    .Y(_07038_));
 NOR2x1_ASAP7_75t_R _21986_ (.A(_06405_),
    .B(_07038_),
    .Y(_07039_));
 OA211x2_ASAP7_75t_R _21987_ (.A1(_06947_),
    .A2(_07038_),
    .B(_06949_),
    .C(_06405_),
    .Y(_07040_));
 OAI22x1_ASAP7_75t_R _21988_ (.A1(_07037_),
    .A2(_06924_),
    .B1(_07039_),
    .B2(_07040_),
    .Y(_02425_));
 OR5x1_ASAP7_75t_R _21989_ (.A(_02108_),
    .B(_02109_),
    .C(_02110_),
    .D(_02111_),
    .E(_02112_),
    .Y(_07041_));
 OR4x1_ASAP7_75t_R _21990_ (.A(_02107_),
    .B(_06914_),
    .C(_07031_),
    .D(_07041_),
    .Y(_07042_));
 AO21x1_ASAP7_75t_R _21991_ (.A1(_06956_),
    .A2(_07042_),
    .B(_06931_),
    .Y(_07043_));
 INVx3_ASAP7_75t_R _21992_ (.A(_06432_),
    .Y(_07044_));
 OAI22x1_ASAP7_75t_R _21993_ (.A1(_07044_),
    .A2(_06924_),
    .B1(_07042_),
    .B2(_06424_),
    .Y(_07045_));
 AO21x1_ASAP7_75t_R _21994_ (.A1(_06424_),
    .A2(_07043_),
    .B(_07045_),
    .Y(_02426_));
 INVx3_ASAP7_75t_R _21995_ (.A(_06454_),
    .Y(_07046_));
 OR3x1_ASAP7_75t_R _21996_ (.A(_02106_),
    .B(_02107_),
    .C(_07041_),
    .Y(_07047_));
 INVx1_ASAP7_75t_R _21997_ (.A(_07047_),
    .Y(_07048_));
 AND3x1_ASAP7_75t_R _21998_ (.A(_06979_),
    .B(_07017_),
    .C(_07048_),
    .Y(_07049_));
 NOR2x1_ASAP7_75t_R _21999_ (.A(_06448_),
    .B(_07049_),
    .Y(_07050_));
 OA211x2_ASAP7_75t_R _22000_ (.A1(_06947_),
    .A2(_07049_),
    .B(_06949_),
    .C(_06448_),
    .Y(_07051_));
 OAI22x1_ASAP7_75t_R _22001_ (.A1(_07046_),
    .A2(_06924_),
    .B1(_07050_),
    .B2(_07051_),
    .Y(_02427_));
 INVx2_ASAP7_75t_R _22002_ (.A(_02232_),
    .Y(_07052_));
 AO21x1_ASAP7_75t_R _22003_ (.A1(_07052_),
    .A2(_06921_),
    .B(_06916_),
    .Y(_07053_));
 NAND2x1_ASAP7_75t_R _22004_ (.A(_06949_),
    .B(_07053_),
    .Y(_07054_));
 AO32x1_ASAP7_75t_R _22005_ (.A1(_02104_),
    .A2(_07052_),
    .A3(_06921_),
    .B1(_06951_),
    .B2(_05850_),
    .Y(_07055_));
 AO21x1_ASAP7_75t_R _22006_ (.A1(_05817_),
    .A2(_07054_),
    .B(_07055_),
    .Y(_02428_));
 AND3x1_ASAP7_75t_R _22007_ (.A(_06448_),
    .B(_07012_),
    .C(_07048_),
    .Y(_07056_));
 AOI211x1_ASAP7_75t_R _22008_ (.A1(_06938_),
    .A2(_07056_),
    .B(_02103_),
    .C(_06906_),
    .Y(_07057_));
 AND3x1_ASAP7_75t_R _22009_ (.A(_02103_),
    .B(_06938_),
    .C(_07056_),
    .Y(_07058_));
 OR2x2_ASAP7_75t_R _22010_ (.A(_07057_),
    .B(_07058_),
    .Y(_07059_));
 AO221x1_ASAP7_75t_R _22011_ (.A1(_06480_),
    .A2(_06986_),
    .B1(_06988_),
    .B2(_06465_),
    .C(_07059_),
    .Y(_02429_));
 OR5x2_ASAP7_75t_R _22012_ (.A(_02103_),
    .B(_02105_),
    .C(_02106_),
    .D(_02107_),
    .E(_07041_),
    .Y(_07060_));
 OR3x1_ASAP7_75t_R _22013_ (.A(_06958_),
    .B(_07011_),
    .C(_07060_),
    .Y(_07061_));
 AO21x1_ASAP7_75t_R _22014_ (.A1(_06956_),
    .A2(_07061_),
    .B(_06918_),
    .Y(_07062_));
 INVx1_ASAP7_75t_R _22015_ (.A(_07061_),
    .Y(_07063_));
 AO32x1_ASAP7_75t_R _22016_ (.A1(_02102_),
    .A2(_06987_),
    .A3(_07063_),
    .B1(_06504_),
    .B2(_06986_),
    .Y(_07064_));
 AO21x1_ASAP7_75t_R _22017_ (.A1(_06489_),
    .A2(_07062_),
    .B(_07064_),
    .Y(_02430_));
 OR3x1_ASAP7_75t_R _22018_ (.A(_06932_),
    .B(_05907_),
    .C(_05937_),
    .Y(_07065_));
 BUFx6f_ASAP7_75t_R _22019_ (.A(_07065_),
    .Y(_07066_));
 AND2x6_ASAP7_75t_R _22020_ (.A(_06914_),
    .B(_07066_),
    .Y(_07067_));
 BUFx6f_ASAP7_75t_R _22021_ (.A(_07067_),
    .Y(_07068_));
 AND3x4_ASAP7_75t_R _22022_ (.A(_06325_),
    .B(_05971_),
    .C(_05768_),
    .Y(_07069_));
 NAND3x2_ASAP7_75t_R _22023_ (.B(_05768_),
    .C(_05901_),
    .Y(_07070_),
    .A(_05897_));
 OR2x6_ASAP7_75t_R _22024_ (.A(_07031_),
    .B(_07060_),
    .Y(_07071_));
 OR3x1_ASAP7_75t_R _22025_ (.A(_02101_),
    .B(_02102_),
    .C(_07071_),
    .Y(_07072_));
 AND2x2_ASAP7_75t_R _22026_ (.A(_07070_),
    .B(_07072_),
    .Y(_07073_));
 AO21x1_ASAP7_75t_R _22027_ (.A1(_05811_),
    .A2(_07069_),
    .B(_07073_),
    .Y(_07074_));
 OA21x2_ASAP7_75t_R _22028_ (.A1(_02102_),
    .A2(_07071_),
    .B(_07070_),
    .Y(_07075_));
 OAI21x1_ASAP7_75t_R _22029_ (.A1(_07075_),
    .A2(_07068_),
    .B(_02101_),
    .Y(_07076_));
 OA21x2_ASAP7_75t_R _22030_ (.A1(_07068_),
    .A2(_07074_),
    .B(_07076_),
    .Y(_02431_));
 OR3x1_ASAP7_75t_R _22031_ (.A(_02101_),
    .B(_02102_),
    .C(_07061_),
    .Y(_07077_));
 AO21x1_ASAP7_75t_R _22032_ (.A1(_06971_),
    .A2(_07077_),
    .B(_07068_),
    .Y(_07078_));
 AO21x2_ASAP7_75t_R _22033_ (.A1(_18560_),
    .A2(_06231_),
    .B(_06234_),
    .Y(_07079_));
 OAI21x1_ASAP7_75t_R _22034_ (.A1(_02100_),
    .A2(_07077_),
    .B(_07070_),
    .Y(_07080_));
 OA21x2_ASAP7_75t_R _22035_ (.A1(_07079_),
    .A2(_07066_),
    .B(_07080_),
    .Y(_07081_));
 NAND2x2_ASAP7_75t_R _22036_ (.A(_06915_),
    .B(_07066_),
    .Y(_07082_));
 AOI22x1_ASAP7_75t_R _22037_ (.A1(_02100_),
    .A2(_07078_),
    .B1(_07081_),
    .B2(_07082_),
    .Y(_02432_));
 AND2x6_ASAP7_75t_R _22038_ (.A(_05768_),
    .B(_06507_),
    .Y(_07083_));
 BUFx6f_ASAP7_75t_R _22039_ (.A(_07083_),
    .Y(_07084_));
 BUFx6f_ASAP7_75t_R _22040_ (.A(_07084_),
    .Y(_07085_));
 OR3x2_ASAP7_75t_R _22041_ (.A(_02100_),
    .B(_02101_),
    .C(_02102_),
    .Y(_07086_));
 OR3x1_ASAP7_75t_R _22042_ (.A(_05818_),
    .B(_07060_),
    .C(_07086_),
    .Y(_07087_));
 INVx1_ASAP7_75t_R _22043_ (.A(_07087_),
    .Y(_07088_));
 OA21x2_ASAP7_75t_R _22044_ (.A1(_07071_),
    .A2(_07086_),
    .B(_07070_),
    .Y(_07089_));
 OA21x2_ASAP7_75t_R _22045_ (.A1(_07067_),
    .A2(_07089_),
    .B(_05818_),
    .Y(_07090_));
 AO221x1_ASAP7_75t_R _22046_ (.A1(_05851_),
    .A2(_07085_),
    .B1(_07088_),
    .B2(_07013_),
    .C(_07090_),
    .Y(_02433_));
 OR5x2_ASAP7_75t_R _22047_ (.A(_02099_),
    .B(_06958_),
    .C(_07011_),
    .D(_07060_),
    .E(_07086_),
    .Y(_07091_));
 OR2x2_ASAP7_75t_R _22048_ (.A(_02098_),
    .B(_07091_),
    .Y(_07092_));
 AO22x1_ASAP7_75t_R _22049_ (.A1(_06556_),
    .A2(_07085_),
    .B1(_07092_),
    .B2(_07070_),
    .Y(_07093_));
 NAND2x1_ASAP7_75t_R _22050_ (.A(_07070_),
    .B(_07091_),
    .Y(_07094_));
 AO21x1_ASAP7_75t_R _22051_ (.A1(_07082_),
    .A2(_07094_),
    .B(_06543_),
    .Y(_07095_));
 OA21x2_ASAP7_75t_R _22052_ (.A1(_07068_),
    .A2(_07093_),
    .B(_07095_),
    .Y(_02434_));
 BUFx6f_ASAP7_75t_R _22053_ (.A(_06934_),
    .Y(_07096_));
 OR4x1_ASAP7_75t_R _22054_ (.A(_02098_),
    .B(_02099_),
    .C(_07071_),
    .D(_07086_),
    .Y(_07097_));
 AOI211x1_ASAP7_75t_R _22055_ (.A1(_06915_),
    .A2(_07066_),
    .B(_07097_),
    .C(_06575_),
    .Y(_07098_));
 AO21x1_ASAP7_75t_R _22056_ (.A1(_06575_),
    .A2(_07097_),
    .B(_07098_),
    .Y(_07099_));
 BUFx6f_ASAP7_75t_R _22057_ (.A(_07067_),
    .Y(_07100_));
 AO22x1_ASAP7_75t_R _22058_ (.A1(_06580_),
    .A2(_07085_),
    .B1(_07100_),
    .B2(_06575_),
    .Y(_07101_));
 AO21x1_ASAP7_75t_R _22059_ (.A1(_07096_),
    .A2(_07099_),
    .B(_07101_),
    .Y(_02435_));
 OR3x2_ASAP7_75t_R _22060_ (.A(_02097_),
    .B(_02098_),
    .C(_07091_),
    .Y(_07102_));
 BUFx6f_ASAP7_75t_R _22061_ (.A(_07067_),
    .Y(_07103_));
 AO21x1_ASAP7_75t_R _22062_ (.A1(_06956_),
    .A2(_07102_),
    .B(_07103_),
    .Y(_07104_));
 INVx1_ASAP7_75t_R _22063_ (.A(_07102_),
    .Y(_07105_));
 BUFx6f_ASAP7_75t_R _22064_ (.A(_07084_),
    .Y(_07106_));
 AO32x1_ASAP7_75t_R _22065_ (.A1(_02096_),
    .A2(_06987_),
    .A3(_07105_),
    .B1(_07106_),
    .B2(_06600_),
    .Y(_07107_));
 AO21x1_ASAP7_75t_R _22066_ (.A1(_06591_),
    .A2(_07104_),
    .B(_07107_),
    .Y(_02436_));
 OR3x1_ASAP7_75t_R _22067_ (.A(_02096_),
    .B(_02097_),
    .C(_07097_),
    .Y(_07108_));
 AO21x1_ASAP7_75t_R _22068_ (.A1(_06956_),
    .A2(_07108_),
    .B(_07103_),
    .Y(_07109_));
 INVx1_ASAP7_75t_R _22069_ (.A(_07108_),
    .Y(_07110_));
 AO32x1_ASAP7_75t_R _22070_ (.A1(_02095_),
    .A2(_06987_),
    .A3(_07110_),
    .B1(_07106_),
    .B2(_06624_),
    .Y(_07111_));
 AO21x1_ASAP7_75t_R _22071_ (.A1(_06614_),
    .A2(_07109_),
    .B(_07111_),
    .Y(_02437_));
 OR2x2_ASAP7_75t_R _22072_ (.A(_02095_),
    .B(_02096_),
    .Y(_07112_));
 NOR2x1_ASAP7_75t_R _22073_ (.A(_07102_),
    .B(_07112_),
    .Y(_07113_));
 INVx1_ASAP7_75t_R _22074_ (.A(_07113_),
    .Y(_07114_));
 OA211x2_ASAP7_75t_R _22075_ (.A1(_06979_),
    .A2(_07084_),
    .B(_07113_),
    .C(_02094_),
    .Y(_07115_));
 AO21x1_ASAP7_75t_R _22076_ (.A1(_06637_),
    .A2(_07114_),
    .B(_07115_),
    .Y(_07116_));
 AO22x1_ASAP7_75t_R _22077_ (.A1(_06650_),
    .A2(_07085_),
    .B1(_07100_),
    .B2(_06637_),
    .Y(_07117_));
 AO21x1_ASAP7_75t_R _22078_ (.A1(_07096_),
    .A2(_07116_),
    .B(_07117_),
    .Y(_02438_));
 OR3x1_ASAP7_75t_R _22079_ (.A(_02104_),
    .B(_06914_),
    .C(_06957_),
    .Y(_07118_));
 NAND2x1_ASAP7_75t_R _22080_ (.A(_02093_),
    .B(_07118_),
    .Y(_07119_));
 AO211x2_ASAP7_75t_R _22081_ (.A1(_06934_),
    .A2(_07118_),
    .B(_06931_),
    .C(_02093_),
    .Y(_07120_));
 AO22x1_ASAP7_75t_R _22082_ (.A1(_06556_),
    .A2(_06951_),
    .B1(_07119_),
    .B2(_07120_),
    .Y(_02439_));
 OR3x2_ASAP7_75t_R _22083_ (.A(_02094_),
    .B(_02095_),
    .C(_07108_),
    .Y(_07121_));
 AO21x1_ASAP7_75t_R _22084_ (.A1(_06956_),
    .A2(_07121_),
    .B(_07103_),
    .Y(_07122_));
 INVx1_ASAP7_75t_R _22085_ (.A(_07121_),
    .Y(_07123_));
 AO32x1_ASAP7_75t_R _22086_ (.A1(_02092_),
    .A2(_06987_),
    .A3(_07123_),
    .B1(_07106_),
    .B2(_06675_),
    .Y(_07124_));
 AO21x1_ASAP7_75t_R _22087_ (.A1(_06670_),
    .A2(_07122_),
    .B(_07124_),
    .Y(_02440_));
 AND3x1_ASAP7_75t_R _22088_ (.A(_06670_),
    .B(_06637_),
    .C(_07113_),
    .Y(_07125_));
 NOR2x1_ASAP7_75t_R _22089_ (.A(_02091_),
    .B(_07125_),
    .Y(_07126_));
 OA211x2_ASAP7_75t_R _22090_ (.A1(_06920_),
    .A2(_07083_),
    .B(_07125_),
    .C(_02091_),
    .Y(_07127_));
 OR2x2_ASAP7_75t_R _22091_ (.A(_07126_),
    .B(_07127_),
    .Y(_07128_));
 INVx3_ASAP7_75t_R _22092_ (.A(_06699_),
    .Y(_07129_));
 OAI22x1_ASAP7_75t_R _22093_ (.A1(_07129_),
    .A2(_07066_),
    .B1(_07082_),
    .B2(_02091_),
    .Y(_07130_));
 AO21x1_ASAP7_75t_R _22094_ (.A1(_07096_),
    .A2(_07128_),
    .B(_07130_),
    .Y(_02441_));
 OR3x1_ASAP7_75t_R _22095_ (.A(_02091_),
    .B(_02092_),
    .C(_07121_),
    .Y(_07131_));
 AO21x1_ASAP7_75t_R _22096_ (.A1(_06956_),
    .A2(_07131_),
    .B(_07103_),
    .Y(_07132_));
 INVx1_ASAP7_75t_R _22097_ (.A(_07131_),
    .Y(_07133_));
 AO32x1_ASAP7_75t_R _22098_ (.A1(_02090_),
    .A2(_06987_),
    .A3(_07133_),
    .B1(_07106_),
    .B2(_05981_),
    .Y(_07134_));
 AO21x1_ASAP7_75t_R _22099_ (.A1(_05968_),
    .A2(_07132_),
    .B(_07134_),
    .Y(_02442_));
 OR5x1_ASAP7_75t_R _22100_ (.A(_02090_),
    .B(_02091_),
    .C(_02092_),
    .D(_02094_),
    .E(_07114_),
    .Y(_07135_));
 AO21x1_ASAP7_75t_R _22101_ (.A1(_06971_),
    .A2(_07135_),
    .B(_07103_),
    .Y(_07136_));
 OR3x1_ASAP7_75t_R _22102_ (.A(_02089_),
    .B(_02090_),
    .C(_02091_),
    .Y(_07137_));
 OR5x2_ASAP7_75t_R _22103_ (.A(_02092_),
    .B(_02094_),
    .C(_07102_),
    .D(_07112_),
    .E(_07137_),
    .Y(_07138_));
 NAND2x1_ASAP7_75t_R _22104_ (.A(_07070_),
    .B(_07138_),
    .Y(_07139_));
 OA21x2_ASAP7_75t_R _22105_ (.A1(_06937_),
    .A2(_07066_),
    .B(_07139_),
    .Y(_07140_));
 AOI22x1_ASAP7_75t_R _22106_ (.A1(_02089_),
    .A2(_07136_),
    .B1(_07140_),
    .B2(_07082_),
    .Y(_02443_));
 OR3x1_ASAP7_75t_R _22107_ (.A(_02092_),
    .B(_07121_),
    .C(_07137_),
    .Y(_07141_));
 AO21x1_ASAP7_75t_R _22108_ (.A1(_06956_),
    .A2(_07141_),
    .B(_07103_),
    .Y(_07142_));
 INVx1_ASAP7_75t_R _22109_ (.A(_07141_),
    .Y(_07143_));
 AO32x1_ASAP7_75t_R _22110_ (.A1(_02088_),
    .A2(_06987_),
    .A3(_07143_),
    .B1(_07106_),
    .B2(_06052_),
    .Y(_07144_));
 AO21x1_ASAP7_75t_R _22111_ (.A1(_06036_),
    .A2(_07142_),
    .B(_07144_),
    .Y(_02444_));
 NOR2x1_ASAP7_75t_R _22112_ (.A(_02088_),
    .B(_07138_),
    .Y(_07145_));
 NOR2x1_ASAP7_75t_R _22113_ (.A(_02087_),
    .B(_07145_),
    .Y(_07146_));
 OA211x2_ASAP7_75t_R _22114_ (.A1(_06920_),
    .A2(_07083_),
    .B(_07145_),
    .C(_02087_),
    .Y(_07147_));
 OR2x2_ASAP7_75t_R _22115_ (.A(_07146_),
    .B(_07147_),
    .Y(_07148_));
 AO22x1_ASAP7_75t_R _22116_ (.A1(_06082_),
    .A2(_07085_),
    .B1(_07100_),
    .B2(_06069_),
    .Y(_07149_));
 AO21x1_ASAP7_75t_R _22117_ (.A1(_07096_),
    .A2(_07148_),
    .B(_07149_),
    .Y(_02445_));
 AND3x1_ASAP7_75t_R _22118_ (.A(_06069_),
    .B(_06036_),
    .C(_07143_),
    .Y(_07150_));
 NOR2x1_ASAP7_75t_R _22119_ (.A(_02086_),
    .B(_07150_),
    .Y(_07151_));
 OA211x2_ASAP7_75t_R _22120_ (.A1(_06920_),
    .A2(_07083_),
    .B(_07150_),
    .C(_02086_),
    .Y(_07152_));
 OR2x2_ASAP7_75t_R _22121_ (.A(_07151_),
    .B(_07152_),
    .Y(_07153_));
 NOR2x1_ASAP7_75t_R _22122_ (.A(_02086_),
    .B(_07082_),
    .Y(_07154_));
 AO221x1_ASAP7_75t_R _22123_ (.A1(_06108_),
    .A2(_07085_),
    .B1(_07153_),
    .B2(_06971_),
    .C(_07154_),
    .Y(_02446_));
 OR4x1_ASAP7_75t_R _22124_ (.A(_02086_),
    .B(_02087_),
    .C(_02088_),
    .D(_07138_),
    .Y(_07155_));
 AO31x2_ASAP7_75t_R _22125_ (.A1(_06857_),
    .A2(_06882_),
    .A3(_06888_),
    .B(_14592_),
    .Y(_07156_));
 AND3x1_ASAP7_75t_R _22126_ (.A(_02228_),
    .B(_14120_),
    .C(_05119_),
    .Y(_07157_));
 INVx1_ASAP7_75t_R _22127_ (.A(_07157_),
    .Y(_07158_));
 NOR2x1_ASAP7_75t_R _22128_ (.A(_05070_),
    .B(_05763_),
    .Y(_07159_));
 OR4x1_ASAP7_75t_R _22129_ (.A(_06903_),
    .B(_05936_),
    .C(_06932_),
    .D(_07159_),
    .Y(_07160_));
 NOR2x1_ASAP7_75t_R _22130_ (.A(_06909_),
    .B(_06910_),
    .Y(_07161_));
 AND5x1_ASAP7_75t_R _22131_ (.A(_05149_),
    .B(_07158_),
    .C(_05192_),
    .D(_07160_),
    .E(_07161_),
    .Y(_07162_));
 OA211x2_ASAP7_75t_R _22132_ (.A1(_06883_),
    .A2(_07156_),
    .B(_07162_),
    .C(_06898_),
    .Y(_07163_));
 INVx1_ASAP7_75t_R _22133_ (.A(_07155_),
    .Y(_07164_));
 OA211x2_ASAP7_75t_R _22134_ (.A1(_07163_),
    .A2(_07069_),
    .B(_07164_),
    .C(_02085_),
    .Y(_07165_));
 AO21x1_ASAP7_75t_R _22135_ (.A1(_06118_),
    .A2(_07155_),
    .B(_07165_),
    .Y(_07166_));
 AO22x1_ASAP7_75t_R _22136_ (.A1(_06131_),
    .A2(_07085_),
    .B1(_07100_),
    .B2(_06118_),
    .Y(_07167_));
 AO21x1_ASAP7_75t_R _22137_ (.A1(_07096_),
    .A2(_07166_),
    .B(_07167_),
    .Y(_02447_));
 OR5x2_ASAP7_75t_R _22138_ (.A(_02085_),
    .B(_02086_),
    .C(_02087_),
    .D(_02088_),
    .E(_07141_),
    .Y(_07168_));
 INVx1_ASAP7_75t_R _22139_ (.A(_07168_),
    .Y(_07169_));
 OA211x2_ASAP7_75t_R _22140_ (.A1(_06979_),
    .A2(_07084_),
    .B(_07169_),
    .C(_02084_),
    .Y(_07170_));
 AO21x1_ASAP7_75t_R _22141_ (.A1(_06147_),
    .A2(_07168_),
    .B(_07170_),
    .Y(_07171_));
 AO22x1_ASAP7_75t_R _22142_ (.A1(_06153_),
    .A2(_07085_),
    .B1(_07100_),
    .B2(_06147_),
    .Y(_07172_));
 AO21x1_ASAP7_75t_R _22143_ (.A1(_07096_),
    .A2(_07171_),
    .B(_07172_),
    .Y(_02448_));
 OR3x1_ASAP7_75t_R _22144_ (.A(_02084_),
    .B(_02085_),
    .C(_07155_),
    .Y(_07173_));
 AOI211x1_ASAP7_75t_R _22145_ (.A1(_06915_),
    .A2(_07066_),
    .B(_07173_),
    .C(_06165_),
    .Y(_07174_));
 AO21x1_ASAP7_75t_R _22146_ (.A1(_06165_),
    .A2(_07173_),
    .B(_07174_),
    .Y(_07175_));
 AO22x1_ASAP7_75t_R _22147_ (.A1(_06179_),
    .A2(_07085_),
    .B1(_07100_),
    .B2(_06165_),
    .Y(_07176_));
 AO21x1_ASAP7_75t_R _22148_ (.A1(_07096_),
    .A2(_07175_),
    .B(_07176_),
    .Y(_02449_));
 INVx2_ASAP7_75t_R _22149_ (.A(_06580_),
    .Y(_07177_));
 AND3x1_ASAP7_75t_R _22150_ (.A(_07052_),
    .B(_06979_),
    .C(_06940_),
    .Y(_07178_));
 NOR2x1_ASAP7_75t_R _22151_ (.A(_06572_),
    .B(_07178_),
    .Y(_07179_));
 OA211x2_ASAP7_75t_R _22152_ (.A1(_06947_),
    .A2(_07178_),
    .B(_06949_),
    .C(_06572_),
    .Y(_07180_));
 OAI22x1_ASAP7_75t_R _22153_ (.A1(_07177_),
    .A2(_06924_),
    .B1(_07179_),
    .B2(_07180_),
    .Y(_02450_));
 OR3x1_ASAP7_75t_R _22154_ (.A(_02083_),
    .B(_02084_),
    .C(_07168_),
    .Y(_07181_));
 AO21x1_ASAP7_75t_R _22155_ (.A1(_06956_),
    .A2(_07181_),
    .B(_07103_),
    .Y(_07182_));
 INVx1_ASAP7_75t_R _22156_ (.A(_07181_),
    .Y(_07183_));
 AO32x1_ASAP7_75t_R _22157_ (.A1(_02081_),
    .A2(_06921_),
    .A3(_07183_),
    .B1(_07106_),
    .B2(_06197_),
    .Y(_07184_));
 AO21x1_ASAP7_75t_R _22158_ (.A1(_06190_),
    .A2(_07182_),
    .B(_07184_),
    .Y(_02451_));
 OR3x1_ASAP7_75t_R _22159_ (.A(_02081_),
    .B(_02083_),
    .C(_07173_),
    .Y(_07185_));
 AOI211x1_ASAP7_75t_R _22160_ (.A1(_06915_),
    .A2(_07066_),
    .B(_07185_),
    .C(_06213_),
    .Y(_07186_));
 AO21x1_ASAP7_75t_R _22161_ (.A1(_06213_),
    .A2(_07185_),
    .B(_07186_),
    .Y(_07187_));
 AO22x1_ASAP7_75t_R _22162_ (.A1(_06219_),
    .A2(_07106_),
    .B1(_07100_),
    .B2(_06213_),
    .Y(_07188_));
 AO21x1_ASAP7_75t_R _22163_ (.A1(_07096_),
    .A2(_07187_),
    .B(_07188_),
    .Y(_02452_));
 AND3x1_ASAP7_75t_R _22164_ (.A(_06213_),
    .B(_06190_),
    .C(_07183_),
    .Y(_07189_));
 INVx1_ASAP7_75t_R _22165_ (.A(_07189_),
    .Y(_07190_));
 OA211x2_ASAP7_75t_R _22166_ (.A1(_06979_),
    .A2(_07084_),
    .B(_07189_),
    .C(_02079_),
    .Y(_07191_));
 AO21x1_ASAP7_75t_R _22167_ (.A1(_06241_),
    .A2(_07190_),
    .B(_07191_),
    .Y(_07192_));
 AO22x1_ASAP7_75t_R _22168_ (.A1(_06254_),
    .A2(_07106_),
    .B1(_07100_),
    .B2(_06241_),
    .Y(_07193_));
 AO21x1_ASAP7_75t_R _22169_ (.A1(_07096_),
    .A2(_07192_),
    .B(_07193_),
    .Y(_02453_));
 OR3x1_ASAP7_75t_R _22170_ (.A(_02079_),
    .B(_02080_),
    .C(_07185_),
    .Y(_07194_));
 AO21x1_ASAP7_75t_R _22171_ (.A1(_06956_),
    .A2(_07194_),
    .B(_07103_),
    .Y(_07195_));
 OR2x6_ASAP7_75t_R _22172_ (.A(_02078_),
    .B(_07194_),
    .Y(_07196_));
 AO21x1_ASAP7_75t_R _22173_ (.A1(_06277_),
    .A2(_06507_),
    .B(_06934_),
    .Y(_07197_));
 OAI21x1_ASAP7_75t_R _22174_ (.A1(_06947_),
    .A2(_07196_),
    .B(_07197_),
    .Y(_07198_));
 AOI22x1_ASAP7_75t_R _22175_ (.A1(_02078_),
    .A2(_07195_),
    .B1(_07198_),
    .B2(_07082_),
    .Y(_02454_));
 OR5x2_ASAP7_75t_R _22176_ (.A(_02078_),
    .B(_02079_),
    .C(_02080_),
    .D(_02081_),
    .E(_07181_),
    .Y(_07199_));
 AO21x1_ASAP7_75t_R _22177_ (.A1(_06934_),
    .A2(_07199_),
    .B(_07103_),
    .Y(_07200_));
 INVx1_ASAP7_75t_R _22178_ (.A(_07199_),
    .Y(_07201_));
 AO32x1_ASAP7_75t_R _22179_ (.A1(_02077_),
    .A2(_06921_),
    .A3(_07201_),
    .B1(_07084_),
    .B2(_06298_),
    .Y(_07202_));
 AO21x1_ASAP7_75t_R _22180_ (.A1(_06291_),
    .A2(_07200_),
    .B(_07202_),
    .Y(_02455_));
 OR3x1_ASAP7_75t_R _22181_ (.A(_02076_),
    .B(_02077_),
    .C(_07196_),
    .Y(_07203_));
 AND2x2_ASAP7_75t_R _22182_ (.A(_07070_),
    .B(_07203_),
    .Y(_07204_));
 AO21x1_ASAP7_75t_R _22183_ (.A1(_06323_),
    .A2(_07069_),
    .B(_07204_),
    .Y(_07205_));
 OA21x2_ASAP7_75t_R _22184_ (.A1(_02077_),
    .A2(_07196_),
    .B(_07070_),
    .Y(_07206_));
 OAI21x1_ASAP7_75t_R _22185_ (.A1(_07068_),
    .A2(_07206_),
    .B(_02076_),
    .Y(_07207_));
 OA21x2_ASAP7_75t_R _22186_ (.A1(_07068_),
    .A2(_07205_),
    .B(_07207_),
    .Y(_02456_));
 OR3x1_ASAP7_75t_R _22187_ (.A(_02076_),
    .B(_02077_),
    .C(_07199_),
    .Y(_07208_));
 AO21x1_ASAP7_75t_R _22188_ (.A1(_06934_),
    .A2(_07208_),
    .B(_07103_),
    .Y(_07209_));
 INVx1_ASAP7_75t_R _22189_ (.A(_07208_),
    .Y(_07210_));
 AO32x1_ASAP7_75t_R _22190_ (.A1(_02075_),
    .A2(_06921_),
    .A3(_07210_),
    .B1(_07084_),
    .B2(_06343_),
    .Y(_07211_));
 AO21x1_ASAP7_75t_R _22191_ (.A1(_06337_),
    .A2(_07209_),
    .B(_07211_),
    .Y(_02457_));
 OR3x1_ASAP7_75t_R _22192_ (.A(_02074_),
    .B(_02075_),
    .C(_07203_),
    .Y(_07212_));
 AND2x2_ASAP7_75t_R _22193_ (.A(_07160_),
    .B(_07212_),
    .Y(_07213_));
 AO21x1_ASAP7_75t_R _22194_ (.A1(_06366_),
    .A2(_07069_),
    .B(_07213_),
    .Y(_07214_));
 OA21x2_ASAP7_75t_R _22195_ (.A1(_02075_),
    .A2(_07203_),
    .B(_07070_),
    .Y(_07215_));
 OAI21x1_ASAP7_75t_R _22196_ (.A1(_07068_),
    .A2(_07215_),
    .B(_02074_),
    .Y(_07216_));
 OA21x2_ASAP7_75t_R _22197_ (.A1(_07068_),
    .A2(_07214_),
    .B(_07216_),
    .Y(_02458_));
 OR3x2_ASAP7_75t_R _22198_ (.A(_02074_),
    .B(_02075_),
    .C(_07208_),
    .Y(_07217_));
 INVx1_ASAP7_75t_R _22199_ (.A(_07217_),
    .Y(_07218_));
 OA211x2_ASAP7_75t_R _22200_ (.A1(_06979_),
    .A2(_07084_),
    .B(_07218_),
    .C(_02073_),
    .Y(_07219_));
 AO21x1_ASAP7_75t_R _22201_ (.A1(_06378_),
    .A2(_07217_),
    .B(_07219_),
    .Y(_07220_));
 AO22x1_ASAP7_75t_R _22202_ (.A1(_06391_),
    .A2(_07106_),
    .B1(_07067_),
    .B2(_06378_),
    .Y(_07221_));
 AO21x1_ASAP7_75t_R _22203_ (.A1(_07096_),
    .A2(_07220_),
    .B(_07221_),
    .Y(_02459_));
 OR3x2_ASAP7_75t_R _22204_ (.A(_02072_),
    .B(_02073_),
    .C(_07212_),
    .Y(_07222_));
 AND2x2_ASAP7_75t_R _22205_ (.A(_07160_),
    .B(_07222_),
    .Y(_07223_));
 AO21x1_ASAP7_75t_R _22206_ (.A1(_06411_),
    .A2(_07069_),
    .B(_07223_),
    .Y(_07224_));
 OA21x2_ASAP7_75t_R _22207_ (.A1(_02073_),
    .A2(_07212_),
    .B(_07160_),
    .Y(_07225_));
 OAI21x1_ASAP7_75t_R _22208_ (.A1(_07068_),
    .A2(_07225_),
    .B(_02072_),
    .Y(_07226_));
 OA21x2_ASAP7_75t_R _22209_ (.A1(_07068_),
    .A2(_07224_),
    .B(_07226_),
    .Y(_02460_));
 INVx2_ASAP7_75t_R _22210_ (.A(_06600_),
    .Y(_07227_));
 AND4x1_ASAP7_75t_R _22211_ (.A(_06572_),
    .B(_06938_),
    .C(_06940_),
    .D(_06944_),
    .Y(_07228_));
 NOR2x1_ASAP7_75t_R _22212_ (.A(_06939_),
    .B(_07228_),
    .Y(_07229_));
 OA211x2_ASAP7_75t_R _22213_ (.A1(_06916_),
    .A2(_07228_),
    .B(_06948_),
    .C(_06939_),
    .Y(_07230_));
 OAI22x1_ASAP7_75t_R _22214_ (.A1(_07227_),
    .A2(_06924_),
    .B1(_07229_),
    .B2(_07230_),
    .Y(_02461_));
 NOR3x1_ASAP7_75t_R _22215_ (.A(_02072_),
    .B(_02073_),
    .C(_07217_),
    .Y(_07231_));
 NOR2x1_ASAP7_75t_R _22216_ (.A(_02070_),
    .B(_07231_),
    .Y(_07232_));
 OA211x2_ASAP7_75t_R _22217_ (.A1(_06920_),
    .A2(_07083_),
    .B(_07231_),
    .C(_02070_),
    .Y(_07233_));
 OR2x2_ASAP7_75t_R _22218_ (.A(_07232_),
    .B(_07233_),
    .Y(_07234_));
 AO22x1_ASAP7_75t_R _22219_ (.A1(_06432_),
    .A2(_07106_),
    .B1(_07067_),
    .B2(_06426_),
    .Y(_07235_));
 AO21x1_ASAP7_75t_R _22220_ (.A1(_06971_),
    .A2(_07234_),
    .B(_07235_),
    .Y(_02462_));
 NOR2x1_ASAP7_75t_R _22221_ (.A(_02070_),
    .B(_07222_),
    .Y(_07236_));
 NOR2x1_ASAP7_75t_R _22222_ (.A(_02069_),
    .B(_07236_),
    .Y(_07237_));
 OA211x2_ASAP7_75t_R _22223_ (.A1(_06920_),
    .A2(_07083_),
    .B(_07236_),
    .C(_02069_),
    .Y(_07238_));
 OR2x2_ASAP7_75t_R _22224_ (.A(_07237_),
    .B(_07238_),
    .Y(_07239_));
 NOR2x1_ASAP7_75t_R _22225_ (.A(_02069_),
    .B(_07082_),
    .Y(_07240_));
 AO221x1_ASAP7_75t_R _22226_ (.A1(_06454_),
    .A2(_07085_),
    .B1(_07239_),
    .B2(_06971_),
    .C(_07240_),
    .Y(_02463_));
 OR5x1_ASAP7_75t_R _22227_ (.A(_02069_),
    .B(_02070_),
    .C(_02072_),
    .D(_02073_),
    .E(_07217_),
    .Y(_07241_));
 AO21x1_ASAP7_75t_R _22228_ (.A1(_06934_),
    .A2(_07241_),
    .B(_07100_),
    .Y(_07242_));
 INVx1_ASAP7_75t_R _22229_ (.A(_07241_),
    .Y(_07243_));
 AO32x1_ASAP7_75t_R _22230_ (.A1(_02068_),
    .A2(_06921_),
    .A3(_07243_),
    .B1(_07084_),
    .B2(_06480_),
    .Y(_07244_));
 AO21x1_ASAP7_75t_R _22231_ (.A1(_06467_),
    .A2(_07242_),
    .B(_07244_),
    .Y(_02464_));
 OR4x1_ASAP7_75t_R _22232_ (.A(_02068_),
    .B(_02069_),
    .C(_02070_),
    .D(_07222_),
    .Y(_07245_));
 AO21x1_ASAP7_75t_R _22233_ (.A1(_06934_),
    .A2(_07245_),
    .B(_07100_),
    .Y(_07246_));
 INVx1_ASAP7_75t_R _22234_ (.A(_07245_),
    .Y(_07247_));
 AO32x1_ASAP7_75t_R _22235_ (.A1(_02067_),
    .A2(_06921_),
    .A3(_07247_),
    .B1(_07084_),
    .B2(_06504_),
    .Y(_07248_));
 AO21x1_ASAP7_75t_R _22236_ (.A1(_06491_),
    .A2(_07246_),
    .B(_07248_),
    .Y(_02465_));
 INVx2_ASAP7_75t_R _22237_ (.A(_06624_),
    .Y(_07249_));
 AND2x2_ASAP7_75t_R _22238_ (.A(_02066_),
    .B(_06928_),
    .Y(_07250_));
 AND3x1_ASAP7_75t_R _22239_ (.A(_07052_),
    .B(_06979_),
    .C(_06941_),
    .Y(_07251_));
 OA211x2_ASAP7_75t_R _22240_ (.A1(_06916_),
    .A2(_07251_),
    .B(_06948_),
    .C(_06611_),
    .Y(_07252_));
 OAI22x1_ASAP7_75t_R _22241_ (.A1(_07249_),
    .A2(_06924_),
    .B1(_07250_),
    .B2(_07252_),
    .Y(_02466_));
 AND3x1_ASAP7_75t_R _22242_ (.A(_06611_),
    .B(_06941_),
    .C(_06944_),
    .Y(_07253_));
 AO21x1_ASAP7_75t_R _22243_ (.A1(_06987_),
    .A2(_07253_),
    .B(_06634_),
    .Y(_07254_));
 AOI21x1_ASAP7_75t_R _22244_ (.A1(_06921_),
    .A2(_07253_),
    .B(_06916_),
    .Y(_07255_));
 OR3x1_ASAP7_75t_R _22245_ (.A(_02065_),
    .B(_06930_),
    .C(_07255_),
    .Y(_07256_));
 AO22x1_ASAP7_75t_R _22246_ (.A1(_06650_),
    .A2(_06951_),
    .B1(_07254_),
    .B2(_07256_),
    .Y(_02467_));
 NOR2x1_ASAP7_75t_R _22247_ (.A(_02065_),
    .B(_02066_),
    .Y(_07257_));
 INVx1_ASAP7_75t_R _22248_ (.A(_02064_),
    .Y(_07258_));
 AO21x1_ASAP7_75t_R _22249_ (.A1(_07257_),
    .A2(_07251_),
    .B(_07258_),
    .Y(_07259_));
 OA33x2_ASAP7_75t_R _22250_ (.A1(_05966_),
    .A2(_05963_),
    .A3(_07030_),
    .B1(_06928_),
    .B2(_02065_),
    .B3(_02066_),
    .Y(_07260_));
 OR3x1_ASAP7_75t_R _22251_ (.A(_02064_),
    .B(_06930_),
    .C(_07260_),
    .Y(_07261_));
 AO22x1_ASAP7_75t_R _22252_ (.A1(_06675_),
    .A2(_06951_),
    .B1(_07259_),
    .B2(_07261_),
    .Y(_02468_));
 INVx1_ASAP7_75t_R _22253_ (.A(_02063_),
    .Y(_07262_));
 AND5x1_ASAP7_75t_R _22254_ (.A(_07258_),
    .B(_06920_),
    .C(_07257_),
    .D(_06941_),
    .E(_06944_),
    .Y(_07263_));
 NOR2x1_ASAP7_75t_R _22255_ (.A(_07262_),
    .B(_07263_),
    .Y(_07264_));
 OA211x2_ASAP7_75t_R _22256_ (.A1(_06916_),
    .A2(_07263_),
    .B(_06948_),
    .C(_07262_),
    .Y(_07265_));
 OAI22x1_ASAP7_75t_R _22257_ (.A1(_07129_),
    .A2(_06924_),
    .B1(_07264_),
    .B2(_07265_),
    .Y(_02469_));
 BUFx6f_ASAP7_75t_R _22258_ (.A(_05504_),
    .Y(_07266_));
 OAI22x1_ASAP7_75t_R _22259_ (.A1(_02061_),
    .A2(_05500_),
    .B1(_07266_),
    .B2(_00331_),
    .Y(_07267_));
 AND2x4_ASAP7_75t_R _22260_ (.A(_05449_),
    .B(_05453_),
    .Y(_07268_));
 OR2x6_ASAP7_75t_R _22261_ (.A(_15274_),
    .B(_05412_),
    .Y(_07269_));
 INVx1_ASAP7_75t_R _22262_ (.A(_05509_),
    .Y(_07270_));
 OA21x2_ASAP7_75t_R _22263_ (.A1(_05416_),
    .A2(_07269_),
    .B(_07270_),
    .Y(_07271_));
 NAND2x1_ASAP7_75t_R _22264_ (.A(_05171_),
    .B(_05402_),
    .Y(_07272_));
 AND2x4_ASAP7_75t_R _22265_ (.A(_05548_),
    .B(_01398_),
    .Y(_07273_));
 INVx1_ASAP7_75t_R _22266_ (.A(_00758_),
    .Y(_07274_));
 OR3x1_ASAP7_75t_R _22267_ (.A(_07274_),
    .B(_05154_),
    .C(_05415_),
    .Y(_07275_));
 OA21x2_ASAP7_75t_R _22268_ (.A1(_05173_),
    .A2(_07273_),
    .B(_07275_),
    .Y(_07276_));
 OR2x6_ASAP7_75t_R _22269_ (.A(_07272_),
    .B(_07276_),
    .Y(_07277_));
 BUFx12f_ASAP7_75t_R _22270_ (.A(_07277_),
    .Y(_07278_));
 INVx5_ASAP7_75t_R _22271_ (.A(_07278_),
    .Y(_07279_));
 OR3x2_ASAP7_75t_R _22272_ (.A(_07268_),
    .B(_07271_),
    .C(_07279_),
    .Y(_07280_));
 OA211x2_ASAP7_75t_R _22273_ (.A1(\cs_registers_i.priv_mode_id_o[0] ),
    .A2(_07280_),
    .B(_07266_),
    .C(_05500_),
    .Y(_07281_));
 OR2x2_ASAP7_75t_R _22274_ (.A(_07267_),
    .B(_07281_),
    .Y(_02470_));
 OAI22x1_ASAP7_75t_R _22275_ (.A1(_02056_),
    .A2(_05500_),
    .B1(_07266_),
    .B2(_00332_),
    .Y(_07282_));
 INVx2_ASAP7_75t_R _22276_ (.A(_18080_),
    .Y(_07283_));
 OA211x2_ASAP7_75t_R _22277_ (.A1(_07283_),
    .A2(_07280_),
    .B(_07266_),
    .C(_05500_),
    .Y(_07284_));
 OR2x2_ASAP7_75t_R _22278_ (.A(_07282_),
    .B(_07284_),
    .Y(_02471_));
 OR3x2_ASAP7_75t_R _22279_ (.A(_05919_),
    .B(_05796_),
    .C(_05937_),
    .Y(_07285_));
 NOR3x1_ASAP7_75t_R _22280_ (.A(_05810_),
    .B(_06235_),
    .C(_07285_),
    .Y(_07286_));
 AOI211x1_ASAP7_75t_R _22281_ (.A1(_02061_),
    .A2(_07285_),
    .B(_07286_),
    .C(_07279_),
    .Y(_07287_));
 AO21x1_ASAP7_75t_R _22282_ (.A1(\cs_registers_i.priv_mode_id_o[0] ),
    .A2(_07279_),
    .B(_07287_),
    .Y(_02472_));
 OR3x1_ASAP7_75t_R _22283_ (.A(_06903_),
    .B(_05936_),
    .C(_06020_),
    .Y(_07288_));
 BUFx6f_ASAP7_75t_R _22284_ (.A(_07288_),
    .Y(_07289_));
 NOR2x1_ASAP7_75t_R _22285_ (.A(_06025_),
    .B(_07289_),
    .Y(_07290_));
 AOI21x1_ASAP7_75t_R _22286_ (.A1(_02060_),
    .A2(_07289_),
    .B(_07290_),
    .Y(_02473_));
 NAND2x1_ASAP7_75t_R _22287_ (.A(_02059_),
    .B(_07289_),
    .Y(_07291_));
 OA21x2_ASAP7_75t_R _22288_ (.A1(_06052_),
    .A2(_07289_),
    .B(_07291_),
    .Y(_02474_));
 NOR2x1_ASAP7_75t_R _22289_ (.A(_06082_),
    .B(_07289_),
    .Y(_07292_));
 AOI21x1_ASAP7_75t_R _22290_ (.A1(_02058_),
    .A2(_07289_),
    .B(_07292_),
    .Y(_02475_));
 NOR2x1_ASAP7_75t_R _22291_ (.A(_06131_),
    .B(_07289_),
    .Y(_07293_));
 AOI21x1_ASAP7_75t_R _22292_ (.A1(_02057_),
    .A2(_07289_),
    .B(_07293_),
    .Y(_02476_));
 AOI211x1_ASAP7_75t_R _22293_ (.A1(_02056_),
    .A2(_07285_),
    .B(_07286_),
    .C(_07279_),
    .Y(_07294_));
 AO21x1_ASAP7_75t_R _22294_ (.A1(_07283_),
    .A2(_07279_),
    .B(_07294_),
    .Y(_02477_));
 NAND2x1_ASAP7_75t_R _22295_ (.A(_01398_),
    .B(_07289_),
    .Y(_07295_));
 OA21x2_ASAP7_75t_R _22296_ (.A1(_05851_),
    .A2(_07289_),
    .B(_07295_),
    .Y(_02478_));
 INVx1_ASAP7_75t_R _22297_ (.A(_02055_),
    .Y(_07296_));
 OR3x2_ASAP7_75t_R _22298_ (.A(_05404_),
    .B(_05173_),
    .C(_05705_),
    .Y(_07297_));
 OR2x2_ASAP7_75t_R _22299_ (.A(_01398_),
    .B(_07297_),
    .Y(_07298_));
 OA21x2_ASAP7_75t_R _22300_ (.A1(_07296_),
    .A2(_07279_),
    .B(_07298_),
    .Y(_02479_));
 NAND2x1_ASAP7_75t_R _22301_ (.A(net81),
    .B(_01398_),
    .Y(_07299_));
 OAI22x1_ASAP7_75t_R _22302_ (.A1(_02054_),
    .A2(_07279_),
    .B1(_07297_),
    .B2(_07299_),
    .Y(_02480_));
 OAI21x1_ASAP7_75t_R _22303_ (.A1(_02053_),
    .A2(_07279_),
    .B(_07298_),
    .Y(_02481_));
 NOR2x2_ASAP7_75t_R _22304_ (.A(_05749_),
    .B(_06010_),
    .Y(_07300_));
 BUFx6f_ASAP7_75t_R _22305_ (.A(_07300_),
    .Y(_07301_));
 OR2x2_ASAP7_75t_R _22306_ (.A(_07279_),
    .B(_07300_),
    .Y(_07302_));
 BUFx6f_ASAP7_75t_R _22307_ (.A(_07302_),
    .Y(_07303_));
 BUFx12f_ASAP7_75t_R _22308_ (.A(_07303_),
    .Y(_07304_));
 OAI21x1_ASAP7_75t_R _22309_ (.A1(_07273_),
    .A2(_07297_),
    .B(_05478_),
    .Y(_07305_));
 BUFx6f_ASAP7_75t_R _22310_ (.A(_07305_),
    .Y(_07306_));
 OA21x2_ASAP7_75t_R _22311_ (.A1(_07273_),
    .A2(_07297_),
    .B(_05478_),
    .Y(_07307_));
 BUFx6f_ASAP7_75t_R _22312_ (.A(_07307_),
    .Y(_07308_));
 AND2x2_ASAP7_75t_R _22313_ (.A(_00019_),
    .B(_07308_),
    .Y(_07309_));
 AO21x2_ASAP7_75t_R _22314_ (.A1(_00022_),
    .A2(_07306_),
    .B(_07309_),
    .Y(_07310_));
 BUFx12f_ASAP7_75t_R _22315_ (.A(_07278_),
    .Y(_07311_));
 OAI22x1_ASAP7_75t_R _22316_ (.A1(_02052_),
    .A2(_07304_),
    .B1(_07310_),
    .B2(_07311_),
    .Y(_07312_));
 AO21x1_ASAP7_75t_R _22317_ (.A1(_05981_),
    .A2(_07301_),
    .B(_07312_),
    .Y(_02482_));
 AND2x2_ASAP7_75t_R _22318_ (.A(_14379_),
    .B(_07308_),
    .Y(_07313_));
 AO21x2_ASAP7_75t_R _22319_ (.A1(_01690_),
    .A2(_07306_),
    .B(_07313_),
    .Y(_07314_));
 OAI22x1_ASAP7_75t_R _22320_ (.A1(_02051_),
    .A2(_07304_),
    .B1(_07314_),
    .B2(_07311_),
    .Y(_07315_));
 AO21x1_ASAP7_75t_R _22321_ (.A1(_06025_),
    .A2(_07301_),
    .B(_07315_),
    .Y(_02483_));
 BUFx6f_ASAP7_75t_R _22322_ (.A(_01689_),
    .Y(_07316_));
 AND2x2_ASAP7_75t_R _22323_ (.A(_01503_),
    .B(_07308_),
    .Y(_07317_));
 AO21x2_ASAP7_75t_R _22324_ (.A1(_07316_),
    .A2(_07306_),
    .B(_07317_),
    .Y(_07318_));
 OAI22x1_ASAP7_75t_R _22325_ (.A1(_02050_),
    .A2(_07304_),
    .B1(_07318_),
    .B2(_07311_),
    .Y(_07319_));
 AO21x1_ASAP7_75t_R _22326_ (.A1(_06052_),
    .A2(_07301_),
    .B(_07319_),
    .Y(_02484_));
 BUFx6f_ASAP7_75t_R _22327_ (.A(_07305_),
    .Y(_07320_));
 BUFx6f_ASAP7_75t_R _22328_ (.A(_07307_),
    .Y(_07321_));
 AND2x2_ASAP7_75t_R _22329_ (.A(_01502_),
    .B(_07321_),
    .Y(_07322_));
 AO21x2_ASAP7_75t_R _22330_ (.A1(_01688_),
    .A2(_07320_),
    .B(_07322_),
    .Y(_07323_));
 OAI22x1_ASAP7_75t_R _22331_ (.A1(_02049_),
    .A2(_07304_),
    .B1(_07323_),
    .B2(_07311_),
    .Y(_07324_));
 AO21x1_ASAP7_75t_R _22332_ (.A1(_06082_),
    .A2(_07301_),
    .B(_07324_),
    .Y(_02485_));
 AND2x2_ASAP7_75t_R _22333_ (.A(_01501_),
    .B(_07321_),
    .Y(_07325_));
 AO21x2_ASAP7_75t_R _22334_ (.A1(_01687_),
    .A2(_07320_),
    .B(_07325_),
    .Y(_07326_));
 OAI22x1_ASAP7_75t_R _22335_ (.A1(_02048_),
    .A2(_07304_),
    .B1(_07326_),
    .B2(_07311_),
    .Y(_07327_));
 AO21x1_ASAP7_75t_R _22336_ (.A1(_06108_),
    .A2(_07301_),
    .B(_07327_),
    .Y(_02486_));
 BUFx3_ASAP7_75t_R _22337_ (.A(_01686_),
    .Y(_07328_));
 AND2x2_ASAP7_75t_R _22338_ (.A(_15708_),
    .B(_07321_),
    .Y(_07329_));
 AO21x2_ASAP7_75t_R _22339_ (.A1(_07328_),
    .A2(_07320_),
    .B(_07329_),
    .Y(_07330_));
 OAI22x1_ASAP7_75t_R _22340_ (.A1(_02047_),
    .A2(_07304_),
    .B1(_07330_),
    .B2(_07311_),
    .Y(_07331_));
 AO21x1_ASAP7_75t_R _22341_ (.A1(_06131_),
    .A2(_07301_),
    .B(_07331_),
    .Y(_02487_));
 AND2x2_ASAP7_75t_R _22342_ (.A(_15832_),
    .B(_07321_),
    .Y(_07332_));
 AO21x2_ASAP7_75t_R _22343_ (.A1(_01685_),
    .A2(_07320_),
    .B(_07332_),
    .Y(_07333_));
 OAI22x1_ASAP7_75t_R _22344_ (.A1(_02046_),
    .A2(_07304_),
    .B1(_07333_),
    .B2(_07311_),
    .Y(_07334_));
 AO21x1_ASAP7_75t_R _22345_ (.A1(_06153_),
    .A2(_07301_),
    .B(_07334_),
    .Y(_02488_));
 BUFx6f_ASAP7_75t_R _22346_ (.A(_01684_),
    .Y(_07335_));
 AND2x2_ASAP7_75t_R _22347_ (.A(_01498_),
    .B(_07321_),
    .Y(_07336_));
 AO21x2_ASAP7_75t_R _22348_ (.A1(_07335_),
    .A2(_07320_),
    .B(_07336_),
    .Y(_07337_));
 OAI22x1_ASAP7_75t_R _22349_ (.A1(_02045_),
    .A2(_07304_),
    .B1(_07337_),
    .B2(_07311_),
    .Y(_07338_));
 AO21x1_ASAP7_75t_R _22350_ (.A1(_06179_),
    .A2(_07301_),
    .B(_07338_),
    .Y(_02489_));
 AND2x2_ASAP7_75t_R _22351_ (.A(_16079_),
    .B(_07321_),
    .Y(_07339_));
 AO21x2_ASAP7_75t_R _22352_ (.A1(_00023_),
    .A2(_07320_),
    .B(_07339_),
    .Y(_07340_));
 OAI22x1_ASAP7_75t_R _22353_ (.A1(_02044_),
    .A2(_07304_),
    .B1(_07340_),
    .B2(_07311_),
    .Y(_07341_));
 AO21x1_ASAP7_75t_R _22354_ (.A1(_06197_),
    .A2(_07301_),
    .B(_07341_),
    .Y(_02490_));
 AND2x2_ASAP7_75t_R _22355_ (.A(_16192_),
    .B(_07321_),
    .Y(_07342_));
 AO21x1_ASAP7_75t_R _22356_ (.A1(_01683_),
    .A2(_07320_),
    .B(_07342_),
    .Y(_07343_));
 OAI22x1_ASAP7_75t_R _22357_ (.A1(_02043_),
    .A2(_07304_),
    .B1(_07343_),
    .B2(_07311_),
    .Y(_07344_));
 AO21x1_ASAP7_75t_R _22358_ (.A1(_06219_),
    .A2(_07301_),
    .B(_07344_),
    .Y(_02491_));
 BUFx6f_ASAP7_75t_R _22359_ (.A(_07300_),
    .Y(_07345_));
 BUFx12f_ASAP7_75t_R _22360_ (.A(_07303_),
    .Y(_07346_));
 BUFx6f_ASAP7_75t_R _22361_ (.A(_05544_),
    .Y(_07347_));
 BUFx6f_ASAP7_75t_R _22362_ (.A(_07347_),
    .Y(_07348_));
 AND2x2_ASAP7_75t_R _22363_ (.A(_01496_),
    .B(_07308_),
    .Y(_07349_));
 AO21x2_ASAP7_75t_R _22364_ (.A1(_07348_),
    .A2(_07306_),
    .B(_07349_),
    .Y(_07350_));
 BUFx12f_ASAP7_75t_R _22365_ (.A(_07278_),
    .Y(_07351_));
 OAI22x1_ASAP7_75t_R _22366_ (.A1(_00749_),
    .A2(_07346_),
    .B1(_07350_),
    .B2(_07351_),
    .Y(_07352_));
 AO21x1_ASAP7_75t_R _22367_ (.A1(_06235_),
    .A2(_07345_),
    .B(_07352_),
    .Y(_02492_));
 AND2x2_ASAP7_75t_R _22368_ (.A(_01495_),
    .B(_07308_),
    .Y(_07353_));
 AO21x2_ASAP7_75t_R _22369_ (.A1(_01682_),
    .A2(_07306_),
    .B(_07353_),
    .Y(_07354_));
 OAI22x1_ASAP7_75t_R _22370_ (.A1(_02042_),
    .A2(_07346_),
    .B1(_07354_),
    .B2(_07351_),
    .Y(_07355_));
 AO21x1_ASAP7_75t_R _22371_ (.A1(_06255_),
    .A2(_07345_),
    .B(_07355_),
    .Y(_02493_));
 AND2x2_ASAP7_75t_R _22372_ (.A(_01494_),
    .B(_07321_),
    .Y(_07356_));
 AO21x2_ASAP7_75t_R _22373_ (.A1(_01681_),
    .A2(_07320_),
    .B(_07356_),
    .Y(_07357_));
 OAI22x1_ASAP7_75t_R _22374_ (.A1(_02041_),
    .A2(_07346_),
    .B1(_07357_),
    .B2(_07351_),
    .Y(_07358_));
 AO21x1_ASAP7_75t_R _22375_ (.A1(_06277_),
    .A2(_07345_),
    .B(_07358_),
    .Y(_02494_));
 AND2x2_ASAP7_75t_R _22376_ (.A(_01493_),
    .B(_07321_),
    .Y(_07359_));
 AO21x2_ASAP7_75t_R _22377_ (.A1(_01680_),
    .A2(_07320_),
    .B(_07359_),
    .Y(_07360_));
 OAI22x1_ASAP7_75t_R _22378_ (.A1(_02040_),
    .A2(_07346_),
    .B1(_07360_),
    .B2(_07351_),
    .Y(_07361_));
 AO21x1_ASAP7_75t_R _22379_ (.A1(_06298_),
    .A2(_07345_),
    .B(_07361_),
    .Y(_02495_));
 AND2x2_ASAP7_75t_R _22380_ (.A(_16698_),
    .B(_07321_),
    .Y(_07362_));
 AO21x2_ASAP7_75t_R _22381_ (.A1(_01679_),
    .A2(_07320_),
    .B(_07362_),
    .Y(_07363_));
 OAI22x1_ASAP7_75t_R _22382_ (.A1(_02039_),
    .A2(_07346_),
    .B1(_07363_),
    .B2(_07351_),
    .Y(_07364_));
 AO21x1_ASAP7_75t_R _22383_ (.A1(_06323_),
    .A2(_07345_),
    .B(_07364_),
    .Y(_02496_));
 BUFx6f_ASAP7_75t_R _22384_ (.A(_07305_),
    .Y(_07365_));
 BUFx6f_ASAP7_75t_R _22385_ (.A(_07307_),
    .Y(_07366_));
 AND2x2_ASAP7_75t_R _22386_ (.A(_01491_),
    .B(_07366_),
    .Y(_07367_));
 AO21x2_ASAP7_75t_R _22387_ (.A1(_01678_),
    .A2(_07365_),
    .B(_07367_),
    .Y(_07368_));
 OAI22x1_ASAP7_75t_R _22388_ (.A1(_02038_),
    .A2(_07346_),
    .B1(_07368_),
    .B2(_07351_),
    .Y(_07369_));
 AO21x1_ASAP7_75t_R _22389_ (.A1(_06343_),
    .A2(_07345_),
    .B(_07369_),
    .Y(_02497_));
 AND2x2_ASAP7_75t_R _22390_ (.A(_01490_),
    .B(_07366_),
    .Y(_07370_));
 AO21x2_ASAP7_75t_R _22391_ (.A1(_01677_),
    .A2(_07365_),
    .B(_07370_),
    .Y(_07371_));
 OAI22x1_ASAP7_75t_R _22392_ (.A1(_02037_),
    .A2(_07346_),
    .B1(_07371_),
    .B2(_07351_),
    .Y(_07372_));
 AO21x1_ASAP7_75t_R _22393_ (.A1(_06366_),
    .A2(_07345_),
    .B(_07372_),
    .Y(_02498_));
 AND2x2_ASAP7_75t_R _22394_ (.A(_04306_),
    .B(_07366_),
    .Y(_07373_));
 AO21x2_ASAP7_75t_R _22395_ (.A1(_01676_),
    .A2(_07365_),
    .B(_07373_),
    .Y(_07374_));
 OAI22x1_ASAP7_75t_R _22396_ (.A1(_02036_),
    .A2(_07346_),
    .B1(_07374_),
    .B2(_07351_),
    .Y(_07375_));
 AO21x1_ASAP7_75t_R _22397_ (.A1(_06391_),
    .A2(_07345_),
    .B(_07375_),
    .Y(_02499_));
 AND2x2_ASAP7_75t_R _22398_ (.A(_04419_),
    .B(_07366_),
    .Y(_07376_));
 AO21x2_ASAP7_75t_R _22399_ (.A1(_01675_),
    .A2(_07365_),
    .B(_07376_),
    .Y(_07377_));
 OAI22x1_ASAP7_75t_R _22400_ (.A1(_02035_),
    .A2(_07346_),
    .B1(_07377_),
    .B2(_07351_),
    .Y(_07378_));
 AO21x1_ASAP7_75t_R _22401_ (.A1(_06411_),
    .A2(_07345_),
    .B(_07378_),
    .Y(_02500_));
 AND2x2_ASAP7_75t_R _22402_ (.A(_01487_),
    .B(_07366_),
    .Y(_07379_));
 AO21x2_ASAP7_75t_R _22403_ (.A1(_01674_),
    .A2(_07365_),
    .B(_07379_),
    .Y(_07380_));
 OAI22x1_ASAP7_75t_R _22404_ (.A1(_02034_),
    .A2(_07346_),
    .B1(_07380_),
    .B2(_07351_),
    .Y(_07381_));
 AO21x1_ASAP7_75t_R _22405_ (.A1(_06432_),
    .A2(_07345_),
    .B(_07381_),
    .Y(_02501_));
 BUFx6f_ASAP7_75t_R _22406_ (.A(_07300_),
    .Y(_07382_));
 BUFx12f_ASAP7_75t_R _22407_ (.A(_07303_),
    .Y(_07383_));
 AND2x2_ASAP7_75t_R _22408_ (.A(_04667_),
    .B(_07366_),
    .Y(_07384_));
 AO21x2_ASAP7_75t_R _22409_ (.A1(_01673_),
    .A2(_07365_),
    .B(_07384_),
    .Y(_07385_));
 BUFx12f_ASAP7_75t_R _22410_ (.A(_07278_),
    .Y(_07386_));
 OAI22x1_ASAP7_75t_R _22411_ (.A1(_02033_),
    .A2(_07383_),
    .B1(_07385_),
    .B2(_07386_),
    .Y(_07387_));
 AO21x1_ASAP7_75t_R _22412_ (.A1(_06454_),
    .A2(_07382_),
    .B(_07387_),
    .Y(_02502_));
 AND2x2_ASAP7_75t_R _22413_ (.A(_00016_),
    .B(_07308_),
    .Y(_07388_));
 AO21x2_ASAP7_75t_R _22414_ (.A1(_17997_),
    .A2(_07306_),
    .B(_07388_),
    .Y(_07389_));
 OAI22x1_ASAP7_75t_R _22415_ (.A1(_02032_),
    .A2(_07383_),
    .B1(_07389_),
    .B2(_07386_),
    .Y(_07390_));
 AO21x1_ASAP7_75t_R _22416_ (.A1(_05851_),
    .A2(_07382_),
    .B(_07390_),
    .Y(_02503_));
 AND2x2_ASAP7_75t_R _22417_ (.A(_01485_),
    .B(_07366_),
    .Y(_07391_));
 AO21x2_ASAP7_75t_R _22418_ (.A1(_01672_),
    .A2(_07365_),
    .B(_07391_),
    .Y(_07392_));
 OAI22x1_ASAP7_75t_R _22419_ (.A1(_02031_),
    .A2(_07383_),
    .B1(_07392_),
    .B2(_07386_),
    .Y(_07393_));
 AO21x1_ASAP7_75t_R _22420_ (.A1(_06480_),
    .A2(_07382_),
    .B(_07393_),
    .Y(_02504_));
 AND2x2_ASAP7_75t_R _22421_ (.A(_01484_),
    .B(_07308_),
    .Y(_07394_));
 AO21x2_ASAP7_75t_R _22422_ (.A1(_01671_),
    .A2(_07306_),
    .B(_07394_),
    .Y(_07395_));
 OAI22x1_ASAP7_75t_R _22423_ (.A1(_02030_),
    .A2(_07383_),
    .B1(_07395_),
    .B2(_07386_),
    .Y(_07396_));
 AO21x1_ASAP7_75t_R _22424_ (.A1(_06504_),
    .A2(_07382_),
    .B(_07396_),
    .Y(_02505_));
 AND2x2_ASAP7_75t_R _22425_ (.A(_14773_),
    .B(_07308_),
    .Y(_07397_));
 AO21x2_ASAP7_75t_R _22426_ (.A1(_00021_),
    .A2(_07306_),
    .B(_07397_),
    .Y(_07398_));
 OAI22x1_ASAP7_75t_R _22427_ (.A1(_01399_),
    .A2(_07383_),
    .B1(_07398_),
    .B2(_07386_),
    .Y(_07399_));
 AO21x1_ASAP7_75t_R _22428_ (.A1(_06556_),
    .A2(_07382_),
    .B(_07399_),
    .Y(_02506_));
 AND2x2_ASAP7_75t_R _22429_ (.A(_14837_),
    .B(_07308_),
    .Y(_07400_));
 AO21x2_ASAP7_75t_R _22430_ (.A1(_01670_),
    .A2(_07306_),
    .B(_07400_),
    .Y(_07401_));
 OAI22x1_ASAP7_75t_R _22431_ (.A1(_01400_),
    .A2(_07383_),
    .B1(_07401_),
    .B2(_07386_),
    .Y(_07402_));
 AO21x1_ASAP7_75t_R _22432_ (.A1(_06580_),
    .A2(_07382_),
    .B(_07402_),
    .Y(_02507_));
 AND2x2_ASAP7_75t_R _22433_ (.A(_14900_),
    .B(_07366_),
    .Y(_07403_));
 AO21x2_ASAP7_75t_R _22434_ (.A1(_01669_),
    .A2(_07365_),
    .B(_07403_),
    .Y(_07404_));
 OAI22x1_ASAP7_75t_R _22435_ (.A1(_01401_),
    .A2(_07383_),
    .B1(_07404_),
    .B2(_07386_),
    .Y(_07405_));
 AO21x1_ASAP7_75t_R _22436_ (.A1(_06600_),
    .A2(_07382_),
    .B(_07405_),
    .Y(_02508_));
 AND2x2_ASAP7_75t_R _22437_ (.A(_14966_),
    .B(_07366_),
    .Y(_07406_));
 AO21x2_ASAP7_75t_R _22438_ (.A1(_01668_),
    .A2(_07365_),
    .B(_07406_),
    .Y(_07407_));
 OAI22x1_ASAP7_75t_R _22439_ (.A1(_01402_),
    .A2(_07383_),
    .B1(_07407_),
    .B2(_07386_),
    .Y(_07408_));
 AO21x1_ASAP7_75t_R _22440_ (.A1(_06624_),
    .A2(_07382_),
    .B(_07408_),
    .Y(_02509_));
 AND2x2_ASAP7_75t_R _22441_ (.A(_01480_),
    .B(_07308_),
    .Y(_07409_));
 AO21x2_ASAP7_75t_R _22442_ (.A1(_01667_),
    .A2(_07306_),
    .B(_07409_),
    .Y(_07410_));
 OAI22x1_ASAP7_75t_R _22443_ (.A1(_02029_),
    .A2(_07383_),
    .B1(_07410_),
    .B2(_07386_),
    .Y(_07411_));
 AO21x1_ASAP7_75t_R _22444_ (.A1(_06650_),
    .A2(_07382_),
    .B(_07411_),
    .Y(_02510_));
 AND2x2_ASAP7_75t_R _22445_ (.A(_15099_),
    .B(_07366_),
    .Y(_07412_));
 AO21x2_ASAP7_75t_R _22446_ (.A1(_01666_),
    .A2(_07365_),
    .B(_07412_),
    .Y(_07413_));
 OAI22x1_ASAP7_75t_R _22447_ (.A1(_02028_),
    .A2(_07383_),
    .B1(_07413_),
    .B2(_07386_),
    .Y(_07414_));
 AO21x1_ASAP7_75t_R _22448_ (.A1(_06675_),
    .A2(_07382_),
    .B(_07414_),
    .Y(_02511_));
 AND2x2_ASAP7_75t_R _22449_ (.A(_15158_),
    .B(_07307_),
    .Y(_07415_));
 AO21x2_ASAP7_75t_R _22450_ (.A1(_01665_),
    .A2(_07305_),
    .B(_07415_),
    .Y(_07416_));
 OAI22x1_ASAP7_75t_R _22451_ (.A1(_02027_),
    .A2(_07303_),
    .B1(_07416_),
    .B2(_07278_),
    .Y(_07417_));
 AO21x1_ASAP7_75t_R _22452_ (.A1(_06699_),
    .A2(_07300_),
    .B(_07417_),
    .Y(_02512_));
 AND2x6_ASAP7_75t_R _22453_ (.A(_04993_),
    .B(_05888_),
    .Y(_07418_));
 NAND3x2_ASAP7_75t_R _22454_ (.B(_05897_),
    .C(_05766_),
    .Y(_07419_),
    .A(_07418_));
 BUFx6f_ASAP7_75t_R _22455_ (.A(_07419_),
    .Y(_07420_));
 BUFx6f_ASAP7_75t_R _22456_ (.A(_07419_),
    .Y(_07421_));
 NAND2x1_ASAP7_75t_R _22457_ (.A(_02026_),
    .B(_07421_),
    .Y(_07422_));
 OA21x2_ASAP7_75t_R _22458_ (.A1(_05811_),
    .A2(_07420_),
    .B(_07422_),
    .Y(_02513_));
 NAND2x1_ASAP7_75t_R _22459_ (.A(_02025_),
    .B(_07421_),
    .Y(_07423_));
 OA21x2_ASAP7_75t_R _22460_ (.A1(_05981_),
    .A2(_07420_),
    .B(_07423_),
    .Y(_02514_));
 NAND2x1_ASAP7_75t_R _22461_ (.A(_02024_),
    .B(_07421_),
    .Y(_07424_));
 OA21x2_ASAP7_75t_R _22462_ (.A1(_06025_),
    .A2(_07420_),
    .B(_07424_),
    .Y(_02515_));
 NAND2x1_ASAP7_75t_R _22463_ (.A(_02023_),
    .B(_07421_),
    .Y(_07425_));
 OA21x2_ASAP7_75t_R _22464_ (.A1(_06052_),
    .A2(_07420_),
    .B(_07425_),
    .Y(_02516_));
 NAND2x1_ASAP7_75t_R _22465_ (.A(_02022_),
    .B(_07421_),
    .Y(_07426_));
 OA21x2_ASAP7_75t_R _22466_ (.A1(_06082_),
    .A2(_07420_),
    .B(_07426_),
    .Y(_02517_));
 NAND2x1_ASAP7_75t_R _22467_ (.A(_02021_),
    .B(_07421_),
    .Y(_07427_));
 OA21x2_ASAP7_75t_R _22468_ (.A1(_06108_),
    .A2(_07420_),
    .B(_07427_),
    .Y(_02518_));
 NAND2x1_ASAP7_75t_R _22469_ (.A(_02020_),
    .B(_07421_),
    .Y(_07428_));
 OA21x2_ASAP7_75t_R _22470_ (.A1(_06131_),
    .A2(_07420_),
    .B(_07428_),
    .Y(_02519_));
 NAND2x1_ASAP7_75t_R _22471_ (.A(_02019_),
    .B(_07421_),
    .Y(_07429_));
 OA21x2_ASAP7_75t_R _22472_ (.A1(_06153_),
    .A2(_07420_),
    .B(_07429_),
    .Y(_02520_));
 BUFx12f_ASAP7_75t_R _22473_ (.A(_07419_),
    .Y(_07430_));
 NAND2x1_ASAP7_75t_R _22474_ (.A(_02018_),
    .B(_07430_),
    .Y(_07431_));
 OA21x2_ASAP7_75t_R _22475_ (.A1(_06179_),
    .A2(_07420_),
    .B(_07431_),
    .Y(_02521_));
 NAND2x1_ASAP7_75t_R _22476_ (.A(_02017_),
    .B(_07430_),
    .Y(_07432_));
 OA21x2_ASAP7_75t_R _22477_ (.A1(_06197_),
    .A2(_07420_),
    .B(_07432_),
    .Y(_02522_));
 BUFx6f_ASAP7_75t_R _22478_ (.A(_07419_),
    .Y(_07433_));
 NAND2x1_ASAP7_75t_R _22479_ (.A(_02016_),
    .B(_07430_),
    .Y(_07434_));
 OA21x2_ASAP7_75t_R _22480_ (.A1(_06219_),
    .A2(_07433_),
    .B(_07434_),
    .Y(_02523_));
 NAND2x1_ASAP7_75t_R _22481_ (.A(_02015_),
    .B(_07430_),
    .Y(_07435_));
 OA21x2_ASAP7_75t_R _22482_ (.A1(_06235_),
    .A2(_07433_),
    .B(_07435_),
    .Y(_02524_));
 NAND2x1_ASAP7_75t_R _22483_ (.A(_02014_),
    .B(_07430_),
    .Y(_07436_));
 OA21x2_ASAP7_75t_R _22484_ (.A1(_06255_),
    .A2(_07433_),
    .B(_07436_),
    .Y(_02525_));
 NAND2x1_ASAP7_75t_R _22485_ (.A(_02013_),
    .B(_07430_),
    .Y(_07437_));
 OA21x2_ASAP7_75t_R _22486_ (.A1(_06277_),
    .A2(_07433_),
    .B(_07437_),
    .Y(_02526_));
 NAND2x1_ASAP7_75t_R _22487_ (.A(_02012_),
    .B(_07430_),
    .Y(_07438_));
 OA21x2_ASAP7_75t_R _22488_ (.A1(_06298_),
    .A2(_07433_),
    .B(_07438_),
    .Y(_02527_));
 NAND2x1_ASAP7_75t_R _22489_ (.A(_02011_),
    .B(_07430_),
    .Y(_07439_));
 OA21x2_ASAP7_75t_R _22490_ (.A1(_06323_),
    .A2(_07433_),
    .B(_07439_),
    .Y(_02528_));
 NAND2x1_ASAP7_75t_R _22491_ (.A(_02010_),
    .B(_07430_),
    .Y(_07440_));
 OA21x2_ASAP7_75t_R _22492_ (.A1(_06343_),
    .A2(_07433_),
    .B(_07440_),
    .Y(_02529_));
 NAND2x1_ASAP7_75t_R _22493_ (.A(_02009_),
    .B(_07430_),
    .Y(_07441_));
 OA21x2_ASAP7_75t_R _22494_ (.A1(_06366_),
    .A2(_07433_),
    .B(_07441_),
    .Y(_02530_));
 BUFx12f_ASAP7_75t_R _22495_ (.A(_07419_),
    .Y(_07442_));
 NAND2x1_ASAP7_75t_R _22496_ (.A(_02008_),
    .B(_07442_),
    .Y(_07443_));
 OA21x2_ASAP7_75t_R _22497_ (.A1(_06391_),
    .A2(_07433_),
    .B(_07443_),
    .Y(_02531_));
 NAND2x1_ASAP7_75t_R _22498_ (.A(_02007_),
    .B(_07442_),
    .Y(_07444_));
 OA21x2_ASAP7_75t_R _22499_ (.A1(_06411_),
    .A2(_07433_),
    .B(_07444_),
    .Y(_02532_));
 BUFx6f_ASAP7_75t_R _22500_ (.A(_07419_),
    .Y(_07445_));
 NAND2x1_ASAP7_75t_R _22501_ (.A(_02006_),
    .B(_07442_),
    .Y(_07446_));
 OA21x2_ASAP7_75t_R _22502_ (.A1(_06432_),
    .A2(_07445_),
    .B(_07446_),
    .Y(_02533_));
 NAND2x1_ASAP7_75t_R _22503_ (.A(_02005_),
    .B(_07442_),
    .Y(_07447_));
 OA21x2_ASAP7_75t_R _22504_ (.A1(_06454_),
    .A2(_07445_),
    .B(_07447_),
    .Y(_02534_));
 NAND2x1_ASAP7_75t_R _22505_ (.A(_02004_),
    .B(_07442_),
    .Y(_07448_));
 OA21x2_ASAP7_75t_R _22506_ (.A1(_05851_),
    .A2(_07445_),
    .B(_07448_),
    .Y(_02535_));
 NAND2x1_ASAP7_75t_R _22507_ (.A(_02003_),
    .B(_07442_),
    .Y(_07449_));
 OA21x2_ASAP7_75t_R _22508_ (.A1(_06480_),
    .A2(_07445_),
    .B(_07449_),
    .Y(_02536_));
 NAND2x1_ASAP7_75t_R _22509_ (.A(_02002_),
    .B(_07442_),
    .Y(_07450_));
 OA21x2_ASAP7_75t_R _22510_ (.A1(_06504_),
    .A2(_07445_),
    .B(_07450_),
    .Y(_02537_));
 NAND2x1_ASAP7_75t_R _22511_ (.A(_02001_),
    .B(_07442_),
    .Y(_07451_));
 OA21x2_ASAP7_75t_R _22512_ (.A1(_06556_),
    .A2(_07445_),
    .B(_07451_),
    .Y(_02538_));
 NAND2x1_ASAP7_75t_R _22513_ (.A(_02000_),
    .B(_07442_),
    .Y(_07452_));
 OA21x2_ASAP7_75t_R _22514_ (.A1(_06580_),
    .A2(_07445_),
    .B(_07452_),
    .Y(_02539_));
 NAND2x1_ASAP7_75t_R _22515_ (.A(_01999_),
    .B(_07442_),
    .Y(_07453_));
 OA21x2_ASAP7_75t_R _22516_ (.A1(_06600_),
    .A2(_07445_),
    .B(_07453_),
    .Y(_02540_));
 NAND2x1_ASAP7_75t_R _22517_ (.A(_01998_),
    .B(_07419_),
    .Y(_07454_));
 OA21x2_ASAP7_75t_R _22518_ (.A1(_06624_),
    .A2(_07445_),
    .B(_07454_),
    .Y(_02541_));
 NAND2x1_ASAP7_75t_R _22519_ (.A(_01997_),
    .B(_07419_),
    .Y(_07455_));
 OA21x2_ASAP7_75t_R _22520_ (.A1(_06650_),
    .A2(_07445_),
    .B(_07455_),
    .Y(_02542_));
 NAND2x1_ASAP7_75t_R _22521_ (.A(_01996_),
    .B(_07419_),
    .Y(_07456_));
 OA21x2_ASAP7_75t_R _22522_ (.A1(_06675_),
    .A2(_07421_),
    .B(_07456_),
    .Y(_02543_));
 NAND2x1_ASAP7_75t_R _22523_ (.A(_01995_),
    .B(_07419_),
    .Y(_07457_));
 OA21x2_ASAP7_75t_R _22524_ (.A1(_06699_),
    .A2(_07421_),
    .B(_07457_),
    .Y(_02544_));
 NAND3x2_ASAP7_75t_R _22525_ (.B(_05072_),
    .C(_05897_),
    .Y(_07458_),
    .A(_07418_));
 BUFx6f_ASAP7_75t_R _22526_ (.A(_07458_),
    .Y(_07459_));
 BUFx6f_ASAP7_75t_R _22527_ (.A(_07458_),
    .Y(_07460_));
 NAND2x1_ASAP7_75t_R _22528_ (.A(_01994_),
    .B(_07460_),
    .Y(_07461_));
 OA21x2_ASAP7_75t_R _22529_ (.A1(_05811_),
    .A2(_07459_),
    .B(_07461_),
    .Y(_02545_));
 NAND2x1_ASAP7_75t_R _22530_ (.A(_01993_),
    .B(_07460_),
    .Y(_07462_));
 OA21x2_ASAP7_75t_R _22531_ (.A1(_05981_),
    .A2(_07459_),
    .B(_07462_),
    .Y(_02546_));
 NAND2x1_ASAP7_75t_R _22532_ (.A(_01992_),
    .B(_07460_),
    .Y(_07463_));
 OA21x2_ASAP7_75t_R _22533_ (.A1(_06025_),
    .A2(_07459_),
    .B(_07463_),
    .Y(_02547_));
 NAND2x1_ASAP7_75t_R _22534_ (.A(_01991_),
    .B(_07460_),
    .Y(_07464_));
 OA21x2_ASAP7_75t_R _22535_ (.A1(_06052_),
    .A2(_07459_),
    .B(_07464_),
    .Y(_02548_));
 NAND2x1_ASAP7_75t_R _22536_ (.A(_01990_),
    .B(_07460_),
    .Y(_07465_));
 OA21x2_ASAP7_75t_R _22537_ (.A1(_06082_),
    .A2(_07459_),
    .B(_07465_),
    .Y(_02549_));
 NAND2x1_ASAP7_75t_R _22538_ (.A(_01989_),
    .B(_07460_),
    .Y(_07466_));
 OA21x2_ASAP7_75t_R _22539_ (.A1(_06108_),
    .A2(_07459_),
    .B(_07466_),
    .Y(_02550_));
 NAND2x1_ASAP7_75t_R _22540_ (.A(_01988_),
    .B(_07460_),
    .Y(_07467_));
 OA21x2_ASAP7_75t_R _22541_ (.A1(_06131_),
    .A2(_07459_),
    .B(_07467_),
    .Y(_02551_));
 NAND2x1_ASAP7_75t_R _22542_ (.A(_01987_),
    .B(_07460_),
    .Y(_07468_));
 OA21x2_ASAP7_75t_R _22543_ (.A1(_06153_),
    .A2(_07459_),
    .B(_07468_),
    .Y(_02552_));
 BUFx6f_ASAP7_75t_R _22544_ (.A(_07458_),
    .Y(_07469_));
 NAND2x1_ASAP7_75t_R _22545_ (.A(_01986_),
    .B(_07469_),
    .Y(_07470_));
 OA21x2_ASAP7_75t_R _22546_ (.A1(_06179_),
    .A2(_07459_),
    .B(_07470_),
    .Y(_02553_));
 NAND2x1_ASAP7_75t_R _22547_ (.A(_01985_),
    .B(_07469_),
    .Y(_07471_));
 OA21x2_ASAP7_75t_R _22548_ (.A1(_06197_),
    .A2(_07459_),
    .B(_07471_),
    .Y(_02554_));
 BUFx6f_ASAP7_75t_R _22549_ (.A(_07458_),
    .Y(_07472_));
 NAND2x1_ASAP7_75t_R _22550_ (.A(_01984_),
    .B(_07469_),
    .Y(_07473_));
 OA21x2_ASAP7_75t_R _22551_ (.A1(_06219_),
    .A2(_07472_),
    .B(_07473_),
    .Y(_02555_));
 NAND2x1_ASAP7_75t_R _22552_ (.A(_01983_),
    .B(_07469_),
    .Y(_07474_));
 OA21x2_ASAP7_75t_R _22553_ (.A1(_06235_),
    .A2(_07472_),
    .B(_07474_),
    .Y(_02556_));
 NAND2x1_ASAP7_75t_R _22554_ (.A(_01982_),
    .B(_07469_),
    .Y(_07475_));
 OA21x2_ASAP7_75t_R _22555_ (.A1(_06255_),
    .A2(_07472_),
    .B(_07475_),
    .Y(_02557_));
 NAND2x1_ASAP7_75t_R _22556_ (.A(_01981_),
    .B(_07469_),
    .Y(_07476_));
 OA21x2_ASAP7_75t_R _22557_ (.A1(_06277_),
    .A2(_07472_),
    .B(_07476_),
    .Y(_02558_));
 NAND2x1_ASAP7_75t_R _22558_ (.A(_01980_),
    .B(_07469_),
    .Y(_07477_));
 OA21x2_ASAP7_75t_R _22559_ (.A1(_06298_),
    .A2(_07472_),
    .B(_07477_),
    .Y(_02559_));
 NAND2x1_ASAP7_75t_R _22560_ (.A(_01979_),
    .B(_07469_),
    .Y(_07478_));
 OA21x2_ASAP7_75t_R _22561_ (.A1(_06323_),
    .A2(_07472_),
    .B(_07478_),
    .Y(_02560_));
 NAND2x1_ASAP7_75t_R _22562_ (.A(_01978_),
    .B(_07469_),
    .Y(_07479_));
 OA21x2_ASAP7_75t_R _22563_ (.A1(_06343_),
    .A2(_07472_),
    .B(_07479_),
    .Y(_02561_));
 NAND2x1_ASAP7_75t_R _22564_ (.A(_01977_),
    .B(_07469_),
    .Y(_07480_));
 OA21x2_ASAP7_75t_R _22565_ (.A1(_06366_),
    .A2(_07472_),
    .B(_07480_),
    .Y(_02562_));
 BUFx12f_ASAP7_75t_R _22566_ (.A(_07458_),
    .Y(_07481_));
 NAND2x1_ASAP7_75t_R _22567_ (.A(_01976_),
    .B(_07481_),
    .Y(_07482_));
 OA21x2_ASAP7_75t_R _22568_ (.A1(_06391_),
    .A2(_07472_),
    .B(_07482_),
    .Y(_02563_));
 NAND2x1_ASAP7_75t_R _22569_ (.A(_01975_),
    .B(_07481_),
    .Y(_07483_));
 OA21x2_ASAP7_75t_R _22570_ (.A1(_06411_),
    .A2(_07472_),
    .B(_07483_),
    .Y(_02564_));
 BUFx6f_ASAP7_75t_R _22571_ (.A(_07458_),
    .Y(_07484_));
 NAND2x1_ASAP7_75t_R _22572_ (.A(_01974_),
    .B(_07481_),
    .Y(_07485_));
 OA21x2_ASAP7_75t_R _22573_ (.A1(_06432_),
    .A2(_07484_),
    .B(_07485_),
    .Y(_02565_));
 NAND2x1_ASAP7_75t_R _22574_ (.A(_01973_),
    .B(_07481_),
    .Y(_07486_));
 OA21x2_ASAP7_75t_R _22575_ (.A1(_06454_),
    .A2(_07484_),
    .B(_07486_),
    .Y(_02566_));
 NAND2x1_ASAP7_75t_R _22576_ (.A(_01972_),
    .B(_07481_),
    .Y(_07487_));
 OA21x2_ASAP7_75t_R _22577_ (.A1(_05851_),
    .A2(_07484_),
    .B(_07487_),
    .Y(_02567_));
 NAND2x1_ASAP7_75t_R _22578_ (.A(_01971_),
    .B(_07481_),
    .Y(_07488_));
 OA21x2_ASAP7_75t_R _22579_ (.A1(_06480_),
    .A2(_07484_),
    .B(_07488_),
    .Y(_02568_));
 NAND2x1_ASAP7_75t_R _22580_ (.A(_01970_),
    .B(_07481_),
    .Y(_07489_));
 OA21x2_ASAP7_75t_R _22581_ (.A1(_06504_),
    .A2(_07484_),
    .B(_07489_),
    .Y(_02569_));
 NAND2x1_ASAP7_75t_R _22582_ (.A(_01969_),
    .B(_07481_),
    .Y(_07490_));
 OA21x2_ASAP7_75t_R _22583_ (.A1(_06556_),
    .A2(_07484_),
    .B(_07490_),
    .Y(_02570_));
 NAND2x1_ASAP7_75t_R _22584_ (.A(_01968_),
    .B(_07481_),
    .Y(_07491_));
 OA21x2_ASAP7_75t_R _22585_ (.A1(_06580_),
    .A2(_07484_),
    .B(_07491_),
    .Y(_02571_));
 NAND2x1_ASAP7_75t_R _22586_ (.A(_01967_),
    .B(_07481_),
    .Y(_07492_));
 OA21x2_ASAP7_75t_R _22587_ (.A1(_06600_),
    .A2(_07484_),
    .B(_07492_),
    .Y(_02572_));
 NAND2x1_ASAP7_75t_R _22588_ (.A(_01966_),
    .B(_07458_),
    .Y(_07493_));
 OA21x2_ASAP7_75t_R _22589_ (.A1(_06624_),
    .A2(_07484_),
    .B(_07493_),
    .Y(_02573_));
 NAND2x1_ASAP7_75t_R _22590_ (.A(_01965_),
    .B(_07458_),
    .Y(_07494_));
 OA21x2_ASAP7_75t_R _22591_ (.A1(_06650_),
    .A2(_07484_),
    .B(_07494_),
    .Y(_02574_));
 NAND2x1_ASAP7_75t_R _22592_ (.A(_01964_),
    .B(_07458_),
    .Y(_07495_));
 OA21x2_ASAP7_75t_R _22593_ (.A1(_06675_),
    .A2(_07460_),
    .B(_07495_),
    .Y(_02575_));
 NAND2x1_ASAP7_75t_R _22594_ (.A(_01963_),
    .B(_07458_),
    .Y(_07496_));
 OA21x2_ASAP7_75t_R _22595_ (.A1(_06699_),
    .A2(_07460_),
    .B(_07496_),
    .Y(_02576_));
 NAND3x1_ASAP7_75t_R _22596_ (.A(_04991_),
    .B(_07278_),
    .C(_07280_),
    .Y(_07497_));
 OR2x6_ASAP7_75t_R _22597_ (.A(_00334_),
    .B(_05504_),
    .Y(_07498_));
 AND2x4_ASAP7_75t_R _22598_ (.A(_07497_),
    .B(_07498_),
    .Y(_07499_));
 BUFx6f_ASAP7_75t_R _22599_ (.A(_07499_),
    .Y(_07500_));
 OA21x2_ASAP7_75t_R _22600_ (.A1(_05749_),
    .A2(_05801_),
    .B(_07500_),
    .Y(_07501_));
 BUFx6f_ASAP7_75t_R _22601_ (.A(_07501_),
    .Y(_07502_));
 BUFx6f_ASAP7_75t_R _22602_ (.A(_07498_),
    .Y(_07503_));
 BUFx12f_ASAP7_75t_R _22603_ (.A(_07503_),
    .Y(_07504_));
 AND2x2_ASAP7_75t_R _22604_ (.A(_01391_),
    .B(_05400_),
    .Y(_07505_));
 AND4x1_ASAP7_75t_R _22605_ (.A(_01758_),
    .B(_01759_),
    .C(_05175_),
    .D(_07505_),
    .Y(_07506_));
 OR2x2_ASAP7_75t_R _22606_ (.A(_05509_),
    .B(_07506_),
    .Y(_07507_));
 AND3x1_ASAP7_75t_R _22607_ (.A(_15594_),
    .B(_07283_),
    .C(\cs_registers_i.priv_mode_id_o[0] ),
    .Y(_07508_));
 AO21x1_ASAP7_75t_R _22608_ (.A1(_16337_),
    .A2(_05416_),
    .B(_07508_),
    .Y(_07509_));
 INVx1_ASAP7_75t_R _22609_ (.A(_07509_),
    .Y(_07510_));
 AO221x1_ASAP7_75t_R _22610_ (.A1(_01758_),
    .A2(_01759_),
    .B1(_14103_),
    .B2(_05164_),
    .C(_05411_),
    .Y(_07511_));
 BUFx6f_ASAP7_75t_R _22611_ (.A(_07511_),
    .Y(_07512_));
 BUFx6f_ASAP7_75t_R _22612_ (.A(_05400_),
    .Y(_07513_));
 OA211x2_ASAP7_75t_R _22613_ (.A1(_05412_),
    .A2(_07510_),
    .B(_07512_),
    .C(_07513_),
    .Y(_07514_));
 OA21x2_ASAP7_75t_R _22614_ (.A1(_07507_),
    .A2(_07514_),
    .B(_05498_),
    .Y(_07515_));
 BUFx12f_ASAP7_75t_R _22615_ (.A(_07497_),
    .Y(_07516_));
 BUFx12f_ASAP7_75t_R _22616_ (.A(_07516_),
    .Y(_07517_));
 OAI22x1_ASAP7_75t_R _22617_ (.A1(_01874_),
    .A2(_07504_),
    .B1(_07515_),
    .B2(_07517_),
    .Y(_07518_));
 AO21x1_ASAP7_75t_R _22618_ (.A1(_05811_),
    .A2(_07500_),
    .B(_07518_),
    .Y(_07519_));
 NAND2x1_ASAP7_75t_R _22619_ (.A(_01962_),
    .B(_07502_),
    .Y(_07520_));
 OA21x2_ASAP7_75t_R _22620_ (.A1(_07502_),
    .A2(_07519_),
    .B(_07520_),
    .Y(_02577_));
 OAI21x1_ASAP7_75t_R _22621_ (.A1(_05749_),
    .A2(_05801_),
    .B(_07500_),
    .Y(_07521_));
 NAND2x1_ASAP7_75t_R _22622_ (.A(_06235_),
    .B(_07500_),
    .Y(_07522_));
 BUFx6f_ASAP7_75t_R _22623_ (.A(_07498_),
    .Y(_07523_));
 NOR2x1_ASAP7_75t_R _22624_ (.A(_13233_),
    .B(_01539_),
    .Y(_07524_));
 NOR2x1_ASAP7_75t_R _22625_ (.A(_05175_),
    .B(_07509_),
    .Y(_07525_));
 AO21x1_ASAP7_75t_R _22626_ (.A1(_01758_),
    .A2(_05175_),
    .B(_07525_),
    .Y(_07526_));
 AO21x1_ASAP7_75t_R _22627_ (.A1(_01391_),
    .A2(_07526_),
    .B(_07507_),
    .Y(_07527_));
 OA21x2_ASAP7_75t_R _22628_ (.A1(_07524_),
    .A2(_07527_),
    .B(_05518_),
    .Y(_07528_));
 BUFx6f_ASAP7_75t_R _22629_ (.A(_07516_),
    .Y(_07529_));
 OA22x2_ASAP7_75t_R _22630_ (.A1(_01873_),
    .A2(_07523_),
    .B1(_07528_),
    .B2(_07529_),
    .Y(_07530_));
 AND3x1_ASAP7_75t_R _22631_ (.A(_07521_),
    .B(_07522_),
    .C(_07530_),
    .Y(_07531_));
 AOI21x1_ASAP7_75t_R _22632_ (.A1(_01961_),
    .A2(_07502_),
    .B(_07531_),
    .Y(_02578_));
 NOR2x1_ASAP7_75t_R _22633_ (.A(_05496_),
    .B(_05445_),
    .Y(_07532_));
 NOR2x1_ASAP7_75t_R _22634_ (.A(_05438_),
    .B(_05441_),
    .Y(_07533_));
 OA21x2_ASAP7_75t_R _22635_ (.A1(_05422_),
    .A2(_05425_),
    .B(_07533_),
    .Y(_07534_));
 OR4x1_ASAP7_75t_R _22636_ (.A(_05435_),
    .B(_05515_),
    .C(_07532_),
    .D(_07534_),
    .Y(_07535_));
 BUFx6f_ASAP7_75t_R _22637_ (.A(_07512_),
    .Y(_07536_));
 INVx1_ASAP7_75t_R _22638_ (.A(_07536_),
    .Y(_07537_));
 AO32x1_ASAP7_75t_R _22639_ (.A1(_05449_),
    .A2(_05453_),
    .A3(_07535_),
    .B1(_07537_),
    .B2(_05406_),
    .Y(_07538_));
 AND3x4_ASAP7_75t_R _22640_ (.A(_04991_),
    .B(_07278_),
    .C(_07280_),
    .Y(_07539_));
 BUFx6f_ASAP7_75t_R _22641_ (.A(_07539_),
    .Y(_07540_));
 NOR2x1_ASAP7_75t_R _22642_ (.A(_01872_),
    .B(_07504_),
    .Y(_07541_));
 AO221x1_ASAP7_75t_R _22643_ (.A1(_05850_),
    .A2(_07500_),
    .B1(_07538_),
    .B2(_07540_),
    .C(_07541_),
    .Y(_07542_));
 NAND2x1_ASAP7_75t_R _22644_ (.A(_01960_),
    .B(_07502_),
    .Y(_07543_));
 OA21x2_ASAP7_75t_R _22645_ (.A1(_07502_),
    .A2(_07542_),
    .B(_07543_),
    .Y(_02579_));
 INVx1_ASAP7_75t_R _22646_ (.A(_01959_),
    .Y(_07544_));
 NAND2x1_ASAP7_75t_R _22647_ (.A(_06555_),
    .B(_07500_),
    .Y(_07545_));
 NOR2x1_ASAP7_75t_R _22648_ (.A(_05442_),
    .B(_05515_),
    .Y(_07546_));
 OR4x1_ASAP7_75t_R _22649_ (.A(_05444_),
    .B(_01918_),
    .C(_05419_),
    .D(_05432_),
    .Y(_07547_));
 AO21x2_ASAP7_75t_R _22650_ (.A1(_07546_),
    .A2(_07547_),
    .B(_05478_),
    .Y(_07548_));
 OR3x1_ASAP7_75t_R _22651_ (.A(_16337_),
    .B(_05412_),
    .C(_05509_),
    .Y(_07549_));
 AO21x1_ASAP7_75t_R _22652_ (.A1(_07548_),
    .A2(_07549_),
    .B(_07516_),
    .Y(_07550_));
 OA211x2_ASAP7_75t_R _22653_ (.A1(_01871_),
    .A2(_07504_),
    .B(_07545_),
    .C(_07550_),
    .Y(_07551_));
 NOR2x1_ASAP7_75t_R _22654_ (.A(_07502_),
    .B(_07551_),
    .Y(_07552_));
 AO21x1_ASAP7_75t_R _22655_ (.A1(_07544_),
    .A2(_07502_),
    .B(_07552_),
    .Y(_02580_));
 NAND2x1_ASAP7_75t_R _22656_ (.A(_06580_),
    .B(_07500_),
    .Y(_07553_));
 INVx1_ASAP7_75t_R _22657_ (.A(_05496_),
    .Y(_07554_));
 AO21x2_ASAP7_75t_R _22658_ (.A1(_07554_),
    .A2(_05495_),
    .B(_05478_),
    .Y(_07555_));
 OA211x2_ASAP7_75t_R _22659_ (.A1(_01870_),
    .A2(_07504_),
    .B(_07521_),
    .C(_07555_),
    .Y(_07556_));
 AOI22x1_ASAP7_75t_R _22660_ (.A1(_01958_),
    .A2(_07502_),
    .B1(_07553_),
    .B2(_07556_),
    .Y(_02581_));
 NAND2x1_ASAP7_75t_R _22661_ (.A(_06504_),
    .B(_07500_),
    .Y(_07557_));
 OA211x2_ASAP7_75t_R _22662_ (.A1(_01869_),
    .A2(_07504_),
    .B(_07521_),
    .C(_05478_),
    .Y(_07558_));
 AOI22x1_ASAP7_75t_R _22663_ (.A1(_01957_),
    .A2(_07502_),
    .B1(_07557_),
    .B2(_07558_),
    .Y(_02582_));
 OAI21x1_ASAP7_75t_R _22664_ (.A1(_05749_),
    .A2(_05791_),
    .B(_07499_),
    .Y(_07559_));
 BUFx6f_ASAP7_75t_R _22665_ (.A(_07559_),
    .Y(_07560_));
 OAI22x1_ASAP7_75t_R _22666_ (.A1(_01865_),
    .A2(_07504_),
    .B1(_07560_),
    .B2(_01956_),
    .Y(_02583_));
 OA21x2_ASAP7_75t_R _22667_ (.A1(_05749_),
    .A2(_05791_),
    .B(_07499_),
    .Y(_07561_));
 BUFx6f_ASAP7_75t_R _22668_ (.A(_07561_),
    .Y(_07562_));
 BUFx12f_ASAP7_75t_R _22669_ (.A(_07562_),
    .Y(_07563_));
 NAND2x2_ASAP7_75t_R _22670_ (.A(_07516_),
    .B(_07498_),
    .Y(_07564_));
 BUFx6f_ASAP7_75t_R _22671_ (.A(_07564_),
    .Y(_07565_));
 BUFx6f_ASAP7_75t_R _22672_ (.A(_07516_),
    .Y(_07566_));
 OA22x2_ASAP7_75t_R _22673_ (.A1(_07310_),
    .A2(_07566_),
    .B1(_07523_),
    .B2(_01864_),
    .Y(_07567_));
 OA211x2_ASAP7_75t_R _22674_ (.A1(_06923_),
    .A2(_07565_),
    .B(_07560_),
    .C(_07567_),
    .Y(_07568_));
 AOI21x1_ASAP7_75t_R _22675_ (.A1(_01955_),
    .A2(_07563_),
    .B(_07568_),
    .Y(_02584_));
 OA22x2_ASAP7_75t_R _22676_ (.A1(_07314_),
    .A2(_07566_),
    .B1(_07523_),
    .B2(_01863_),
    .Y(_07569_));
 OA211x2_ASAP7_75t_R _22677_ (.A1(_06937_),
    .A2(_07565_),
    .B(_07560_),
    .C(_07569_),
    .Y(_07570_));
 AOI21x1_ASAP7_75t_R _22678_ (.A1(_01954_),
    .A2(_07563_),
    .B(_07570_),
    .Y(_02585_));
 INVx1_ASAP7_75t_R _22679_ (.A(_06051_),
    .Y(_07571_));
 OA22x2_ASAP7_75t_R _22680_ (.A1(_07318_),
    .A2(_07566_),
    .B1(_07523_),
    .B2(_01862_),
    .Y(_07572_));
 OA211x2_ASAP7_75t_R _22681_ (.A1(_07571_),
    .A2(_07565_),
    .B(_07560_),
    .C(_07572_),
    .Y(_07573_));
 AOI21x1_ASAP7_75t_R _22682_ (.A1(_01953_),
    .A2(_07563_),
    .B(_07573_),
    .Y(_02586_));
 OA22x2_ASAP7_75t_R _22683_ (.A1(_07323_),
    .A2(_07566_),
    .B1(_07523_),
    .B2(_01861_),
    .Y(_07574_));
 OA211x2_ASAP7_75t_R _22684_ (.A1(_06961_),
    .A2(_07565_),
    .B(_07560_),
    .C(_07574_),
    .Y(_07575_));
 AOI21x1_ASAP7_75t_R _22685_ (.A1(_01952_),
    .A2(_07563_),
    .B(_07575_),
    .Y(_02587_));
 INVx1_ASAP7_75t_R _22686_ (.A(_06108_),
    .Y(_07576_));
 BUFx6f_ASAP7_75t_R _22687_ (.A(_07516_),
    .Y(_07577_));
 OA22x2_ASAP7_75t_R _22688_ (.A1(_07326_),
    .A2(_07577_),
    .B1(_07523_),
    .B2(_01860_),
    .Y(_07578_));
 OA211x2_ASAP7_75t_R _22689_ (.A1(_07576_),
    .A2(_07565_),
    .B(_07560_),
    .C(_07578_),
    .Y(_07579_));
 AOI21x1_ASAP7_75t_R _22690_ (.A1(_01951_),
    .A2(_07563_),
    .B(_07579_),
    .Y(_02588_));
 BUFx3_ASAP7_75t_R _22691_ (.A(_07559_),
    .Y(_07580_));
 BUFx6f_ASAP7_75t_R _22692_ (.A(_07498_),
    .Y(_07581_));
 OA22x2_ASAP7_75t_R _22693_ (.A1(_07330_),
    .A2(_07577_),
    .B1(_07581_),
    .B2(_01859_),
    .Y(_07582_));
 OA211x2_ASAP7_75t_R _22694_ (.A1(_06968_),
    .A2(_07565_),
    .B(_07580_),
    .C(_07582_),
    .Y(_07583_));
 AOI21x1_ASAP7_75t_R _22695_ (.A1(_01950_),
    .A2(_07563_),
    .B(_07583_),
    .Y(_02589_));
 OA22x2_ASAP7_75t_R _22696_ (.A1(_07333_),
    .A2(_07577_),
    .B1(_07581_),
    .B2(_01858_),
    .Y(_07584_));
 OA211x2_ASAP7_75t_R _22697_ (.A1(_06973_),
    .A2(_07565_),
    .B(_07580_),
    .C(_07584_),
    .Y(_07585_));
 AOI21x1_ASAP7_75t_R _22698_ (.A1(_01949_),
    .A2(_07563_),
    .B(_07585_),
    .Y(_02590_));
 OA22x2_ASAP7_75t_R _22699_ (.A1(_07337_),
    .A2(_07577_),
    .B1(_07581_),
    .B2(_01857_),
    .Y(_07586_));
 OA211x2_ASAP7_75t_R _22700_ (.A1(_06978_),
    .A2(_07565_),
    .B(_07580_),
    .C(_07586_),
    .Y(_07587_));
 AOI21x1_ASAP7_75t_R _22701_ (.A1(_01948_),
    .A2(_07563_),
    .B(_07587_),
    .Y(_02591_));
 INVx2_ASAP7_75t_R _22702_ (.A(_06196_),
    .Y(_07588_));
 OA22x2_ASAP7_75t_R _22703_ (.A1(_07340_),
    .A2(_07577_),
    .B1(_07581_),
    .B2(_01856_),
    .Y(_07589_));
 OA211x2_ASAP7_75t_R _22704_ (.A1(_07588_),
    .A2(_07565_),
    .B(_07580_),
    .C(_07589_),
    .Y(_07590_));
 AOI21x1_ASAP7_75t_R _22705_ (.A1(_01947_),
    .A2(_07563_),
    .B(_07590_),
    .Y(_02592_));
 OA22x2_ASAP7_75t_R _22706_ (.A1(_07343_),
    .A2(_07577_),
    .B1(_07581_),
    .B2(_01855_),
    .Y(_07591_));
 OA211x2_ASAP7_75t_R _22707_ (.A1(_06995_),
    .A2(_07565_),
    .B(_07580_),
    .C(_07591_),
    .Y(_07592_));
 AOI21x1_ASAP7_75t_R _22708_ (.A1(_01946_),
    .A2(_07563_),
    .B(_07592_),
    .Y(_02593_));
 BUFx12f_ASAP7_75t_R _22709_ (.A(_07562_),
    .Y(_07593_));
 OA22x2_ASAP7_75t_R _22710_ (.A1(_07350_),
    .A2(_07517_),
    .B1(_07523_),
    .B2(_01854_),
    .Y(_07594_));
 AND3x1_ASAP7_75t_R _22711_ (.A(_07522_),
    .B(_07560_),
    .C(_07594_),
    .Y(_07595_));
 AOI21x1_ASAP7_75t_R _22712_ (.A1(_01945_),
    .A2(_07593_),
    .B(_07595_),
    .Y(_02594_));
 BUFx12f_ASAP7_75t_R _22713_ (.A(_07562_),
    .Y(_07596_));
 OAI22x1_ASAP7_75t_R _22714_ (.A1(_07354_),
    .A2(_07517_),
    .B1(_07504_),
    .B2(_01853_),
    .Y(_07597_));
 AO21x1_ASAP7_75t_R _22715_ (.A1(_06255_),
    .A2(_07500_),
    .B(_07597_),
    .Y(_07598_));
 NAND2x1_ASAP7_75t_R _22716_ (.A(_01944_),
    .B(_07562_),
    .Y(_07599_));
 OA21x2_ASAP7_75t_R _22717_ (.A1(_07596_),
    .A2(_07598_),
    .B(_07599_),
    .Y(_02595_));
 BUFx6f_ASAP7_75t_R _22718_ (.A(_07564_),
    .Y(_07600_));
 OA22x2_ASAP7_75t_R _22719_ (.A1(_07357_),
    .A2(_07577_),
    .B1(_07581_),
    .B2(_01852_),
    .Y(_07601_));
 OA211x2_ASAP7_75t_R _22720_ (.A1(_07006_),
    .A2(_07600_),
    .B(_07580_),
    .C(_07601_),
    .Y(_07602_));
 AOI21x1_ASAP7_75t_R _22721_ (.A1(_01943_),
    .A2(_07593_),
    .B(_07602_),
    .Y(_02596_));
 INVx2_ASAP7_75t_R _22722_ (.A(_06297_),
    .Y(_07603_));
 OA22x2_ASAP7_75t_R _22723_ (.A1(_07360_),
    .A2(_07577_),
    .B1(_07581_),
    .B2(_01851_),
    .Y(_07604_));
 OA211x2_ASAP7_75t_R _22724_ (.A1(_07603_),
    .A2(_07600_),
    .B(_07580_),
    .C(_07604_),
    .Y(_07605_));
 AOI21x1_ASAP7_75t_R _22725_ (.A1(_01942_),
    .A2(_07593_),
    .B(_07605_),
    .Y(_02597_));
 OA22x2_ASAP7_75t_R _22726_ (.A1(_07363_),
    .A2(_07577_),
    .B1(_07581_),
    .B2(_01850_),
    .Y(_07606_));
 OA211x2_ASAP7_75t_R _22727_ (.A1(_07016_),
    .A2(_07600_),
    .B(_07580_),
    .C(_07606_),
    .Y(_07607_));
 AOI21x1_ASAP7_75t_R _22728_ (.A1(_01941_),
    .A2(_07593_),
    .B(_07607_),
    .Y(_02598_));
 OA22x2_ASAP7_75t_R _22729_ (.A1(_07368_),
    .A2(_07577_),
    .B1(_07581_),
    .B2(_01849_),
    .Y(_07608_));
 OA211x2_ASAP7_75t_R _22730_ (.A1(_06344_),
    .A2(_07600_),
    .B(_07580_),
    .C(_07608_),
    .Y(_07609_));
 AOI21x1_ASAP7_75t_R _22731_ (.A1(_01940_),
    .A2(_07593_),
    .B(_07609_),
    .Y(_02599_));
 BUFx6f_ASAP7_75t_R _22732_ (.A(_07516_),
    .Y(_07610_));
 OA22x2_ASAP7_75t_R _22733_ (.A1(_07371_),
    .A2(_07610_),
    .B1(_07581_),
    .B2(_01848_),
    .Y(_07611_));
 OA211x2_ASAP7_75t_R _22734_ (.A1(_07026_),
    .A2(_07600_),
    .B(_07580_),
    .C(_07611_),
    .Y(_07612_));
 AOI21x1_ASAP7_75t_R _22735_ (.A1(_01939_),
    .A2(_07593_),
    .B(_07612_),
    .Y(_02600_));
 INVx2_ASAP7_75t_R _22736_ (.A(_06390_),
    .Y(_07613_));
 BUFx6f_ASAP7_75t_R _22737_ (.A(_07559_),
    .Y(_07614_));
 OA22x2_ASAP7_75t_R _22738_ (.A1(_07374_),
    .A2(_07610_),
    .B1(_07503_),
    .B2(_01847_),
    .Y(_07615_));
 OA211x2_ASAP7_75t_R _22739_ (.A1(_07613_),
    .A2(_07600_),
    .B(_07614_),
    .C(_07615_),
    .Y(_07616_));
 AOI21x1_ASAP7_75t_R _22740_ (.A1(_01938_),
    .A2(_07593_),
    .B(_07616_),
    .Y(_02601_));
 OA22x2_ASAP7_75t_R _22741_ (.A1(_07377_),
    .A2(_07610_),
    .B1(_07503_),
    .B2(_01846_),
    .Y(_07617_));
 OA211x2_ASAP7_75t_R _22742_ (.A1(_07037_),
    .A2(_07600_),
    .B(_07614_),
    .C(_07617_),
    .Y(_07618_));
 AOI21x1_ASAP7_75t_R _22743_ (.A1(_01937_),
    .A2(_07593_),
    .B(_07618_),
    .Y(_02602_));
 OA22x2_ASAP7_75t_R _22744_ (.A1(_07380_),
    .A2(_07610_),
    .B1(_07503_),
    .B2(_01845_),
    .Y(_07619_));
 OA211x2_ASAP7_75t_R _22745_ (.A1(_07044_),
    .A2(_07600_),
    .B(_07614_),
    .C(_07619_),
    .Y(_07620_));
 AOI21x1_ASAP7_75t_R _22746_ (.A1(_01936_),
    .A2(_07593_),
    .B(_07620_),
    .Y(_02603_));
 OA22x2_ASAP7_75t_R _22747_ (.A1(_07385_),
    .A2(_07610_),
    .B1(_07503_),
    .B2(_01844_),
    .Y(_07621_));
 OA211x2_ASAP7_75t_R _22748_ (.A1(_07046_),
    .A2(_07600_),
    .B(_07614_),
    .C(_07621_),
    .Y(_07622_));
 AOI21x1_ASAP7_75t_R _22749_ (.A1(_01935_),
    .A2(_07593_),
    .B(_07622_),
    .Y(_02604_));
 OAI22x1_ASAP7_75t_R _22750_ (.A1(_07389_),
    .A2(_07517_),
    .B1(_07504_),
    .B2(_01843_),
    .Y(_07623_));
 AO21x1_ASAP7_75t_R _22751_ (.A1(_05851_),
    .A2(_07500_),
    .B(_07623_),
    .Y(_07624_));
 NAND2x1_ASAP7_75t_R _22752_ (.A(_01934_),
    .B(_07562_),
    .Y(_07625_));
 OA21x2_ASAP7_75t_R _22753_ (.A1(_07562_),
    .A2(_07624_),
    .B(_07625_),
    .Y(_02605_));
 INVx2_ASAP7_75t_R _22754_ (.A(_06479_),
    .Y(_07626_));
 OA22x2_ASAP7_75t_R _22755_ (.A1(_07392_),
    .A2(_07610_),
    .B1(_07503_),
    .B2(_01842_),
    .Y(_07627_));
 OA211x2_ASAP7_75t_R _22756_ (.A1(_07626_),
    .A2(_07600_),
    .B(_07614_),
    .C(_07627_),
    .Y(_07628_));
 AOI21x1_ASAP7_75t_R _22757_ (.A1(_01933_),
    .A2(_07596_),
    .B(_07628_),
    .Y(_02606_));
 OA22x2_ASAP7_75t_R _22758_ (.A1(_07395_),
    .A2(_07517_),
    .B1(_07523_),
    .B2(_01841_),
    .Y(_07629_));
 AND3x1_ASAP7_75t_R _22759_ (.A(_07557_),
    .B(_07560_),
    .C(_07629_),
    .Y(_07630_));
 AOI21x1_ASAP7_75t_R _22760_ (.A1(_01932_),
    .A2(_07596_),
    .B(_07630_),
    .Y(_02607_));
 OA22x2_ASAP7_75t_R _22761_ (.A1(_07398_),
    .A2(_07529_),
    .B1(_07523_),
    .B2(_01840_),
    .Y(_07631_));
 AND3x1_ASAP7_75t_R _22762_ (.A(_07545_),
    .B(_07560_),
    .C(_07631_),
    .Y(_07632_));
 AOI21x1_ASAP7_75t_R _22763_ (.A1(_01931_),
    .A2(_07596_),
    .B(_07632_),
    .Y(_02608_));
 OA22x2_ASAP7_75t_R _22764_ (.A1(_07401_),
    .A2(_07529_),
    .B1(_07523_),
    .B2(_01839_),
    .Y(_07633_));
 AND3x1_ASAP7_75t_R _22765_ (.A(_07553_),
    .B(_07560_),
    .C(_07633_),
    .Y(_07634_));
 AOI21x1_ASAP7_75t_R _22766_ (.A1(_01930_),
    .A2(_07596_),
    .B(_07634_),
    .Y(_02609_));
 OA22x2_ASAP7_75t_R _22767_ (.A1(_07404_),
    .A2(_07610_),
    .B1(_07503_),
    .B2(_01838_),
    .Y(_07635_));
 OA211x2_ASAP7_75t_R _22768_ (.A1(_07227_),
    .A2(_07564_),
    .B(_07614_),
    .C(_07635_),
    .Y(_07636_));
 AOI21x1_ASAP7_75t_R _22769_ (.A1(_01929_),
    .A2(_07596_),
    .B(_07636_),
    .Y(_02610_));
 OA22x2_ASAP7_75t_R _22770_ (.A1(_07407_),
    .A2(_07610_),
    .B1(_07503_),
    .B2(_01837_),
    .Y(_07637_));
 OA211x2_ASAP7_75t_R _22771_ (.A1(_07249_),
    .A2(_07564_),
    .B(_07614_),
    .C(_07637_),
    .Y(_07638_));
 AOI21x1_ASAP7_75t_R _22772_ (.A1(_01928_),
    .A2(_07596_),
    .B(_07638_),
    .Y(_02611_));
 INVx2_ASAP7_75t_R _22773_ (.A(_00334_),
    .Y(_07639_));
 NOR2x1_ASAP7_75t_R _22774_ (.A(_07639_),
    .B(_06649_),
    .Y(_07640_));
 AO21x1_ASAP7_75t_R _22775_ (.A1(_07639_),
    .A2(_01836_),
    .B(_07640_),
    .Y(_07641_));
 AND2x4_ASAP7_75t_R _22776_ (.A(_07266_),
    .B(_07516_),
    .Y(_07642_));
 NAND2x1_ASAP7_75t_R _22777_ (.A(_06649_),
    .B(_07642_),
    .Y(_07643_));
 OA21x2_ASAP7_75t_R _22778_ (.A1(_07410_),
    .A2(_07529_),
    .B(_07643_),
    .Y(_07644_));
 OA211x2_ASAP7_75t_R _22779_ (.A1(_07266_),
    .A2(_07641_),
    .B(_07644_),
    .C(_07614_),
    .Y(_07645_));
 AOI21x1_ASAP7_75t_R _22780_ (.A1(_01927_),
    .A2(_07596_),
    .B(_07645_),
    .Y(_02612_));
 INVx1_ASAP7_75t_R _22781_ (.A(_06675_),
    .Y(_07646_));
 OA22x2_ASAP7_75t_R _22782_ (.A1(_07413_),
    .A2(_07610_),
    .B1(_07503_),
    .B2(_01835_),
    .Y(_07647_));
 OA211x2_ASAP7_75t_R _22783_ (.A1(_07646_),
    .A2(_07564_),
    .B(_07614_),
    .C(_07647_),
    .Y(_07648_));
 AOI21x1_ASAP7_75t_R _22784_ (.A1(_01926_),
    .A2(_07596_),
    .B(_07648_),
    .Y(_02613_));
 OA22x2_ASAP7_75t_R _22785_ (.A1(_07416_),
    .A2(_07610_),
    .B1(_07503_),
    .B2(_01834_),
    .Y(_07649_));
 OA211x2_ASAP7_75t_R _22786_ (.A1(_07129_),
    .A2(_07564_),
    .B(_07614_),
    .C(_07649_),
    .Y(_07650_));
 AOI21x1_ASAP7_75t_R _22787_ (.A1(_01925_),
    .A2(_07596_),
    .B(_07650_),
    .Y(_02614_));
 NAND2x1_ASAP7_75t_R _22788_ (.A(_05123_),
    .B(_05912_),
    .Y(_07651_));
 NOR2x2_ASAP7_75t_R _22789_ (.A(_05937_),
    .B(_07651_),
    .Y(_07652_));
 BUFx6f_ASAP7_75t_R _22790_ (.A(_07652_),
    .Y(_07653_));
 BUFx6f_ASAP7_75t_R _22791_ (.A(_07652_),
    .Y(_07654_));
 NOR2x1_ASAP7_75t_R _22792_ (.A(_01924_),
    .B(_07654_),
    .Y(_07655_));
 AO21x1_ASAP7_75t_R _22793_ (.A1(_06153_),
    .A2(_07653_),
    .B(_07655_),
    .Y(_02615_));
 NOR2x1_ASAP7_75t_R _22794_ (.A(_01923_),
    .B(_07654_),
    .Y(_07656_));
 AO21x1_ASAP7_75t_R _22795_ (.A1(_06391_),
    .A2(_07653_),
    .B(_07656_),
    .Y(_02616_));
 BUFx12f_ASAP7_75t_R _22796_ (.A(_07652_),
    .Y(_07657_));
 NOR2x1_ASAP7_75t_R _22797_ (.A(_01922_),
    .B(_07657_),
    .Y(_07658_));
 AO21x1_ASAP7_75t_R _22798_ (.A1(_06411_),
    .A2(_07653_),
    .B(_07658_),
    .Y(_02617_));
 NOR2x1_ASAP7_75t_R _22799_ (.A(_01921_),
    .B(_07657_),
    .Y(_07659_));
 AO21x1_ASAP7_75t_R _22800_ (.A1(_06432_),
    .A2(_07653_),
    .B(_07659_),
    .Y(_02618_));
 NOR2x1_ASAP7_75t_R _22801_ (.A(_01920_),
    .B(_07657_),
    .Y(_07660_));
 AO21x1_ASAP7_75t_R _22802_ (.A1(_06454_),
    .A2(_07653_),
    .B(_07660_),
    .Y(_02619_));
 NOR2x1_ASAP7_75t_R _22803_ (.A(_01919_),
    .B(_07657_),
    .Y(_07661_));
 AO21x1_ASAP7_75t_R _22804_ (.A1(_06480_),
    .A2(_07653_),
    .B(_07661_),
    .Y(_02620_));
 NOR2x1_ASAP7_75t_R _22805_ (.A(_01918_),
    .B(_07657_),
    .Y(_07662_));
 AO21x1_ASAP7_75t_R _22806_ (.A1(_06025_),
    .A2(_07653_),
    .B(_07662_),
    .Y(_02621_));
 NOR2x1_ASAP7_75t_R _22807_ (.A(_01917_),
    .B(_07657_),
    .Y(_07663_));
 AO21x1_ASAP7_75t_R _22808_ (.A1(_06650_),
    .A2(_07653_),
    .B(_07663_),
    .Y(_02622_));
 NOR2x1_ASAP7_75t_R _22809_ (.A(_01916_),
    .B(_07657_),
    .Y(_07664_));
 AO21x1_ASAP7_75t_R _22810_ (.A1(_06556_),
    .A2(_07653_),
    .B(_07664_),
    .Y(_02623_));
 NOR2x1_ASAP7_75t_R _22811_ (.A(_01915_),
    .B(_07657_),
    .Y(_07665_));
 AO21x1_ASAP7_75t_R _22812_ (.A1(_06179_),
    .A2(_07653_),
    .B(_07665_),
    .Y(_02624_));
 NOR2x1_ASAP7_75t_R _22813_ (.A(_01914_),
    .B(_07657_),
    .Y(_07666_));
 AO21x1_ASAP7_75t_R _22814_ (.A1(_06197_),
    .A2(_07654_),
    .B(_07666_),
    .Y(_02625_));
 NOR2x1_ASAP7_75t_R _22815_ (.A(_01913_),
    .B(_07657_),
    .Y(_07667_));
 AO21x1_ASAP7_75t_R _22816_ (.A1(_06219_),
    .A2(_07654_),
    .B(_07667_),
    .Y(_02626_));
 NOR2x1_ASAP7_75t_R _22817_ (.A(_01912_),
    .B(_07652_),
    .Y(_07668_));
 AO21x1_ASAP7_75t_R _22818_ (.A1(_06255_),
    .A2(_07654_),
    .B(_07668_),
    .Y(_02627_));
 NOR2x1_ASAP7_75t_R _22819_ (.A(_01911_),
    .B(_07652_),
    .Y(_07669_));
 AO21x1_ASAP7_75t_R _22820_ (.A1(_06277_),
    .A2(_07654_),
    .B(_07669_),
    .Y(_02628_));
 NOR2x1_ASAP7_75t_R _22821_ (.A(_01910_),
    .B(_07652_),
    .Y(_07670_));
 AO21x1_ASAP7_75t_R _22822_ (.A1(_06298_),
    .A2(_07654_),
    .B(_07670_),
    .Y(_02629_));
 NOR2x1_ASAP7_75t_R _22823_ (.A(_01909_),
    .B(_07652_),
    .Y(_07671_));
 AO21x1_ASAP7_75t_R _22824_ (.A1(_06323_),
    .A2(_07654_),
    .B(_07671_),
    .Y(_02630_));
 NOR2x1_ASAP7_75t_R _22825_ (.A(_01908_),
    .B(_07652_),
    .Y(_07672_));
 AO21x1_ASAP7_75t_R _22826_ (.A1(_06343_),
    .A2(_07654_),
    .B(_07672_),
    .Y(_02631_));
 NOR2x1_ASAP7_75t_R _22827_ (.A(_01907_),
    .B(_07652_),
    .Y(_07673_));
 AO21x1_ASAP7_75t_R _22828_ (.A1(_06366_),
    .A2(_07654_),
    .B(_07673_),
    .Y(_02632_));
 NAND3x2_ASAP7_75t_R _22829_ (.B(_05897_),
    .C(_05777_),
    .Y(_07674_),
    .A(_05867_));
 BUFx6f_ASAP7_75t_R _22830_ (.A(_07674_),
    .Y(_07675_));
 BUFx6f_ASAP7_75t_R _22831_ (.A(_07674_),
    .Y(_07676_));
 NAND2x1_ASAP7_75t_R _22832_ (.A(_01906_),
    .B(_07676_),
    .Y(_07677_));
 OA21x2_ASAP7_75t_R _22833_ (.A1(_05811_),
    .A2(_07675_),
    .B(_07677_),
    .Y(_02633_));
 NAND2x1_ASAP7_75t_R _22834_ (.A(_01905_),
    .B(_07676_),
    .Y(_07678_));
 OA21x2_ASAP7_75t_R _22835_ (.A1(_05981_),
    .A2(_07675_),
    .B(_07678_),
    .Y(_02634_));
 NAND2x1_ASAP7_75t_R _22836_ (.A(_01904_),
    .B(_07676_),
    .Y(_07679_));
 OA21x2_ASAP7_75t_R _22837_ (.A1(_06025_),
    .A2(_07675_),
    .B(_07679_),
    .Y(_02635_));
 NAND2x1_ASAP7_75t_R _22838_ (.A(_01903_),
    .B(_07676_),
    .Y(_07680_));
 OA21x2_ASAP7_75t_R _22839_ (.A1(_06052_),
    .A2(_07675_),
    .B(_07680_),
    .Y(_02636_));
 NAND2x1_ASAP7_75t_R _22840_ (.A(_01902_),
    .B(_07676_),
    .Y(_07681_));
 OA21x2_ASAP7_75t_R _22841_ (.A1(_06082_),
    .A2(_07675_),
    .B(_07681_),
    .Y(_02637_));
 NAND2x1_ASAP7_75t_R _22842_ (.A(_01901_),
    .B(_07676_),
    .Y(_07682_));
 OA21x2_ASAP7_75t_R _22843_ (.A1(_06108_),
    .A2(_07675_),
    .B(_07682_),
    .Y(_02638_));
 NAND2x1_ASAP7_75t_R _22844_ (.A(_01900_),
    .B(_07676_),
    .Y(_07683_));
 OA21x2_ASAP7_75t_R _22845_ (.A1(_06131_),
    .A2(_07675_),
    .B(_07683_),
    .Y(_02639_));
 NAND2x1_ASAP7_75t_R _22846_ (.A(_01899_),
    .B(_07676_),
    .Y(_07684_));
 OA21x2_ASAP7_75t_R _22847_ (.A1(_06153_),
    .A2(_07675_),
    .B(_07684_),
    .Y(_02640_));
 BUFx12f_ASAP7_75t_R _22848_ (.A(_07674_),
    .Y(_07685_));
 NAND2x1_ASAP7_75t_R _22849_ (.A(_01898_),
    .B(_07685_),
    .Y(_07686_));
 OA21x2_ASAP7_75t_R _22850_ (.A1(_06179_),
    .A2(_07675_),
    .B(_07686_),
    .Y(_02641_));
 NAND2x1_ASAP7_75t_R _22851_ (.A(_01897_),
    .B(_07685_),
    .Y(_07687_));
 OA21x2_ASAP7_75t_R _22852_ (.A1(_06197_),
    .A2(_07675_),
    .B(_07687_),
    .Y(_02642_));
 BUFx6f_ASAP7_75t_R _22853_ (.A(_07674_),
    .Y(_07688_));
 NAND2x1_ASAP7_75t_R _22854_ (.A(_01896_),
    .B(_07685_),
    .Y(_07689_));
 OA21x2_ASAP7_75t_R _22855_ (.A1(_06219_),
    .A2(_07688_),
    .B(_07689_),
    .Y(_02643_));
 NAND2x1_ASAP7_75t_R _22856_ (.A(_01895_),
    .B(_07685_),
    .Y(_07690_));
 OA21x2_ASAP7_75t_R _22857_ (.A1(_06235_),
    .A2(_07688_),
    .B(_07690_),
    .Y(_02644_));
 NAND2x1_ASAP7_75t_R _22858_ (.A(_01894_),
    .B(_07685_),
    .Y(_07691_));
 OA21x2_ASAP7_75t_R _22859_ (.A1(_06255_),
    .A2(_07688_),
    .B(_07691_),
    .Y(_02645_));
 NAND2x1_ASAP7_75t_R _22860_ (.A(_01893_),
    .B(_07685_),
    .Y(_07692_));
 OA21x2_ASAP7_75t_R _22861_ (.A1(_06277_),
    .A2(_07688_),
    .B(_07692_),
    .Y(_02646_));
 NAND2x1_ASAP7_75t_R _22862_ (.A(_01892_),
    .B(_07685_),
    .Y(_07693_));
 OA21x2_ASAP7_75t_R _22863_ (.A1(_06298_),
    .A2(_07688_),
    .B(_07693_),
    .Y(_02647_));
 NAND2x1_ASAP7_75t_R _22864_ (.A(_01891_),
    .B(_07685_),
    .Y(_07694_));
 OA21x2_ASAP7_75t_R _22865_ (.A1(_06323_),
    .A2(_07688_),
    .B(_07694_),
    .Y(_02648_));
 NAND2x1_ASAP7_75t_R _22866_ (.A(_01890_),
    .B(_07685_),
    .Y(_07695_));
 OA21x2_ASAP7_75t_R _22867_ (.A1(_06343_),
    .A2(_07688_),
    .B(_07695_),
    .Y(_02649_));
 NAND2x1_ASAP7_75t_R _22868_ (.A(_01889_),
    .B(_07685_),
    .Y(_07696_));
 OA21x2_ASAP7_75t_R _22869_ (.A1(_06366_),
    .A2(_07688_),
    .B(_07696_),
    .Y(_02650_));
 BUFx12f_ASAP7_75t_R _22870_ (.A(_07674_),
    .Y(_07697_));
 NAND2x1_ASAP7_75t_R _22871_ (.A(_01888_),
    .B(_07697_),
    .Y(_07698_));
 OA21x2_ASAP7_75t_R _22872_ (.A1(_06391_),
    .A2(_07688_),
    .B(_07698_),
    .Y(_02651_));
 NAND2x1_ASAP7_75t_R _22873_ (.A(_01887_),
    .B(_07697_),
    .Y(_07699_));
 OA21x2_ASAP7_75t_R _22874_ (.A1(_06411_),
    .A2(_07688_),
    .B(_07699_),
    .Y(_02652_));
 BUFx6f_ASAP7_75t_R _22875_ (.A(_07674_),
    .Y(_07700_));
 NAND2x1_ASAP7_75t_R _22876_ (.A(_01886_),
    .B(_07697_),
    .Y(_07701_));
 OA21x2_ASAP7_75t_R _22877_ (.A1(_06432_),
    .A2(_07700_),
    .B(_07701_),
    .Y(_02653_));
 NAND2x1_ASAP7_75t_R _22878_ (.A(_01885_),
    .B(_07697_),
    .Y(_07702_));
 OA21x2_ASAP7_75t_R _22879_ (.A1(_06454_),
    .A2(_07700_),
    .B(_07702_),
    .Y(_02654_));
 NAND2x1_ASAP7_75t_R _22880_ (.A(_01884_),
    .B(_07697_),
    .Y(_07703_));
 OA21x2_ASAP7_75t_R _22881_ (.A1(_05851_),
    .A2(_07700_),
    .B(_07703_),
    .Y(_02655_));
 NAND2x1_ASAP7_75t_R _22882_ (.A(_01883_),
    .B(_07697_),
    .Y(_07704_));
 OA21x2_ASAP7_75t_R _22883_ (.A1(_06480_),
    .A2(_07700_),
    .B(_07704_),
    .Y(_02656_));
 NAND2x1_ASAP7_75t_R _22884_ (.A(_01882_),
    .B(_07697_),
    .Y(_07705_));
 OA21x2_ASAP7_75t_R _22885_ (.A1(_06504_),
    .A2(_07700_),
    .B(_07705_),
    .Y(_02657_));
 NAND2x1_ASAP7_75t_R _22886_ (.A(_01881_),
    .B(_07697_),
    .Y(_07706_));
 OA21x2_ASAP7_75t_R _22887_ (.A1(_06556_),
    .A2(_07700_),
    .B(_07706_),
    .Y(_02658_));
 NAND2x1_ASAP7_75t_R _22888_ (.A(_01880_),
    .B(_07697_),
    .Y(_07707_));
 OA21x2_ASAP7_75t_R _22889_ (.A1(_06580_),
    .A2(_07700_),
    .B(_07707_),
    .Y(_02659_));
 NAND2x1_ASAP7_75t_R _22890_ (.A(_01879_),
    .B(_07697_),
    .Y(_07708_));
 OA21x2_ASAP7_75t_R _22891_ (.A1(_06600_),
    .A2(_07700_),
    .B(_07708_),
    .Y(_02660_));
 NAND2x1_ASAP7_75t_R _22892_ (.A(_01878_),
    .B(_07674_),
    .Y(_07709_));
 OA21x2_ASAP7_75t_R _22893_ (.A1(_06624_),
    .A2(_07700_),
    .B(_07709_),
    .Y(_02661_));
 NAND2x1_ASAP7_75t_R _22894_ (.A(_01877_),
    .B(_07674_),
    .Y(_07710_));
 OA21x2_ASAP7_75t_R _22895_ (.A1(_06650_),
    .A2(_07700_),
    .B(_07710_),
    .Y(_02662_));
 NAND2x1_ASAP7_75t_R _22896_ (.A(_01876_),
    .B(_07674_),
    .Y(_07711_));
 OA21x2_ASAP7_75t_R _22897_ (.A1(_06675_),
    .A2(_07676_),
    .B(_07711_),
    .Y(_02663_));
 NAND2x1_ASAP7_75t_R _22898_ (.A(_01875_),
    .B(_07674_),
    .Y(_07712_));
 OA21x2_ASAP7_75t_R _22899_ (.A1(_06699_),
    .A2(_07676_),
    .B(_07712_),
    .Y(_02664_));
 BUFx12f_ASAP7_75t_R _22900_ (.A(_07529_),
    .Y(_07713_));
 BUFx12f_ASAP7_75t_R _22901_ (.A(_07713_),
    .Y(_07714_));
 BUFx6f_ASAP7_75t_R _22902_ (.A(_07539_),
    .Y(_07715_));
 AND2x2_ASAP7_75t_R _22903_ (.A(_01962_),
    .B(_07715_),
    .Y(_07716_));
 AOI21x1_ASAP7_75t_R _22904_ (.A1(_01874_),
    .A2(_07714_),
    .B(_07716_),
    .Y(_02665_));
 AND2x2_ASAP7_75t_R _22905_ (.A(_01961_),
    .B(_07715_),
    .Y(_07717_));
 AOI21x1_ASAP7_75t_R _22906_ (.A1(_01873_),
    .A2(_07714_),
    .B(_07717_),
    .Y(_02666_));
 AND2x2_ASAP7_75t_R _22907_ (.A(_01960_),
    .B(_07715_),
    .Y(_07718_));
 AOI21x1_ASAP7_75t_R _22908_ (.A1(_01872_),
    .A2(_07714_),
    .B(_07718_),
    .Y(_02667_));
 NAND2x1_ASAP7_75t_R _22909_ (.A(_01871_),
    .B(_07713_),
    .Y(_07719_));
 OA21x2_ASAP7_75t_R _22910_ (.A1(_07544_),
    .A2(_07713_),
    .B(_07719_),
    .Y(_02668_));
 AND2x2_ASAP7_75t_R _22911_ (.A(_01958_),
    .B(_07715_),
    .Y(_07720_));
 AOI21x1_ASAP7_75t_R _22912_ (.A1(_01870_),
    .A2(_07714_),
    .B(_07720_),
    .Y(_02669_));
 AND2x2_ASAP7_75t_R _22913_ (.A(_01957_),
    .B(_07715_),
    .Y(_07721_));
 AOI21x1_ASAP7_75t_R _22914_ (.A1(_01869_),
    .A2(_07714_),
    .B(_07721_),
    .Y(_02670_));
 AND2x2_ASAP7_75t_R _22915_ (.A(_00331_),
    .B(_07715_),
    .Y(_07722_));
 AOI21x1_ASAP7_75t_R _22916_ (.A1(_01868_),
    .A2(_07714_),
    .B(_07722_),
    .Y(_02671_));
 AND2x2_ASAP7_75t_R _22917_ (.A(_00332_),
    .B(_07715_),
    .Y(_07723_));
 AOI21x1_ASAP7_75t_R _22918_ (.A1(_01867_),
    .A2(_07714_),
    .B(_07723_),
    .Y(_02672_));
 AND2x2_ASAP7_75t_R _22919_ (.A(_00333_),
    .B(_07715_),
    .Y(_07724_));
 AOI21x1_ASAP7_75t_R _22920_ (.A1(_01866_),
    .A2(_07714_),
    .B(_07724_),
    .Y(_02673_));
 AND2x2_ASAP7_75t_R _22921_ (.A(_01956_),
    .B(_07715_),
    .Y(_07725_));
 AOI21x1_ASAP7_75t_R _22922_ (.A1(_01865_),
    .A2(_07714_),
    .B(_07725_),
    .Y(_02674_));
 BUFx6f_ASAP7_75t_R _22923_ (.A(_07540_),
    .Y(_07726_));
 AND2x2_ASAP7_75t_R _22924_ (.A(_01955_),
    .B(_07726_),
    .Y(_07727_));
 AOI21x1_ASAP7_75t_R _22925_ (.A1(_01864_),
    .A2(_07714_),
    .B(_07727_),
    .Y(_02675_));
 BUFx12f_ASAP7_75t_R _22926_ (.A(_07713_),
    .Y(_07728_));
 AND2x2_ASAP7_75t_R _22927_ (.A(_01954_),
    .B(_07726_),
    .Y(_07729_));
 AOI21x1_ASAP7_75t_R _22928_ (.A1(_01863_),
    .A2(_07728_),
    .B(_07729_),
    .Y(_02676_));
 AND2x2_ASAP7_75t_R _22929_ (.A(_01953_),
    .B(_07726_),
    .Y(_07730_));
 AOI21x1_ASAP7_75t_R _22930_ (.A1(_01862_),
    .A2(_07728_),
    .B(_07730_),
    .Y(_02677_));
 AND2x2_ASAP7_75t_R _22931_ (.A(_01952_),
    .B(_07726_),
    .Y(_07731_));
 AOI21x1_ASAP7_75t_R _22932_ (.A1(_01861_),
    .A2(_07728_),
    .B(_07731_),
    .Y(_02678_));
 AND2x2_ASAP7_75t_R _22933_ (.A(_01951_),
    .B(_07726_),
    .Y(_07732_));
 AOI21x1_ASAP7_75t_R _22934_ (.A1(_01860_),
    .A2(_07728_),
    .B(_07732_),
    .Y(_02679_));
 AND2x2_ASAP7_75t_R _22935_ (.A(_01950_),
    .B(_07726_),
    .Y(_07733_));
 AOI21x1_ASAP7_75t_R _22936_ (.A1(_01859_),
    .A2(_07728_),
    .B(_07733_),
    .Y(_02680_));
 AND2x2_ASAP7_75t_R _22937_ (.A(_01949_),
    .B(_07726_),
    .Y(_07734_));
 AOI21x1_ASAP7_75t_R _22938_ (.A1(_01858_),
    .A2(_07728_),
    .B(_07734_),
    .Y(_02681_));
 AND2x2_ASAP7_75t_R _22939_ (.A(_01948_),
    .B(_07726_),
    .Y(_07735_));
 AOI21x1_ASAP7_75t_R _22940_ (.A1(_01857_),
    .A2(_07728_),
    .B(_07735_),
    .Y(_02682_));
 AND2x2_ASAP7_75t_R _22941_ (.A(_01947_),
    .B(_07726_),
    .Y(_07736_));
 AOI21x1_ASAP7_75t_R _22942_ (.A1(_01856_),
    .A2(_07728_),
    .B(_07736_),
    .Y(_02683_));
 AND2x2_ASAP7_75t_R _22943_ (.A(_01946_),
    .B(_07726_),
    .Y(_07737_));
 AOI21x1_ASAP7_75t_R _22944_ (.A1(_01855_),
    .A2(_07728_),
    .B(_07737_),
    .Y(_02684_));
 BUFx6f_ASAP7_75t_R _22945_ (.A(_07540_),
    .Y(_07738_));
 AND2x2_ASAP7_75t_R _22946_ (.A(_01945_),
    .B(_07738_),
    .Y(_07739_));
 AOI21x1_ASAP7_75t_R _22947_ (.A1(_01854_),
    .A2(_07728_),
    .B(_07739_),
    .Y(_02685_));
 BUFx12f_ASAP7_75t_R _22948_ (.A(_07713_),
    .Y(_07740_));
 AND2x2_ASAP7_75t_R _22949_ (.A(_01944_),
    .B(_07738_),
    .Y(_07741_));
 AOI21x1_ASAP7_75t_R _22950_ (.A1(_01853_),
    .A2(_07740_),
    .B(_07741_),
    .Y(_02686_));
 AND2x2_ASAP7_75t_R _22951_ (.A(_01943_),
    .B(_07738_),
    .Y(_07742_));
 AOI21x1_ASAP7_75t_R _22952_ (.A1(_01852_),
    .A2(_07740_),
    .B(_07742_),
    .Y(_02687_));
 AND2x2_ASAP7_75t_R _22953_ (.A(_01942_),
    .B(_07738_),
    .Y(_07743_));
 AOI21x1_ASAP7_75t_R _22954_ (.A1(_01851_),
    .A2(_07740_),
    .B(_07743_),
    .Y(_02688_));
 AND2x2_ASAP7_75t_R _22955_ (.A(_01941_),
    .B(_07738_),
    .Y(_07744_));
 AOI21x1_ASAP7_75t_R _22956_ (.A1(_01850_),
    .A2(_07740_),
    .B(_07744_),
    .Y(_02689_));
 AND2x2_ASAP7_75t_R _22957_ (.A(_01940_),
    .B(_07738_),
    .Y(_07745_));
 AOI21x1_ASAP7_75t_R _22958_ (.A1(_01849_),
    .A2(_07740_),
    .B(_07745_),
    .Y(_02690_));
 AND2x2_ASAP7_75t_R _22959_ (.A(_01939_),
    .B(_07738_),
    .Y(_07746_));
 AOI21x1_ASAP7_75t_R _22960_ (.A1(_01848_),
    .A2(_07740_),
    .B(_07746_),
    .Y(_02691_));
 AND2x2_ASAP7_75t_R _22961_ (.A(_01938_),
    .B(_07738_),
    .Y(_07747_));
 AOI21x1_ASAP7_75t_R _22962_ (.A1(_01847_),
    .A2(_07740_),
    .B(_07747_),
    .Y(_02692_));
 AND2x2_ASAP7_75t_R _22963_ (.A(_01937_),
    .B(_07738_),
    .Y(_07748_));
 AOI21x1_ASAP7_75t_R _22964_ (.A1(_01846_),
    .A2(_07740_),
    .B(_07748_),
    .Y(_02693_));
 AND2x2_ASAP7_75t_R _22965_ (.A(_01936_),
    .B(_07738_),
    .Y(_07749_));
 AOI21x1_ASAP7_75t_R _22966_ (.A1(_01845_),
    .A2(_07740_),
    .B(_07749_),
    .Y(_02694_));
 BUFx6f_ASAP7_75t_R _22967_ (.A(_07540_),
    .Y(_07750_));
 AND2x2_ASAP7_75t_R _22968_ (.A(_01935_),
    .B(_07750_),
    .Y(_07751_));
 AOI21x1_ASAP7_75t_R _22969_ (.A1(_01844_),
    .A2(_07740_),
    .B(_07751_),
    .Y(_02695_));
 BUFx12f_ASAP7_75t_R _22970_ (.A(_07713_),
    .Y(_07752_));
 AND2x2_ASAP7_75t_R _22971_ (.A(_01934_),
    .B(_07750_),
    .Y(_07753_));
 AOI21x1_ASAP7_75t_R _22972_ (.A1(_01843_),
    .A2(_07752_),
    .B(_07753_),
    .Y(_02696_));
 AND2x2_ASAP7_75t_R _22973_ (.A(_01933_),
    .B(_07750_),
    .Y(_07754_));
 AOI21x1_ASAP7_75t_R _22974_ (.A1(_01842_),
    .A2(_07752_),
    .B(_07754_),
    .Y(_02697_));
 AND2x2_ASAP7_75t_R _22975_ (.A(_01932_),
    .B(_07750_),
    .Y(_07755_));
 AOI21x1_ASAP7_75t_R _22976_ (.A1(_01841_),
    .A2(_07752_),
    .B(_07755_),
    .Y(_02698_));
 AND2x2_ASAP7_75t_R _22977_ (.A(_01931_),
    .B(_07750_),
    .Y(_07756_));
 AOI21x1_ASAP7_75t_R _22978_ (.A1(_01840_),
    .A2(_07752_),
    .B(_07756_),
    .Y(_02699_));
 AND2x2_ASAP7_75t_R _22979_ (.A(_01930_),
    .B(_07750_),
    .Y(_07757_));
 AOI21x1_ASAP7_75t_R _22980_ (.A1(_01839_),
    .A2(_07752_),
    .B(_07757_),
    .Y(_02700_));
 AND2x2_ASAP7_75t_R _22981_ (.A(_01929_),
    .B(_07750_),
    .Y(_07758_));
 AOI21x1_ASAP7_75t_R _22982_ (.A1(_01838_),
    .A2(_07752_),
    .B(_07758_),
    .Y(_02701_));
 AND2x2_ASAP7_75t_R _22983_ (.A(_01928_),
    .B(_07750_),
    .Y(_07759_));
 AOI21x1_ASAP7_75t_R _22984_ (.A1(_01837_),
    .A2(_07752_),
    .B(_07759_),
    .Y(_02702_));
 AND2x2_ASAP7_75t_R _22985_ (.A(_01927_),
    .B(_07750_),
    .Y(_07760_));
 AOI21x1_ASAP7_75t_R _22986_ (.A1(_01836_),
    .A2(_07752_),
    .B(_07760_),
    .Y(_02703_));
 AND2x2_ASAP7_75t_R _22987_ (.A(_01926_),
    .B(_07750_),
    .Y(_07761_));
 AOI21x1_ASAP7_75t_R _22988_ (.A1(_01835_),
    .A2(_07752_),
    .B(_07761_),
    .Y(_02704_));
 BUFx6f_ASAP7_75t_R _22989_ (.A(_07539_),
    .Y(_07762_));
 AND2x2_ASAP7_75t_R _22990_ (.A(_01925_),
    .B(_07762_),
    .Y(_07763_));
 AOI21x1_ASAP7_75t_R _22991_ (.A1(_01834_),
    .A2(_07752_),
    .B(_07763_),
    .Y(_02705_));
 NAND2x1_ASAP7_75t_R _22992_ (.A(_05912_),
    .B(_05777_),
    .Y(_07764_));
 OR2x6_ASAP7_75t_R _22993_ (.A(_05937_),
    .B(_07764_),
    .Y(_07765_));
 INVx2_ASAP7_75t_R _22994_ (.A(_07765_),
    .Y(_07766_));
 NAND2x1_ASAP7_75t_R _22995_ (.A(_06277_),
    .B(_07766_),
    .Y(_07767_));
 OAI21x1_ASAP7_75t_R _22996_ (.A1(_01833_),
    .A2(_07766_),
    .B(_07767_),
    .Y(_02706_));
 NAND2x1_ASAP7_75t_R _22997_ (.A(_06179_),
    .B(_07766_),
    .Y(_07768_));
 OAI21x1_ASAP7_75t_R _22998_ (.A1(_01832_),
    .A2(_07766_),
    .B(_07768_),
    .Y(_02707_));
 INVx1_ASAP7_75t_R _22999_ (.A(_01831_),
    .Y(_07769_));
 OAI21x1_ASAP7_75t_R _23000_ (.A1(_05749_),
    .A2(_06004_),
    .B(_07516_),
    .Y(_07770_));
 BUFx6f_ASAP7_75t_R _23001_ (.A(_07770_),
    .Y(_07771_));
 OR2x6_ASAP7_75t_R _23002_ (.A(_01391_),
    .B(_07524_),
    .Y(_07772_));
 BUFx6f_ASAP7_75t_R _23003_ (.A(_07772_),
    .Y(_07773_));
 BUFx6f_ASAP7_75t_R _23004_ (.A(_13534_),
    .Y(_07774_));
 BUFx3_ASAP7_75t_R _23005_ (.A(_13533_),
    .Y(_07775_));
 AND2x2_ASAP7_75t_R _23006_ (.A(_07775_),
    .B(_13238_),
    .Y(_07776_));
 AO21x1_ASAP7_75t_R _23007_ (.A1(_07774_),
    .A2(_01537_),
    .B(_07776_),
    .Y(_07777_));
 OAI22x1_ASAP7_75t_R _23008_ (.A1(_01477_),
    .A2(_07536_),
    .B1(_07773_),
    .B2(_07777_),
    .Y(_07778_));
 AO21x2_ASAP7_75t_R _23009_ (.A1(_07505_),
    .A2(_07512_),
    .B(_05509_),
    .Y(_07779_));
 OR2x2_ASAP7_75t_R _23010_ (.A(_07497_),
    .B(_07779_),
    .Y(_07780_));
 BUFx6f_ASAP7_75t_R _23011_ (.A(_07780_),
    .Y(_07781_));
 INVx1_ASAP7_75t_R _23012_ (.A(_07781_),
    .Y(_07782_));
 INVx3_ASAP7_75t_R _23013_ (.A(_07770_),
    .Y(_07783_));
 AO221x1_ASAP7_75t_R _23014_ (.A1(_05811_),
    .A2(_07517_),
    .B1(_07778_),
    .B2(_07782_),
    .C(_07783_),
    .Y(_07784_));
 OA21x2_ASAP7_75t_R _23015_ (.A1(_07769_),
    .A2(_07771_),
    .B(_07784_),
    .Y(_02712_));
 BUFx12f_ASAP7_75t_R _23016_ (.A(_07783_),
    .Y(_07785_));
 BUFx12f_ASAP7_75t_R _23017_ (.A(_07785_),
    .Y(_07786_));
 BUFx6f_ASAP7_75t_R _23018_ (.A(_07779_),
    .Y(_07787_));
 AND2x2_ASAP7_75t_R _23019_ (.A(_07775_),
    .B(_13685_),
    .Y(_07788_));
 AO21x1_ASAP7_75t_R _23020_ (.A1(_07774_),
    .A2(_01536_),
    .B(_07788_),
    .Y(_07789_));
 BUFx6f_ASAP7_75t_R _23021_ (.A(_01538_),
    .Y(_07790_));
 OR4x1_ASAP7_75t_R _23022_ (.A(_00016_),
    .B(_07790_),
    .C(_14773_),
    .D(_01496_),
    .Y(_07791_));
 OR4x1_ASAP7_75t_R _23023_ (.A(_01480_),
    .B(_14966_),
    .C(_14900_),
    .D(_14837_),
    .Y(_07792_));
 OR4x1_ASAP7_75t_R _23024_ (.A(_15158_),
    .B(_15099_),
    .C(_07791_),
    .D(_07792_),
    .Y(_07793_));
 XNOR2x2_ASAP7_75t_R _23025_ (.A(_00019_),
    .B(_07793_),
    .Y(_07794_));
 BUFx6f_ASAP7_75t_R _23026_ (.A(_05400_),
    .Y(_07795_));
 OA222x2_ASAP7_75t_R _23027_ (.A1(_01476_),
    .A2(_07536_),
    .B1(_07773_),
    .B2(_07789_),
    .C1(_07794_),
    .C2(_07795_),
    .Y(_07796_));
 OR3x1_ASAP7_75t_R _23028_ (.A(_07529_),
    .B(_07787_),
    .C(_07796_),
    .Y(_07797_));
 OA211x2_ASAP7_75t_R _23029_ (.A1(_06923_),
    .A2(_07762_),
    .B(_07771_),
    .C(_07797_),
    .Y(_07798_));
 AOI21x1_ASAP7_75t_R _23030_ (.A1(_01830_),
    .A2(_07786_),
    .B(_07798_),
    .Y(_02713_));
 BUFx12f_ASAP7_75t_R _23031_ (.A(_00339_),
    .Y(_07799_));
 AND2x2_ASAP7_75t_R _23032_ (.A(_07775_),
    .B(_07799_),
    .Y(_07800_));
 AO21x1_ASAP7_75t_R _23033_ (.A1(_07774_),
    .A2(_01535_),
    .B(_07800_),
    .Y(_07801_));
 OR3x2_ASAP7_75t_R _23034_ (.A(_07790_),
    .B(_14773_),
    .C(_02236_),
    .Y(_07802_));
 BUFx6f_ASAP7_75t_R _23035_ (.A(_07802_),
    .Y(_07803_));
 OR4x1_ASAP7_75t_R _23036_ (.A(_00019_),
    .B(_15158_),
    .C(_15099_),
    .D(_07792_),
    .Y(_07804_));
 OR2x2_ASAP7_75t_R _23037_ (.A(_07803_),
    .B(_07804_),
    .Y(_07805_));
 XNOR2x2_ASAP7_75t_R _23038_ (.A(_14379_),
    .B(_07805_),
    .Y(_07806_));
 OA222x2_ASAP7_75t_R _23039_ (.A1(_01475_),
    .A2(_07536_),
    .B1(_07773_),
    .B2(_07801_),
    .C1(_07806_),
    .C2(_07795_),
    .Y(_07807_));
 OR3x1_ASAP7_75t_R _23040_ (.A(_07529_),
    .B(_07787_),
    .C(_07807_),
    .Y(_07808_));
 OA211x2_ASAP7_75t_R _23041_ (.A1(_06937_),
    .A2(_07762_),
    .B(_07771_),
    .C(_07808_),
    .Y(_07809_));
 AOI21x1_ASAP7_75t_R _23042_ (.A1(_01829_),
    .A2(_07786_),
    .B(_07809_),
    .Y(_02714_));
 BUFx6f_ASAP7_75t_R _23043_ (.A(_07512_),
    .Y(_07810_));
 AND2x2_ASAP7_75t_R _23044_ (.A(_07775_),
    .B(_14272_),
    .Y(_07811_));
 AO21x1_ASAP7_75t_R _23045_ (.A1(_07774_),
    .A2(_01534_),
    .B(_07811_),
    .Y(_07812_));
 BUFx6f_ASAP7_75t_R _23046_ (.A(_07791_),
    .Y(_07813_));
 OR3x1_ASAP7_75t_R _23047_ (.A(_14379_),
    .B(_07813_),
    .C(_07804_),
    .Y(_07814_));
 XNOR2x2_ASAP7_75t_R _23048_ (.A(_01503_),
    .B(_07814_),
    .Y(_07815_));
 OA222x2_ASAP7_75t_R _23049_ (.A1(_01474_),
    .A2(_07810_),
    .B1(_07773_),
    .B2(_07812_),
    .C1(_07815_),
    .C2(_07795_),
    .Y(_07816_));
 OR3x1_ASAP7_75t_R _23050_ (.A(_07529_),
    .B(_07787_),
    .C(_07816_),
    .Y(_07817_));
 OA211x2_ASAP7_75t_R _23051_ (.A1(_07571_),
    .A2(_07762_),
    .B(_07771_),
    .C(_07817_),
    .Y(_07818_));
 AOI21x1_ASAP7_75t_R _23052_ (.A1(_01828_),
    .A2(_07786_),
    .B(_07818_),
    .Y(_02715_));
 AND2x2_ASAP7_75t_R _23053_ (.A(_14112_),
    .B(_13533_),
    .Y(_07819_));
 AO21x1_ASAP7_75t_R _23054_ (.A1(_07774_),
    .A2(_01533_),
    .B(_07819_),
    .Y(_07820_));
 OR4x1_ASAP7_75t_R _23055_ (.A(_01503_),
    .B(_14379_),
    .C(_07803_),
    .D(_07804_),
    .Y(_07821_));
 XNOR2x2_ASAP7_75t_R _23056_ (.A(_01502_),
    .B(_07821_),
    .Y(_07822_));
 OA222x2_ASAP7_75t_R _23057_ (.A1(_01473_),
    .A2(_07810_),
    .B1(_07773_),
    .B2(_07820_),
    .C1(_07822_),
    .C2(_07795_),
    .Y(_07823_));
 OR3x1_ASAP7_75t_R _23058_ (.A(_07529_),
    .B(_07787_),
    .C(_07823_),
    .Y(_07824_));
 OA211x2_ASAP7_75t_R _23059_ (.A1(_06961_),
    .A2(_07762_),
    .B(_07771_),
    .C(_07824_),
    .Y(_07825_));
 AOI21x1_ASAP7_75t_R _23060_ (.A1(_01827_),
    .A2(_07786_),
    .B(_07825_),
    .Y(_02716_));
 AND2x2_ASAP7_75t_R _23061_ (.A(_14533_),
    .B(_13533_),
    .Y(_07826_));
 AO21x1_ASAP7_75t_R _23062_ (.A1(_13534_),
    .A2(_01532_),
    .B(_07826_),
    .Y(_07827_));
 OR5x1_ASAP7_75t_R _23063_ (.A(_01502_),
    .B(_01503_),
    .C(_14379_),
    .D(_07791_),
    .E(_07804_),
    .Y(_07828_));
 XNOR2x2_ASAP7_75t_R _23064_ (.A(_01501_),
    .B(_07828_),
    .Y(_07829_));
 OA222x2_ASAP7_75t_R _23065_ (.A1(_01472_),
    .A2(_07810_),
    .B1(_07773_),
    .B2(_07827_),
    .C1(_07829_),
    .C2(_07795_),
    .Y(_07830_));
 OR3x1_ASAP7_75t_R _23066_ (.A(_07529_),
    .B(_07787_),
    .C(_07830_),
    .Y(_07831_));
 OA211x2_ASAP7_75t_R _23067_ (.A1(_07576_),
    .A2(_07762_),
    .B(_07771_),
    .C(_07831_),
    .Y(_07832_));
 AOI21x1_ASAP7_75t_R _23068_ (.A1(_01826_),
    .A2(_07786_),
    .B(_07832_),
    .Y(_02717_));
 BUFx3_ASAP7_75t_R _23069_ (.A(_07770_),
    .Y(_07833_));
 BUFx6f_ASAP7_75t_R _23070_ (.A(_07516_),
    .Y(_07834_));
 AND2x2_ASAP7_75t_R _23071_ (.A(_14289_),
    .B(_13533_),
    .Y(_07835_));
 AO21x1_ASAP7_75t_R _23072_ (.A1(_13534_),
    .A2(_01531_),
    .B(_07835_),
    .Y(_07836_));
 OR5x2_ASAP7_75t_R _23073_ (.A(_01501_),
    .B(_01502_),
    .C(_01503_),
    .D(_14379_),
    .E(_07804_),
    .Y(_07837_));
 OR2x6_ASAP7_75t_R _23074_ (.A(_07802_),
    .B(_07837_),
    .Y(_07838_));
 XNOR2x2_ASAP7_75t_R _23075_ (.A(_15708_),
    .B(_07838_),
    .Y(_07839_));
 OA222x2_ASAP7_75t_R _23076_ (.A1(_01471_),
    .A2(_07810_),
    .B1(_07772_),
    .B2(_07836_),
    .C1(_07839_),
    .C2(_07513_),
    .Y(_07840_));
 OR3x1_ASAP7_75t_R _23077_ (.A(_07834_),
    .B(_07787_),
    .C(_07840_),
    .Y(_07841_));
 OA211x2_ASAP7_75t_R _23078_ (.A1(_06968_),
    .A2(_07762_),
    .B(_07833_),
    .C(_07841_),
    .Y(_07842_));
 AOI21x1_ASAP7_75t_R _23079_ (.A1(_01825_),
    .A2(_07786_),
    .B(_07842_),
    .Y(_02718_));
 OR3x1_ASAP7_75t_R _23080_ (.A(_15708_),
    .B(_07813_),
    .C(_07837_),
    .Y(_07843_));
 XNOR2x2_ASAP7_75t_R _23081_ (.A(_15832_),
    .B(_07843_),
    .Y(_07844_));
 BUFx6f_ASAP7_75t_R _23082_ (.A(_05400_),
    .Y(_07845_));
 OR3x2_ASAP7_75t_R _23083_ (.A(_13534_),
    .B(_01391_),
    .C(_07524_),
    .Y(_07846_));
 BUFx6f_ASAP7_75t_R _23084_ (.A(_07846_),
    .Y(_07847_));
 OA222x2_ASAP7_75t_R _23085_ (.A1(_01470_),
    .A2(_07810_),
    .B1(_07844_),
    .B2(_07845_),
    .C1(_07847_),
    .C2(_14278_),
    .Y(_07848_));
 OR3x1_ASAP7_75t_R _23086_ (.A(_07834_),
    .B(_07787_),
    .C(_07848_),
    .Y(_07849_));
 OA211x2_ASAP7_75t_R _23087_ (.A1(_06973_),
    .A2(_07762_),
    .B(_07833_),
    .C(_07849_),
    .Y(_07850_));
 AOI21x1_ASAP7_75t_R _23088_ (.A1(_01824_),
    .A2(_07786_),
    .B(_07850_),
    .Y(_02719_));
 OR3x1_ASAP7_75t_R _23089_ (.A(_15832_),
    .B(_15708_),
    .C(_07838_),
    .Y(_07851_));
 XNOR2x2_ASAP7_75t_R _23090_ (.A(_01498_),
    .B(_07851_),
    .Y(_07852_));
 OA222x2_ASAP7_75t_R _23091_ (.A1(_01469_),
    .A2(_07810_),
    .B1(_07852_),
    .B2(_07845_),
    .C1(_07847_),
    .C2(_14778_),
    .Y(_07853_));
 OR3x1_ASAP7_75t_R _23092_ (.A(_07834_),
    .B(_07787_),
    .C(_07853_),
    .Y(_07854_));
 OA211x2_ASAP7_75t_R _23093_ (.A1(_06978_),
    .A2(_07762_),
    .B(_07833_),
    .C(_07854_),
    .Y(_07855_));
 AOI21x1_ASAP7_75t_R _23094_ (.A1(_01823_),
    .A2(_07786_),
    .B(_07855_),
    .Y(_02720_));
 OR3x2_ASAP7_75t_R _23095_ (.A(_01498_),
    .B(_15832_),
    .C(_15708_),
    .Y(_07856_));
 OR3x1_ASAP7_75t_R _23096_ (.A(_07813_),
    .B(_07837_),
    .C(_07856_),
    .Y(_07857_));
 XNOR2x2_ASAP7_75t_R _23097_ (.A(_16079_),
    .B(_07857_),
    .Y(_07858_));
 OA222x2_ASAP7_75t_R _23098_ (.A1(_01468_),
    .A2(_07810_),
    .B1(_07858_),
    .B2(_07845_),
    .C1(_07847_),
    .C2(_14354_),
    .Y(_07859_));
 OR3x1_ASAP7_75t_R _23099_ (.A(_07834_),
    .B(_07787_),
    .C(_07859_),
    .Y(_07860_));
 OA211x2_ASAP7_75t_R _23100_ (.A1(_07588_),
    .A2(_07762_),
    .B(_07833_),
    .C(_07860_),
    .Y(_07861_));
 AOI21x1_ASAP7_75t_R _23101_ (.A1(_01822_),
    .A2(_07786_),
    .B(_07861_),
    .Y(_02721_));
 BUFx6f_ASAP7_75t_R _23102_ (.A(_07539_),
    .Y(_07862_));
 OR3x1_ASAP7_75t_R _23103_ (.A(_16079_),
    .B(_07838_),
    .C(_07856_),
    .Y(_07863_));
 XNOR2x2_ASAP7_75t_R _23104_ (.A(_16192_),
    .B(_07863_),
    .Y(_07864_));
 OA222x2_ASAP7_75t_R _23105_ (.A1(_01467_),
    .A2(_07810_),
    .B1(_07864_),
    .B2(_07845_),
    .C1(_07847_),
    .C2(_14339_),
    .Y(_07865_));
 OR3x1_ASAP7_75t_R _23106_ (.A(_07834_),
    .B(_07787_),
    .C(_07865_),
    .Y(_07866_));
 OA211x2_ASAP7_75t_R _23107_ (.A1(_06995_),
    .A2(_07862_),
    .B(_07833_),
    .C(_07866_),
    .Y(_07867_));
 AOI21x1_ASAP7_75t_R _23108_ (.A1(_01821_),
    .A2(_07786_),
    .B(_07867_),
    .Y(_02722_));
 AND2x2_ASAP7_75t_R _23109_ (.A(_07775_),
    .B(_13237_),
    .Y(_07868_));
 AO21x1_ASAP7_75t_R _23110_ (.A1(_07774_),
    .A2(_01530_),
    .B(_07868_),
    .Y(_07869_));
 XNOR2x2_ASAP7_75t_R _23111_ (.A(_07790_),
    .B(_01496_),
    .Y(_07870_));
 OA222x2_ASAP7_75t_R _23112_ (.A1(_01466_),
    .A2(_07536_),
    .B1(_07773_),
    .B2(_07869_),
    .C1(_07870_),
    .C2(_07845_),
    .Y(_07871_));
 OAI22x1_ASAP7_75t_R _23113_ (.A1(_07079_),
    .A2(_07715_),
    .B1(_07781_),
    .B2(_07871_),
    .Y(_07872_));
 NOR2x1_ASAP7_75t_R _23114_ (.A(_01820_),
    .B(_07771_),
    .Y(_07873_));
 AO21x1_ASAP7_75t_R _23115_ (.A1(_07771_),
    .A2(_07872_),
    .B(_07873_),
    .Y(_02723_));
 OR5x1_ASAP7_75t_R _23116_ (.A(_16079_),
    .B(_16192_),
    .C(_07813_),
    .D(_07837_),
    .E(_07856_),
    .Y(_07874_));
 XNOR2x2_ASAP7_75t_R _23117_ (.A(_01495_),
    .B(_07874_),
    .Y(_07875_));
 OA222x2_ASAP7_75t_R _23118_ (.A1(_01465_),
    .A2(_07536_),
    .B1(_07875_),
    .B2(_07845_),
    .C1(_07847_),
    .C2(_15594_),
    .Y(_07876_));
 NOR2x1_ASAP7_75t_R _23119_ (.A(_07781_),
    .B(_07876_),
    .Y(_07877_));
 AO21x1_ASAP7_75t_R _23120_ (.A1(_06254_),
    .A2(_07713_),
    .B(_07877_),
    .Y(_07878_));
 NOR2x1_ASAP7_75t_R _23121_ (.A(_01819_),
    .B(_07771_),
    .Y(_07879_));
 AO21x1_ASAP7_75t_R _23122_ (.A1(_07771_),
    .A2(_07878_),
    .B(_07879_),
    .Y(_02724_));
 BUFx12f_ASAP7_75t_R _23123_ (.A(_07783_),
    .Y(_07880_));
 BUFx6f_ASAP7_75t_R _23124_ (.A(_07779_),
    .Y(_07881_));
 OR5x1_ASAP7_75t_R _23125_ (.A(_16079_),
    .B(_01495_),
    .C(_16192_),
    .D(_07838_),
    .E(_07856_),
    .Y(_07882_));
 XNOR2x2_ASAP7_75t_R _23126_ (.A(_01494_),
    .B(_07882_),
    .Y(_07883_));
 OA222x2_ASAP7_75t_R _23127_ (.A1(_01464_),
    .A2(_07810_),
    .B1(_07883_),
    .B2(_07795_),
    .C1(_07847_),
    .C2(_16332_),
    .Y(_07884_));
 OR3x1_ASAP7_75t_R _23128_ (.A(_07834_),
    .B(_07881_),
    .C(_07884_),
    .Y(_07885_));
 OA211x2_ASAP7_75t_R _23129_ (.A1(_07006_),
    .A2(_07862_),
    .B(_07833_),
    .C(_07885_),
    .Y(_07886_));
 AOI21x1_ASAP7_75t_R _23130_ (.A1(_01818_),
    .A2(_07880_),
    .B(_07886_),
    .Y(_02725_));
 OR5x1_ASAP7_75t_R _23131_ (.A(_16079_),
    .B(_01494_),
    .C(_01495_),
    .D(_16192_),
    .E(_07856_),
    .Y(_07887_));
 OR3x1_ASAP7_75t_R _23132_ (.A(_07813_),
    .B(_07837_),
    .C(_07887_),
    .Y(_07888_));
 XNOR2x2_ASAP7_75t_R _23133_ (.A(_01493_),
    .B(_07888_),
    .Y(_07889_));
 OA222x2_ASAP7_75t_R _23134_ (.A1(_01463_),
    .A2(_07810_),
    .B1(_07889_),
    .B2(_07795_),
    .C1(_07847_),
    .C2(_15587_),
    .Y(_07890_));
 OR3x1_ASAP7_75t_R _23135_ (.A(_07834_),
    .B(_07881_),
    .C(_07890_),
    .Y(_07891_));
 OA211x2_ASAP7_75t_R _23136_ (.A1(_07603_),
    .A2(_07862_),
    .B(_07833_),
    .C(_07891_),
    .Y(_07892_));
 AOI21x1_ASAP7_75t_R _23137_ (.A1(_01817_),
    .A2(_07880_),
    .B(_07892_),
    .Y(_02726_));
 BUFx6f_ASAP7_75t_R _23138_ (.A(_07512_),
    .Y(_07893_));
 OR3x1_ASAP7_75t_R _23139_ (.A(_01493_),
    .B(_07837_),
    .C(_07887_),
    .Y(_07894_));
 OR2x2_ASAP7_75t_R _23140_ (.A(_07803_),
    .B(_07894_),
    .Y(_07895_));
 XNOR2x2_ASAP7_75t_R _23141_ (.A(_16698_),
    .B(_07895_),
    .Y(_07896_));
 OA222x2_ASAP7_75t_R _23142_ (.A1(_01462_),
    .A2(_07893_),
    .B1(_07896_),
    .B2(_07795_),
    .C1(_07847_),
    .C2(_15482_),
    .Y(_07897_));
 OR3x1_ASAP7_75t_R _23143_ (.A(_07834_),
    .B(_07881_),
    .C(_07897_),
    .Y(_07898_));
 OA211x2_ASAP7_75t_R _23144_ (.A1(_07016_),
    .A2(_07862_),
    .B(_07833_),
    .C(_07898_),
    .Y(_07899_));
 AOI21x1_ASAP7_75t_R _23145_ (.A1(_01816_),
    .A2(_07880_),
    .B(_07899_),
    .Y(_02727_));
 OR3x1_ASAP7_75t_R _23146_ (.A(_16698_),
    .B(_07813_),
    .C(_07894_),
    .Y(_07900_));
 XNOR2x2_ASAP7_75t_R _23147_ (.A(_01491_),
    .B(_07900_),
    .Y(_07901_));
 OA222x2_ASAP7_75t_R _23148_ (.A1(_01461_),
    .A2(_07893_),
    .B1(_07901_),
    .B2(_07795_),
    .C1(_07846_),
    .C2(_15466_),
    .Y(_07902_));
 OR3x1_ASAP7_75t_R _23149_ (.A(_07834_),
    .B(_07881_),
    .C(_07902_),
    .Y(_07903_));
 OA211x2_ASAP7_75t_R _23150_ (.A1(_06344_),
    .A2(_07862_),
    .B(_07833_),
    .C(_07903_),
    .Y(_07904_));
 AOI21x1_ASAP7_75t_R _23151_ (.A1(_01815_),
    .A2(_07880_),
    .B(_07904_),
    .Y(_02728_));
 OR3x1_ASAP7_75t_R _23152_ (.A(_01491_),
    .B(_16698_),
    .C(_07894_),
    .Y(_07905_));
 OR2x2_ASAP7_75t_R _23153_ (.A(_07803_),
    .B(_07905_),
    .Y(_07906_));
 XNOR2x2_ASAP7_75t_R _23154_ (.A(_01490_),
    .B(_07906_),
    .Y(_07907_));
 OA222x2_ASAP7_75t_R _23155_ (.A1(_01460_),
    .A2(_07893_),
    .B1(_07847_),
    .B2(_13831_),
    .C1(_07907_),
    .C2(_07513_),
    .Y(_07908_));
 OR3x1_ASAP7_75t_R _23156_ (.A(_07834_),
    .B(_07881_),
    .C(_07908_),
    .Y(_07909_));
 OA211x2_ASAP7_75t_R _23157_ (.A1(_07026_),
    .A2(_07862_),
    .B(_07833_),
    .C(_07909_),
    .Y(_07910_));
 AOI21x1_ASAP7_75t_R _23158_ (.A1(_01814_),
    .A2(_07880_),
    .B(_07910_),
    .Y(_02729_));
 BUFx3_ASAP7_75t_R _23159_ (.A(_07770_),
    .Y(_07911_));
 OR3x1_ASAP7_75t_R _23160_ (.A(_01490_),
    .B(_07813_),
    .C(_07905_),
    .Y(_07912_));
 XNOR2x2_ASAP7_75t_R _23161_ (.A(_04306_),
    .B(_07912_),
    .Y(_07913_));
 OA222x2_ASAP7_75t_R _23162_ (.A1(_01459_),
    .A2(_07893_),
    .B1(_07913_),
    .B2(_07795_),
    .C1(_07846_),
    .C2(_13837_),
    .Y(_07914_));
 OR3x1_ASAP7_75t_R _23163_ (.A(_07566_),
    .B(_07881_),
    .C(_07914_),
    .Y(_07915_));
 OA211x2_ASAP7_75t_R _23164_ (.A1(_07613_),
    .A2(_07862_),
    .B(_07911_),
    .C(_07915_),
    .Y(_07916_));
 AOI21x1_ASAP7_75t_R _23165_ (.A1(_01813_),
    .A2(_07880_),
    .B(_07916_),
    .Y(_02730_));
 OR2x2_ASAP7_75t_R _23166_ (.A(_01490_),
    .B(_07905_),
    .Y(_07917_));
 OR3x1_ASAP7_75t_R _23167_ (.A(_04306_),
    .B(_07803_),
    .C(_07917_),
    .Y(_07918_));
 XNOR2x2_ASAP7_75t_R _23168_ (.A(_04419_),
    .B(_07918_),
    .Y(_07919_));
 OA222x2_ASAP7_75t_R _23169_ (.A1(_01458_),
    .A2(_07893_),
    .B1(_07846_),
    .B2(_13909_),
    .C1(_07919_),
    .C2(_07513_),
    .Y(_07920_));
 OR2x2_ASAP7_75t_R _23170_ (.A(_07781_),
    .B(_07920_),
    .Y(_07921_));
 OA211x2_ASAP7_75t_R _23171_ (.A1(_07037_),
    .A2(_07862_),
    .B(_07911_),
    .C(_07921_),
    .Y(_07922_));
 AOI21x1_ASAP7_75t_R _23172_ (.A1(_01812_),
    .A2(_07880_),
    .B(_07922_),
    .Y(_02731_));
 OR4x1_ASAP7_75t_R _23173_ (.A(_04419_),
    .B(_04306_),
    .C(_07791_),
    .D(_07917_),
    .Y(_07923_));
 XNOR2x2_ASAP7_75t_R _23174_ (.A(_01487_),
    .B(_07923_),
    .Y(_07924_));
 OA222x2_ASAP7_75t_R _23175_ (.A1(_01457_),
    .A2(_07512_),
    .B1(_07846_),
    .B2(_01513_),
    .C1(_07924_),
    .C2(_07513_),
    .Y(_07925_));
 OR2x2_ASAP7_75t_R _23176_ (.A(_07781_),
    .B(_07925_),
    .Y(_07926_));
 OA211x2_ASAP7_75t_R _23177_ (.A1(_07044_),
    .A2(_07862_),
    .B(_07911_),
    .C(_07926_),
    .Y(_07927_));
 AOI21x1_ASAP7_75t_R _23178_ (.A1(_01811_),
    .A2(_07880_),
    .B(_07927_),
    .Y(_02732_));
 OR4x1_ASAP7_75t_R _23179_ (.A(_01487_),
    .B(_04419_),
    .C(_04306_),
    .D(_07917_),
    .Y(_07928_));
 OR2x2_ASAP7_75t_R _23180_ (.A(_07803_),
    .B(_07928_),
    .Y(_07929_));
 XNOR2x2_ASAP7_75t_R _23181_ (.A(_04667_),
    .B(_07929_),
    .Y(_07930_));
 OA222x2_ASAP7_75t_R _23182_ (.A1(_01456_),
    .A2(_07512_),
    .B1(_07846_),
    .B2(_01512_),
    .C1(_07930_),
    .C2(_05400_),
    .Y(_07931_));
 OR2x2_ASAP7_75t_R _23183_ (.A(_07781_),
    .B(_07931_),
    .Y(_07932_));
 OA211x2_ASAP7_75t_R _23184_ (.A1(_07046_),
    .A2(_07862_),
    .B(_07911_),
    .C(_07932_),
    .Y(_07933_));
 AOI21x1_ASAP7_75t_R _23185_ (.A1(_01810_),
    .A2(_07880_),
    .B(_07933_),
    .Y(_02733_));
 AND2x2_ASAP7_75t_R _23186_ (.A(_07775_),
    .B(_13217_),
    .Y(_07934_));
 AO21x1_ASAP7_75t_R _23187_ (.A1(_07774_),
    .A2(_01529_),
    .B(_07934_),
    .Y(_07935_));
 NAND2x1_ASAP7_75t_R _23188_ (.A(\cs_registers_i.pc_id_i[2] ),
    .B(_07790_),
    .Y(_07936_));
 OA21x2_ASAP7_75t_R _23189_ (.A1(_00017_),
    .A2(_07790_),
    .B(_07936_),
    .Y(_07937_));
 OA222x2_ASAP7_75t_R _23190_ (.A1(_01455_),
    .A2(_07536_),
    .B1(_07773_),
    .B2(_07935_),
    .C1(_07937_),
    .C2(_07845_),
    .Y(_07938_));
 NAND2x1_ASAP7_75t_R _23191_ (.A(_05850_),
    .B(_07517_),
    .Y(_07939_));
 OA211x2_ASAP7_75t_R _23192_ (.A1(_07781_),
    .A2(_07938_),
    .B(_07939_),
    .C(_07770_),
    .Y(_07940_));
 AOI21x1_ASAP7_75t_R _23193_ (.A1(_01809_),
    .A2(_07880_),
    .B(_07940_),
    .Y(_02734_));
 OR3x1_ASAP7_75t_R _23194_ (.A(_04667_),
    .B(_07791_),
    .C(_07928_),
    .Y(_07941_));
 XNOR2x2_ASAP7_75t_R _23195_ (.A(_01485_),
    .B(_07941_),
    .Y(_07942_));
 OA222x2_ASAP7_75t_R _23196_ (.A1(_01454_),
    .A2(_07512_),
    .B1(_07846_),
    .B2(_14122_),
    .C1(_07942_),
    .C2(_05400_),
    .Y(_07943_));
 OR2x2_ASAP7_75t_R _23197_ (.A(_07780_),
    .B(_07943_),
    .Y(_07944_));
 OA211x2_ASAP7_75t_R _23198_ (.A1(_07626_),
    .A2(_07540_),
    .B(_07911_),
    .C(_07944_),
    .Y(_07945_));
 AOI21x1_ASAP7_75t_R _23199_ (.A1(_01808_),
    .A2(_07785_),
    .B(_07945_),
    .Y(_02735_));
 OR3x1_ASAP7_75t_R _23200_ (.A(_01485_),
    .B(_04667_),
    .C(_07929_),
    .Y(_07946_));
 XNOR2x2_ASAP7_75t_R _23201_ (.A(_01484_),
    .B(_07946_),
    .Y(_07947_));
 OA222x2_ASAP7_75t_R _23202_ (.A1(_01453_),
    .A2(_07536_),
    .B1(_07947_),
    .B2(_07845_),
    .C1(_07847_),
    .C2(_14099_),
    .Y(_07948_));
 NAND2x1_ASAP7_75t_R _23203_ (.A(_06503_),
    .B(_07517_),
    .Y(_07949_));
 OA211x2_ASAP7_75t_R _23204_ (.A1(_07781_),
    .A2(_07948_),
    .B(_07949_),
    .C(_07770_),
    .Y(_07950_));
 AOI21x1_ASAP7_75t_R _23205_ (.A1(_01807_),
    .A2(_07785_),
    .B(_07950_),
    .Y(_02736_));
 AND2x2_ASAP7_75t_R _23206_ (.A(_07775_),
    .B(_13263_),
    .Y(_07951_));
 AO21x1_ASAP7_75t_R _23207_ (.A1(_07774_),
    .A2(_01528_),
    .B(_07951_),
    .Y(_07952_));
 OAI21x1_ASAP7_75t_R _23208_ (.A1(_07790_),
    .A2(_02236_),
    .B(_14773_),
    .Y(_07953_));
 NAND2x1_ASAP7_75t_R _23209_ (.A(_07803_),
    .B(_07953_),
    .Y(_07954_));
 OA222x2_ASAP7_75t_R _23210_ (.A1(_01452_),
    .A2(_07536_),
    .B1(_07773_),
    .B2(_07952_),
    .C1(_07954_),
    .C2(_07845_),
    .Y(_07955_));
 NAND2x1_ASAP7_75t_R _23211_ (.A(_06556_),
    .B(_07517_),
    .Y(_07956_));
 OA211x2_ASAP7_75t_R _23212_ (.A1(_07781_),
    .A2(_07955_),
    .B(_07956_),
    .C(_07770_),
    .Y(_07957_));
 AOI21x1_ASAP7_75t_R _23213_ (.A1(_01806_),
    .A2(_07785_),
    .B(_07957_),
    .Y(_02737_));
 AND2x2_ASAP7_75t_R _23214_ (.A(_07775_),
    .B(_13280_),
    .Y(_07958_));
 AO21x1_ASAP7_75t_R _23215_ (.A1(_13534_),
    .A2(_01527_),
    .B(_07958_),
    .Y(_07959_));
 XNOR2x2_ASAP7_75t_R _23216_ (.A(_14837_),
    .B(_07813_),
    .Y(_07960_));
 OA222x2_ASAP7_75t_R _23217_ (.A1(_01451_),
    .A2(_07893_),
    .B1(_07772_),
    .B2(_07959_),
    .C1(_07960_),
    .C2(_07513_),
    .Y(_07961_));
 OR3x1_ASAP7_75t_R _23218_ (.A(_07566_),
    .B(_07881_),
    .C(_07961_),
    .Y(_07962_));
 OA211x2_ASAP7_75t_R _23219_ (.A1(_07177_),
    .A2(_07540_),
    .B(_07911_),
    .C(_07962_),
    .Y(_07963_));
 AOI21x1_ASAP7_75t_R _23220_ (.A1(_01805_),
    .A2(_07785_),
    .B(_07963_),
    .Y(_02738_));
 AND2x2_ASAP7_75t_R _23221_ (.A(_07775_),
    .B(_13242_),
    .Y(_07964_));
 AO21x1_ASAP7_75t_R _23222_ (.A1(_13534_),
    .A2(_01526_),
    .B(_07964_),
    .Y(_07965_));
 OR2x2_ASAP7_75t_R _23223_ (.A(_14837_),
    .B(_07803_),
    .Y(_07966_));
 XNOR2x2_ASAP7_75t_R _23224_ (.A(_14900_),
    .B(_07966_),
    .Y(_07967_));
 OA222x2_ASAP7_75t_R _23225_ (.A1(_01450_),
    .A2(_07893_),
    .B1(_07772_),
    .B2(_07965_),
    .C1(_07967_),
    .C2(_07513_),
    .Y(_07968_));
 OR3x1_ASAP7_75t_R _23226_ (.A(_07566_),
    .B(_07881_),
    .C(_07968_),
    .Y(_07969_));
 OA211x2_ASAP7_75t_R _23227_ (.A1(_07227_),
    .A2(_07540_),
    .B(_07911_),
    .C(_07969_),
    .Y(_07970_));
 AOI21x1_ASAP7_75t_R _23228_ (.A1(_01804_),
    .A2(_07785_),
    .B(_07970_),
    .Y(_02739_));
 AND2x2_ASAP7_75t_R _23229_ (.A(_13277_),
    .B(_13533_),
    .Y(_07971_));
 AO21x1_ASAP7_75t_R _23230_ (.A1(_13534_),
    .A2(_01525_),
    .B(_07971_),
    .Y(_07972_));
 OR3x1_ASAP7_75t_R _23231_ (.A(_14900_),
    .B(_14837_),
    .C(_07813_),
    .Y(_07973_));
 XNOR2x2_ASAP7_75t_R _23232_ (.A(_14966_),
    .B(_07973_),
    .Y(_07974_));
 OA222x2_ASAP7_75t_R _23233_ (.A1(_01449_),
    .A2(_07893_),
    .B1(_07772_),
    .B2(_07972_),
    .C1(_07974_),
    .C2(_07513_),
    .Y(_07975_));
 OR3x1_ASAP7_75t_R _23234_ (.A(_07566_),
    .B(_07881_),
    .C(_07975_),
    .Y(_07976_));
 OA211x2_ASAP7_75t_R _23235_ (.A1(_07249_),
    .A2(_07540_),
    .B(_07911_),
    .C(_07976_),
    .Y(_07977_));
 AOI21x1_ASAP7_75t_R _23236_ (.A1(_01803_),
    .A2(_07785_),
    .B(_07977_),
    .Y(_02740_));
 AND2x2_ASAP7_75t_R _23237_ (.A(_07775_),
    .B(_13430_),
    .Y(_07978_));
 AO21x1_ASAP7_75t_R _23238_ (.A1(_07774_),
    .A2(_01524_),
    .B(_07978_),
    .Y(_07979_));
 OR4x1_ASAP7_75t_R _23239_ (.A(_14966_),
    .B(_14900_),
    .C(_14837_),
    .D(_07803_),
    .Y(_07980_));
 XNOR2x2_ASAP7_75t_R _23240_ (.A(_01480_),
    .B(_07980_),
    .Y(_07981_));
 OA222x2_ASAP7_75t_R _23241_ (.A1(_01448_),
    .A2(_07536_),
    .B1(_07773_),
    .B2(_07979_),
    .C1(_07981_),
    .C2(_07845_),
    .Y(_07982_));
 NAND2x1_ASAP7_75t_R _23242_ (.A(_06650_),
    .B(_07517_),
    .Y(_07983_));
 OA211x2_ASAP7_75t_R _23243_ (.A1(_07781_),
    .A2(_07982_),
    .B(_07983_),
    .C(_07770_),
    .Y(_07984_));
 AOI21x1_ASAP7_75t_R _23244_ (.A1(_01802_),
    .A2(_07785_),
    .B(_07984_),
    .Y(_02741_));
 AND2x2_ASAP7_75t_R _23245_ (.A(_13533_),
    .B(_13455_),
    .Y(_07985_));
 AO21x1_ASAP7_75t_R _23246_ (.A1(_13534_),
    .A2(_01523_),
    .B(_07985_),
    .Y(_07986_));
 OR2x2_ASAP7_75t_R _23247_ (.A(_07813_),
    .B(_07792_),
    .Y(_07987_));
 XNOR2x2_ASAP7_75t_R _23248_ (.A(_15099_),
    .B(_07987_),
    .Y(_07988_));
 OA222x2_ASAP7_75t_R _23249_ (.A1(_01447_),
    .A2(_07893_),
    .B1(_07772_),
    .B2(_07986_),
    .C1(_07988_),
    .C2(_07513_),
    .Y(_07989_));
 OR3x1_ASAP7_75t_R _23250_ (.A(_07566_),
    .B(_07881_),
    .C(_07989_),
    .Y(_07990_));
 OA211x2_ASAP7_75t_R _23251_ (.A1(_07646_),
    .A2(_07540_),
    .B(_07911_),
    .C(_07990_),
    .Y(_07991_));
 AOI21x1_ASAP7_75t_R _23252_ (.A1(_01801_),
    .A2(_07785_),
    .B(_07991_),
    .Y(_02742_));
 AND2x2_ASAP7_75t_R _23253_ (.A(_13533_),
    .B(_13602_),
    .Y(_07992_));
 AO21x1_ASAP7_75t_R _23254_ (.A1(_13534_),
    .A2(_01522_),
    .B(_07992_),
    .Y(_07993_));
 OR3x1_ASAP7_75t_R _23255_ (.A(_15099_),
    .B(_07792_),
    .C(_07803_),
    .Y(_07994_));
 XNOR2x2_ASAP7_75t_R _23256_ (.A(_15158_),
    .B(_07994_),
    .Y(_07995_));
 OA222x2_ASAP7_75t_R _23257_ (.A1(_01446_),
    .A2(_07893_),
    .B1(_07772_),
    .B2(_07993_),
    .C1(_07995_),
    .C2(_07513_),
    .Y(_07996_));
 OR3x1_ASAP7_75t_R _23258_ (.A(_07566_),
    .B(_07779_),
    .C(_07996_),
    .Y(_07997_));
 OA211x2_ASAP7_75t_R _23259_ (.A1(_07129_),
    .A2(_07540_),
    .B(_07911_),
    .C(_07997_),
    .Y(_07998_));
 AOI21x1_ASAP7_75t_R _23260_ (.A1(_01800_),
    .A2(_07785_),
    .B(_07998_),
    .Y(_02743_));
 NAND2x1_ASAP7_75t_R _23261_ (.A(_05121_),
    .B(_05916_),
    .Y(_07999_));
 OR2x2_ASAP7_75t_R _23262_ (.A(_07999_),
    .B(_05937_),
    .Y(_08000_));
 BUFx6f_ASAP7_75t_R _23263_ (.A(_08000_),
    .Y(_08001_));
 BUFx6f_ASAP7_75t_R _23264_ (.A(_08001_),
    .Y(_08002_));
 INVx1_ASAP7_75t_R _23265_ (.A(net1),
    .Y(_08003_));
 AND3x4_ASAP7_75t_R _23266_ (.A(_05404_),
    .B(_05172_),
    .C(_05704_),
    .Y(_08004_));
 BUFx12f_ASAP7_75t_R _23267_ (.A(_08004_),
    .Y(_08005_));
 BUFx12f_ASAP7_75t_R _23268_ (.A(_08005_),
    .Y(_08006_));
 OA21x2_ASAP7_75t_R _23269_ (.A1(_05171_),
    .A2(_05705_),
    .B(_08001_),
    .Y(_08007_));
 BUFx6f_ASAP7_75t_R _23270_ (.A(_08007_),
    .Y(_08008_));
 BUFx12f_ASAP7_75t_R _23271_ (.A(_08008_),
    .Y(_08009_));
 AOI22x1_ASAP7_75t_R _23272_ (.A1(_08003_),
    .A2(_08006_),
    .B1(_08009_),
    .B2(_01405_),
    .Y(_08010_));
 OA21x2_ASAP7_75t_R _23273_ (.A1(_05981_),
    .A2(_08002_),
    .B(_08010_),
    .Y(_02744_));
 INVx1_ASAP7_75t_R _23274_ (.A(net2),
    .Y(_08011_));
 AOI22x1_ASAP7_75t_R _23275_ (.A1(_08011_),
    .A2(_08006_),
    .B1(_08009_),
    .B2(_00746_),
    .Y(_08012_));
 OA21x2_ASAP7_75t_R _23276_ (.A1(_06025_),
    .A2(_08002_),
    .B(_08012_),
    .Y(_02745_));
 INVx1_ASAP7_75t_R _23277_ (.A(net3),
    .Y(_08013_));
 AOI22x1_ASAP7_75t_R _23278_ (.A1(_08013_),
    .A2(_08006_),
    .B1(_08009_),
    .B2(_00745_),
    .Y(_08014_));
 OA21x2_ASAP7_75t_R _23279_ (.A1(_06052_),
    .A2(_08002_),
    .B(_08014_),
    .Y(_02746_));
 INVx1_ASAP7_75t_R _23280_ (.A(net4),
    .Y(_08015_));
 AOI22x1_ASAP7_75t_R _23281_ (.A1(_08015_),
    .A2(_08006_),
    .B1(_08009_),
    .B2(_01406_),
    .Y(_08016_));
 OA21x2_ASAP7_75t_R _23282_ (.A1(_06082_),
    .A2(_08002_),
    .B(_08016_),
    .Y(_02747_));
 INVx1_ASAP7_75t_R _23283_ (.A(net5),
    .Y(_08017_));
 AOI22x1_ASAP7_75t_R _23284_ (.A1(_08017_),
    .A2(_08006_),
    .B1(_08009_),
    .B2(_01407_),
    .Y(_08018_));
 OA21x2_ASAP7_75t_R _23285_ (.A1(_06108_),
    .A2(_08002_),
    .B(_08018_),
    .Y(_02748_));
 INVx1_ASAP7_75t_R _23286_ (.A(net6),
    .Y(_08019_));
 AOI22x1_ASAP7_75t_R _23287_ (.A1(_08019_),
    .A2(_08006_),
    .B1(_08009_),
    .B2(_01408_),
    .Y(_08020_));
 OA21x2_ASAP7_75t_R _23288_ (.A1(_06131_),
    .A2(_08002_),
    .B(_08020_),
    .Y(_02749_));
 INVx1_ASAP7_75t_R _23289_ (.A(net7),
    .Y(_08021_));
 AOI22x1_ASAP7_75t_R _23290_ (.A1(_08021_),
    .A2(_08006_),
    .B1(_08009_),
    .B2(_01409_),
    .Y(_08022_));
 OA21x2_ASAP7_75t_R _23291_ (.A1(_06153_),
    .A2(_08002_),
    .B(_08022_),
    .Y(_02750_));
 INVx1_ASAP7_75t_R _23292_ (.A(net8),
    .Y(_08023_));
 AOI22x1_ASAP7_75t_R _23293_ (.A1(_08023_),
    .A2(_08006_),
    .B1(_08009_),
    .B2(_01410_),
    .Y(_08024_));
 OA21x2_ASAP7_75t_R _23294_ (.A1(_06179_),
    .A2(_08002_),
    .B(_08024_),
    .Y(_02751_));
 INVx1_ASAP7_75t_R _23295_ (.A(net9),
    .Y(_08025_));
 AOI22x1_ASAP7_75t_R _23296_ (.A1(_08025_),
    .A2(_08006_),
    .B1(_08009_),
    .B2(_01411_),
    .Y(_08026_));
 OA21x2_ASAP7_75t_R _23297_ (.A1(_06197_),
    .A2(_08002_),
    .B(_08026_),
    .Y(_02752_));
 INVx1_ASAP7_75t_R _23298_ (.A(net10),
    .Y(_08027_));
 AOI22x1_ASAP7_75t_R _23299_ (.A1(_08027_),
    .A2(_08006_),
    .B1(_08009_),
    .B2(_01412_),
    .Y(_08028_));
 OA21x2_ASAP7_75t_R _23300_ (.A1(_06219_),
    .A2(_08002_),
    .B(_08028_),
    .Y(_02753_));
 BUFx6f_ASAP7_75t_R _23301_ (.A(_08001_),
    .Y(_08029_));
 INVx1_ASAP7_75t_R _23302_ (.A(net11),
    .Y(_08030_));
 BUFx12f_ASAP7_75t_R _23303_ (.A(_08005_),
    .Y(_08031_));
 BUFx12f_ASAP7_75t_R _23304_ (.A(_08008_),
    .Y(_08032_));
 AOI22x1_ASAP7_75t_R _23305_ (.A1(_08030_),
    .A2(_08031_),
    .B1(_08032_),
    .B2(_01413_),
    .Y(_08033_));
 OA21x2_ASAP7_75t_R _23306_ (.A1(_06255_),
    .A2(_08029_),
    .B(_08033_),
    .Y(_02754_));
 INVx1_ASAP7_75t_R _23307_ (.A(net12),
    .Y(_08034_));
 AOI22x1_ASAP7_75t_R _23308_ (.A1(_08034_),
    .A2(_08031_),
    .B1(_08032_),
    .B2(_01414_),
    .Y(_08035_));
 OA21x2_ASAP7_75t_R _23309_ (.A1(_06277_),
    .A2(_08029_),
    .B(_08035_),
    .Y(_02755_));
 INVx1_ASAP7_75t_R _23310_ (.A(net13),
    .Y(_08036_));
 AOI22x1_ASAP7_75t_R _23311_ (.A1(_08036_),
    .A2(_08031_),
    .B1(_08032_),
    .B2(_01415_),
    .Y(_08037_));
 OA21x2_ASAP7_75t_R _23312_ (.A1(_06298_),
    .A2(_08029_),
    .B(_08037_),
    .Y(_02756_));
 INVx1_ASAP7_75t_R _23313_ (.A(net14),
    .Y(_08038_));
 AOI22x1_ASAP7_75t_R _23314_ (.A1(_08038_),
    .A2(_08031_),
    .B1(_08032_),
    .B2(_00007_),
    .Y(_08039_));
 OA21x2_ASAP7_75t_R _23315_ (.A1(_06323_),
    .A2(_08029_),
    .B(_08039_),
    .Y(_02757_));
 INVx1_ASAP7_75t_R _23316_ (.A(net15),
    .Y(_08040_));
 AOI22x1_ASAP7_75t_R _23317_ (.A1(_08040_),
    .A2(_08031_),
    .B1(_08032_),
    .B2(_00008_),
    .Y(_08041_));
 OA21x2_ASAP7_75t_R _23318_ (.A1(_06343_),
    .A2(_08029_),
    .B(_08041_),
    .Y(_02758_));
 INVx1_ASAP7_75t_R _23319_ (.A(net16),
    .Y(_08042_));
 AOI22x1_ASAP7_75t_R _23320_ (.A1(_08042_),
    .A2(_08031_),
    .B1(_08032_),
    .B2(_00009_),
    .Y(_08043_));
 OA21x2_ASAP7_75t_R _23321_ (.A1(_06366_),
    .A2(_08029_),
    .B(_08043_),
    .Y(_02759_));
 INVx1_ASAP7_75t_R _23322_ (.A(net17),
    .Y(_08044_));
 AOI22x1_ASAP7_75t_R _23323_ (.A1(_08044_),
    .A2(_08031_),
    .B1(_08032_),
    .B2(_00010_),
    .Y(_08045_));
 OA21x2_ASAP7_75t_R _23324_ (.A1(_06391_),
    .A2(_08029_),
    .B(_08045_),
    .Y(_02760_));
 INVx1_ASAP7_75t_R _23325_ (.A(net18),
    .Y(_08046_));
 AOI22x1_ASAP7_75t_R _23326_ (.A1(_08046_),
    .A2(_08031_),
    .B1(_08032_),
    .B2(_00011_),
    .Y(_08047_));
 OA21x2_ASAP7_75t_R _23327_ (.A1(_06411_),
    .A2(_08029_),
    .B(_08047_),
    .Y(_02761_));
 INVx1_ASAP7_75t_R _23328_ (.A(net19),
    .Y(_08048_));
 AOI22x1_ASAP7_75t_R _23329_ (.A1(_08048_),
    .A2(_08031_),
    .B1(_08032_),
    .B2(_00012_),
    .Y(_08049_));
 OA21x2_ASAP7_75t_R _23330_ (.A1(_06432_),
    .A2(_08029_),
    .B(_08049_),
    .Y(_02762_));
 INVx1_ASAP7_75t_R _23331_ (.A(net20),
    .Y(_08050_));
 AOI22x1_ASAP7_75t_R _23332_ (.A1(_08050_),
    .A2(_08031_),
    .B1(_08032_),
    .B2(_00013_),
    .Y(_08051_));
 OA21x2_ASAP7_75t_R _23333_ (.A1(_06454_),
    .A2(_08029_),
    .B(_08051_),
    .Y(_02763_));
 INVx1_ASAP7_75t_R _23334_ (.A(net21),
    .Y(_08052_));
 AOI22x1_ASAP7_75t_R _23335_ (.A1(_08052_),
    .A2(_08005_),
    .B1(_08008_),
    .B2(_00014_),
    .Y(_08053_));
 OA21x2_ASAP7_75t_R _23336_ (.A1(_06480_),
    .A2(_08001_),
    .B(_08053_),
    .Y(_02764_));
 INVx1_ASAP7_75t_R _23337_ (.A(net22),
    .Y(_08054_));
 AOI22x1_ASAP7_75t_R _23338_ (.A1(_08054_),
    .A2(_08005_),
    .B1(_08008_),
    .B2(_00015_),
    .Y(_08055_));
 OA21x2_ASAP7_75t_R _23339_ (.A1(_06504_),
    .A2(_08001_),
    .B(_08055_),
    .Y(_02765_));
 INVx1_ASAP7_75t_R _23340_ (.A(net23),
    .Y(_08056_));
 AOI22x1_ASAP7_75t_R _23341_ (.A1(_08056_),
    .A2(_08005_),
    .B1(_08008_),
    .B2(_01403_),
    .Y(_08057_));
 OA21x2_ASAP7_75t_R _23342_ (.A1(_06675_),
    .A2(_08001_),
    .B(_08057_),
    .Y(_02766_));
 INVx1_ASAP7_75t_R _23343_ (.A(net24),
    .Y(_08058_));
 AOI22x1_ASAP7_75t_R _23344_ (.A1(_08058_),
    .A2(_08005_),
    .B1(_08008_),
    .B2(_01404_),
    .Y(_08059_));
 OA21x2_ASAP7_75t_R _23345_ (.A1(_06699_),
    .A2(_08001_),
    .B(_08059_),
    .Y(_02767_));
 OA21x2_ASAP7_75t_R _23346_ (.A1(_13837_),
    .A2(_14272_),
    .B(_14112_),
    .Y(_08060_));
 AND3x4_ASAP7_75t_R _23347_ (.A(_14541_),
    .B(_14623_),
    .C(_08060_),
    .Y(_08061_));
 BUFx6f_ASAP7_75t_R _23348_ (.A(_08061_),
    .Y(_08062_));
 INVx1_ASAP7_75t_R _23349_ (.A(_08062_),
    .Y(_08063_));
 OR3x1_ASAP7_75t_R _23350_ (.A(_02192_),
    .B(_05205_),
    .C(_08063_),
    .Y(_08064_));
 NAND2x1_ASAP7_75t_R _23351_ (.A(_01799_),
    .B(_08064_),
    .Y(_08065_));
 OA21x2_ASAP7_75t_R _23352_ (.A1(_05233_),
    .A2(_08064_),
    .B(_08065_),
    .Y(_02768_));
 AND3x4_ASAP7_75t_R _23353_ (.A(_14634_),
    .B(_02192_),
    .C(_02193_),
    .Y(_08066_));
 AND3x1_ASAP7_75t_R _23354_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_05196_),
    .C(_08066_),
    .Y(_08067_));
 AOI21x1_ASAP7_75t_R _23355_ (.A1(_05254_),
    .A2(_05206_),
    .B(_08067_),
    .Y(_02769_));
 BUFx6f_ASAP7_75t_R _23356_ (.A(_02237_),
    .Y(_08068_));
 INVx2_ASAP7_75t_R _23357_ (.A(_08068_),
    .Y(_08069_));
 AND3x1_ASAP7_75t_R _23358_ (.A(_08069_),
    .B(_05196_),
    .C(_08066_),
    .Y(_08070_));
 AOI21x1_ASAP7_75t_R _23359_ (.A1(_18084_),
    .A2(_05206_),
    .B(_08070_),
    .Y(_02770_));
 XNOR2x2_ASAP7_75t_R _23360_ (.A(_05186_),
    .B(_02238_),
    .Y(_08071_));
 AND3x1_ASAP7_75t_R _23361_ (.A(_05196_),
    .B(_08066_),
    .C(_08071_),
    .Y(_08072_));
 AOI21x1_ASAP7_75t_R _23362_ (.A1(_05186_),
    .A2(_05206_),
    .B(_08072_),
    .Y(_02771_));
 INVx2_ASAP7_75t_R _23363_ (.A(_05187_),
    .Y(_08073_));
 AND3x1_ASAP7_75t_R _23364_ (.A(_05186_),
    .B(_18083_),
    .C(_18084_),
    .Y(_08074_));
 XNOR2x2_ASAP7_75t_R _23365_ (.A(_08073_),
    .B(_08074_),
    .Y(_08075_));
 AND3x1_ASAP7_75t_R _23366_ (.A(_05196_),
    .B(_08066_),
    .C(_08075_),
    .Y(_08076_));
 AOI21x1_ASAP7_75t_R _23367_ (.A1(_05187_),
    .A2(_05206_),
    .B(_08076_),
    .Y(_02772_));
 NAND2x1_ASAP7_75t_R _23368_ (.A(_05186_),
    .B(_05187_),
    .Y(_08077_));
 BUFx6f_ASAP7_75t_R _23369_ (.A(_08077_),
    .Y(_08078_));
 OA21x2_ASAP7_75t_R _23370_ (.A1(_02238_),
    .A2(_08078_),
    .B(_08066_),
    .Y(_08079_));
 OA21x2_ASAP7_75t_R _23371_ (.A1(_05205_),
    .A2(_08079_),
    .B(_01394_),
    .Y(_08080_));
 INVx2_ASAP7_75t_R _23372_ (.A(_01394_),
    .Y(_08081_));
 NOR2x1_ASAP7_75t_R _23373_ (.A(_02238_),
    .B(_08078_),
    .Y(_08082_));
 AND5x1_ASAP7_75t_R _23374_ (.A(_08081_),
    .B(_05193_),
    .C(_05722_),
    .D(_08066_),
    .E(_08082_),
    .Y(_08083_));
 NOR2x1_ASAP7_75t_R _23375_ (.A(_08080_),
    .B(_08083_),
    .Y(_02773_));
 NAND2x2_ASAP7_75t_R _23376_ (.A(_14640_),
    .B(_05195_),
    .Y(_08084_));
 BUFx6f_ASAP7_75t_R _23377_ (.A(_08084_),
    .Y(_08085_));
 INVx1_ASAP7_75t_R _23378_ (.A(_05350_),
    .Y(_08086_));
 BUFx6f_ASAP7_75t_R _23379_ (.A(_08086_),
    .Y(_08087_));
 BUFx6f_ASAP7_75t_R _23380_ (.A(_08087_),
    .Y(_08088_));
 AND2x2_ASAP7_75t_R _23381_ (.A(_14624_),
    .B(_05348_),
    .Y(_08089_));
 AND3x1_ASAP7_75t_R _23382_ (.A(_05255_),
    .B(_04962_),
    .C(_08089_),
    .Y(_08090_));
 AO21x1_ASAP7_75t_R _23383_ (.A1(_14635_),
    .A2(_08088_),
    .B(_08090_),
    .Y(_08091_));
 BUFx6f_ASAP7_75t_R _23384_ (.A(_14640_),
    .Y(_08092_));
 INVx1_ASAP7_75t_R _23385_ (.A(_00066_),
    .Y(_08093_));
 AO21x1_ASAP7_75t_R _23386_ (.A1(_08092_),
    .A2(_05204_),
    .B(_08093_),
    .Y(_08094_));
 OA21x2_ASAP7_75t_R _23387_ (.A1(_08085_),
    .A2(_08091_),
    .B(_08094_),
    .Y(_02774_));
 BUFx6f_ASAP7_75t_R _23388_ (.A(_05350_),
    .Y(_08095_));
 AND2x2_ASAP7_75t_R _23389_ (.A(_05324_),
    .B(_08087_),
    .Y(_08096_));
 AO21x1_ASAP7_75t_R _23390_ (.A1(\alu_adder_result_ex[10] ),
    .A2(_08095_),
    .B(_08096_),
    .Y(_08097_));
 BUFx6f_ASAP7_75t_R _23391_ (.A(_08084_),
    .Y(_08098_));
 NAND2x1_ASAP7_75t_R _23392_ (.A(_00076_),
    .B(_08098_),
    .Y(_08099_));
 OA21x2_ASAP7_75t_R _23393_ (.A1(_08085_),
    .A2(_08097_),
    .B(_08099_),
    .Y(_02775_));
 BUFx6f_ASAP7_75t_R _23394_ (.A(_05350_),
    .Y(_08100_));
 OR2x2_ASAP7_75t_R _23395_ (.A(_05328_),
    .B(_08100_),
    .Y(_08101_));
 OA21x2_ASAP7_75t_R _23396_ (.A1(\alu_adder_result_ex[11] ),
    .A2(_08088_),
    .B(_08101_),
    .Y(_08102_));
 NAND2x1_ASAP7_75t_R _23397_ (.A(_00075_),
    .B(_08098_),
    .Y(_08103_));
 OA21x2_ASAP7_75t_R _23398_ (.A1(_08085_),
    .A2(_08102_),
    .B(_08103_),
    .Y(_02776_));
 NOR2x1_ASAP7_75t_R _23399_ (.A(_05618_),
    .B(_08095_),
    .Y(_08104_));
 AO21x1_ASAP7_75t_R _23400_ (.A1(\alu_adder_result_ex[12] ),
    .A2(_08095_),
    .B(_08104_),
    .Y(_08105_));
 INVx1_ASAP7_75t_R _23401_ (.A(_00078_),
    .Y(_08106_));
 AO21x1_ASAP7_75t_R _23402_ (.A1(_08092_),
    .A2(_05204_),
    .B(_08106_),
    .Y(_08107_));
 OA21x2_ASAP7_75t_R _23403_ (.A1(_08085_),
    .A2(_08105_),
    .B(_08107_),
    .Y(_02777_));
 OR2x2_ASAP7_75t_R _23404_ (.A(_05624_),
    .B(_08100_),
    .Y(_08108_));
 OA21x2_ASAP7_75t_R _23405_ (.A1(\alu_adder_result_ex[13] ),
    .A2(_08088_),
    .B(_08108_),
    .Y(_08109_));
 INVx1_ASAP7_75t_R _23406_ (.A(_00077_),
    .Y(_08110_));
 AO21x1_ASAP7_75t_R _23407_ (.A1(_08092_),
    .A2(_05204_),
    .B(_08110_),
    .Y(_08111_));
 OA21x2_ASAP7_75t_R _23408_ (.A1(_08085_),
    .A2(_08109_),
    .B(_08111_),
    .Y(_02778_));
 AO21x1_ASAP7_75t_R _23409_ (.A1(_15551_),
    .A2(_15582_),
    .B(_08100_),
    .Y(_08112_));
 OA21x2_ASAP7_75t_R _23410_ (.A1(\alu_adder_result_ex[14] ),
    .A2(_08088_),
    .B(_08112_),
    .Y(_08113_));
 NAND2x1_ASAP7_75t_R _23411_ (.A(_00080_),
    .B(_08098_),
    .Y(_08114_));
 OA21x2_ASAP7_75t_R _23412_ (.A1(_08085_),
    .A2(_08113_),
    .B(_08114_),
    .Y(_02779_));
 OR2x2_ASAP7_75t_R _23413_ (.A(_15707_),
    .B(_08100_),
    .Y(_08115_));
 OA21x2_ASAP7_75t_R _23414_ (.A1(\alu_adder_result_ex[15] ),
    .A2(_08088_),
    .B(_08115_),
    .Y(_08116_));
 NAND2x1_ASAP7_75t_R _23415_ (.A(_00079_),
    .B(_08098_),
    .Y(_08117_));
 OA21x2_ASAP7_75t_R _23416_ (.A1(_08085_),
    .A2(_08116_),
    .B(_08117_),
    .Y(_02780_));
 OR2x2_ASAP7_75t_R _23417_ (.A(_15831_),
    .B(_08100_),
    .Y(_08118_));
 OA21x2_ASAP7_75t_R _23418_ (.A1(\alu_adder_result_ex[16] ),
    .A2(_08088_),
    .B(_08118_),
    .Y(_08119_));
 NAND2x1_ASAP7_75t_R _23419_ (.A(_00082_),
    .B(_08098_),
    .Y(_08120_));
 OA21x2_ASAP7_75t_R _23420_ (.A1(_08085_),
    .A2(_08119_),
    .B(_08120_),
    .Y(_02781_));
 OR2x2_ASAP7_75t_R _23421_ (.A(_05281_),
    .B(_08100_),
    .Y(_08121_));
 OA21x2_ASAP7_75t_R _23422_ (.A1(\alu_adder_result_ex[17] ),
    .A2(_08088_),
    .B(_08121_),
    .Y(_08122_));
 INVx1_ASAP7_75t_R _23423_ (.A(_00081_),
    .Y(_08123_));
 AO21x1_ASAP7_75t_R _23424_ (.A1(_08092_),
    .A2(_05204_),
    .B(_08123_),
    .Y(_08124_));
 OA21x2_ASAP7_75t_R _23425_ (.A1(_08085_),
    .A2(_08122_),
    .B(_08124_),
    .Y(_02782_));
 OR2x2_ASAP7_75t_R _23426_ (.A(_16078_),
    .B(_08100_),
    .Y(_08125_));
 OA21x2_ASAP7_75t_R _23427_ (.A1(\alu_adder_result_ex[18] ),
    .A2(_08088_),
    .B(_08125_),
    .Y(_08126_));
 NAND2x1_ASAP7_75t_R _23428_ (.A(_00084_),
    .B(_08098_),
    .Y(_08127_));
 OA21x2_ASAP7_75t_R _23429_ (.A1(_08085_),
    .A2(_08126_),
    .B(_08127_),
    .Y(_02783_));
 BUFx6f_ASAP7_75t_R _23430_ (.A(_08084_),
    .Y(_08128_));
 OR2x2_ASAP7_75t_R _23431_ (.A(_05650_),
    .B(_08100_),
    .Y(_08129_));
 OA21x2_ASAP7_75t_R _23432_ (.A1(\alu_adder_result_ex[19] ),
    .A2(_08088_),
    .B(_08129_),
    .Y(_08130_));
 NAND2x1_ASAP7_75t_R _23433_ (.A(_00083_),
    .B(_08098_),
    .Y(_08131_));
 OA21x2_ASAP7_75t_R _23434_ (.A1(_08128_),
    .A2(_08130_),
    .B(_08131_),
    .Y(_02784_));
 NOR2x1_ASAP7_75t_R _23435_ (.A(_14528_),
    .B(_08095_),
    .Y(_08132_));
 AO21x1_ASAP7_75t_R _23436_ (.A1(\alu_adder_result_ex[1] ),
    .A2(_08095_),
    .B(_08132_),
    .Y(_08133_));
 INVx1_ASAP7_75t_R _23437_ (.A(_00065_),
    .Y(_08134_));
 AO21x1_ASAP7_75t_R _23438_ (.A1(_08092_),
    .A2(_05204_),
    .B(_08134_),
    .Y(_08135_));
 OA21x2_ASAP7_75t_R _23439_ (.A1(_08128_),
    .A2(_08133_),
    .B(_08135_),
    .Y(_02785_));
 OR2x2_ASAP7_75t_R _23440_ (.A(_05654_),
    .B(_08100_),
    .Y(_08136_));
 OA21x2_ASAP7_75t_R _23441_ (.A1(\alu_adder_result_ex[20] ),
    .A2(_08088_),
    .B(_08136_),
    .Y(_08137_));
 NAND2x1_ASAP7_75t_R _23442_ (.A(_00086_),
    .B(_08098_),
    .Y(_08138_));
 OA21x2_ASAP7_75t_R _23443_ (.A1(_08128_),
    .A2(_08137_),
    .B(_08138_),
    .Y(_02786_));
 BUFx6f_ASAP7_75t_R _23444_ (.A(_08087_),
    .Y(_08139_));
 OR2x2_ASAP7_75t_R _23445_ (.A(_05295_),
    .B(_08100_),
    .Y(_08140_));
 OA21x2_ASAP7_75t_R _23446_ (.A1(\alu_adder_result_ex[21] ),
    .A2(_08139_),
    .B(_08140_),
    .Y(_08141_));
 INVx1_ASAP7_75t_R _23447_ (.A(_00085_),
    .Y(_08142_));
 AO21x1_ASAP7_75t_R _23448_ (.A1(_08092_),
    .A2(_05204_),
    .B(_08142_),
    .Y(_08143_));
 OA21x2_ASAP7_75t_R _23449_ (.A1(_08128_),
    .A2(_08141_),
    .B(_08143_),
    .Y(_02787_));
 BUFx3_ASAP7_75t_R _23450_ (.A(_05350_),
    .Y(_08144_));
 OR2x2_ASAP7_75t_R _23451_ (.A(_16587_),
    .B(_08144_),
    .Y(_08145_));
 OA21x2_ASAP7_75t_R _23452_ (.A1(\alu_adder_result_ex[22] ),
    .A2(_08139_),
    .B(_08145_),
    .Y(_08146_));
 BUFx12f_ASAP7_75t_R _23453_ (.A(_08084_),
    .Y(_08147_));
 NAND2x1_ASAP7_75t_R _23454_ (.A(_00088_),
    .B(_08147_),
    .Y(_08148_));
 OA21x2_ASAP7_75t_R _23455_ (.A1(_08128_),
    .A2(_08146_),
    .B(_08148_),
    .Y(_02788_));
 OR2x2_ASAP7_75t_R _23456_ (.A(_05308_),
    .B(_08144_),
    .Y(_08149_));
 OA21x2_ASAP7_75t_R _23457_ (.A1(\alu_adder_result_ex[23] ),
    .A2(_08139_),
    .B(_08149_),
    .Y(_08150_));
 NAND2x1_ASAP7_75t_R _23458_ (.A(_00087_),
    .B(_08147_),
    .Y(_08151_));
 OA21x2_ASAP7_75t_R _23459_ (.A1(_08128_),
    .A2(_08150_),
    .B(_08151_),
    .Y(_02789_));
 OR2x2_ASAP7_75t_R _23460_ (.A(_05672_),
    .B(_08144_),
    .Y(_08152_));
 OA21x2_ASAP7_75t_R _23461_ (.A1(\alu_adder_result_ex[24] ),
    .A2(_08139_),
    .B(_08152_),
    .Y(_08153_));
 NAND2x1_ASAP7_75t_R _23462_ (.A(_00090_),
    .B(_08147_),
    .Y(_08154_));
 OA21x2_ASAP7_75t_R _23463_ (.A1(_08128_),
    .A2(_08153_),
    .B(_08154_),
    .Y(_02790_));
 OR2x2_ASAP7_75t_R _23464_ (.A(_16931_),
    .B(_08144_),
    .Y(_08155_));
 OA21x2_ASAP7_75t_R _23465_ (.A1(\alu_adder_result_ex[25] ),
    .A2(_08139_),
    .B(_08155_),
    .Y(_08156_));
 INVx1_ASAP7_75t_R _23466_ (.A(_00089_),
    .Y(_08157_));
 AO21x1_ASAP7_75t_R _23467_ (.A1(_08092_),
    .A2(_05204_),
    .B(_08157_),
    .Y(_08158_));
 OA21x2_ASAP7_75t_R _23468_ (.A1(_08128_),
    .A2(_08156_),
    .B(_08158_),
    .Y(_02791_));
 OR2x2_ASAP7_75t_R _23469_ (.A(_04305_),
    .B(_08144_),
    .Y(_08159_));
 OA21x2_ASAP7_75t_R _23470_ (.A1(\alu_adder_result_ex[26] ),
    .A2(_08139_),
    .B(_08159_),
    .Y(_08160_));
 NAND2x1_ASAP7_75t_R _23471_ (.A(_00092_),
    .B(_08147_),
    .Y(_08161_));
 OA21x2_ASAP7_75t_R _23472_ (.A1(_08128_),
    .A2(_08160_),
    .B(_08161_),
    .Y(_02792_));
 NOR2x1_ASAP7_75t_R _23473_ (.A(_05685_),
    .B(_08095_),
    .Y(_08162_));
 AO21x1_ASAP7_75t_R _23474_ (.A1(\alu_adder_result_ex[27] ),
    .A2(_08095_),
    .B(_08162_),
    .Y(_08163_));
 NAND2x1_ASAP7_75t_R _23475_ (.A(_00091_),
    .B(_08147_),
    .Y(_08164_));
 OA21x2_ASAP7_75t_R _23476_ (.A1(_08128_),
    .A2(_08163_),
    .B(_08164_),
    .Y(_02793_));
 BUFx6f_ASAP7_75t_R _23477_ (.A(_08084_),
    .Y(_08165_));
 OR2x2_ASAP7_75t_R _23478_ (.A(_04554_),
    .B(_08144_),
    .Y(_08166_));
 OA21x2_ASAP7_75t_R _23479_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_08139_),
    .B(_08166_),
    .Y(_08167_));
 NAND2x1_ASAP7_75t_R _23480_ (.A(_00094_),
    .B(_08147_),
    .Y(_08168_));
 OA21x2_ASAP7_75t_R _23481_ (.A1(_08165_),
    .A2(_08167_),
    .B(_08168_),
    .Y(_02794_));
 OR2x2_ASAP7_75t_R _23482_ (.A(_05343_),
    .B(_08144_),
    .Y(_08169_));
 OA21x2_ASAP7_75t_R _23483_ (.A1(\alu_adder_result_ex[29] ),
    .A2(_08139_),
    .B(_08169_),
    .Y(_08170_));
 BUFx6f_ASAP7_75t_R _23484_ (.A(_05196_),
    .Y(_08171_));
 INVx1_ASAP7_75t_R _23485_ (.A(_00093_),
    .Y(_08172_));
 AO21x1_ASAP7_75t_R _23486_ (.A1(_08092_),
    .A2(_08171_),
    .B(_08172_),
    .Y(_08173_));
 OA21x2_ASAP7_75t_R _23487_ (.A1(_08165_),
    .A2(_08170_),
    .B(_08173_),
    .Y(_02795_));
 OR2x2_ASAP7_75t_R _23488_ (.A(_14703_),
    .B(_08144_),
    .Y(_08174_));
 OA21x2_ASAP7_75t_R _23489_ (.A1(\alu_adder_result_ex[2] ),
    .A2(_08139_),
    .B(_08174_),
    .Y(_08175_));
 NAND2x1_ASAP7_75t_R _23490_ (.A(_00068_),
    .B(_08147_),
    .Y(_08176_));
 OA21x2_ASAP7_75t_R _23491_ (.A1(_08165_),
    .A2(_08175_),
    .B(_08176_),
    .Y(_02796_));
 OR2x2_ASAP7_75t_R _23492_ (.A(_05358_),
    .B(_08144_),
    .Y(_08177_));
 OA21x2_ASAP7_75t_R _23493_ (.A1(\alu_adder_result_ex[30] ),
    .A2(_08139_),
    .B(_08177_),
    .Y(_08178_));
 NAND2x1_ASAP7_75t_R _23494_ (.A(_00096_),
    .B(_08147_),
    .Y(_08179_));
 OA21x2_ASAP7_75t_R _23495_ (.A1(_08165_),
    .A2(_08178_),
    .B(_08179_),
    .Y(_02797_));
 AOI21x1_ASAP7_75t_R _23496_ (.A1(_04971_),
    .A2(_08089_),
    .B(_04900_),
    .Y(_08180_));
 NAND2x1_ASAP7_75t_R _23497_ (.A(_00095_),
    .B(_08147_),
    .Y(_08181_));
 OA21x2_ASAP7_75t_R _23498_ (.A1(_08165_),
    .A2(_08180_),
    .B(_08181_),
    .Y(_02798_));
 OR2x2_ASAP7_75t_R _23499_ (.A(_14770_),
    .B(_08144_),
    .Y(_08182_));
 OA21x2_ASAP7_75t_R _23500_ (.A1(\alu_adder_result_ex[3] ),
    .A2(_08087_),
    .B(_08182_),
    .Y(_08183_));
 NAND2x1_ASAP7_75t_R _23501_ (.A(_00067_),
    .B(_08147_),
    .Y(_08184_));
 OA21x2_ASAP7_75t_R _23502_ (.A1(_08165_),
    .A2(_08183_),
    .B(_08184_),
    .Y(_02799_));
 AND2x2_ASAP7_75t_R _23503_ (.A(_14835_),
    .B(_08087_),
    .Y(_08185_));
 AO21x1_ASAP7_75t_R _23504_ (.A1(\alu_adder_result_ex[4] ),
    .A2(_08095_),
    .B(_08185_),
    .Y(_08186_));
 INVx1_ASAP7_75t_R _23505_ (.A(_00070_),
    .Y(_08187_));
 AO21x1_ASAP7_75t_R _23506_ (.A1(_08092_),
    .A2(_08171_),
    .B(_08187_),
    .Y(_08188_));
 OA21x2_ASAP7_75t_R _23507_ (.A1(_08165_),
    .A2(_08186_),
    .B(_08188_),
    .Y(_02800_));
 OR2x2_ASAP7_75t_R _23508_ (.A(_05583_),
    .B(_05350_),
    .Y(_08189_));
 OA21x2_ASAP7_75t_R _23509_ (.A1(\alu_adder_result_ex[5] ),
    .A2(_08087_),
    .B(_08189_),
    .Y(_08190_));
 INVx1_ASAP7_75t_R _23510_ (.A(_00069_),
    .Y(_08191_));
 AO21x1_ASAP7_75t_R _23511_ (.A1(_08092_),
    .A2(_08171_),
    .B(_08191_),
    .Y(_08192_));
 OA21x2_ASAP7_75t_R _23512_ (.A1(_08165_),
    .A2(_08190_),
    .B(_08192_),
    .Y(_02801_));
 AND2x2_ASAP7_75t_R _23513_ (.A(_05303_),
    .B(_08087_),
    .Y(_08193_));
 AO21x1_ASAP7_75t_R _23514_ (.A1(\alu_adder_result_ex[6] ),
    .A2(_08095_),
    .B(_08193_),
    .Y(_08194_));
 NAND2x1_ASAP7_75t_R _23515_ (.A(_00072_),
    .B(_08084_),
    .Y(_08195_));
 OA21x2_ASAP7_75t_R _23516_ (.A1(_08165_),
    .A2(_08194_),
    .B(_08195_),
    .Y(_02802_));
 OR2x2_ASAP7_75t_R _23517_ (.A(_05595_),
    .B(_05350_),
    .Y(_08196_));
 OA21x2_ASAP7_75t_R _23518_ (.A1(\alu_adder_result_ex[7] ),
    .A2(_08087_),
    .B(_08196_),
    .Y(_08197_));
 NAND2x1_ASAP7_75t_R _23519_ (.A(_00071_),
    .B(_08084_),
    .Y(_08198_));
 OA21x2_ASAP7_75t_R _23520_ (.A1(_08165_),
    .A2(_08197_),
    .B(_08198_),
    .Y(_02803_));
 AND2x2_ASAP7_75t_R _23521_ (.A(_15098_),
    .B(_08087_),
    .Y(_08199_));
 AO21x1_ASAP7_75t_R _23522_ (.A1(\alu_adder_result_ex[8] ),
    .A2(_08095_),
    .B(_08199_),
    .Y(_08200_));
 INVx1_ASAP7_75t_R _23523_ (.A(_00074_),
    .Y(_08201_));
 AO21x1_ASAP7_75t_R _23524_ (.A1(_14640_),
    .A2(_08171_),
    .B(_08201_),
    .Y(_08202_));
 OA21x2_ASAP7_75t_R _23525_ (.A1(_08098_),
    .A2(_08200_),
    .B(_08202_),
    .Y(_02804_));
 OR2x2_ASAP7_75t_R _23526_ (.A(_05605_),
    .B(_05350_),
    .Y(_08203_));
 OA21x2_ASAP7_75t_R _23527_ (.A1(\alu_adder_result_ex[9] ),
    .A2(_08087_),
    .B(_08203_),
    .Y(_08204_));
 INVx1_ASAP7_75t_R _23528_ (.A(_00073_),
    .Y(_08205_));
 AO21x1_ASAP7_75t_R _23529_ (.A1(_14640_),
    .A2(_08171_),
    .B(_08205_),
    .Y(_08206_));
 OA21x2_ASAP7_75t_R _23530_ (.A1(_08098_),
    .A2(_08204_),
    .B(_08206_),
    .Y(_02805_));
 INVx1_ASAP7_75t_R _23531_ (.A(_01732_),
    .Y(_08207_));
 MAJx3_ASAP7_75t_R _23532_ (.A(_04959_),
    .B(_08207_),
    .C(net1961),
    .Y(_08208_));
 OR3x1_ASAP7_75t_R _23533_ (.A(_08081_),
    .B(_00025_),
    .C(_08208_),
    .Y(_08209_));
 BUFx6f_ASAP7_75t_R _23534_ (.A(_08209_),
    .Y(_08210_));
 OR3x2_ASAP7_75t_R _23535_ (.A(_05197_),
    .B(_08078_),
    .C(_05205_),
    .Y(_08211_));
 OA21x2_ASAP7_75t_R _23536_ (.A1(_08210_),
    .A2(_08211_),
    .B(_00028_),
    .Y(_08212_));
 AND3x4_ASAP7_75t_R _23537_ (.A(_14640_),
    .B(_05197_),
    .C(_05195_),
    .Y(_08213_));
 BUFx6f_ASAP7_75t_R _23538_ (.A(_08213_),
    .Y(_08214_));
 BUFx12f_ASAP7_75t_R _23539_ (.A(_08214_),
    .Y(_08215_));
 NOR2x1_ASAP7_75t_R _23540_ (.A(_08212_),
    .B(_08215_),
    .Y(_02806_));
 BUFx12f_ASAP7_75t_R _23541_ (.A(_08214_),
    .Y(_08216_));
 OR3x1_ASAP7_75t_R _23542_ (.A(_08081_),
    .B(_00032_),
    .C(_08208_),
    .Y(_08217_));
 BUFx6f_ASAP7_75t_R _23543_ (.A(_08217_),
    .Y(_08218_));
 BUFx6f_ASAP7_75t_R _23544_ (.A(_05197_),
    .Y(_08219_));
 NAND2x2_ASAP7_75t_R _23545_ (.A(_05186_),
    .B(_08073_),
    .Y(_08220_));
 OR3x1_ASAP7_75t_R _23546_ (.A(_08219_),
    .B(_05205_),
    .C(_08220_),
    .Y(_08221_));
 BUFx6f_ASAP7_75t_R _23547_ (.A(_08221_),
    .Y(_08222_));
 OAI22x1_ASAP7_75t_R _23548_ (.A1(_00040_),
    .A2(_08216_),
    .B1(_08218_),
    .B2(_08222_),
    .Y(_02807_));
 BUFx6f_ASAP7_75t_R _23549_ (.A(_08208_),
    .Y(_08223_));
 OR3x1_ASAP7_75t_R _23550_ (.A(_08081_),
    .B(_00024_),
    .C(_08223_),
    .Y(_08224_));
 BUFx6f_ASAP7_75t_R _23551_ (.A(_08224_),
    .Y(_08225_));
 OAI22x1_ASAP7_75t_R _23552_ (.A1(_00041_),
    .A2(_08216_),
    .B1(_08222_),
    .B2(_08225_),
    .Y(_02808_));
 OR2x2_ASAP7_75t_R _23553_ (.A(_05186_),
    .B(_05187_),
    .Y(_08226_));
 BUFx6f_ASAP7_75t_R _23554_ (.A(_08226_),
    .Y(_08227_));
 OR3x1_ASAP7_75t_R _23555_ (.A(_08219_),
    .B(_05205_),
    .C(_08227_),
    .Y(_08228_));
 BUFx6f_ASAP7_75t_R _23556_ (.A(_08228_),
    .Y(_08229_));
 OAI22x1_ASAP7_75t_R _23557_ (.A1(_00042_),
    .A2(_08216_),
    .B1(_08229_),
    .B2(_08210_),
    .Y(_02809_));
 OR3x2_ASAP7_75t_R _23558_ (.A(_01395_),
    .B(_08081_),
    .C(_08223_),
    .Y(_08230_));
 OAI22x1_ASAP7_75t_R _23559_ (.A1(_00043_),
    .A2(_08216_),
    .B1(_08229_),
    .B2(_08230_),
    .Y(_02810_));
 OAI22x1_ASAP7_75t_R _23560_ (.A1(_00044_),
    .A2(_08216_),
    .B1(_08218_),
    .B2(_08229_),
    .Y(_02811_));
 OAI22x1_ASAP7_75t_R _23561_ (.A1(_00045_),
    .A2(_08216_),
    .B1(_08225_),
    .B2(_08229_),
    .Y(_02812_));
 OR3x1_ASAP7_75t_R _23562_ (.A(_01394_),
    .B(_00025_),
    .C(_08208_),
    .Y(_08231_));
 BUFx6f_ASAP7_75t_R _23563_ (.A(_08231_),
    .Y(_08232_));
 OA21x2_ASAP7_75t_R _23564_ (.A1(_08211_),
    .A2(_08232_),
    .B(_00046_),
    .Y(_08233_));
 NOR2x1_ASAP7_75t_R _23565_ (.A(_08215_),
    .B(_08233_),
    .Y(_02813_));
 OR3x1_ASAP7_75t_R _23566_ (.A(_01395_),
    .B(_01394_),
    .C(_08208_),
    .Y(_08234_));
 BUFx6f_ASAP7_75t_R _23567_ (.A(_08234_),
    .Y(_08235_));
 OA21x2_ASAP7_75t_R _23568_ (.A1(_08211_),
    .A2(_08235_),
    .B(_00047_),
    .Y(_08236_));
 NOR2x1_ASAP7_75t_R _23569_ (.A(_08215_),
    .B(_08236_),
    .Y(_02814_));
 OR3x1_ASAP7_75t_R _23570_ (.A(_01394_),
    .B(_00032_),
    .C(_08208_),
    .Y(_08237_));
 BUFx6f_ASAP7_75t_R _23571_ (.A(_08237_),
    .Y(_08238_));
 OA21x2_ASAP7_75t_R _23572_ (.A1(_08211_),
    .A2(_08238_),
    .B(_00048_),
    .Y(_08239_));
 NOR2x1_ASAP7_75t_R _23573_ (.A(_08215_),
    .B(_08239_),
    .Y(_02815_));
 OR3x1_ASAP7_75t_R _23574_ (.A(_01394_),
    .B(_00024_),
    .C(_08208_),
    .Y(_08240_));
 BUFx6f_ASAP7_75t_R _23575_ (.A(_08240_),
    .Y(_08241_));
 OA21x2_ASAP7_75t_R _23576_ (.A1(_08211_),
    .A2(_08241_),
    .B(_00049_),
    .Y(_08242_));
 NOR2x1_ASAP7_75t_R _23577_ (.A(_08215_),
    .B(_08242_),
    .Y(_02816_));
 OR4x1_ASAP7_75t_R _23578_ (.A(_01395_),
    .B(_08081_),
    .C(_08077_),
    .D(_08223_),
    .Y(_08243_));
 OR3x1_ASAP7_75t_R _23579_ (.A(_05198_),
    .B(_05206_),
    .C(_08243_),
    .Y(_08244_));
 OAI21x1_ASAP7_75t_R _23580_ (.A1(_00030_),
    .A2(_08216_),
    .B(_08244_),
    .Y(_02817_));
 OR2x2_ASAP7_75t_R _23581_ (.A(_05186_),
    .B(_08073_),
    .Y(_08245_));
 BUFx6f_ASAP7_75t_R _23582_ (.A(_08245_),
    .Y(_08246_));
 OR3x1_ASAP7_75t_R _23583_ (.A(_08219_),
    .B(_05205_),
    .C(_08246_),
    .Y(_08247_));
 BUFx6f_ASAP7_75t_R _23584_ (.A(_08247_),
    .Y(_08248_));
 OAI22x1_ASAP7_75t_R _23585_ (.A1(_00050_),
    .A2(_08216_),
    .B1(_08232_),
    .B2(_08248_),
    .Y(_02818_));
 OAI22x1_ASAP7_75t_R _23586_ (.A1(_00051_),
    .A2(_08216_),
    .B1(_08235_),
    .B2(_08248_),
    .Y(_02819_));
 OAI22x1_ASAP7_75t_R _23587_ (.A1(_00052_),
    .A2(_08216_),
    .B1(_08238_),
    .B2(_08248_),
    .Y(_02820_));
 BUFx12f_ASAP7_75t_R _23588_ (.A(_08214_),
    .Y(_08249_));
 OAI22x1_ASAP7_75t_R _23589_ (.A1(_00053_),
    .A2(_08249_),
    .B1(_08241_),
    .B2(_08248_),
    .Y(_02821_));
 OAI22x1_ASAP7_75t_R _23590_ (.A1(_00054_),
    .A2(_08249_),
    .B1(_08222_),
    .B2(_08232_),
    .Y(_02822_));
 OAI22x1_ASAP7_75t_R _23591_ (.A1(_00055_),
    .A2(_08249_),
    .B1(_08222_),
    .B2(_08235_),
    .Y(_02823_));
 OAI22x1_ASAP7_75t_R _23592_ (.A1(_00056_),
    .A2(_08249_),
    .B1(_08222_),
    .B2(_08238_),
    .Y(_02824_));
 OAI22x1_ASAP7_75t_R _23593_ (.A1(_00057_),
    .A2(_08249_),
    .B1(_08222_),
    .B2(_08241_),
    .Y(_02825_));
 OAI22x1_ASAP7_75t_R _23594_ (.A1(_00058_),
    .A2(_08249_),
    .B1(_08229_),
    .B2(_08232_),
    .Y(_02826_));
 OAI22x1_ASAP7_75t_R _23595_ (.A1(_00059_),
    .A2(_08249_),
    .B1(_08229_),
    .B2(_08235_),
    .Y(_02827_));
 OA21x2_ASAP7_75t_R _23596_ (.A1(_08211_),
    .A2(_08218_),
    .B(_00031_),
    .Y(_08250_));
 NOR2x1_ASAP7_75t_R _23597_ (.A(_08214_),
    .B(_08250_),
    .Y(_02828_));
 OAI22x1_ASAP7_75t_R _23598_ (.A1(_00060_),
    .A2(_08249_),
    .B1(_08229_),
    .B2(_08238_),
    .Y(_02829_));
 OAI22x1_ASAP7_75t_R _23599_ (.A1(_00061_),
    .A2(_08249_),
    .B1(_08229_),
    .B2(_08241_),
    .Y(_02830_));
 OA21x2_ASAP7_75t_R _23600_ (.A1(_08211_),
    .A2(_08225_),
    .B(_00033_),
    .Y(_08251_));
 NOR2x1_ASAP7_75t_R _23601_ (.A(_08214_),
    .B(_08251_),
    .Y(_02831_));
 OAI22x1_ASAP7_75t_R _23602_ (.A1(_00034_),
    .A2(_08249_),
    .B1(_08248_),
    .B2(_08210_),
    .Y(_02832_));
 OAI22x1_ASAP7_75t_R _23603_ (.A1(_00035_),
    .A2(_08215_),
    .B1(_08230_),
    .B2(_08248_),
    .Y(_02833_));
 OAI22x1_ASAP7_75t_R _23604_ (.A1(_00036_),
    .A2(_08215_),
    .B1(_08218_),
    .B2(_08248_),
    .Y(_02834_));
 OAI22x1_ASAP7_75t_R _23605_ (.A1(_00037_),
    .A2(_08215_),
    .B1(_08225_),
    .B2(_08248_),
    .Y(_02835_));
 OAI22x1_ASAP7_75t_R _23606_ (.A1(_00038_),
    .A2(_08215_),
    .B1(_08222_),
    .B2(_08210_),
    .Y(_02836_));
 OAI22x1_ASAP7_75t_R _23607_ (.A1(_00039_),
    .A2(_08215_),
    .B1(_08222_),
    .B2(_08230_),
    .Y(_02837_));
 INVx1_ASAP7_75t_R _23608_ (.A(net82),
    .Y(_08252_));
 NAND2x1_ASAP7_75t_R _23609_ (.A(_01797_),
    .B(_08252_),
    .Y(_02838_));
 OR2x6_ASAP7_75t_R _23610_ (.A(_13685_),
    .B(_13602_),
    .Y(_08253_));
 BUFx12f_ASAP7_75t_R _23611_ (.A(_08253_),
    .Y(_08254_));
 AND4x1_ASAP7_75t_R _23612_ (.A(_05182_),
    .B(_05178_),
    .C(_01442_),
    .D(_05181_),
    .Y(_08255_));
 INVx3_ASAP7_75t_R _23613_ (.A(_08255_),
    .Y(_08256_));
 AO32x1_ASAP7_75t_R _23614_ (.A1(_13277_),
    .A2(_13220_),
    .A3(_13263_),
    .B1(_14124_),
    .B2(_13296_),
    .Y(_08257_));
 AO21x1_ASAP7_75t_R _23615_ (.A1(_13240_),
    .A2(_08257_),
    .B(_14120_),
    .Y(_08258_));
 NAND2x1_ASAP7_75t_R _23616_ (.A(_06891_),
    .B(_08258_),
    .Y(_08259_));
 OR4x1_ASAP7_75t_R _23617_ (.A(_06904_),
    .B(_06905_),
    .C(_06912_),
    .D(_08259_),
    .Y(_08260_));
 BUFx6f_ASAP7_75t_R _23618_ (.A(_08260_),
    .Y(_08261_));
 OR2x2_ASAP7_75t_R _23619_ (.A(_13455_),
    .B(_13430_),
    .Y(_08262_));
 AO211x2_ASAP7_75t_R _23620_ (.A1(_08256_),
    .A2(_08261_),
    .B(_07799_),
    .C(_08262_),
    .Y(_08263_));
 NOR2x2_ASAP7_75t_R _23621_ (.A(_08254_),
    .B(_08263_),
    .Y(_08264_));
 BUFx12f_ASAP7_75t_R _23622_ (.A(_08264_),
    .Y(_08265_));
 NOR2x1_ASAP7_75t_R _23623_ (.A(_06905_),
    .B(_06912_),
    .Y(_08266_));
 INVx1_ASAP7_75t_R _23624_ (.A(_08259_),
    .Y(_08267_));
 AND3x4_ASAP7_75t_R _23625_ (.A(_05149_),
    .B(_08266_),
    .C(_08267_),
    .Y(_08268_));
 BUFx6f_ASAP7_75t_R _23626_ (.A(_01440_),
    .Y(_08269_));
 BUFx6f_ASAP7_75t_R _23627_ (.A(_08269_),
    .Y(_08270_));
 BUFx6f_ASAP7_75t_R _23628_ (.A(_08270_),
    .Y(_08271_));
 BUFx6f_ASAP7_75t_R _23629_ (.A(_01441_),
    .Y(_08272_));
 BUFx6f_ASAP7_75t_R _23630_ (.A(_08272_),
    .Y(_08273_));
 BUFx6f_ASAP7_75t_R _23631_ (.A(_08273_),
    .Y(_08274_));
 BUFx6f_ASAP7_75t_R _23632_ (.A(_08274_),
    .Y(_08275_));
 BUFx6f_ASAP7_75t_R _23633_ (.A(_08273_),
    .Y(_08276_));
 NAND2x1_ASAP7_75t_R _23634_ (.A(net78),
    .B(_08276_),
    .Y(_08277_));
 OAI21x1_ASAP7_75t_R _23635_ (.A1(_01417_),
    .A2(_08275_),
    .B(_08277_),
    .Y(_08278_));
 BUFx6f_ASAP7_75t_R _23636_ (.A(_08273_),
    .Y(_08279_));
 NAND2x1_ASAP7_75t_R _23637_ (.A(_01432_),
    .B(_08279_),
    .Y(_08280_));
 INVx2_ASAP7_75t_R _23638_ (.A(_08269_),
    .Y(_08281_));
 BUFx6f_ASAP7_75t_R _23639_ (.A(_08281_),
    .Y(_08282_));
 OA211x2_ASAP7_75t_R _23640_ (.A1(net27),
    .A2(_08275_),
    .B(_08280_),
    .C(_08282_),
    .Y(_08283_));
 AOI21x1_ASAP7_75t_R _23641_ (.A1(_08271_),
    .A2(_08278_),
    .B(_08283_),
    .Y(_08284_));
 NAND2x2_ASAP7_75t_R _23642_ (.A(_02191_),
    .B(_02196_),
    .Y(_08285_));
 BUFx6f_ASAP7_75t_R _23643_ (.A(_08285_),
    .Y(_08286_));
 BUFx6f_ASAP7_75t_R _23644_ (.A(_08282_),
    .Y(_08287_));
 INVx3_ASAP7_75t_R _23645_ (.A(_08272_),
    .Y(_08288_));
 BUFx6f_ASAP7_75t_R _23646_ (.A(_08288_),
    .Y(_08289_));
 BUFx6f_ASAP7_75t_R _23647_ (.A(_08289_),
    .Y(_08290_));
 AND2x2_ASAP7_75t_R _23648_ (.A(net64),
    .B(_08274_),
    .Y(_08291_));
 AOI21x1_ASAP7_75t_R _23649_ (.A1(net27),
    .A2(_08290_),
    .B(_08291_),
    .Y(_08292_));
 INVx1_ASAP7_75t_R _23650_ (.A(net55),
    .Y(_08293_));
 BUFx6f_ASAP7_75t_R _23651_ (.A(_08269_),
    .Y(_08294_));
 OA211x2_ASAP7_75t_R _23652_ (.A1(_08293_),
    .A2(_08279_),
    .B(_08277_),
    .C(_08294_),
    .Y(_08295_));
 BUFx6f_ASAP7_75t_R _23653_ (.A(_02191_),
    .Y(_08296_));
 AO211x2_ASAP7_75t_R _23654_ (.A1(_08287_),
    .A2(_08292_),
    .B(_08295_),
    .C(_08296_),
    .Y(_08297_));
 BUFx12f_ASAP7_75t_R _23655_ (.A(_02196_),
    .Y(_08298_));
 OR2x2_ASAP7_75t_R _23656_ (.A(net77),
    .B(_08288_),
    .Y(_08299_));
 OA211x2_ASAP7_75t_R _23657_ (.A1(net54),
    .A2(_08272_),
    .B(_08299_),
    .C(_08269_),
    .Y(_08300_));
 OR2x2_ASAP7_75t_R _23658_ (.A(net63),
    .B(_08288_),
    .Y(_08301_));
 OA211x2_ASAP7_75t_R _23659_ (.A1(net72),
    .A2(_08272_),
    .B(_08301_),
    .C(_08281_),
    .Y(_08302_));
 NOR2x1_ASAP7_75t_R _23660_ (.A(_08300_),
    .B(_08302_),
    .Y(_08303_));
 OR3x2_ASAP7_75t_R _23661_ (.A(_01445_),
    .B(_08298_),
    .C(_08303_),
    .Y(_08304_));
 OA211x2_ASAP7_75t_R _23662_ (.A1(_08284_),
    .A2(_08286_),
    .B(_08297_),
    .C(_08304_),
    .Y(_08305_));
 OA21x2_ASAP7_75t_R _23663_ (.A1(_02291_),
    .A2(_05795_),
    .B(_14591_),
    .Y(_08306_));
 XNOR2x1_ASAP7_75t_R _23664_ (.B(_08306_),
    .Y(_08307_),
    .A(_18575_));
 BUFx6f_ASAP7_75t_R _23665_ (.A(_08307_),
    .Y(_08308_));
 OA31x2_ASAP7_75t_R _23666_ (.A1(_13449_),
    .A2(_18559_),
    .A3(_18563_),
    .B1(_14591_),
    .Y(_08309_));
 XNOR2x1_ASAP7_75t_R _23667_ (.B(_08309_),
    .Y(_08310_),
    .A(_18570_));
 BUFx6f_ASAP7_75t_R _23668_ (.A(_08310_),
    .Y(_08311_));
 BUFx6f_ASAP7_75t_R _23669_ (.A(_08311_),
    .Y(_08312_));
 AND2x4_ASAP7_75t_R _23670_ (.A(_02291_),
    .B(_14591_),
    .Y(_08313_));
 XNOR2x1_ASAP7_75t_R _23671_ (.B(_08313_),
    .Y(_08314_),
    .A(_18565_));
 BUFx6f_ASAP7_75t_R _23672_ (.A(_08314_),
    .Y(_08315_));
 BUFx6f_ASAP7_75t_R _23673_ (.A(_08315_),
    .Y(_08316_));
 NAND2x1_ASAP7_75t_R _23674_ (.A(_00268_),
    .B(_14591_),
    .Y(_08317_));
 OA21x2_ASAP7_75t_R _23675_ (.A1(_14591_),
    .A2(_13543_),
    .B(_08317_),
    .Y(_08318_));
 BUFx6f_ASAP7_75t_R _23676_ (.A(_08318_),
    .Y(_08319_));
 BUFx6f_ASAP7_75t_R _23677_ (.A(_08319_),
    .Y(_08320_));
 OR4x1_ASAP7_75t_R _23678_ (.A(_14544_),
    .B(_14576_),
    .C(_14609_),
    .D(_14610_),
    .Y(_08321_));
 OR3x2_ASAP7_75t_R _23679_ (.A(_01389_),
    .B(_14603_),
    .C(_08321_),
    .Y(_08322_));
 BUFx6f_ASAP7_75t_R _23680_ (.A(_08322_),
    .Y(_08323_));
 INVx1_ASAP7_75t_R _23681_ (.A(_01389_),
    .Y(_08324_));
 AND3x4_ASAP7_75t_R _23682_ (.A(_08324_),
    .B(_14615_),
    .C(_06865_),
    .Y(_08325_));
 BUFx6f_ASAP7_75t_R _23683_ (.A(_08325_),
    .Y(_08326_));
 AND3x1_ASAP7_75t_R _23684_ (.A(_15430_),
    .B(_15432_),
    .C(_08326_),
    .Y(_08327_));
 BUFx6f_ASAP7_75t_R _23685_ (.A(_13449_),
    .Y(_08328_));
 AO211x2_ASAP7_75t_R _23686_ (.A1(_18645_),
    .A2(_08323_),
    .B(_08327_),
    .C(_08328_),
    .Y(_08329_));
 AND3x1_ASAP7_75t_R _23687_ (.A(_13269_),
    .B(_13293_),
    .C(_08326_),
    .Y(_08330_));
 BUFx6f_ASAP7_75t_R _23688_ (.A(_08322_),
    .Y(_08331_));
 AND3x1_ASAP7_75t_R _23689_ (.A(_16191_),
    .B(_16194_),
    .C(_08331_),
    .Y(_08332_));
 OR3x1_ASAP7_75t_R _23690_ (.A(_05829_),
    .B(_08330_),
    .C(_08332_),
    .Y(_08333_));
 AND3x1_ASAP7_75t_R _23691_ (.A(_08320_),
    .B(_08329_),
    .C(_08333_),
    .Y(_08334_));
 OAI21x1_ASAP7_75t_R _23692_ (.A1(_14591_),
    .A2(_18559_),
    .B(_08317_),
    .Y(_08335_));
 BUFx6f_ASAP7_75t_R _23693_ (.A(_08335_),
    .Y(_08336_));
 BUFx6f_ASAP7_75t_R _23694_ (.A(_08336_),
    .Y(_08337_));
 AOI221x1_ASAP7_75t_R _23695_ (.A1(_14446_),
    .A2(_15583_),
    .B1(_15584_),
    .B2(_15585_),
    .C(_08323_),
    .Y(_08338_));
 AND3x1_ASAP7_75t_R _23696_ (.A(_15944_),
    .B(_15946_),
    .C(_08331_),
    .Y(_08339_));
 OR3x1_ASAP7_75t_R _23697_ (.A(_05829_),
    .B(_08338_),
    .C(_08339_),
    .Y(_08340_));
 BUFx6f_ASAP7_75t_R _23698_ (.A(_08325_),
    .Y(_08341_));
 OA211x2_ASAP7_75t_R _23699_ (.A1(_14709_),
    .A2(_15707_),
    .B(_15710_),
    .C(_08341_),
    .Y(_08342_));
 AO211x2_ASAP7_75t_R _23700_ (.A1(_18635_),
    .A2(_08323_),
    .B(_08342_),
    .C(_13450_),
    .Y(_08343_));
 AND3x1_ASAP7_75t_R _23701_ (.A(_08337_),
    .B(_08340_),
    .C(_08343_),
    .Y(_08344_));
 OR3x1_ASAP7_75t_R _23702_ (.A(_08316_),
    .B(_08334_),
    .C(_08344_),
    .Y(_08345_));
 XNOR2x1_ASAP7_75t_R _23703_ (.B(_08313_),
    .Y(_08346_),
    .A(_18563_));
 BUFx6f_ASAP7_75t_R _23704_ (.A(_08346_),
    .Y(_08347_));
 BUFx6f_ASAP7_75t_R _23705_ (.A(_08319_),
    .Y(_08348_));
 BUFx6f_ASAP7_75t_R _23706_ (.A(_08331_),
    .Y(_08349_));
 AND3x1_ASAP7_75t_R _23707_ (.A(_15157_),
    .B(_15160_),
    .C(_08326_),
    .Y(_08350_));
 AO211x2_ASAP7_75t_R _23708_ (.A1(_18665_),
    .A2(_08349_),
    .B(_08350_),
    .C(_08328_),
    .Y(_08351_));
 BUFx6f_ASAP7_75t_R _23709_ (.A(_08326_),
    .Y(_08352_));
 BUFx6f_ASAP7_75t_R _23710_ (.A(_08322_),
    .Y(_08353_));
 AND3x1_ASAP7_75t_R _23711_ (.A(_16697_),
    .B(_16700_),
    .C(_08353_),
    .Y(_08354_));
 AO211x2_ASAP7_75t_R _23712_ (.A1(_18592_),
    .A2(_08352_),
    .B(_08354_),
    .C(_13452_),
    .Y(_08355_));
 AND3x1_ASAP7_75t_R _23713_ (.A(_08348_),
    .B(_08351_),
    .C(_08355_),
    .Y(_08356_));
 BUFx6f_ASAP7_75t_R _23714_ (.A(_08335_),
    .Y(_08357_));
 AND3x1_ASAP7_75t_R _23715_ (.A(_14378_),
    .B(_14387_),
    .C(_08326_),
    .Y(_08358_));
 AND3x1_ASAP7_75t_R _23716_ (.A(_16326_),
    .B(_16328_),
    .C(_08331_),
    .Y(_08359_));
 OR3x1_ASAP7_75t_R _23717_ (.A(_13450_),
    .B(_08358_),
    .C(_08359_),
    .Y(_08360_));
 AND3x1_ASAP7_75t_R _23718_ (.A(_15228_),
    .B(_15230_),
    .C(_08341_),
    .Y(_08361_));
 AND3x1_ASAP7_75t_R _23719_ (.A(_16449_),
    .B(_16451_),
    .C(_08331_),
    .Y(_08362_));
 OR3x1_ASAP7_75t_R _23720_ (.A(_05829_),
    .B(_08361_),
    .C(_08362_),
    .Y(_08363_));
 AND3x1_ASAP7_75t_R _23721_ (.A(_08357_),
    .B(_08360_),
    .C(_08363_),
    .Y(_08364_));
 OR3x1_ASAP7_75t_R _23722_ (.A(_08347_),
    .B(_08356_),
    .C(_08364_),
    .Y(_08365_));
 AND3x1_ASAP7_75t_R _23723_ (.A(_08312_),
    .B(_08345_),
    .C(_08365_),
    .Y(_08366_));
 XNOR2x1_ASAP7_75t_R _23724_ (.B(_08309_),
    .Y(_08367_),
    .A(_18568_));
 BUFx6f_ASAP7_75t_R _23725_ (.A(_08367_),
    .Y(_08368_));
 AND3x1_ASAP7_75t_R _23726_ (.A(_15944_),
    .B(_15946_),
    .C(_08341_),
    .Y(_08369_));
 AO21x2_ASAP7_75t_R _23727_ (.A1(_18625_),
    .A2(_08323_),
    .B(_08369_),
    .Y(_08370_));
 BUFx6f_ASAP7_75t_R _23728_ (.A(_08341_),
    .Y(_08371_));
 OA211x2_ASAP7_75t_R _23729_ (.A1(_14709_),
    .A2(_15707_),
    .B(_15710_),
    .C(_08353_),
    .Y(_08372_));
 AO211x2_ASAP7_75t_R _23730_ (.A1(_18635_),
    .A2(_08371_),
    .B(_08372_),
    .C(_05829_),
    .Y(_08373_));
 OA21x2_ASAP7_75t_R _23731_ (.A1(_18555_),
    .A2(_08370_),
    .B(_08373_),
    .Y(_08374_));
 AND3x1_ASAP7_75t_R _23732_ (.A(_16191_),
    .B(_16194_),
    .C(_08341_),
    .Y(_08375_));
 AND3x1_ASAP7_75t_R _23733_ (.A(_13269_),
    .B(_13293_),
    .C(_08331_),
    .Y(_08376_));
 OR3x1_ASAP7_75t_R _23734_ (.A(_13450_),
    .B(_08375_),
    .C(_08376_),
    .Y(_08377_));
 AND3x1_ASAP7_75t_R _23735_ (.A(_15430_),
    .B(_15432_),
    .C(_08331_),
    .Y(_08378_));
 AO211x2_ASAP7_75t_R _23736_ (.A1(_18645_),
    .A2(_08371_),
    .B(_08378_),
    .C(_05829_),
    .Y(_08379_));
 AND3x1_ASAP7_75t_R _23737_ (.A(_08357_),
    .B(_08377_),
    .C(_08379_),
    .Y(_08380_));
 AO21x1_ASAP7_75t_R _23738_ (.A1(_08320_),
    .A2(_08374_),
    .B(_08380_),
    .Y(_08381_));
 AND3x1_ASAP7_75t_R _23739_ (.A(_16449_),
    .B(_16451_),
    .C(_08341_),
    .Y(_08382_));
 AND3x1_ASAP7_75t_R _23740_ (.A(_15228_),
    .B(_15230_),
    .C(_08353_),
    .Y(_08383_));
 OR3x1_ASAP7_75t_R _23741_ (.A(_13450_),
    .B(_08382_),
    .C(_08383_),
    .Y(_08384_));
 AND3x1_ASAP7_75t_R _23742_ (.A(_16326_),
    .B(_16328_),
    .C(_08341_),
    .Y(_08385_));
 AND3x1_ASAP7_75t_R _23743_ (.A(_14378_),
    .B(_14387_),
    .C(_08353_),
    .Y(_08386_));
 OR3x1_ASAP7_75t_R _23744_ (.A(_05829_),
    .B(_08385_),
    .C(_08386_),
    .Y(_08387_));
 AND3x1_ASAP7_75t_R _23745_ (.A(_08348_),
    .B(_08384_),
    .C(_08387_),
    .Y(_08388_));
 AND3x1_ASAP7_75t_R _23746_ (.A(_16697_),
    .B(_16700_),
    .C(_08326_),
    .Y(_08389_));
 AO21x1_ASAP7_75t_R _23747_ (.A1(_18592_),
    .A2(_08323_),
    .B(_08389_),
    .Y(_08390_));
 AND3x1_ASAP7_75t_R _23748_ (.A(_15157_),
    .B(_15160_),
    .C(_08353_),
    .Y(_08391_));
 AO211x2_ASAP7_75t_R _23749_ (.A1(_18665_),
    .A2(_08371_),
    .B(_08391_),
    .C(_05829_),
    .Y(_08392_));
 OA211x2_ASAP7_75t_R _23750_ (.A1(_18555_),
    .A2(_08390_),
    .B(_08392_),
    .C(_08336_),
    .Y(_08393_));
 OR3x1_ASAP7_75t_R _23751_ (.A(_08315_),
    .B(_08388_),
    .C(_08393_),
    .Y(_08394_));
 OA21x2_ASAP7_75t_R _23752_ (.A1(_08347_),
    .A2(_08381_),
    .B(_08394_),
    .Y(_08395_));
 AND2x2_ASAP7_75t_R _23753_ (.A(_08368_),
    .B(_08395_),
    .Y(_08396_));
 OR3x1_ASAP7_75t_R _23754_ (.A(_08308_),
    .B(_08366_),
    .C(_08396_),
    .Y(_08397_));
 AND3x1_ASAP7_75t_R _23755_ (.A(_14965_),
    .B(_14970_),
    .C(_08325_),
    .Y(_08398_));
 OA211x2_ASAP7_75t_R _23756_ (.A1(_14709_),
    .A2(_16931_),
    .B(_16933_),
    .C(_08353_),
    .Y(_08399_));
 OR2x2_ASAP7_75t_R _23757_ (.A(_08398_),
    .B(_08399_),
    .Y(_08400_));
 AND3x4_ASAP7_75t_R _23758_ (.A(_04418_),
    .B(_04421_),
    .C(_08353_),
    .Y(_08401_));
 AO211x2_ASAP7_75t_R _23759_ (.A1(_18572_),
    .A2(_08371_),
    .B(_08335_),
    .C(_08401_),
    .Y(_08402_));
 OA21x2_ASAP7_75t_R _23760_ (.A1(_08348_),
    .A2(_08400_),
    .B(_08402_),
    .Y(_08403_));
 AND3x1_ASAP7_75t_R _23761_ (.A(_14899_),
    .B(_14902_),
    .C(_08341_),
    .Y(_08404_));
 AO21x1_ASAP7_75t_R _23762_ (.A1(_18685_),
    .A2(_08323_),
    .B(_08404_),
    .Y(_08405_));
 AND3x1_ASAP7_75t_R _23763_ (.A(_15024_),
    .B(_15026_),
    .C(_08341_),
    .Y(_08406_));
 AND3x1_ASAP7_75t_R _23764_ (.A(_16820_),
    .B(_16822_),
    .C(_08353_),
    .Y(_08407_));
 OR3x1_ASAP7_75t_R _23765_ (.A(_08319_),
    .B(_08406_),
    .C(_08407_),
    .Y(_08408_));
 BUFx6f_ASAP7_75t_R _23766_ (.A(_13451_),
    .Y(_08409_));
 OA211x2_ASAP7_75t_R _23767_ (.A1(_08357_),
    .A2(_08405_),
    .B(_08408_),
    .C(_08409_),
    .Y(_08410_));
 AO21x1_ASAP7_75t_R _23768_ (.A1(_18555_),
    .A2(_08403_),
    .B(_08410_),
    .Y(_08411_));
 AND3x1_ASAP7_75t_R _23769_ (.A(_04788_),
    .B(_04790_),
    .C(_08353_),
    .Y(_08412_));
 AO21x2_ASAP7_75t_R _23770_ (.A1(_18558_),
    .A2(_08371_),
    .B(_08412_),
    .Y(_08413_));
 OA211x2_ASAP7_75t_R _23771_ (.A1(_14709_),
    .A2(_14770_),
    .B(_14775_),
    .C(_08325_),
    .Y(_08414_));
 OA211x2_ASAP7_75t_R _23772_ (.A1(_14709_),
    .A2(_04554_),
    .B(_04556_),
    .C(_08322_),
    .Y(_08415_));
 OR3x1_ASAP7_75t_R _23773_ (.A(_08319_),
    .B(_08414_),
    .C(_08415_),
    .Y(_08416_));
 OA211x2_ASAP7_75t_R _23774_ (.A1(_08357_),
    .A2(_08413_),
    .B(_08416_),
    .C(_13453_),
    .Y(_08417_));
 AND3x4_ASAP7_75t_R _23775_ (.A(_14390_),
    .B(_14444_),
    .C(_08325_),
    .Y(_08418_));
 AND2x6_ASAP7_75t_R _23776_ (.A(_18072_),
    .B(_08322_),
    .Y(_08419_));
 OR2x6_ASAP7_75t_R _23777_ (.A(_08418_),
    .B(_08419_),
    .Y(_08420_));
 AND3x4_ASAP7_75t_R _23778_ (.A(_04666_),
    .B(_04669_),
    .C(_08353_),
    .Y(_08421_));
 AO211x2_ASAP7_75t_R _23779_ (.A1(_18562_),
    .A2(_08371_),
    .B(_08319_),
    .C(_08421_),
    .Y(_08422_));
 OA211x2_ASAP7_75t_R _23780_ (.A1(_08357_),
    .A2(_08420_),
    .B(_08422_),
    .C(_05930_),
    .Y(_08423_));
 OR3x1_ASAP7_75t_R _23781_ (.A(_08347_),
    .B(_08417_),
    .C(_08423_),
    .Y(_08424_));
 OA21x2_ASAP7_75t_R _23782_ (.A1(_08316_),
    .A2(_08411_),
    .B(_08424_),
    .Y(_08425_));
 NAND2x1_ASAP7_75t_R _23783_ (.A(_08307_),
    .B(_08367_),
    .Y(_08426_));
 XNOR2x1_ASAP7_75t_R _23784_ (.B(_08306_),
    .Y(_08427_),
    .A(_18573_));
 AND2x6_ASAP7_75t_R _23785_ (.A(_06865_),
    .B(_06880_),
    .Y(_08428_));
 OA21x2_ASAP7_75t_R _23786_ (.A1(_08418_),
    .A2(_08419_),
    .B(_08428_),
    .Y(_08429_));
 BUFx6f_ASAP7_75t_R _23787_ (.A(_08429_),
    .Y(_08430_));
 OR3x1_ASAP7_75t_R _23788_ (.A(_08427_),
    .B(_08368_),
    .C(_08430_),
    .Y(_08431_));
 OA21x2_ASAP7_75t_R _23789_ (.A1(_08425_),
    .A2(_08426_),
    .B(_08431_),
    .Y(_08432_));
 NAND2x1_ASAP7_75t_R _23790_ (.A(_08397_),
    .B(_08432_),
    .Y(_08433_));
 BUFx6f_ASAP7_75t_R _23791_ (.A(_08349_),
    .Y(_08434_));
 AND2x2_ASAP7_75t_R _23792_ (.A(_02222_),
    .B(net1974),
    .Y(_08435_));
 AOI211x1_ASAP7_75t_R _23793_ (.A1(_06858_),
    .A2(_08435_),
    .B(_08321_),
    .C(_14603_),
    .Y(_08436_));
 BUFx6f_ASAP7_75t_R _23794_ (.A(_08436_),
    .Y(_08437_));
 NAND2x1_ASAP7_75t_R _23795_ (.A(_08434_),
    .B(_08437_),
    .Y(_08438_));
 BUFx6f_ASAP7_75t_R _23796_ (.A(_08352_),
    .Y(_08439_));
 BUFx6f_ASAP7_75t_R _23797_ (.A(_08439_),
    .Y(_08440_));
 AO211x2_ASAP7_75t_R _23798_ (.A1(_18592_),
    .A2(_08371_),
    .B(_08354_),
    .C(_13450_),
    .Y(_08441_));
 OR3x1_ASAP7_75t_R _23799_ (.A(_05829_),
    .B(_08406_),
    .C(_08407_),
    .Y(_08442_));
 AND3x1_ASAP7_75t_R _23800_ (.A(_08336_),
    .B(_08441_),
    .C(_08442_),
    .Y(_08443_));
 OR3x1_ASAP7_75t_R _23801_ (.A(_13450_),
    .B(_08398_),
    .C(_08399_),
    .Y(_08444_));
 BUFx6f_ASAP7_75t_R _23802_ (.A(_08319_),
    .Y(_08445_));
 OA211x2_ASAP7_75t_R _23803_ (.A1(_08409_),
    .A2(_08405_),
    .B(_08444_),
    .C(_08445_),
    .Y(_08446_));
 OR3x1_ASAP7_75t_R _23804_ (.A(_08314_),
    .B(_08443_),
    .C(_08446_),
    .Y(_08447_));
 BUFx6f_ASAP7_75t_R _23805_ (.A(_08346_),
    .Y(_08448_));
 AO211x2_ASAP7_75t_R _23806_ (.A1(_18562_),
    .A2(_08371_),
    .B(_08335_),
    .C(_08421_),
    .Y(_08449_));
 AO211x2_ASAP7_75t_R _23807_ (.A1(_18572_),
    .A2(_08371_),
    .B(_08319_),
    .C(_08401_),
    .Y(_08450_));
 AND3x1_ASAP7_75t_R _23808_ (.A(_08409_),
    .B(_08449_),
    .C(_08450_),
    .Y(_08451_));
 OA211x2_ASAP7_75t_R _23809_ (.A1(_08336_),
    .A2(_08413_),
    .B(_08416_),
    .C(_05930_),
    .Y(_08452_));
 OR3x1_ASAP7_75t_R _23810_ (.A(_08448_),
    .B(_08451_),
    .C(_08452_),
    .Y(_08453_));
 AND2x4_ASAP7_75t_R _23811_ (.A(_08447_),
    .B(_08453_),
    .Y(_08454_));
 AND2x2_ASAP7_75t_R _23812_ (.A(_08427_),
    .B(_08367_),
    .Y(_08455_));
 BUFx6f_ASAP7_75t_R _23813_ (.A(_08455_),
    .Y(_08456_));
 INVx1_ASAP7_75t_R _23814_ (.A(_08456_),
    .Y(_08457_));
 NAND2x2_ASAP7_75t_R _23815_ (.A(_08420_),
    .B(_08428_),
    .Y(_08458_));
 NAND2x1_ASAP7_75t_R _23816_ (.A(_08307_),
    .B(_08458_),
    .Y(_08459_));
 BUFx6f_ASAP7_75t_R _23817_ (.A(_08459_),
    .Y(_08460_));
 OA211x2_ASAP7_75t_R _23818_ (.A1(_08418_),
    .A2(_08419_),
    .B(_13452_),
    .C(_08335_),
    .Y(_08461_));
 AND2x2_ASAP7_75t_R _23819_ (.A(_08448_),
    .B(_08461_),
    .Y(_08462_));
 OR3x1_ASAP7_75t_R _23820_ (.A(_08367_),
    .B(_08430_),
    .C(_08462_),
    .Y(_08463_));
 OA211x2_ASAP7_75t_R _23821_ (.A1(_08454_),
    .A2(_08457_),
    .B(_08460_),
    .C(_08463_),
    .Y(_08464_));
 NAND2x1_ASAP7_75t_R _23822_ (.A(_08440_),
    .B(_08464_),
    .Y(_08465_));
 INVx1_ASAP7_75t_R _23823_ (.A(_08436_),
    .Y(_08466_));
 AOI21x1_ASAP7_75t_R _23824_ (.A1(net1975),
    .A2(_02222_),
    .B(_08321_),
    .Y(_08467_));
 NAND2x2_ASAP7_75t_R _23825_ (.A(_14604_),
    .B(_08467_),
    .Y(_08468_));
 INVx1_ASAP7_75t_R _23826_ (.A(_06880_),
    .Y(_08469_));
 AO21x1_ASAP7_75t_R _23827_ (.A1(net1974),
    .A2(_06858_),
    .B(_06860_),
    .Y(_08470_));
 AO21x1_ASAP7_75t_R _23828_ (.A1(_08469_),
    .A2(_08470_),
    .B(_06855_),
    .Y(_08471_));
 NOR2x1_ASAP7_75t_R _23829_ (.A(net1975),
    .B(_06860_),
    .Y(_08472_));
 AND3x1_ASAP7_75t_R _23830_ (.A(_08324_),
    .B(_06860_),
    .C(_14603_),
    .Y(_08473_));
 OA21x2_ASAP7_75t_R _23831_ (.A1(_08472_),
    .A2(_08473_),
    .B(_06865_),
    .Y(_08474_));
 OR3x2_ASAP7_75t_R _23832_ (.A(_06860_),
    .B(_08321_),
    .C(_08435_),
    .Y(_08475_));
 OA21x2_ASAP7_75t_R _23833_ (.A1(_01389_),
    .A2(_06860_),
    .B(_06872_),
    .Y(_08476_));
 OR2x2_ASAP7_75t_R _23834_ (.A(_08321_),
    .B(_08476_),
    .Y(_08477_));
 BUFx6f_ASAP7_75t_R _23835_ (.A(_08477_),
    .Y(_08478_));
 NAND2x1_ASAP7_75t_R _23836_ (.A(_08475_),
    .B(_08478_),
    .Y(_08479_));
 NOR2x1_ASAP7_75t_R _23837_ (.A(_08474_),
    .B(_08479_),
    .Y(_08480_));
 AND5x1_ASAP7_75t_R _23838_ (.A(_06874_),
    .B(_08466_),
    .C(_08468_),
    .D(_08471_),
    .E(_08480_),
    .Y(_08481_));
 OR2x6_ASAP7_75t_R _23839_ (.A(_15234_),
    .B(_08481_),
    .Y(_08482_));
 BUFx6f_ASAP7_75t_R _23840_ (.A(_08482_),
    .Y(_08483_));
 BUFx6f_ASAP7_75t_R _23841_ (.A(_08468_),
    .Y(_08484_));
 BUFx6f_ASAP7_75t_R _23842_ (.A(_08475_),
    .Y(_08485_));
 BUFx6f_ASAP7_75t_R _23843_ (.A(_08478_),
    .Y(_08486_));
 INVx1_ASAP7_75t_R _23844_ (.A(_02301_),
    .Y(_08487_));
 NAND3x1_ASAP7_75t_R _23845_ (.A(_08474_),
    .B(_08475_),
    .C(_08478_),
    .Y(_08488_));
 BUFx6f_ASAP7_75t_R _23846_ (.A(_08488_),
    .Y(_08489_));
 OA222x2_ASAP7_75t_R _23847_ (.A1(_00285_),
    .A2(_08485_),
    .B1(_08486_),
    .B2(_08487_),
    .C1(_08489_),
    .C2(_00284_),
    .Y(_08490_));
 OA21x2_ASAP7_75t_R _23848_ (.A1(_15179_),
    .A2(_08484_),
    .B(_08490_),
    .Y(_08491_));
 AND2x2_ASAP7_75t_R _23849_ (.A(_13262_),
    .B(_00135_),
    .Y(_08492_));
 AND2x2_ASAP7_75t_R _23850_ (.A(_14119_),
    .B(_14623_),
    .Y(_08493_));
 NAND2x1_ASAP7_75t_R _23851_ (.A(_05237_),
    .B(_02197_),
    .Y(_08494_));
 NOR2x2_ASAP7_75t_R _23852_ (.A(_08493_),
    .B(_08494_),
    .Y(_08495_));
 XOR2x1_ASAP7_75t_R _23853_ (.A(_00142_),
    .Y(_08496_),
    .B(_00174_));
 AO21x1_ASAP7_75t_R _23854_ (.A1(_14119_),
    .A2(_15234_),
    .B(_08494_),
    .Y(_08497_));
 BUFx6f_ASAP7_75t_R _23855_ (.A(_08497_),
    .Y(_08498_));
 OR2x2_ASAP7_75t_R _23856_ (.A(_00135_),
    .B(_08498_),
    .Y(_08499_));
 OA211x2_ASAP7_75t_R _23857_ (.A1(_08495_),
    .A2(_08496_),
    .B(_08499_),
    .C(_14533_),
    .Y(_08500_));
 OR3x1_ASAP7_75t_R _23858_ (.A(_14626_),
    .B(_08492_),
    .C(_08500_),
    .Y(_08501_));
 OA211x2_ASAP7_75t_R _23859_ (.A1(_08483_),
    .A2(_08491_),
    .B(_08501_),
    .C(_14388_),
    .Y(_08502_));
 OA211x2_ASAP7_75t_R _23860_ (.A1(_08433_),
    .A2(_08438_),
    .B(_08465_),
    .C(_08502_),
    .Y(_08503_));
 BUFx6f_ASAP7_75t_R _23861_ (.A(_08261_),
    .Y(_08504_));
 AO21x1_ASAP7_75t_R _23862_ (.A1(_14120_),
    .A2(_06674_),
    .B(_08504_),
    .Y(_08505_));
 OAI22x1_ASAP7_75t_R _23863_ (.A1(_08268_),
    .A2(_08305_),
    .B1(_08503_),
    .B2(_08505_),
    .Y(_08506_));
 OR2x6_ASAP7_75t_R _23864_ (.A(_08254_),
    .B(_08263_),
    .Y(_08507_));
 BUFx12f_ASAP7_75t_R _23865_ (.A(_08507_),
    .Y(_08508_));
 BUFx12f_ASAP7_75t_R _23866_ (.A(_08508_),
    .Y(_08509_));
 AND2x2_ASAP7_75t_R _23867_ (.A(_13981_),
    .B(_08509_),
    .Y(_08510_));
 AO21x1_ASAP7_75t_R _23868_ (.A1(_08265_),
    .A2(_08506_),
    .B(_08510_),
    .Y(_02839_));
 AND2x6_ASAP7_75t_R _23869_ (.A(_08349_),
    .B(_08436_),
    .Y(_08511_));
 BUFx6f_ASAP7_75t_R _23870_ (.A(_08511_),
    .Y(_08512_));
 BUFx6f_ASAP7_75t_R _23871_ (.A(_08427_),
    .Y(_08513_));
 BUFx6f_ASAP7_75t_R _23872_ (.A(_08448_),
    .Y(_08514_));
 AO21x1_ASAP7_75t_R _23873_ (.A1(_18665_),
    .A2(_08352_),
    .B(_08391_),
    .Y(_08515_));
 OR3x1_ASAP7_75t_R _23874_ (.A(_08409_),
    .B(_08382_),
    .C(_08383_),
    .Y(_08516_));
 OA21x2_ASAP7_75t_R _23875_ (.A1(_18555_),
    .A2(_08515_),
    .B(_08516_),
    .Y(_08517_));
 OR3x1_ASAP7_75t_R _23876_ (.A(_05930_),
    .B(_08385_),
    .C(_08386_),
    .Y(_08518_));
 OR3x1_ASAP7_75t_R _23877_ (.A(_08409_),
    .B(_08375_),
    .C(_08376_),
    .Y(_08519_));
 AND3x1_ASAP7_75t_R _23878_ (.A(_08320_),
    .B(_08518_),
    .C(_08519_),
    .Y(_08520_));
 AOI21x1_ASAP7_75t_R _23879_ (.A1(_08337_),
    .A2(_08517_),
    .B(_08520_),
    .Y(_08521_));
 AO211x2_ASAP7_75t_R _23880_ (.A1(_18645_),
    .A2(_08352_),
    .B(_08378_),
    .C(_08328_),
    .Y(_08522_));
 OAI21x1_ASAP7_75t_R _23881_ (.A1(_13453_),
    .A2(_08370_),
    .B(_08522_),
    .Y(_08523_));
 XNOR2x2_ASAP7_75t_R _23882_ (.A(_13451_),
    .B(_08326_),
    .Y(_08524_));
 NOR2x1_ASAP7_75t_R _23883_ (.A(_18628_),
    .B(_08524_),
    .Y(_08525_));
 AND2x2_ASAP7_75t_R _23884_ (.A(_18635_),
    .B(_08524_),
    .Y(_08526_));
 OAI21x1_ASAP7_75t_R _23885_ (.A1(_08525_),
    .A2(_08526_),
    .B(_08320_),
    .Y(_08527_));
 BUFx6f_ASAP7_75t_R _23886_ (.A(_08314_),
    .Y(_08528_));
 OA211x2_ASAP7_75t_R _23887_ (.A1(_08320_),
    .A2(_08523_),
    .B(_08527_),
    .C(_08528_),
    .Y(_08529_));
 AOI21x1_ASAP7_75t_R _23888_ (.A1(_08514_),
    .A2(_08521_),
    .B(_08529_),
    .Y(_08530_));
 OA211x2_ASAP7_75t_R _23889_ (.A1(_08445_),
    .A2(_08400_),
    .B(_08402_),
    .C(_08409_),
    .Y(_08531_));
 OR3x1_ASAP7_75t_R _23890_ (.A(_08335_),
    .B(_08414_),
    .C(_08415_),
    .Y(_08532_));
 AO211x2_ASAP7_75t_R _23891_ (.A1(_18685_),
    .A2(_08323_),
    .B(_08319_),
    .C(_08404_),
    .Y(_08533_));
 AND3x1_ASAP7_75t_R _23892_ (.A(_05930_),
    .B(_08532_),
    .C(_08533_),
    .Y(_08534_));
 AND2x4_ASAP7_75t_R _23893_ (.A(_08445_),
    .B(_08430_),
    .Y(_08535_));
 OA211x2_ASAP7_75t_R _23894_ (.A1(_08336_),
    .A2(_08420_),
    .B(_08422_),
    .C(_08409_),
    .Y(_08536_));
 AND2x2_ASAP7_75t_R _23895_ (.A(_13450_),
    .B(_08335_),
    .Y(_08537_));
 AO21x1_ASAP7_75t_R _23896_ (.A1(_08413_),
    .A2(_08537_),
    .B(_08346_),
    .Y(_08538_));
 OA33x2_ASAP7_75t_R _23897_ (.A1(_08315_),
    .A2(_08531_),
    .A3(_08534_),
    .B1(_08535_),
    .B2(_08536_),
    .B3(_08538_),
    .Y(_08539_));
 AND2x2_ASAP7_75t_R _23898_ (.A(_08307_),
    .B(_08539_),
    .Y(_08540_));
 AO211x2_ASAP7_75t_R _23899_ (.A1(_08513_),
    .A2(_08530_),
    .B(_08540_),
    .C(_08312_),
    .Y(_08541_));
 OR3x1_ASAP7_75t_R _23900_ (.A(_08328_),
    .B(_08330_),
    .C(_08332_),
    .Y(_08542_));
 OR3x1_ASAP7_75t_R _23901_ (.A(_13452_),
    .B(_08358_),
    .C(_08359_),
    .Y(_08543_));
 AND3x1_ASAP7_75t_R _23902_ (.A(_08348_),
    .B(_08542_),
    .C(_08543_),
    .Y(_08544_));
 OR3x1_ASAP7_75t_R _23903_ (.A(_08328_),
    .B(_08338_),
    .C(_08339_),
    .Y(_08545_));
 AO211x2_ASAP7_75t_R _23904_ (.A1(_18645_),
    .A2(_08349_),
    .B(_08327_),
    .C(_13452_),
    .Y(_08546_));
 AND3x1_ASAP7_75t_R _23905_ (.A(_08357_),
    .B(_08545_),
    .C(_08546_),
    .Y(_08547_));
 OR3x1_ASAP7_75t_R _23906_ (.A(_08315_),
    .B(_08544_),
    .C(_08547_),
    .Y(_08548_));
 AND3x1_ASAP7_75t_R _23907_ (.A(_08445_),
    .B(_08441_),
    .C(_08442_),
    .Y(_08549_));
 OR3x1_ASAP7_75t_R _23908_ (.A(_13450_),
    .B(_08361_),
    .C(_08362_),
    .Y(_08550_));
 AO211x2_ASAP7_75t_R _23909_ (.A1(_18665_),
    .A2(_08323_),
    .B(_08350_),
    .C(_13452_),
    .Y(_08551_));
 AND3x1_ASAP7_75t_R _23910_ (.A(_08336_),
    .B(_08550_),
    .C(_08551_),
    .Y(_08552_));
 OR3x1_ASAP7_75t_R _23911_ (.A(_08448_),
    .B(_08549_),
    .C(_08552_),
    .Y(_08553_));
 AO21x1_ASAP7_75t_R _23912_ (.A1(_08548_),
    .A2(_08553_),
    .B(_08308_),
    .Y(_08554_));
 BUFx6f_ASAP7_75t_R _23913_ (.A(_08368_),
    .Y(_08555_));
 AO21x1_ASAP7_75t_R _23914_ (.A1(_08460_),
    .A2(_08554_),
    .B(_08555_),
    .Y(_08556_));
 AND2x2_ASAP7_75t_R _23915_ (.A(_08541_),
    .B(_08556_),
    .Y(_08557_));
 BUFx6f_ASAP7_75t_R _23916_ (.A(_08489_),
    .Y(_08558_));
 BUFx6f_ASAP7_75t_R _23917_ (.A(_08475_),
    .Y(_08559_));
 INVx1_ASAP7_75t_R _23918_ (.A(_02302_),
    .Y(_08560_));
 OA222x2_ASAP7_75t_R _23919_ (.A1(_00287_),
    .A2(_08559_),
    .B1(_08486_),
    .B2(_08560_),
    .C1(_15166_),
    .C2(_08484_),
    .Y(_08561_));
 OA21x2_ASAP7_75t_R _23920_ (.A1(_00286_),
    .A2(_08558_),
    .B(_08561_),
    .Y(_08562_));
 OA21x2_ASAP7_75t_R _23921_ (.A1(_00134_),
    .A2(_17089_),
    .B(_00143_),
    .Y(_08563_));
 OA21x2_ASAP7_75t_R _23922_ (.A1(_00142_),
    .A2(_08563_),
    .B(_00151_),
    .Y(_08564_));
 XNOR2x1_ASAP7_75t_R _23923_ (.B(_08564_),
    .Y(_08565_),
    .A(_00150_));
 NAND2x1_ASAP7_75t_R _23924_ (.A(_05240_),
    .B(_08498_),
    .Y(_08566_));
 BUFx6f_ASAP7_75t_R _23925_ (.A(_08566_),
    .Y(_08567_));
 BUFx6f_ASAP7_75t_R _23926_ (.A(_14620_),
    .Y(_08568_));
 AO21x2_ASAP7_75t_R _23927_ (.A1(_14533_),
    .A2(_08498_),
    .B(_08568_),
    .Y(_08569_));
 BUFx6f_ASAP7_75t_R _23928_ (.A(_08569_),
    .Y(_08570_));
 OA22x2_ASAP7_75t_R _23929_ (.A1(_08565_),
    .A2(_08567_),
    .B1(_08570_),
    .B2(_00144_),
    .Y(_08571_));
 OA21x2_ASAP7_75t_R _23930_ (.A1(_08483_),
    .A2(_08562_),
    .B(_08571_),
    .Y(_08572_));
 NAND2x1_ASAP7_75t_R _23931_ (.A(_06698_),
    .B(_08572_),
    .Y(_08573_));
 AO21x1_ASAP7_75t_R _23932_ (.A1(_08512_),
    .A2(_08557_),
    .B(_08573_),
    .Y(_08574_));
 AND3x1_ASAP7_75t_R _23933_ (.A(_08409_),
    .B(_08532_),
    .C(_08533_),
    .Y(_08575_));
 AND3x1_ASAP7_75t_R _23934_ (.A(_05930_),
    .B(_08449_),
    .C(_08450_),
    .Y(_08576_));
 OR2x2_ASAP7_75t_R _23935_ (.A(_08575_),
    .B(_08576_),
    .Y(_08577_));
 AND3x1_ASAP7_75t_R _23936_ (.A(_08357_),
    .B(_08351_),
    .C(_08355_),
    .Y(_08578_));
 OR3x1_ASAP7_75t_R _23937_ (.A(_08328_),
    .B(_08406_),
    .C(_08407_),
    .Y(_08579_));
 OA211x2_ASAP7_75t_R _23938_ (.A1(_13453_),
    .A2(_08400_),
    .B(_08579_),
    .C(_08445_),
    .Y(_08580_));
 OR3x1_ASAP7_75t_R _23939_ (.A(_08315_),
    .B(_08578_),
    .C(_08580_),
    .Y(_08581_));
 OA21x2_ASAP7_75t_R _23940_ (.A1(_08514_),
    .A2(_08577_),
    .B(_08581_),
    .Y(_08582_));
 OR3x1_ASAP7_75t_R _23941_ (.A(_13451_),
    .B(_08418_),
    .C(_08419_),
    .Y(_08583_));
 OA211x2_ASAP7_75t_R _23942_ (.A1(_05930_),
    .A2(_08413_),
    .B(_08583_),
    .C(_08336_),
    .Y(_08584_));
 OR2x2_ASAP7_75t_R _23943_ (.A(_08535_),
    .B(_08584_),
    .Y(_08585_));
 OR2x2_ASAP7_75t_R _23944_ (.A(_08346_),
    .B(_08430_),
    .Y(_08586_));
 OA211x2_ASAP7_75t_R _23945_ (.A1(_08316_),
    .A2(_08585_),
    .B(_08586_),
    .C(_08311_),
    .Y(_08587_));
 AO21x2_ASAP7_75t_R _23946_ (.A1(_08368_),
    .A2(_08582_),
    .B(_08587_),
    .Y(_08588_));
 OR2x2_ASAP7_75t_R _23947_ (.A(_08308_),
    .B(_08588_),
    .Y(_08589_));
 AND2x4_ASAP7_75t_R _23948_ (.A(_08439_),
    .B(_08460_),
    .Y(_08590_));
 OR4x1_ASAP7_75t_R _23949_ (.A(_06904_),
    .B(_07157_),
    .C(_06905_),
    .D(_08259_),
    .Y(_08591_));
 BUFx6f_ASAP7_75t_R _23950_ (.A(_08591_),
    .Y(_08592_));
 BUFx6f_ASAP7_75t_R _23951_ (.A(_08592_),
    .Y(_08593_));
 AO21x1_ASAP7_75t_R _23952_ (.A1(_08589_),
    .A2(_08590_),
    .B(_08593_),
    .Y(_08594_));
 AND2x4_ASAP7_75t_R _23953_ (.A(_02191_),
    .B(_08298_),
    .Y(_08595_));
 BUFx6f_ASAP7_75t_R _23954_ (.A(_08595_),
    .Y(_08596_));
 BUFx6f_ASAP7_75t_R _23955_ (.A(_08596_),
    .Y(_08597_));
 NOR2x1_ASAP7_75t_R _23956_ (.A(net59),
    .B(_08276_),
    .Y(_08598_));
 AOI21x1_ASAP7_75t_R _23957_ (.A1(_01431_),
    .A2(_08275_),
    .B(_08598_),
    .Y(_08599_));
 INVx1_ASAP7_75t_R _23958_ (.A(_01416_),
    .Y(_08600_));
 OR2x2_ASAP7_75t_R _23959_ (.A(net79),
    .B(_08289_),
    .Y(_08601_));
 BUFx6f_ASAP7_75t_R _23960_ (.A(_08269_),
    .Y(_08602_));
 OA211x2_ASAP7_75t_R _23961_ (.A1(_08600_),
    .A2(_08279_),
    .B(_08601_),
    .C(_08602_),
    .Y(_08603_));
 AO21x1_ASAP7_75t_R _23962_ (.A1(_08287_),
    .A2(_08599_),
    .B(_08603_),
    .Y(_08604_));
 BUFx6f_ASAP7_75t_R _23963_ (.A(_08602_),
    .Y(_08605_));
 BUFx6f_ASAP7_75t_R _23964_ (.A(_08276_),
    .Y(_08606_));
 OA21x2_ASAP7_75t_R _23965_ (.A1(net56),
    .A2(_08606_),
    .B(_08601_),
    .Y(_08607_));
 INVx1_ASAP7_75t_R _23966_ (.A(net65),
    .Y(_08608_));
 BUFx6f_ASAP7_75t_R _23967_ (.A(_08273_),
    .Y(_08609_));
 AO21x1_ASAP7_75t_R _23968_ (.A1(_08608_),
    .A2(_08609_),
    .B(_08598_),
    .Y(_08610_));
 NOR2x1_ASAP7_75t_R _23969_ (.A(_08270_),
    .B(_08610_),
    .Y(_08611_));
 AO21x1_ASAP7_75t_R _23970_ (.A1(_08605_),
    .A2(_08607_),
    .B(_08611_),
    .Y(_08612_));
 NAND2x1_ASAP7_75t_R _23971_ (.A(_08504_),
    .B(_08304_),
    .Y(_08613_));
 AO221x1_ASAP7_75t_R _23972_ (.A1(_08597_),
    .A2(_08604_),
    .B1(_08612_),
    .B2(_05727_),
    .C(_08613_),
    .Y(_08614_));
 OA21x2_ASAP7_75t_R _23973_ (.A1(_08574_),
    .A2(_08594_),
    .B(_08614_),
    .Y(_08615_));
 AND2x2_ASAP7_75t_R _23974_ (.A(_14079_),
    .B(_08509_),
    .Y(_08616_));
 AO21x1_ASAP7_75t_R _23975_ (.A1(_08265_),
    .A2(_08615_),
    .B(_08616_),
    .Y(_02840_));
 BUFx6f_ASAP7_75t_R _23976_ (.A(_08308_),
    .Y(_08617_));
 OR3x1_ASAP7_75t_R _23977_ (.A(_08315_),
    .B(_08549_),
    .C(_08552_),
    .Y(_08618_));
 OR3x1_ASAP7_75t_R _23978_ (.A(_08448_),
    .B(_08531_),
    .C(_08534_),
    .Y(_08619_));
 AND2x4_ASAP7_75t_R _23979_ (.A(_08618_),
    .B(_08619_),
    .Y(_08620_));
 AO221x1_ASAP7_75t_R _23980_ (.A1(_08445_),
    .A2(_08430_),
    .B1(_08537_),
    .B2(_08413_),
    .C(_08314_),
    .Y(_08621_));
 OA21x2_ASAP7_75t_R _23981_ (.A1(_08536_),
    .A2(_08621_),
    .B(_08586_),
    .Y(_08622_));
 AND2x2_ASAP7_75t_R _23982_ (.A(_08311_),
    .B(_08622_),
    .Y(_08623_));
 AO21x1_ASAP7_75t_R _23983_ (.A1(_08368_),
    .A2(_08620_),
    .B(_08623_),
    .Y(_08624_));
 OA21x2_ASAP7_75t_R _23984_ (.A1(_08617_),
    .A2(_08624_),
    .B(_08460_),
    .Y(_08625_));
 AND3x1_ASAP7_75t_R _23985_ (.A(_08445_),
    .B(_08360_),
    .C(_08363_),
    .Y(_08626_));
 AND3x1_ASAP7_75t_R _23986_ (.A(_08336_),
    .B(_08329_),
    .C(_08333_),
    .Y(_08627_));
 OR2x6_ASAP7_75t_R _23987_ (.A(_08626_),
    .B(_08627_),
    .Y(_08628_));
 OR3x1_ASAP7_75t_R _23988_ (.A(_08448_),
    .B(_08578_),
    .C(_08580_),
    .Y(_08629_));
 OA21x2_ASAP7_75t_R _23989_ (.A1(_08316_),
    .A2(_08628_),
    .B(_08629_),
    .Y(_08630_));
 AND3x1_ASAP7_75t_R _23990_ (.A(_08445_),
    .B(_08377_),
    .C(_08379_),
    .Y(_08631_));
 AND3x1_ASAP7_75t_R _23991_ (.A(_08336_),
    .B(_08384_),
    .C(_08387_),
    .Y(_08632_));
 OR3x1_ASAP7_75t_R _23992_ (.A(_08315_),
    .B(_08631_),
    .C(_08632_),
    .Y(_08633_));
 AND3x1_ASAP7_75t_R _23993_ (.A(_08445_),
    .B(_08340_),
    .C(_08343_),
    .Y(_08634_));
 OA211x2_ASAP7_75t_R _23994_ (.A1(_05930_),
    .A2(_08370_),
    .B(_08373_),
    .C(_08336_),
    .Y(_08635_));
 OR3x1_ASAP7_75t_R _23995_ (.A(_08448_),
    .B(_08634_),
    .C(_08635_),
    .Y(_08636_));
 AND3x1_ASAP7_75t_R _23996_ (.A(_08368_),
    .B(_08633_),
    .C(_08636_),
    .Y(_08637_));
 AO21x1_ASAP7_75t_R _23997_ (.A1(_08312_),
    .A2(_08630_),
    .B(_08637_),
    .Y(_08638_));
 OR3x1_ASAP7_75t_R _23998_ (.A(_08528_),
    .B(_08575_),
    .C(_08576_),
    .Y(_08639_));
 OA21x2_ASAP7_75t_R _23999_ (.A1(_08514_),
    .A2(_08585_),
    .B(_08639_),
    .Y(_08640_));
 OA21x2_ASAP7_75t_R _24000_ (.A1(_08426_),
    .A2(_08640_),
    .B(_08431_),
    .Y(_08641_));
 OA21x2_ASAP7_75t_R _24001_ (.A1(_08308_),
    .A2(_08638_),
    .B(_08641_),
    .Y(_08642_));
 INVx1_ASAP7_75t_R _24002_ (.A(_02303_),
    .Y(_08643_));
 OA222x2_ASAP7_75t_R _24003_ (.A1(_00289_),
    .A2(_08559_),
    .B1(_08486_),
    .B2(_08643_),
    .C1(_08489_),
    .C2(_00288_),
    .Y(_08644_));
 OA21x2_ASAP7_75t_R _24004_ (.A1(_15248_),
    .A2(_08484_),
    .B(_08644_),
    .Y(_08645_));
 INVx1_ASAP7_75t_R _24005_ (.A(_00174_),
    .Y(_08646_));
 OA21x2_ASAP7_75t_R _24006_ (.A1(_00142_),
    .A2(_08646_),
    .B(_00151_),
    .Y(_08647_));
 OA21x2_ASAP7_75t_R _24007_ (.A1(_00150_),
    .A2(_08647_),
    .B(_00159_),
    .Y(_08648_));
 XOR2x1_ASAP7_75t_R _24008_ (.A(_00158_),
    .Y(_08649_),
    .B(_08648_));
 NAND3x1_ASAP7_75t_R _24009_ (.A(_05241_),
    .B(_08498_),
    .C(_08649_),
    .Y(_08650_));
 OA21x2_ASAP7_75t_R _24010_ (.A1(_00152_),
    .A2(_08569_),
    .B(_08650_),
    .Y(_08651_));
 OA21x2_ASAP7_75t_R _24011_ (.A1(_08483_),
    .A2(_08645_),
    .B(_08651_),
    .Y(_08652_));
 NAND2x1_ASAP7_75t_R _24012_ (.A(_05980_),
    .B(_08652_),
    .Y(_08653_));
 AO221x1_ASAP7_75t_R _24013_ (.A1(_08440_),
    .A2(_08625_),
    .B1(_08642_),
    .B2(_08512_),
    .C(_08653_),
    .Y(_08654_));
 INVx1_ASAP7_75t_R _24014_ (.A(net66),
    .Y(_08655_));
 NOR2x1_ASAP7_75t_R _24015_ (.A(net70),
    .B(_08276_),
    .Y(_08656_));
 AO21x1_ASAP7_75t_R _24016_ (.A1(_08655_),
    .A2(_08609_),
    .B(_08656_),
    .Y(_08657_));
 INVx1_ASAP7_75t_R _24017_ (.A(net28),
    .Y(_08658_));
 NAND2x1_ASAP7_75t_R _24018_ (.A(_08658_),
    .B(_08276_),
    .Y(_08659_));
 OA21x2_ASAP7_75t_R _24019_ (.A1(net57),
    .A2(_08274_),
    .B(_08659_),
    .Y(_08660_));
 NOR2x1_ASAP7_75t_R _24020_ (.A(_08282_),
    .B(_08660_),
    .Y(_08661_));
 AO21x1_ASAP7_75t_R _24021_ (.A1(_08287_),
    .A2(_08657_),
    .B(_08661_),
    .Y(_08662_));
 AOI211x1_ASAP7_75t_R _24022_ (.A1(_01430_),
    .A2(_08606_),
    .B(_08656_),
    .C(_08270_),
    .Y(_08663_));
 INVx1_ASAP7_75t_R _24023_ (.A(_01438_),
    .Y(_08664_));
 OA211x2_ASAP7_75t_R _24024_ (.A1(_08664_),
    .A2(_08279_),
    .B(_08659_),
    .C(_08294_),
    .Y(_08665_));
 OAI21x1_ASAP7_75t_R _24025_ (.A1(_08663_),
    .A2(_08665_),
    .B(_08596_),
    .Y(_08666_));
 OA211x2_ASAP7_75t_R _24026_ (.A1(_08296_),
    .A2(_08662_),
    .B(_08666_),
    .C(_08304_),
    .Y(_08667_));
 NAND2x1_ASAP7_75t_R _24027_ (.A(_08504_),
    .B(_08667_),
    .Y(_08668_));
 OA21x2_ASAP7_75t_R _24028_ (.A1(_08593_),
    .A2(_08654_),
    .B(_08668_),
    .Y(_08669_));
 AND2x2_ASAP7_75t_R _24029_ (.A(_14160_),
    .B(_08509_),
    .Y(_08670_));
 AO21x1_ASAP7_75t_R _24030_ (.A1(_08265_),
    .A2(_08669_),
    .B(_08670_),
    .Y(_02841_));
 OR3x1_ASAP7_75t_R _24031_ (.A(_08315_),
    .B(_08356_),
    .C(_08364_),
    .Y(_08671_));
 OA21x2_ASAP7_75t_R _24032_ (.A1(_08347_),
    .A2(_08411_),
    .B(_08671_),
    .Y(_08672_));
 OA31x2_ASAP7_75t_R _24033_ (.A1(_08315_),
    .A2(_08417_),
    .A3(_08423_),
    .B1(_08586_),
    .Y(_08673_));
 AND2x2_ASAP7_75t_R _24034_ (.A(_08311_),
    .B(_08673_),
    .Y(_08674_));
 AO21x1_ASAP7_75t_R _24035_ (.A1(_08368_),
    .A2(_08672_),
    .B(_08674_),
    .Y(_08675_));
 OA21x2_ASAP7_75t_R _24036_ (.A1(_08617_),
    .A2(_08675_),
    .B(_08460_),
    .Y(_08676_));
 OR3x1_ASAP7_75t_R _24037_ (.A(_08346_),
    .B(_08430_),
    .C(_08461_),
    .Y(_08677_));
 OA31x2_ASAP7_75t_R _24038_ (.A1(_08528_),
    .A2(_08451_),
    .A3(_08452_),
    .B1(_08677_),
    .Y(_08678_));
 AND2x2_ASAP7_75t_R _24039_ (.A(_08312_),
    .B(_08430_),
    .Y(_08679_));
 AO21x2_ASAP7_75t_R _24040_ (.A1(_08555_),
    .A2(_08678_),
    .B(_08679_),
    .Y(_08680_));
 AND3x1_ASAP7_75t_R _24041_ (.A(_08320_),
    .B(_08550_),
    .C(_08551_),
    .Y(_08681_));
 AND3x1_ASAP7_75t_R _24042_ (.A(_08337_),
    .B(_08542_),
    .C(_08543_),
    .Y(_08682_));
 OR3x1_ASAP7_75t_R _24043_ (.A(_08528_),
    .B(_08681_),
    .C(_08682_),
    .Y(_08683_));
 OR3x1_ASAP7_75t_R _24044_ (.A(_08347_),
    .B(_08443_),
    .C(_08446_),
    .Y(_08684_));
 AND2x4_ASAP7_75t_R _24045_ (.A(_08683_),
    .B(_08684_),
    .Y(_08685_));
 OA211x2_ASAP7_75t_R _24046_ (.A1(_13453_),
    .A2(_08370_),
    .B(_08522_),
    .C(_08348_),
    .Y(_08686_));
 AND3x1_ASAP7_75t_R _24047_ (.A(_08337_),
    .B(_08518_),
    .C(_08519_),
    .Y(_08687_));
 OA21x2_ASAP7_75t_R _24048_ (.A1(_08686_),
    .A2(_08687_),
    .B(_08347_),
    .Y(_08688_));
 AO21x1_ASAP7_75t_R _24049_ (.A1(_08545_),
    .A2(_08546_),
    .B(_08337_),
    .Y(_08689_));
 OR3x1_ASAP7_75t_R _24050_ (.A(_08348_),
    .B(_08525_),
    .C(_08526_),
    .Y(_08690_));
 AND3x1_ASAP7_75t_R _24051_ (.A(_08528_),
    .B(_08689_),
    .C(_08690_),
    .Y(_08691_));
 OR3x1_ASAP7_75t_R _24052_ (.A(_08312_),
    .B(_08688_),
    .C(_08691_),
    .Y(_08692_));
 OA211x2_ASAP7_75t_R _24053_ (.A1(_08555_),
    .A2(_08685_),
    .B(_08692_),
    .C(_08513_),
    .Y(_08693_));
 AO21x1_ASAP7_75t_R _24054_ (.A1(_08617_),
    .A2(_08680_),
    .B(_08693_),
    .Y(_08694_));
 BUFx6f_ASAP7_75t_R _24055_ (.A(_08488_),
    .Y(_08695_));
 INVx1_ASAP7_75t_R _24056_ (.A(_02304_),
    .Y(_08696_));
 OA222x2_ASAP7_75t_R _24057_ (.A1(_00291_),
    .A2(_08559_),
    .B1(_08486_),
    .B2(_08696_),
    .C1(_15240_),
    .C2(_08468_),
    .Y(_08697_));
 OA21x2_ASAP7_75t_R _24058_ (.A1(_00290_),
    .A2(_08695_),
    .B(_08697_),
    .Y(_08698_));
 OA21x2_ASAP7_75t_R _24059_ (.A1(_00150_),
    .A2(_08564_),
    .B(_00159_),
    .Y(_08699_));
 OA21x2_ASAP7_75t_R _24060_ (.A1(_00158_),
    .A2(_08699_),
    .B(_00167_),
    .Y(_08700_));
 XNOR2x1_ASAP7_75t_R _24061_ (.B(_08700_),
    .Y(_08701_),
    .A(_00166_));
 OA22x2_ASAP7_75t_R _24062_ (.A1(_00160_),
    .A2(_08569_),
    .B1(_08701_),
    .B2(_08566_),
    .Y(_08702_));
 OA21x2_ASAP7_75t_R _24063_ (.A1(_08483_),
    .A2(_08698_),
    .B(_08702_),
    .Y(_08703_));
 NAND2x1_ASAP7_75t_R _24064_ (.A(_06023_),
    .B(_08703_),
    .Y(_08704_));
 AO221x1_ASAP7_75t_R _24065_ (.A1(_08440_),
    .A2(_08676_),
    .B1(_08694_),
    .B2(_08512_),
    .C(_08704_),
    .Y(_08705_));
 INVx1_ASAP7_75t_R _24066_ (.A(net67),
    .Y(_08706_));
 NOR2x1_ASAP7_75t_R _24067_ (.A(net73),
    .B(_08276_),
    .Y(_08707_));
 AO21x1_ASAP7_75t_R _24068_ (.A1(_08706_),
    .A2(_08609_),
    .B(_08707_),
    .Y(_08708_));
 OR2x2_ASAP7_75t_R _24069_ (.A(net29),
    .B(_08288_),
    .Y(_08709_));
 OA21x2_ASAP7_75t_R _24070_ (.A1(net58),
    .A2(_08274_),
    .B(_08709_),
    .Y(_08710_));
 NOR2x1_ASAP7_75t_R _24071_ (.A(_08282_),
    .B(_08710_),
    .Y(_08711_));
 AO21x1_ASAP7_75t_R _24072_ (.A1(_08287_),
    .A2(_08708_),
    .B(_08711_),
    .Y(_08712_));
 AOI211x1_ASAP7_75t_R _24073_ (.A1(_01429_),
    .A2(_08606_),
    .B(_08707_),
    .C(_08270_),
    .Y(_08713_));
 INVx1_ASAP7_75t_R _24074_ (.A(_01437_),
    .Y(_08714_));
 OA211x2_ASAP7_75t_R _24075_ (.A1(_08714_),
    .A2(_08609_),
    .B(_08709_),
    .C(_08294_),
    .Y(_08715_));
 OAI21x1_ASAP7_75t_R _24076_ (.A1(_08713_),
    .A2(_08715_),
    .B(_08596_),
    .Y(_08716_));
 OA211x2_ASAP7_75t_R _24077_ (.A1(_08296_),
    .A2(_08712_),
    .B(_08716_),
    .C(_08304_),
    .Y(_08717_));
 NAND2x1_ASAP7_75t_R _24078_ (.A(_08504_),
    .B(_08717_),
    .Y(_08718_));
 OA21x2_ASAP7_75t_R _24079_ (.A1(_08593_),
    .A2(_08705_),
    .B(_08718_),
    .Y(_08719_));
 AND2x2_ASAP7_75t_R _24080_ (.A(_14251_),
    .B(_08509_),
    .Y(_08720_));
 AO21x1_ASAP7_75t_R _24081_ (.A1(_08265_),
    .A2(_08719_),
    .B(_08720_),
    .Y(_02842_));
 INVx3_ASAP7_75t_R _24082_ (.A(_08482_),
    .Y(_08721_));
 AND2x4_ASAP7_75t_R _24083_ (.A(_08427_),
    .B(_08310_),
    .Y(_08722_));
 INVx1_ASAP7_75t_R _24084_ (.A(_08722_),
    .Y(_08723_));
 OA22x2_ASAP7_75t_R _24085_ (.A1(_08723_),
    .A2(_08678_),
    .B1(_08685_),
    .B2(_08457_),
    .Y(_08724_));
 AND2x4_ASAP7_75t_R _24086_ (.A(_08307_),
    .B(_08367_),
    .Y(_08725_));
 OR3x1_ASAP7_75t_R _24087_ (.A(_08347_),
    .B(_08334_),
    .C(_08344_),
    .Y(_08726_));
 OA21x2_ASAP7_75t_R _24088_ (.A1(_08316_),
    .A2(_08381_),
    .B(_08726_),
    .Y(_08727_));
 OA211x2_ASAP7_75t_R _24089_ (.A1(_08307_),
    .A2(_08672_),
    .B(_08459_),
    .C(_08311_),
    .Y(_08728_));
 AO221x1_ASAP7_75t_R _24090_ (.A1(_08725_),
    .A2(_08673_),
    .B1(_08727_),
    .B2(_08456_),
    .C(_08728_),
    .Y(_08729_));
 BUFx6f_ASAP7_75t_R _24091_ (.A(_08484_),
    .Y(_08730_));
 BUFx6f_ASAP7_75t_R _24092_ (.A(_08559_),
    .Y(_08731_));
 BUFx6f_ASAP7_75t_R _24093_ (.A(_08486_),
    .Y(_08732_));
 INVx1_ASAP7_75t_R _24094_ (.A(_02305_),
    .Y(_08733_));
 OA222x2_ASAP7_75t_R _24095_ (.A1(_00293_),
    .A2(_08731_),
    .B1(_08732_),
    .B2(_08733_),
    .C1(_08558_),
    .C2(_00292_),
    .Y(_08734_));
 OAI21x1_ASAP7_75t_R _24096_ (.A1(_15524_),
    .A2(_08730_),
    .B(_08734_),
    .Y(_08735_));
 AO221x1_ASAP7_75t_R _24097_ (.A1(_08590_),
    .A2(_08724_),
    .B1(_08729_),
    .B2(_08512_),
    .C(_08735_),
    .Y(_08736_));
 NAND2x1_ASAP7_75t_R _24098_ (.A(_08721_),
    .B(_08736_),
    .Y(_08737_));
 AND4x1_ASAP7_75t_R _24099_ (.A(_05149_),
    .B(_07158_),
    .C(_05192_),
    .D(_08267_),
    .Y(_08738_));
 OA21x2_ASAP7_75t_R _24100_ (.A1(_00158_),
    .A2(_08648_),
    .B(_00167_),
    .Y(_08739_));
 OA21x2_ASAP7_75t_R _24101_ (.A1(_00166_),
    .A2(_08739_),
    .B(_00173_),
    .Y(_08740_));
 XOR2x1_ASAP7_75t_R _24102_ (.A(_00172_),
    .Y(_08741_),
    .B(_08740_));
 INVx1_ASAP7_75t_R _24103_ (.A(_08741_),
    .Y(_08742_));
 OA22x2_ASAP7_75t_R _24104_ (.A1(_00168_),
    .A2(_08570_),
    .B1(_08742_),
    .B2(_08567_),
    .Y(_08743_));
 AND3x1_ASAP7_75t_R _24105_ (.A(_06050_),
    .B(_08738_),
    .C(_08743_),
    .Y(_08744_));
 NAND2x1_ASAP7_75t_R _24106_ (.A(net74),
    .B(_08289_),
    .Y(_08745_));
 OA211x2_ASAP7_75t_R _24107_ (.A1(_01427_),
    .A2(_08289_),
    .B(_08745_),
    .C(_08282_),
    .Y(_08746_));
 NAND2x1_ASAP7_75t_R _24108_ (.A(net30),
    .B(_08273_),
    .Y(_08747_));
 OA211x2_ASAP7_75t_R _24109_ (.A1(_01436_),
    .A2(_08279_),
    .B(_08747_),
    .C(_08294_),
    .Y(_08748_));
 INVx1_ASAP7_75t_R _24110_ (.A(net68),
    .Y(_08749_));
 OAI21x1_ASAP7_75t_R _24111_ (.A1(_08749_),
    .A2(_08289_),
    .B(_08745_),
    .Y(_08750_));
 NOR2x1_ASAP7_75t_R _24112_ (.A(_08270_),
    .B(_08750_),
    .Y(_08751_));
 INVx1_ASAP7_75t_R _24113_ (.A(net60),
    .Y(_08752_));
 OA21x2_ASAP7_75t_R _24114_ (.A1(_08752_),
    .A2(_08276_),
    .B(_08747_),
    .Y(_08753_));
 AND2x2_ASAP7_75t_R _24115_ (.A(_08602_),
    .B(_08753_),
    .Y(_08754_));
 OA33x2_ASAP7_75t_R _24116_ (.A1(_08286_),
    .A2(_08746_),
    .A3(_08748_),
    .B1(_08751_),
    .B2(_08754_),
    .B3(_08296_),
    .Y(_08755_));
 AND3x4_ASAP7_75t_R _24117_ (.A(_08504_),
    .B(_08304_),
    .C(_08755_),
    .Y(_08756_));
 AOI21x1_ASAP7_75t_R _24118_ (.A1(_08737_),
    .A2(_08744_),
    .B(_08756_),
    .Y(_08757_));
 AND2x2_ASAP7_75t_R _24119_ (.A(_13177_),
    .B(_08509_),
    .Y(_08758_));
 AO21x1_ASAP7_75t_R _24120_ (.A1(_08265_),
    .A2(_08757_),
    .B(_08758_),
    .Y(_02843_));
 INVx1_ASAP7_75t_R _24121_ (.A(_02306_),
    .Y(_08759_));
 OA222x2_ASAP7_75t_R _24122_ (.A1(_00295_),
    .A2(_08731_),
    .B1(_08732_),
    .B2(_08759_),
    .C1(_15518_),
    .C2(_08730_),
    .Y(_08760_));
 OAI21x1_ASAP7_75t_R _24123_ (.A1(_00294_),
    .A2(_08558_),
    .B(_08760_),
    .Y(_08761_));
 AND2x2_ASAP7_75t_R _24124_ (.A(_08312_),
    .B(_08640_),
    .Y(_08762_));
 AND2x2_ASAP7_75t_R _24125_ (.A(_08555_),
    .B(_08630_),
    .Y(_08763_));
 OR3x1_ASAP7_75t_R _24126_ (.A(_08617_),
    .B(_08762_),
    .C(_08763_),
    .Y(_08764_));
 OA21x2_ASAP7_75t_R _24127_ (.A1(_08308_),
    .A2(_08620_),
    .B(_08460_),
    .Y(_08765_));
 OR2x2_ASAP7_75t_R _24128_ (.A(_08544_),
    .B(_08547_),
    .Y(_08766_));
 OA211x2_ASAP7_75t_R _24129_ (.A1(_08320_),
    .A2(_08523_),
    .B(_08527_),
    .C(_08448_),
    .Y(_08767_));
 INVx1_ASAP7_75t_R _24130_ (.A(_08767_),
    .Y(_08768_));
 OA21x2_ASAP7_75t_R _24131_ (.A1(_08514_),
    .A2(_08766_),
    .B(_08768_),
    .Y(_08769_));
 AND2x2_ASAP7_75t_R _24132_ (.A(_08307_),
    .B(_08622_),
    .Y(_08770_));
 AO211x2_ASAP7_75t_R _24133_ (.A1(_08513_),
    .A2(_08769_),
    .B(_08770_),
    .C(_08312_),
    .Y(_08771_));
 OA211x2_ASAP7_75t_R _24134_ (.A1(_08555_),
    .A2(_08765_),
    .B(_08771_),
    .C(_08511_),
    .Y(_08772_));
 AO221x1_ASAP7_75t_R _24135_ (.A1(_08721_),
    .A2(_08761_),
    .B1(_08764_),
    .B2(_08590_),
    .C(_08772_),
    .Y(_08773_));
 AND3x1_ASAP7_75t_R _24136_ (.A(_00159_),
    .B(_00167_),
    .C(_00173_),
    .Y(_08774_));
 OA21x2_ASAP7_75t_R _24137_ (.A1(_00150_),
    .A2(_08564_),
    .B(_08774_),
    .Y(_08775_));
 AND3x1_ASAP7_75t_R _24138_ (.A(_00158_),
    .B(_00167_),
    .C(_00173_),
    .Y(_08776_));
 AO21x1_ASAP7_75t_R _24139_ (.A1(_00166_),
    .A2(_00173_),
    .B(_08776_),
    .Y(_08777_));
 OR3x1_ASAP7_75t_R _24140_ (.A(_00172_),
    .B(_08775_),
    .C(_08777_),
    .Y(_08778_));
 AND2x4_ASAP7_75t_R _24141_ (.A(_00179_),
    .B(_08778_),
    .Y(_08779_));
 XNOR2x1_ASAP7_75t_R _24142_ (.B(_08779_),
    .Y(_08780_),
    .A(_00178_));
 AND2x2_ASAP7_75t_R _24143_ (.A(_00175_),
    .B(_08495_),
    .Y(_08781_));
 AO21x1_ASAP7_75t_R _24144_ (.A1(_08498_),
    .A2(_08780_),
    .B(_08781_),
    .Y(_08782_));
 AO21x1_ASAP7_75t_R _24145_ (.A1(_14533_),
    .A2(_08782_),
    .B(_08568_),
    .Y(_08783_));
 AO21x2_ASAP7_75t_R _24146_ (.A1(_00175_),
    .A2(_05720_),
    .B(_08783_),
    .Y(_08784_));
 AND3x1_ASAP7_75t_R _24147_ (.A(_06081_),
    .B(_08738_),
    .C(_08784_),
    .Y(_08785_));
 INVx1_ASAP7_75t_R _24148_ (.A(_08785_),
    .Y(_08786_));
 AND2x6_ASAP7_75t_R _24149_ (.A(_08269_),
    .B(_08288_),
    .Y(_08787_));
 AO221x1_ASAP7_75t_R _24150_ (.A1(net69),
    .A2(_08272_),
    .B1(_08787_),
    .B2(net61),
    .C(_08296_),
    .Y(_08788_));
 INVx1_ASAP7_75t_R _24151_ (.A(_01426_),
    .Y(_08789_));
 AND2x4_ASAP7_75t_R _24152_ (.A(_08281_),
    .B(_08272_),
    .Y(_08790_));
 INVx1_ASAP7_75t_R _24153_ (.A(_01435_),
    .Y(_08791_));
 AO221x1_ASAP7_75t_R _24154_ (.A1(_08789_),
    .A2(_08790_),
    .B1(_08787_),
    .B2(_08791_),
    .C(_05727_),
    .Y(_08792_));
 NAND2x1_ASAP7_75t_R _24155_ (.A(_08788_),
    .B(_08792_),
    .Y(_08793_));
 NAND2x1_ASAP7_75t_R _24156_ (.A(net75),
    .B(_08289_),
    .Y(_08794_));
 AO21x1_ASAP7_75t_R _24157_ (.A1(_08793_),
    .A2(_08794_),
    .B(_08294_),
    .Y(_08795_));
 AND2x6_ASAP7_75t_R _24158_ (.A(_08269_),
    .B(_08273_),
    .Y(_08796_));
 NAND2x1_ASAP7_75t_R _24159_ (.A(net31),
    .B(_08796_),
    .Y(_08797_));
 OA211x2_ASAP7_75t_R _24160_ (.A1(_08275_),
    .A2(_08793_),
    .B(_08795_),
    .C(_08797_),
    .Y(_08798_));
 AND2x6_ASAP7_75t_R _24161_ (.A(_08296_),
    .B(_05738_),
    .Y(_08799_));
 OA211x2_ASAP7_75t_R _24162_ (.A1(_08798_),
    .A2(_08799_),
    .B(_08504_),
    .C(_08304_),
    .Y(_08800_));
 INVx1_ASAP7_75t_R _24163_ (.A(_08800_),
    .Y(_08801_));
 OA21x2_ASAP7_75t_R _24164_ (.A1(_08773_),
    .A2(_08786_),
    .B(_08801_),
    .Y(_08802_));
 AND2x2_ASAP7_75t_R _24165_ (.A(_15406_),
    .B(_08509_),
    .Y(_08803_));
 AO21x1_ASAP7_75t_R _24166_ (.A1(_08265_),
    .A2(_08802_),
    .B(_08803_),
    .Y(_02844_));
 BUFx6f_ASAP7_75t_R _24167_ (.A(_08508_),
    .Y(_08804_));
 AND2x2_ASAP7_75t_R _24168_ (.A(_00180_),
    .B(_08495_),
    .Y(_08805_));
 AND3x1_ASAP7_75t_R _24169_ (.A(_00173_),
    .B(_00179_),
    .C(_00186_),
    .Y(_08806_));
 OA21x2_ASAP7_75t_R _24170_ (.A1(_00166_),
    .A2(_08739_),
    .B(_08806_),
    .Y(_08807_));
 AND3x1_ASAP7_75t_R _24171_ (.A(_00172_),
    .B(_00179_),
    .C(_00186_),
    .Y(_08808_));
 AO21x2_ASAP7_75t_R _24172_ (.A1(_00178_),
    .A2(_00186_),
    .B(_08808_),
    .Y(_08809_));
 NOR2x1_ASAP7_75t_R _24173_ (.A(_08807_),
    .B(_08809_),
    .Y(_08810_));
 XNOR2x1_ASAP7_75t_R _24174_ (.B(_08810_),
    .Y(_08811_),
    .A(net1967));
 NOR2x1_ASAP7_75t_R _24175_ (.A(_08495_),
    .B(_08811_),
    .Y(_08812_));
 OR3x2_ASAP7_75t_R _24176_ (.A(_14541_),
    .B(_08805_),
    .C(_08812_),
    .Y(_08813_));
 OA21x2_ASAP7_75t_R _24177_ (.A1(_14533_),
    .A2(_00180_),
    .B(_08813_),
    .Y(_08814_));
 BUFx6f_ASAP7_75t_R _24178_ (.A(_08478_),
    .Y(_08815_));
 INVx1_ASAP7_75t_R _24179_ (.A(_02307_),
    .Y(_08816_));
 OA222x2_ASAP7_75t_R _24180_ (.A1(_00297_),
    .A2(_08485_),
    .B1(_08815_),
    .B2(_08816_),
    .C1(_08489_),
    .C2(_00296_),
    .Y(_08817_));
 AND2x6_ASAP7_75t_R _24181_ (.A(_14604_),
    .B(_08467_),
    .Y(_08818_));
 NAND2x1_ASAP7_75t_R _24182_ (.A(\alu_adder_result_ex[14] ),
    .B(_08818_),
    .Y(_08819_));
 AO21x1_ASAP7_75t_R _24183_ (.A1(_08817_),
    .A2(_08819_),
    .B(_08483_),
    .Y(_08820_));
 OA211x2_ASAP7_75t_R _24184_ (.A1(_14627_),
    .A2(_08814_),
    .B(_08820_),
    .C(_06107_),
    .Y(_08821_));
 OA211x2_ASAP7_75t_R _24185_ (.A1(_08514_),
    .A2(_08577_),
    .B(_08581_),
    .C(_08311_),
    .Y(_08822_));
 OR3x1_ASAP7_75t_R _24186_ (.A(_08528_),
    .B(_08634_),
    .C(_08635_),
    .Y(_08823_));
 OA211x2_ASAP7_75t_R _24187_ (.A1(_08514_),
    .A2(_08628_),
    .B(_08823_),
    .C(_08368_),
    .Y(_08824_));
 NAND2x1_ASAP7_75t_R _24188_ (.A(_08346_),
    .B(_08367_),
    .Y(_08825_));
 AO21x1_ASAP7_75t_R _24189_ (.A1(_08346_),
    .A2(_08367_),
    .B(_08430_),
    .Y(_08826_));
 OA31x2_ASAP7_75t_R _24190_ (.A1(_08535_),
    .A2(_08584_),
    .A3(_08825_),
    .B1(_08826_),
    .Y(_08827_));
 OR2x2_ASAP7_75t_R _24191_ (.A(_08427_),
    .B(_08827_),
    .Y(_08828_));
 OA31x2_ASAP7_75t_R _24192_ (.A1(_08308_),
    .A2(_08822_),
    .A3(_08824_),
    .B1(_08828_),
    .Y(_08829_));
 AND2x2_ASAP7_75t_R _24193_ (.A(_08548_),
    .B(_08553_),
    .Y(_08830_));
 AND2x2_ASAP7_75t_R _24194_ (.A(_08311_),
    .B(_08539_),
    .Y(_08831_));
 AO21x1_ASAP7_75t_R _24195_ (.A1(_08555_),
    .A2(_08830_),
    .B(_08831_),
    .Y(_08832_));
 BUFx6f_ASAP7_75t_R _24196_ (.A(_08439_),
    .Y(_08833_));
 OA211x2_ASAP7_75t_R _24197_ (.A1(_08617_),
    .A2(_08832_),
    .B(_08460_),
    .C(_08833_),
    .Y(_08834_));
 BUFx6f_ASAP7_75t_R _24198_ (.A(_08592_),
    .Y(_08835_));
 AOI211x1_ASAP7_75t_R _24199_ (.A1(_08512_),
    .A2(_08829_),
    .B(_08834_),
    .C(_08835_),
    .Y(_08836_));
 NOR2x1_ASAP7_75t_R _24200_ (.A(net76),
    .B(_08272_),
    .Y(_08837_));
 AOI211x1_ASAP7_75t_R _24201_ (.A1(_01425_),
    .A2(_08279_),
    .B(_08837_),
    .C(_08602_),
    .Y(_08838_));
 INVx1_ASAP7_75t_R _24202_ (.A(_01434_),
    .Y(_08839_));
 OR2x2_ASAP7_75t_R _24203_ (.A(net53),
    .B(_08288_),
    .Y(_08840_));
 OA211x2_ASAP7_75t_R _24204_ (.A1(_08839_),
    .A2(_08274_),
    .B(_08840_),
    .C(_08294_),
    .Y(_08841_));
 OAI21x1_ASAP7_75t_R _24205_ (.A1(_08838_),
    .A2(_08841_),
    .B(_08596_),
    .Y(_08842_));
 INVx1_ASAP7_75t_R _24206_ (.A(net71),
    .Y(_08843_));
 AO21x1_ASAP7_75t_R _24207_ (.A1(_08843_),
    .A2(_08273_),
    .B(_08837_),
    .Y(_08844_));
 AND2x2_ASAP7_75t_R _24208_ (.A(_08282_),
    .B(_08844_),
    .Y(_08845_));
 OA21x2_ASAP7_75t_R _24209_ (.A1(net62),
    .A2(_08273_),
    .B(_08840_),
    .Y(_08846_));
 NOR2x1_ASAP7_75t_R _24210_ (.A(_08282_),
    .B(_08846_),
    .Y(_08847_));
 OR3x1_ASAP7_75t_R _24211_ (.A(_08296_),
    .B(_08845_),
    .C(_08847_),
    .Y(_08848_));
 AND4x1_ASAP7_75t_R _24212_ (.A(_08261_),
    .B(_08304_),
    .C(_08842_),
    .D(_08848_),
    .Y(_08849_));
 AO21x2_ASAP7_75t_R _24213_ (.A1(_08821_),
    .A2(_08836_),
    .B(_08849_),
    .Y(_08850_));
 BUFx12f_ASAP7_75t_R _24214_ (.A(_08850_),
    .Y(_08851_));
 NOR2x1_ASAP7_75t_R _24215_ (.A(_08804_),
    .B(_08851_),
    .Y(_08852_));
 AO21x1_ASAP7_75t_R _24216_ (.A1(_15559_),
    .A2(_08804_),
    .B(_08852_),
    .Y(_02845_));
 BUFx12f_ASAP7_75t_R _24217_ (.A(_08738_),
    .Y(_08853_));
 NOR2x1_ASAP7_75t_R _24218_ (.A(net77),
    .B(_08272_),
    .Y(_08854_));
 AO21x1_ASAP7_75t_R _24219_ (.A1(_01424_),
    .A2(_08275_),
    .B(_08854_),
    .Y(_08855_));
 INVx1_ASAP7_75t_R _24220_ (.A(_01433_),
    .Y(_08856_));
 OR2x2_ASAP7_75t_R _24221_ (.A(net54),
    .B(_08288_),
    .Y(_08857_));
 OA211x2_ASAP7_75t_R _24222_ (.A1(_08856_),
    .A2(_08279_),
    .B(_08857_),
    .C(_08294_),
    .Y(_08858_));
 INVx1_ASAP7_75t_R _24223_ (.A(_08858_),
    .Y(_08859_));
 OA21x2_ASAP7_75t_R _24224_ (.A1(_08605_),
    .A2(_08855_),
    .B(_08859_),
    .Y(_08860_));
 OA21x2_ASAP7_75t_R _24225_ (.A1(net63),
    .A2(_08272_),
    .B(_08857_),
    .Y(_08861_));
 NAND2x1_ASAP7_75t_R _24226_ (.A(_08269_),
    .B(_08861_),
    .Y(_08862_));
 INVx1_ASAP7_75t_R _24227_ (.A(net72),
    .Y(_08863_));
 AO21x1_ASAP7_75t_R _24228_ (.A1(_08863_),
    .A2(_08272_),
    .B(_08854_),
    .Y(_08864_));
 OR2x2_ASAP7_75t_R _24229_ (.A(_08269_),
    .B(_08864_),
    .Y(_08865_));
 AO21x1_ASAP7_75t_R _24230_ (.A1(_08862_),
    .A2(_08865_),
    .B(_08296_),
    .Y(_08866_));
 OA211x2_ASAP7_75t_R _24231_ (.A1(_08286_),
    .A2(_08860_),
    .B(_08866_),
    .C(_08304_),
    .Y(_08867_));
 NAND2x1_ASAP7_75t_R _24232_ (.A(_08312_),
    .B(_08425_),
    .Y(_08868_));
 AND2x4_ASAP7_75t_R _24233_ (.A(_08345_),
    .B(_08365_),
    .Y(_08869_));
 NAND2x1_ASAP7_75t_R _24234_ (.A(_08555_),
    .B(_08869_),
    .Y(_08870_));
 INVx1_ASAP7_75t_R _24235_ (.A(_08460_),
    .Y(_08871_));
 AO31x2_ASAP7_75t_R _24236_ (.A1(_08513_),
    .A2(_08868_),
    .A3(_08870_),
    .B(_08871_),
    .Y(_08872_));
 AO21x2_ASAP7_75t_R _24237_ (.A1(_08367_),
    .A2(_08462_),
    .B(_08430_),
    .Y(_08873_));
 OA21x2_ASAP7_75t_R _24238_ (.A1(_08681_),
    .A2(_08682_),
    .B(_08528_),
    .Y(_08874_));
 AND3x1_ASAP7_75t_R _24239_ (.A(_08347_),
    .B(_08689_),
    .C(_08690_),
    .Y(_08875_));
 OR3x1_ASAP7_75t_R _24240_ (.A(_08312_),
    .B(_08874_),
    .C(_08875_),
    .Y(_08876_));
 OA211x2_ASAP7_75t_R _24241_ (.A1(_08454_),
    .A2(_08555_),
    .B(_08876_),
    .C(_08513_),
    .Y(_08877_));
 AOI211x1_ASAP7_75t_R _24242_ (.A1(_08617_),
    .A2(_08873_),
    .B(_08877_),
    .C(_08440_),
    .Y(_08878_));
 AO21x1_ASAP7_75t_R _24243_ (.A1(_08440_),
    .A2(_08872_),
    .B(_08878_),
    .Y(_08879_));
 BUFx6f_ASAP7_75t_R _24244_ (.A(_08482_),
    .Y(_08880_));
 INVx1_ASAP7_75t_R _24245_ (.A(_02308_),
    .Y(_08881_));
 OA222x2_ASAP7_75t_R _24246_ (.A1(_00299_),
    .A2(_08731_),
    .B1(_08732_),
    .B2(_08881_),
    .C1(_08695_),
    .C2(_00298_),
    .Y(_08882_));
 OA21x2_ASAP7_75t_R _24247_ (.A1(_15764_),
    .A2(_08730_),
    .B(_08882_),
    .Y(_08883_));
 OA21x2_ASAP7_75t_R _24248_ (.A1(_00178_),
    .A2(_08779_),
    .B(_00186_),
    .Y(_08884_));
 OA21x2_ASAP7_75t_R _24249_ (.A1(net1967),
    .A2(_08884_),
    .B(_00195_),
    .Y(_08885_));
 XNOR2x1_ASAP7_75t_R _24250_ (.B(_08885_),
    .Y(_08886_),
    .A(_00194_));
 OA21x2_ASAP7_75t_R _24251_ (.A1(_00187_),
    .A2(_08570_),
    .B(_14388_),
    .Y(_08887_));
 OA21x2_ASAP7_75t_R _24252_ (.A1(_08567_),
    .A2(_08886_),
    .B(_08887_),
    .Y(_08888_));
 OA21x2_ASAP7_75t_R _24253_ (.A1(_08880_),
    .A2(_08883_),
    .B(_08888_),
    .Y(_08889_));
 OA21x2_ASAP7_75t_R _24254_ (.A1(_08466_),
    .A2(_08879_),
    .B(_08889_),
    .Y(_08890_));
 AO21x1_ASAP7_75t_R _24255_ (.A1(_14120_),
    .A2(_06130_),
    .B(_08593_),
    .Y(_08891_));
 OAI22x1_ASAP7_75t_R _24256_ (.A1(_08853_),
    .A2(_08867_),
    .B1(_08890_),
    .B2(_08891_),
    .Y(_08892_));
 NAND2x1_ASAP7_75t_R _24257_ (.A(_00876_),
    .B(_08804_),
    .Y(_08893_));
 OA21x2_ASAP7_75t_R _24258_ (.A1(_08804_),
    .A2(_08892_),
    .B(_08893_),
    .Y(_02846_));
 AO21x1_ASAP7_75t_R _24259_ (.A1(_08617_),
    .A2(_08873_),
    .B(_08434_),
    .Y(_08894_));
 OAI21x1_ASAP7_75t_R _24260_ (.A1(_08877_),
    .A2(_08894_),
    .B(_08437_),
    .Y(_08895_));
 AO21x1_ASAP7_75t_R _24261_ (.A1(_08434_),
    .A2(_08872_),
    .B(_08895_),
    .Y(_08896_));
 INVx1_ASAP7_75t_R _24262_ (.A(_02309_),
    .Y(_08897_));
 OA222x2_ASAP7_75t_R _24263_ (.A1(_00301_),
    .A2(_08485_),
    .B1(_08815_),
    .B2(_08897_),
    .C1(_08695_),
    .C2(_00300_),
    .Y(_08898_));
 OR2x2_ASAP7_75t_R _24264_ (.A(_16019_),
    .B(_08484_),
    .Y(_08899_));
 AO21x1_ASAP7_75t_R _24265_ (.A1(_08898_),
    .A2(_08899_),
    .B(_08483_),
    .Y(_08900_));
 NAND2x2_ASAP7_75t_R _24266_ (.A(_14541_),
    .B(_15234_),
    .Y(_08901_));
 BUFx6f_ASAP7_75t_R _24267_ (.A(_08498_),
    .Y(_08902_));
 OR3x1_ASAP7_75t_R _24268_ (.A(net1967),
    .B(_08807_),
    .C(_08809_),
    .Y(_08903_));
 AO21x1_ASAP7_75t_R _24269_ (.A1(_00195_),
    .A2(_08903_),
    .B(_00194_),
    .Y(_08904_));
 AND2x2_ASAP7_75t_R _24270_ (.A(_00200_),
    .B(_08904_),
    .Y(_08905_));
 XNOR2x2_ASAP7_75t_R _24271_ (.A(_00199_),
    .B(_08905_),
    .Y(_08906_));
 AND2x2_ASAP7_75t_R _24272_ (.A(_00064_),
    .B(_08495_),
    .Y(_08907_));
 AO21x1_ASAP7_75t_R _24273_ (.A1(_08902_),
    .A2(_08906_),
    .B(_08907_),
    .Y(_08908_));
 AOI21x1_ASAP7_75t_R _24274_ (.A1(_14533_),
    .A2(_08908_),
    .B(_08568_),
    .Y(_08909_));
 OAI21x1_ASAP7_75t_R _24275_ (.A1(_05636_),
    .A2(_08901_),
    .B(_08909_),
    .Y(_08910_));
 AND4x1_ASAP7_75t_R _24276_ (.A(_06152_),
    .B(_08738_),
    .C(_08900_),
    .D(_08910_),
    .Y(_08911_));
 OA21x2_ASAP7_75t_R _24277_ (.A1(_01445_),
    .A2(_08866_),
    .B(_08304_),
    .Y(_08912_));
 OR2x2_ASAP7_75t_R _24278_ (.A(_01432_),
    .B(_08273_),
    .Y(_08913_));
 OA211x2_ASAP7_75t_R _24279_ (.A1(_08293_),
    .A2(_08289_),
    .B(_08913_),
    .C(_08294_),
    .Y(_08914_));
 INVx1_ASAP7_75t_R _24280_ (.A(net78),
    .Y(_08915_));
 NAND2x1_ASAP7_75t_R _24281_ (.A(net27),
    .B(_08273_),
    .Y(_08916_));
 OA211x2_ASAP7_75t_R _24282_ (.A1(_08915_),
    .A2(_08276_),
    .B(_08916_),
    .C(_08282_),
    .Y(_08917_));
 OR3x1_ASAP7_75t_R _24283_ (.A(_08285_),
    .B(_08914_),
    .C(_08917_),
    .Y(_08918_));
 AND3x2_ASAP7_75t_R _24284_ (.A(_08261_),
    .B(_08912_),
    .C(_08918_),
    .Y(_08919_));
 AOI21x1_ASAP7_75t_R _24285_ (.A1(_08896_),
    .A2(_08911_),
    .B(_08919_),
    .Y(_08920_));
 AND2x2_ASAP7_75t_R _24286_ (.A(_08264_),
    .B(_08920_),
    .Y(_08921_));
 AO21x1_ASAP7_75t_R _24287_ (.A1(_15795_),
    .A2(_08804_),
    .B(_08921_),
    .Y(_02847_));
 NAND2x2_ASAP7_75t_R _24288_ (.A(_08592_),
    .B(_08912_),
    .Y(_08922_));
 AND2x2_ASAP7_75t_R _24289_ (.A(net59),
    .B(_08274_),
    .Y(_08923_));
 AO21x1_ASAP7_75t_R _24290_ (.A1(net79),
    .A2(_08290_),
    .B(_08923_),
    .Y(_08924_));
 NAND2x1_ASAP7_75t_R _24291_ (.A(net56),
    .B(_08276_),
    .Y(_08925_));
 OA211x2_ASAP7_75t_R _24292_ (.A1(_01431_),
    .A2(_08274_),
    .B(_08925_),
    .C(_08294_),
    .Y(_08926_));
 INVx1_ASAP7_75t_R _24293_ (.A(_08926_),
    .Y(_08927_));
 OA211x2_ASAP7_75t_R _24294_ (.A1(_08605_),
    .A2(_08924_),
    .B(_08927_),
    .C(_08596_),
    .Y(_08928_));
 AND2x2_ASAP7_75t_R _24295_ (.A(_08439_),
    .B(_08829_),
    .Y(_08929_));
 OA211x2_ASAP7_75t_R _24296_ (.A1(_08617_),
    .A2(_08832_),
    .B(_08511_),
    .C(_08460_),
    .Y(_08930_));
 INVx1_ASAP7_75t_R _24297_ (.A(_02310_),
    .Y(_08931_));
 OA222x2_ASAP7_75t_R _24298_ (.A1(_00303_),
    .A2(_08475_),
    .B1(_08478_),
    .B2(_08931_),
    .C1(_08488_),
    .C2(_00302_),
    .Y(_08932_));
 OA21x2_ASAP7_75t_R _24299_ (.A1(_16004_),
    .A2(_08484_),
    .B(_08932_),
    .Y(_08933_));
 OR5x1_ASAP7_75t_R _24300_ (.A(_00172_),
    .B(_00178_),
    .C(net1967),
    .D(_08775_),
    .E(_08777_),
    .Y(_08934_));
 OA21x2_ASAP7_75t_R _24301_ (.A1(_00179_),
    .A2(_00178_),
    .B(_00186_),
    .Y(_08935_));
 OA211x2_ASAP7_75t_R _24302_ (.A1(net1967),
    .A2(_08935_),
    .B(_00200_),
    .C(_00195_),
    .Y(_08936_));
 AO221x1_ASAP7_75t_R _24303_ (.A1(_00194_),
    .A2(_00200_),
    .B1(_08934_),
    .B2(_08936_),
    .C(_00199_),
    .Y(_08937_));
 AND3x1_ASAP7_75t_R _24304_ (.A(_00204_),
    .B(_00203_),
    .C(_08937_),
    .Y(_08938_));
 AOI21x1_ASAP7_75t_R _24305_ (.A1(_00204_),
    .A2(_08937_),
    .B(_00203_),
    .Y(_08939_));
 OA21x2_ASAP7_75t_R _24306_ (.A1(_08938_),
    .A2(_08939_),
    .B(_08498_),
    .Y(_08940_));
 AO21x1_ASAP7_75t_R _24307_ (.A1(_00099_),
    .A2(_08495_),
    .B(_08940_),
    .Y(_08941_));
 AO21x1_ASAP7_75t_R _24308_ (.A1(_14533_),
    .A2(_08941_),
    .B(_08568_),
    .Y(_08942_));
 AO21x1_ASAP7_75t_R _24309_ (.A1(_15947_),
    .A2(_05720_),
    .B(_08942_),
    .Y(_08943_));
 OA21x2_ASAP7_75t_R _24310_ (.A1(_08482_),
    .A2(_08933_),
    .B(_08943_),
    .Y(_08944_));
 NAND2x1_ASAP7_75t_R _24311_ (.A(_06177_),
    .B(_08944_),
    .Y(_08945_));
 OR4x1_ASAP7_75t_R _24312_ (.A(_08592_),
    .B(_08929_),
    .C(_08930_),
    .D(_08945_),
    .Y(_08946_));
 OAI21x1_ASAP7_75t_R _24313_ (.A1(_08922_),
    .A2(_08928_),
    .B(_08946_),
    .Y(_08947_));
 BUFx12f_ASAP7_75t_R _24314_ (.A(_08947_),
    .Y(_08948_));
 NOR2x1_ASAP7_75t_R _24315_ (.A(_08804_),
    .B(_08948_),
    .Y(_08949_));
 AO21x1_ASAP7_75t_R _24316_ (.A1(_15920_),
    .A2(_08804_),
    .B(_08949_),
    .Y(_02848_));
 BUFx12f_ASAP7_75t_R _24317_ (.A(_14094_),
    .Y(_08950_));
 INVx1_ASAP7_75t_R _24318_ (.A(_08262_),
    .Y(_08951_));
 OA211x2_ASAP7_75t_R _24319_ (.A1(_08255_),
    .A2(_08268_),
    .B(_00339_),
    .C(_08951_),
    .Y(_08952_));
 BUFx6f_ASAP7_75t_R _24320_ (.A(_08952_),
    .Y(_08953_));
 BUFx6f_ASAP7_75t_R _24321_ (.A(_08953_),
    .Y(_08954_));
 AND2x6_ASAP7_75t_R _24322_ (.A(_08950_),
    .B(_08954_),
    .Y(_08955_));
 BUFx6f_ASAP7_75t_R _24323_ (.A(_08955_),
    .Y(_08956_));
 OA211x2_ASAP7_75t_R _24324_ (.A1(_14709_),
    .A2(_16931_),
    .B(_16933_),
    .C(_08341_),
    .Y(_08957_));
 AND3x1_ASAP7_75t_R _24325_ (.A(_14965_),
    .B(_14970_),
    .C(_08331_),
    .Y(_08958_));
 OR3x1_ASAP7_75t_R _24326_ (.A(_08328_),
    .B(_08957_),
    .C(_08958_),
    .Y(_08959_));
 AND3x1_ASAP7_75t_R _24327_ (.A(_16820_),
    .B(_16822_),
    .C(_08326_),
    .Y(_08960_));
 AND3x1_ASAP7_75t_R _24328_ (.A(_15024_),
    .B(_15026_),
    .C(_08331_),
    .Y(_08961_));
 OR3x1_ASAP7_75t_R _24329_ (.A(_05829_),
    .B(_08960_),
    .C(_08961_),
    .Y(_08962_));
 AND3x1_ASAP7_75t_R _24330_ (.A(_08348_),
    .B(_08959_),
    .C(_08962_),
    .Y(_08963_));
 AND3x1_ASAP7_75t_R _24331_ (.A(_04418_),
    .B(_04421_),
    .C(_08326_),
    .Y(_08964_));
 AO211x2_ASAP7_75t_R _24332_ (.A1(_18572_),
    .A2(_08349_),
    .B(_08964_),
    .C(_08328_),
    .Y(_08965_));
 AND3x1_ASAP7_75t_R _24333_ (.A(_14899_),
    .B(_14902_),
    .C(_08331_),
    .Y(_08966_));
 AO211x2_ASAP7_75t_R _24334_ (.A1(_18685_),
    .A2(_08352_),
    .B(_08966_),
    .C(_13452_),
    .Y(_08967_));
 AND3x1_ASAP7_75t_R _24335_ (.A(_08337_),
    .B(_08965_),
    .C(_08967_),
    .Y(_08968_));
 OR3x1_ASAP7_75t_R _24336_ (.A(_08528_),
    .B(_08963_),
    .C(_08968_),
    .Y(_08969_));
 OR3x1_ASAP7_75t_R _24337_ (.A(_08448_),
    .B(_08388_),
    .C(_08393_),
    .Y(_08970_));
 AND3x1_ASAP7_75t_R _24338_ (.A(_08368_),
    .B(_08969_),
    .C(_08970_),
    .Y(_08971_));
 AO211x2_ASAP7_75t_R _24339_ (.A1(_08312_),
    .A2(_08727_),
    .B(_08971_),
    .C(_08308_),
    .Y(_08972_));
 OA21x2_ASAP7_75t_R _24340_ (.A1(_08513_),
    .A2(_08675_),
    .B(_08972_),
    .Y(_08973_));
 OA21x2_ASAP7_75t_R _24341_ (.A1(_08617_),
    .A2(_08680_),
    .B(_08590_),
    .Y(_08974_));
 INVx1_ASAP7_75t_R _24342_ (.A(_02297_),
    .Y(_08975_));
 OA222x2_ASAP7_75t_R _24343_ (.A1(_00277_),
    .A2(_08731_),
    .B1(_08732_),
    .B2(_08975_),
    .C1(_08558_),
    .C2(_00276_),
    .Y(_08976_));
 OAI21x1_ASAP7_75t_R _24344_ (.A1(_05226_),
    .A2(_08730_),
    .B(_08976_),
    .Y(_08977_));
 AOI211x1_ASAP7_75t_R _24345_ (.A1(_08512_),
    .A2(_08973_),
    .B(_08974_),
    .C(_08977_),
    .Y(_08978_));
 OA22x2_ASAP7_75t_R _24346_ (.A1(_00113_),
    .A2(_08567_),
    .B1(_08570_),
    .B2(_00109_),
    .Y(_08979_));
 OA211x2_ASAP7_75t_R _24347_ (.A1(_08880_),
    .A2(_08978_),
    .B(_08979_),
    .C(_06579_),
    .Y(_08980_));
 BUFx3_ASAP7_75t_R _24348_ (.A(_08790_),
    .Y(_08981_));
 BUFx6f_ASAP7_75t_R _24349_ (.A(_08787_),
    .Y(_08982_));
 AO221x1_ASAP7_75t_R _24350_ (.A1(net60),
    .A2(_08981_),
    .B1(_08982_),
    .B2(net30),
    .C(_08596_),
    .Y(_08983_));
 INVx1_ASAP7_75t_R _24351_ (.A(_01436_),
    .Y(_08984_));
 INVx1_ASAP7_75t_R _24352_ (.A(_01421_),
    .Y(_08985_));
 AO221x1_ASAP7_75t_R _24353_ (.A1(_08984_),
    .A2(_08981_),
    .B1(_08982_),
    .B2(_08985_),
    .C(_08286_),
    .Y(_08986_));
 NOR2x1_ASAP7_75t_R _24354_ (.A(_08602_),
    .B(_08279_),
    .Y(_08987_));
 NOR2x1_ASAP7_75t_R _24355_ (.A(_01427_),
    .B(_08799_),
    .Y(_08988_));
 AO21x1_ASAP7_75t_R _24356_ (.A1(net68),
    .A2(_05738_),
    .B(_08988_),
    .Y(_08989_));
 AO222x2_ASAP7_75t_R _24357_ (.A1(net74),
    .A2(_08796_),
    .B1(_08983_),
    .B2(_08986_),
    .C1(_08987_),
    .C2(_08989_),
    .Y(_08990_));
 NAND2x1_ASAP7_75t_R _24358_ (.A(_08504_),
    .B(_08990_),
    .Y(_08991_));
 OAI21x1_ASAP7_75t_R _24359_ (.A1(_08593_),
    .A2(_08980_),
    .B(_08991_),
    .Y(_08992_));
 BUFx12f_ASAP7_75t_R _24360_ (.A(_08992_),
    .Y(_08993_));
 BUFx6f_ASAP7_75t_R _24361_ (.A(_08955_),
    .Y(_08994_));
 NOR2x1_ASAP7_75t_R _24362_ (.A(_00506_),
    .B(_08994_),
    .Y(_08995_));
 AO21x1_ASAP7_75t_R _24363_ (.A1(_08956_),
    .A2(_08993_),
    .B(_08995_),
    .Y(_02849_));
 AND2x4_ASAP7_75t_R _24364_ (.A(_08460_),
    .B(_08511_),
    .Y(_08996_));
 OA211x2_ASAP7_75t_R _24365_ (.A1(_08555_),
    .A2(_08765_),
    .B(_08771_),
    .C(_08440_),
    .Y(_08997_));
 AOI21x1_ASAP7_75t_R _24366_ (.A1(_08764_),
    .A2(_08996_),
    .B(_08997_),
    .Y(_08998_));
 INVx1_ASAP7_75t_R _24367_ (.A(_02311_),
    .Y(_08999_));
 OA222x2_ASAP7_75t_R _24368_ (.A1(_00305_),
    .A2(_08731_),
    .B1(_08732_),
    .B2(_08999_),
    .C1(_08558_),
    .C2(_00304_),
    .Y(_09000_));
 NAND2x1_ASAP7_75t_R _24369_ (.A(\alu_adder_result_ex[18] ),
    .B(_08818_),
    .Y(_09001_));
 AO21x1_ASAP7_75t_R _24370_ (.A1(_09000_),
    .A2(_09001_),
    .B(_08880_),
    .Y(_09002_));
 OR3x1_ASAP7_75t_R _24371_ (.A(net1967),
    .B(_00194_),
    .C(_00199_),
    .Y(_09003_));
 OR2x2_ASAP7_75t_R _24372_ (.A(_00195_),
    .B(_00194_),
    .Y(_09004_));
 AO21x1_ASAP7_75t_R _24373_ (.A1(_00200_),
    .A2(_09004_),
    .B(_00199_),
    .Y(_09005_));
 OA31x2_ASAP7_75t_R _24374_ (.A1(_08807_),
    .A2(_08809_),
    .A3(_09003_),
    .B1(_09005_),
    .Y(_09006_));
 AO21x1_ASAP7_75t_R _24375_ (.A1(_00204_),
    .A2(_09006_),
    .B(_00203_),
    .Y(_09007_));
 AND2x2_ASAP7_75t_R _24376_ (.A(_00208_),
    .B(_09007_),
    .Y(_09008_));
 XNOR2x2_ASAP7_75t_R _24377_ (.A(_00207_),
    .B(_09008_),
    .Y(_09009_));
 AND2x2_ASAP7_75t_R _24378_ (.A(_00103_),
    .B(_08495_),
    .Y(_09010_));
 AO21x1_ASAP7_75t_R _24379_ (.A1(_08902_),
    .A2(_09009_),
    .B(_09010_),
    .Y(_09011_));
 AO21x1_ASAP7_75t_R _24380_ (.A1(_14534_),
    .A2(_09011_),
    .B(_08568_),
    .Y(_09012_));
 AO21x2_ASAP7_75t_R _24381_ (.A1(_16083_),
    .A2(_05721_),
    .B(_09012_),
    .Y(_09013_));
 AND4x1_ASAP7_75t_R _24382_ (.A(_06195_),
    .B(_08738_),
    .C(_09002_),
    .D(_09013_),
    .Y(_09014_));
 NAND2x1_ASAP7_75t_R _24383_ (.A(net57),
    .B(_08609_),
    .Y(_09015_));
 OA211x2_ASAP7_75t_R _24384_ (.A1(_01430_),
    .A2(_08606_),
    .B(_09015_),
    .C(_08602_),
    .Y(_09016_));
 NAND2x1_ASAP7_75t_R _24385_ (.A(net70),
    .B(_08274_),
    .Y(_09017_));
 OA211x2_ASAP7_75t_R _24386_ (.A1(_08658_),
    .A2(_08606_),
    .B(_09017_),
    .C(_08282_),
    .Y(_09018_));
 OR3x1_ASAP7_75t_R _24387_ (.A(_08286_),
    .B(_09016_),
    .C(_09018_),
    .Y(_09019_));
 AND3x4_ASAP7_75t_R _24388_ (.A(_08504_),
    .B(_08912_),
    .C(_09019_),
    .Y(_09020_));
 AOI21x1_ASAP7_75t_R _24389_ (.A1(_08998_),
    .A2(_09014_),
    .B(_09020_),
    .Y(_09021_));
 BUFx6f_ASAP7_75t_R _24390_ (.A(_09021_),
    .Y(_09022_));
 AND2x2_ASAP7_75t_R _24391_ (.A(_16042_),
    .B(_08509_),
    .Y(_09023_));
 AO21x1_ASAP7_75t_R _24392_ (.A1(_08265_),
    .A2(_09022_),
    .B(_09023_),
    .Y(_02850_));
 BUFx6f_ASAP7_75t_R _24393_ (.A(_08922_),
    .Y(_09024_));
 AND2x2_ASAP7_75t_R _24394_ (.A(net73),
    .B(_08606_),
    .Y(_09025_));
 AO21x1_ASAP7_75t_R _24395_ (.A1(net29),
    .A2(_08290_),
    .B(_09025_),
    .Y(_09026_));
 NAND2x1_ASAP7_75t_R _24396_ (.A(net58),
    .B(_08609_),
    .Y(_09027_));
 OA211x2_ASAP7_75t_R _24397_ (.A1(_01429_),
    .A2(_08606_),
    .B(_09027_),
    .C(_08602_),
    .Y(_09028_));
 INVx1_ASAP7_75t_R _24398_ (.A(_09028_),
    .Y(_09029_));
 OA211x2_ASAP7_75t_R _24399_ (.A1(_08271_),
    .A2(_09026_),
    .B(_09029_),
    .C(_08597_),
    .Y(_09030_));
 INVx1_ASAP7_75t_R _24400_ (.A(_02312_),
    .Y(_09031_));
 OA22x2_ASAP7_75t_R _24401_ (.A1(_00307_),
    .A2(_08559_),
    .B1(_08486_),
    .B2(_09031_),
    .Y(_09032_));
 OA21x2_ASAP7_75t_R _24402_ (.A1(_00306_),
    .A2(_08479_),
    .B(_09032_),
    .Y(_09033_));
 OAI22x1_ASAP7_75t_R _24403_ (.A1(_16253_),
    .A2(_08730_),
    .B1(_08480_),
    .B2(_09033_),
    .Y(_09034_));
 AO221x1_ASAP7_75t_R _24404_ (.A1(_08833_),
    .A2(_08729_),
    .B1(_08996_),
    .B2(_08724_),
    .C(_09034_),
    .Y(_09035_));
 AND2x2_ASAP7_75t_R _24405_ (.A(_08721_),
    .B(_09035_),
    .Y(_09036_));
 BUFx12f_ASAP7_75t_R _24406_ (.A(_08901_),
    .Y(_09037_));
 AND3x4_ASAP7_75t_R _24407_ (.A(_00204_),
    .B(_00208_),
    .C(_00211_),
    .Y(_09038_));
 AND3x1_ASAP7_75t_R _24408_ (.A(_00203_),
    .B(_00208_),
    .C(_00211_),
    .Y(_09039_));
 AO21x2_ASAP7_75t_R _24409_ (.A1(_00207_),
    .A2(_00211_),
    .B(_09039_),
    .Y(_09040_));
 AO21x1_ASAP7_75t_R _24410_ (.A1(_08937_),
    .A2(_09038_),
    .B(_09040_),
    .Y(_09041_));
 XOR2x2_ASAP7_75t_R _24411_ (.A(_00210_),
    .B(_09041_),
    .Y(_09042_));
 NOR2x1_ASAP7_75t_R _24412_ (.A(_00108_),
    .B(_08902_),
    .Y(_09043_));
 AO21x1_ASAP7_75t_R _24413_ (.A1(_08902_),
    .A2(_09042_),
    .B(_09043_),
    .Y(_09044_));
 NAND2x1_ASAP7_75t_R _24414_ (.A(_05241_),
    .B(_09044_),
    .Y(_09045_));
 OA211x2_ASAP7_75t_R _24415_ (.A1(_16195_),
    .A2(_09037_),
    .B(_06218_),
    .C(_09045_),
    .Y(_09046_));
 NAND2x1_ASAP7_75t_R _24416_ (.A(_08853_),
    .B(_09046_),
    .Y(_09047_));
 OA22x2_ASAP7_75t_R _24417_ (.A1(_09024_),
    .A2(_09030_),
    .B1(_09036_),
    .B2(_09047_),
    .Y(_09048_));
 BUFx6f_ASAP7_75t_R _24418_ (.A(_09048_),
    .Y(_09049_));
 BUFx6f_ASAP7_75t_R _24419_ (.A(_08508_),
    .Y(_09050_));
 AND2x2_ASAP7_75t_R _24420_ (.A(_16167_),
    .B(_09050_),
    .Y(_09051_));
 AO21x1_ASAP7_75t_R _24421_ (.A1(_08265_),
    .A2(_09049_),
    .B(_09051_),
    .Y(_02851_));
 BUFx6f_ASAP7_75t_R _24422_ (.A(_08264_),
    .Y(_09052_));
 INVx1_ASAP7_75t_R _24423_ (.A(_02313_),
    .Y(_09053_));
 OA222x2_ASAP7_75t_R _24424_ (.A1(_00309_),
    .A2(_08731_),
    .B1(_08732_),
    .B2(_09053_),
    .C1(_08558_),
    .C2(_00308_),
    .Y(_09054_));
 NAND2x1_ASAP7_75t_R _24425_ (.A(\alu_adder_result_ex[20] ),
    .B(_08818_),
    .Y(_09055_));
 AO21x1_ASAP7_75t_R _24426_ (.A1(_09054_),
    .A2(_09055_),
    .B(_08880_),
    .Y(_09056_));
 OR3x1_ASAP7_75t_R _24427_ (.A(_14534_),
    .B(_16329_),
    .C(_08568_),
    .Y(_09057_));
 AND4x1_ASAP7_75t_R _24428_ (.A(_06253_),
    .B(_08738_),
    .C(_09056_),
    .D(_09057_),
    .Y(_09058_));
 BUFx6f_ASAP7_75t_R _24429_ (.A(_08495_),
    .Y(_09059_));
 BUFx6f_ASAP7_75t_R _24430_ (.A(_09059_),
    .Y(_09060_));
 AO21x1_ASAP7_75t_R _24431_ (.A1(_09006_),
    .A2(_09038_),
    .B(_09040_),
    .Y(_09061_));
 OA21x2_ASAP7_75t_R _24432_ (.A1(_00210_),
    .A2(_09061_),
    .B(_00214_),
    .Y(_09062_));
 XOR2x2_ASAP7_75t_R _24433_ (.A(_00213_),
    .B(_09062_),
    .Y(_09063_));
 NAND2x1_ASAP7_75t_R _24434_ (.A(_00113_),
    .B(_09059_),
    .Y(_09064_));
 OA211x2_ASAP7_75t_R _24435_ (.A1(_09060_),
    .A2(_09063_),
    .B(_09064_),
    .C(_05242_),
    .Y(_09065_));
 AOI221x1_ASAP7_75t_R _24436_ (.A1(_08512_),
    .A2(_08676_),
    .B1(_08694_),
    .B2(_08440_),
    .C(_09065_),
    .Y(_09066_));
 OR2x2_ASAP7_75t_R _24437_ (.A(_01427_),
    .B(_08276_),
    .Y(_09067_));
 OA211x2_ASAP7_75t_R _24438_ (.A1(_08752_),
    .A2(_08289_),
    .B(_09067_),
    .C(_08602_),
    .Y(_09068_));
 INVx1_ASAP7_75t_R _24439_ (.A(net30),
    .Y(_09069_));
 NAND2x1_ASAP7_75t_R _24440_ (.A(net74),
    .B(_08274_),
    .Y(_09070_));
 OA211x2_ASAP7_75t_R _24441_ (.A1(_09069_),
    .A2(_08606_),
    .B(_09070_),
    .C(_08282_),
    .Y(_09071_));
 OR3x1_ASAP7_75t_R _24442_ (.A(_08286_),
    .B(_09068_),
    .C(_09071_),
    .Y(_09072_));
 AND3x4_ASAP7_75t_R _24443_ (.A(_08504_),
    .B(_08912_),
    .C(_09072_),
    .Y(_09073_));
 AOI21x1_ASAP7_75t_R _24444_ (.A1(_09058_),
    .A2(_09066_),
    .B(_09073_),
    .Y(_09074_));
 BUFx6f_ASAP7_75t_R _24445_ (.A(_09074_),
    .Y(_09075_));
 AND2x2_ASAP7_75t_R _24446_ (.A(_16302_),
    .B(_09050_),
    .Y(_09076_));
 AO21x1_ASAP7_75t_R _24447_ (.A1(_09052_),
    .A2(_09075_),
    .B(_09076_),
    .Y(_02852_));
 AND2x2_ASAP7_75t_R _24448_ (.A(net75),
    .B(_08606_),
    .Y(_09077_));
 AO21x1_ASAP7_75t_R _24449_ (.A1(net31),
    .A2(_08290_),
    .B(_09077_),
    .Y(_09078_));
 NAND2x1_ASAP7_75t_R _24450_ (.A(net61),
    .B(_08609_),
    .Y(_09079_));
 OA211x2_ASAP7_75t_R _24451_ (.A1(_01426_),
    .A2(_08606_),
    .B(_09079_),
    .C(_08602_),
    .Y(_09080_));
 INVx1_ASAP7_75t_R _24452_ (.A(_09080_),
    .Y(_09081_));
 OA211x2_ASAP7_75t_R _24453_ (.A1(_08271_),
    .A2(_09078_),
    .B(_09081_),
    .C(_08597_),
    .Y(_09082_));
 INVx1_ASAP7_75t_R _24454_ (.A(_06275_),
    .Y(_09083_));
 AND2x2_ASAP7_75t_R _24455_ (.A(_08833_),
    .B(_08642_),
    .Y(_09084_));
 INVx1_ASAP7_75t_R _24456_ (.A(_02314_),
    .Y(_09085_));
 OA222x2_ASAP7_75t_R _24457_ (.A1(_00311_),
    .A2(_08559_),
    .B1(_08486_),
    .B2(_09085_),
    .C1(_08489_),
    .C2(_00310_),
    .Y(_09086_));
 OAI21x1_ASAP7_75t_R _24458_ (.A1(_16515_),
    .A2(_08730_),
    .B(_09086_),
    .Y(_09087_));
 AO32x1_ASAP7_75t_R _24459_ (.A1(_14541_),
    .A2(_16452_),
    .A3(_14623_),
    .B1(_08721_),
    .B2(_09087_),
    .Y(_09088_));
 OR4x1_ASAP7_75t_R _24460_ (.A(_09083_),
    .B(_08835_),
    .C(_09084_),
    .D(_09088_),
    .Y(_09089_));
 OR2x2_ASAP7_75t_R _24461_ (.A(_00210_),
    .B(_00213_),
    .Y(_09090_));
 AO211x2_ASAP7_75t_R _24462_ (.A1(_08937_),
    .A2(_09038_),
    .B(_09040_),
    .C(_09090_),
    .Y(_09091_));
 OR2x2_ASAP7_75t_R _24463_ (.A(_00214_),
    .B(_00213_),
    .Y(_09092_));
 AND2x2_ASAP7_75t_R _24464_ (.A(_00217_),
    .B(_09092_),
    .Y(_09093_));
 NAND2x1_ASAP7_75t_R _24465_ (.A(_09091_),
    .B(_09093_),
    .Y(_09094_));
 XNOR2x2_ASAP7_75t_R _24466_ (.A(_00216_),
    .B(_09094_),
    .Y(_09095_));
 NAND2x1_ASAP7_75t_R _24467_ (.A(_00120_),
    .B(_09059_),
    .Y(_09096_));
 OA211x2_ASAP7_75t_R _24468_ (.A1(_09059_),
    .A2(_09095_),
    .B(_09096_),
    .C(_05241_),
    .Y(_09097_));
 AO21x1_ASAP7_75t_R _24469_ (.A1(_08512_),
    .A2(_08625_),
    .B(_09097_),
    .Y(_09098_));
 OA22x2_ASAP7_75t_R _24470_ (.A1(_09024_),
    .A2(_09082_),
    .B1(_09089_),
    .B2(_09098_),
    .Y(_09099_));
 BUFx6f_ASAP7_75t_R _24471_ (.A(_09099_),
    .Y(_09100_));
 AND2x2_ASAP7_75t_R _24472_ (.A(_16425_),
    .B(_09050_),
    .Y(_09101_));
 AO21x1_ASAP7_75t_R _24473_ (.A1(_09052_),
    .A2(_09100_),
    .B(_09101_),
    .Y(_02853_));
 AND2x2_ASAP7_75t_R _24474_ (.A(net76),
    .B(_08609_),
    .Y(_09102_));
 AO21x1_ASAP7_75t_R _24475_ (.A1(net53),
    .A2(_08290_),
    .B(_09102_),
    .Y(_09103_));
 NAND2x1_ASAP7_75t_R _24476_ (.A(net62),
    .B(_08609_),
    .Y(_09104_));
 OA211x2_ASAP7_75t_R _24477_ (.A1(_01425_),
    .A2(_08275_),
    .B(_09104_),
    .C(_08270_),
    .Y(_09105_));
 INVx1_ASAP7_75t_R _24478_ (.A(_09105_),
    .Y(_09106_));
 OA211x2_ASAP7_75t_R _24479_ (.A1(_08271_),
    .A2(_09103_),
    .B(_09106_),
    .C(_08597_),
    .Y(_09107_));
 OR3x1_ASAP7_75t_R _24480_ (.A(_00210_),
    .B(_00213_),
    .C(_00216_),
    .Y(_09108_));
 AO21x1_ASAP7_75t_R _24481_ (.A1(_00217_),
    .A2(_09092_),
    .B(_00216_),
    .Y(_09109_));
 OA21x2_ASAP7_75t_R _24482_ (.A1(_09061_),
    .A2(_09108_),
    .B(_09109_),
    .Y(_09110_));
 NAND2x1_ASAP7_75t_R _24483_ (.A(_00220_),
    .B(_09110_),
    .Y(_09111_));
 XNOR2x2_ASAP7_75t_R _24484_ (.A(_00219_),
    .B(_09111_),
    .Y(_09112_));
 NAND2x1_ASAP7_75t_R _24485_ (.A(_00127_),
    .B(_09059_),
    .Y(_09113_));
 OA211x2_ASAP7_75t_R _24486_ (.A1(_09059_),
    .A2(_09112_),
    .B(_09113_),
    .C(_05241_),
    .Y(_09114_));
 INVx1_ASAP7_75t_R _24487_ (.A(_02315_),
    .Y(_09115_));
 OA222x2_ASAP7_75t_R _24488_ (.A1(_00313_),
    .A2(_08485_),
    .B1(_08815_),
    .B2(_09115_),
    .C1(_08695_),
    .C2(_00312_),
    .Y(_09116_));
 OA21x2_ASAP7_75t_R _24489_ (.A1(_16761_),
    .A2(_08730_),
    .B(_09116_),
    .Y(_09117_));
 NOR2x1_ASAP7_75t_R _24490_ (.A(_08880_),
    .B(_09117_),
    .Y(_09118_));
 AO21x1_ASAP7_75t_R _24491_ (.A1(_08589_),
    .A2(_08996_),
    .B(_08592_),
    .Y(_09119_));
 AND3x1_ASAP7_75t_R _24492_ (.A(_08833_),
    .B(_08541_),
    .C(_08556_),
    .Y(_09120_));
 OAI21x1_ASAP7_75t_R _24493_ (.A1(_16591_),
    .A2(_09037_),
    .B(_06296_),
    .Y(_09121_));
 OR5x1_ASAP7_75t_R _24494_ (.A(_09114_),
    .B(_09118_),
    .C(_09119_),
    .D(_09120_),
    .E(_09121_),
    .Y(_09122_));
 OA21x2_ASAP7_75t_R _24495_ (.A1(_09024_),
    .A2(_09107_),
    .B(_09122_),
    .Y(_09123_));
 BUFx6f_ASAP7_75t_R _24496_ (.A(_09123_),
    .Y(_09124_));
 AND2x2_ASAP7_75t_R _24497_ (.A(_16563_),
    .B(_09050_),
    .Y(_09125_));
 AO21x1_ASAP7_75t_R _24498_ (.A1(_09052_),
    .A2(_09124_),
    .B(_09125_),
    .Y(_02854_));
 OA211x2_ASAP7_75t_R _24499_ (.A1(net54),
    .A2(_08275_),
    .B(_08299_),
    .C(_08287_),
    .Y(_09126_));
 INVx1_ASAP7_75t_R _24500_ (.A(_01424_),
    .Y(_09127_));
 OA211x2_ASAP7_75t_R _24501_ (.A1(_09127_),
    .A2(_08275_),
    .B(_08301_),
    .C(_08270_),
    .Y(_09128_));
 OA21x2_ASAP7_75t_R _24502_ (.A1(_09126_),
    .A2(_09128_),
    .B(_08597_),
    .Y(_09129_));
 AO21x1_ASAP7_75t_R _24503_ (.A1(_09091_),
    .A2(_09093_),
    .B(_00216_),
    .Y(_09130_));
 AO21x1_ASAP7_75t_R _24504_ (.A1(_00220_),
    .A2(_09130_),
    .B(_00219_),
    .Y(_09131_));
 NAND2x1_ASAP7_75t_R _24505_ (.A(_00223_),
    .B(_09131_),
    .Y(_09132_));
 XNOR2x2_ASAP7_75t_R _24506_ (.A(_00222_),
    .B(_09132_),
    .Y(_09133_));
 OR2x2_ASAP7_75t_R _24507_ (.A(_02209_),
    .B(_08498_),
    .Y(_09134_));
 OA211x2_ASAP7_75t_R _24508_ (.A1(_09059_),
    .A2(_09133_),
    .B(_09134_),
    .C(_05241_),
    .Y(_09135_));
 INVx1_ASAP7_75t_R _24509_ (.A(_02316_),
    .Y(_09136_));
 OA222x2_ASAP7_75t_R _24510_ (.A1(_00315_),
    .A2(_08485_),
    .B1(_08815_),
    .B2(_09136_),
    .C1(_08695_),
    .C2(_00314_),
    .Y(_09137_));
 OA21x2_ASAP7_75t_R _24511_ (.A1(_16753_),
    .A2(_08730_),
    .B(_09137_),
    .Y(_09138_));
 OAI22x1_ASAP7_75t_R _24512_ (.A1(_16701_),
    .A2(_09037_),
    .B1(_08880_),
    .B2(_09138_),
    .Y(_09139_));
 AND3x1_ASAP7_75t_R _24513_ (.A(_08833_),
    .B(_08397_),
    .C(_08432_),
    .Y(_09140_));
 NAND2x1_ASAP7_75t_R _24514_ (.A(_08464_),
    .B(_08511_),
    .Y(_09141_));
 NAND2x1_ASAP7_75t_R _24515_ (.A(_06322_),
    .B(_09141_),
    .Y(_09142_));
 OR5x1_ASAP7_75t_R _24516_ (.A(_08593_),
    .B(_09135_),
    .C(_09139_),
    .D(_09140_),
    .E(_09142_),
    .Y(_09143_));
 OA21x2_ASAP7_75t_R _24517_ (.A1(_09024_),
    .A2(_09129_),
    .B(_09143_),
    .Y(_09144_));
 BUFx6f_ASAP7_75t_R _24518_ (.A(_09144_),
    .Y(_09145_));
 AND2x2_ASAP7_75t_R _24519_ (.A(_16673_),
    .B(_09050_),
    .Y(_09146_));
 AO21x1_ASAP7_75t_R _24520_ (.A1(_09052_),
    .A2(_09145_),
    .B(_09146_),
    .Y(_02855_));
 OA211x2_ASAP7_75t_R _24521_ (.A1(_08293_),
    .A2(_08275_),
    .B(_08277_),
    .C(_08287_),
    .Y(_09147_));
 AOI211x1_ASAP7_75t_R _24522_ (.A1(_08271_),
    .A2(_08292_),
    .B(_08286_),
    .C(_09147_),
    .Y(_09148_));
 AND3x1_ASAP7_75t_R _24523_ (.A(_00220_),
    .B(_00223_),
    .C(_00226_),
    .Y(_09149_));
 AND3x1_ASAP7_75t_R _24524_ (.A(_00219_),
    .B(_00223_),
    .C(_00226_),
    .Y(_09150_));
 AO21x1_ASAP7_75t_R _24525_ (.A1(_00222_),
    .A2(_00226_),
    .B(_09150_),
    .Y(_09151_));
 AO21x2_ASAP7_75t_R _24526_ (.A1(_09110_),
    .A2(_09149_),
    .B(_09151_),
    .Y(_09152_));
 XOR2x2_ASAP7_75t_R _24527_ (.A(_00225_),
    .B(_09152_),
    .Y(_09153_));
 NAND2x1_ASAP7_75t_R _24528_ (.A(_08495_),
    .B(_08496_),
    .Y(_09154_));
 OA211x2_ASAP7_75t_R _24529_ (.A1(_09059_),
    .A2(_09153_),
    .B(_09154_),
    .C(_05241_),
    .Y(_09155_));
 OR3x1_ASAP7_75t_R _24530_ (.A(_08328_),
    .B(_08960_),
    .C(_08961_),
    .Y(_09156_));
 AO211x2_ASAP7_75t_R _24531_ (.A1(_18592_),
    .A2(_08349_),
    .B(_08389_),
    .C(_13452_),
    .Y(_09157_));
 AND3x1_ASAP7_75t_R _24532_ (.A(_08337_),
    .B(_09156_),
    .C(_09157_),
    .Y(_09158_));
 AO21x1_ASAP7_75t_R _24533_ (.A1(_08320_),
    .A2(_08517_),
    .B(_09158_),
    .Y(_09159_));
 OR3x1_ASAP7_75t_R _24534_ (.A(_08347_),
    .B(_08686_),
    .C(_08687_),
    .Y(_09160_));
 OA21x2_ASAP7_75t_R _24535_ (.A1(_08316_),
    .A2(_09159_),
    .B(_09160_),
    .Y(_09161_));
 OR3x1_ASAP7_75t_R _24536_ (.A(_08723_),
    .B(_08874_),
    .C(_08875_),
    .Y(_09162_));
 OA22x2_ASAP7_75t_R _24537_ (.A1(_08427_),
    .A2(_08463_),
    .B1(_08426_),
    .B2(_08454_),
    .Y(_09163_));
 OA211x2_ASAP7_75t_R _24538_ (.A1(_08457_),
    .A2(_09161_),
    .B(_09162_),
    .C(_09163_),
    .Y(_09164_));
 NOR2x2_ASAP7_75t_R _24539_ (.A(_08456_),
    .B(_08458_),
    .Y(_09165_));
 AOI21x1_ASAP7_75t_R _24540_ (.A1(_08456_),
    .A2(_08425_),
    .B(_09165_),
    .Y(_09166_));
 NAND2x1_ASAP7_75t_R _24541_ (.A(_08434_),
    .B(_09166_),
    .Y(_09167_));
 OA211x2_ASAP7_75t_R _24542_ (.A1(_08434_),
    .A2(_09164_),
    .B(_09167_),
    .C(_08437_),
    .Y(_09168_));
 NAND2x2_ASAP7_75t_R _24543_ (.A(_08568_),
    .B(_08818_),
    .Y(_09169_));
 NOR2x1_ASAP7_75t_R _24544_ (.A(_04246_),
    .B(_09169_),
    .Y(_09170_));
 INVx1_ASAP7_75t_R _24545_ (.A(_02317_),
    .Y(_09171_));
 OA222x2_ASAP7_75t_R _24546_ (.A1(_00317_),
    .A2(_08485_),
    .B1(_08815_),
    .B2(_09171_),
    .C1(_08489_),
    .C2(_00316_),
    .Y(_09172_));
 OA22x2_ASAP7_75t_R _24547_ (.A1(_16823_),
    .A2(_08901_),
    .B1(_08482_),
    .B2(_09172_),
    .Y(_09173_));
 NAND2x1_ASAP7_75t_R _24548_ (.A(_06342_),
    .B(_09173_),
    .Y(_09174_));
 OR5x1_ASAP7_75t_R _24549_ (.A(_08593_),
    .B(_09155_),
    .C(_09168_),
    .D(_09170_),
    .E(_09174_),
    .Y(_09175_));
 OA21x2_ASAP7_75t_R _24550_ (.A1(_09024_),
    .A2(_09148_),
    .B(_09175_),
    .Y(_09176_));
 BUFx6f_ASAP7_75t_R _24551_ (.A(_09176_),
    .Y(_09177_));
 AND2x2_ASAP7_75t_R _24552_ (.A(_16796_),
    .B(_09050_),
    .Y(_09178_));
 AO21x1_ASAP7_75t_R _24553_ (.A1(_09052_),
    .A2(_09177_),
    .B(_09178_),
    .Y(_02856_));
 NAND2x1_ASAP7_75t_R _24554_ (.A(_08605_),
    .B(_08610_),
    .Y(_09179_));
 OA211x2_ASAP7_75t_R _24555_ (.A1(_08271_),
    .A2(_08607_),
    .B(_09179_),
    .C(_08597_),
    .Y(_09180_));
 AO21x1_ASAP7_75t_R _24556_ (.A1(_09130_),
    .A2(_09149_),
    .B(_09151_),
    .Y(_09181_));
 OA21x2_ASAP7_75t_R _24557_ (.A1(_00225_),
    .A2(_09181_),
    .B(_00229_),
    .Y(_09182_));
 XOR2x2_ASAP7_75t_R _24558_ (.A(_00228_),
    .B(_09182_),
    .Y(_09183_));
 NAND2x1_ASAP7_75t_R _24559_ (.A(_08495_),
    .B(_08565_),
    .Y(_09184_));
 OA211x2_ASAP7_75t_R _24560_ (.A1(_09059_),
    .A2(_09183_),
    .B(_09184_),
    .C(_05241_),
    .Y(_09185_));
 OA211x2_ASAP7_75t_R _24561_ (.A1(_08514_),
    .A2(_08628_),
    .B(_08823_),
    .C(_08311_),
    .Y(_09186_));
 OA211x2_ASAP7_75t_R _24562_ (.A1(_05930_),
    .A2(_08390_),
    .B(_08392_),
    .C(_08445_),
    .Y(_09187_));
 AND3x1_ASAP7_75t_R _24563_ (.A(_08357_),
    .B(_08959_),
    .C(_08962_),
    .Y(_09188_));
 OR3x1_ASAP7_75t_R _24564_ (.A(_08316_),
    .B(_09187_),
    .C(_09188_),
    .Y(_09189_));
 OR3x1_ASAP7_75t_R _24565_ (.A(_08514_),
    .B(_08631_),
    .C(_08632_),
    .Y(_09190_));
 AND3x1_ASAP7_75t_R _24566_ (.A(_08368_),
    .B(_09189_),
    .C(_09190_),
    .Y(_09191_));
 OR3x1_ASAP7_75t_R _24567_ (.A(_08308_),
    .B(_09186_),
    .C(_09191_),
    .Y(_09192_));
 OAI21x1_ASAP7_75t_R _24568_ (.A1(_08513_),
    .A2(_08588_),
    .B(_09192_),
    .Y(_09193_));
 AO21x1_ASAP7_75t_R _24569_ (.A1(_08456_),
    .A2(_08539_),
    .B(_09165_),
    .Y(_09194_));
 OAI21x1_ASAP7_75t_R _24570_ (.A1(_08833_),
    .A2(_09194_),
    .B(_08437_),
    .Y(_09195_));
 AOI21x1_ASAP7_75t_R _24571_ (.A1(_08440_),
    .A2(_09193_),
    .B(_09195_),
    .Y(_09196_));
 INVx1_ASAP7_75t_R _24572_ (.A(_02318_),
    .Y(_09197_));
 OA222x2_ASAP7_75t_R _24573_ (.A1(_00319_),
    .A2(_08559_),
    .B1(_08478_),
    .B2(_09197_),
    .C1(_08488_),
    .C2(_00318_),
    .Y(_09198_));
 OA21x2_ASAP7_75t_R _24574_ (.A1(_16995_),
    .A2(_08484_),
    .B(_09198_),
    .Y(_09199_));
 OA22x2_ASAP7_75t_R _24575_ (.A1(_16935_),
    .A2(_08901_),
    .B1(_08483_),
    .B2(_09199_),
    .Y(_09200_));
 NAND2x1_ASAP7_75t_R _24576_ (.A(_06365_),
    .B(_09200_),
    .Y(_09201_));
 OR4x1_ASAP7_75t_R _24577_ (.A(_08593_),
    .B(_09185_),
    .C(_09196_),
    .D(_09201_),
    .Y(_09202_));
 OA21x2_ASAP7_75t_R _24578_ (.A1(_09024_),
    .A2(_09180_),
    .B(_09202_),
    .Y(_09203_));
 BUFx6f_ASAP7_75t_R _24579_ (.A(_09203_),
    .Y(_09204_));
 AND2x2_ASAP7_75t_R _24580_ (.A(_16895_),
    .B(_09050_),
    .Y(_09205_));
 AO21x1_ASAP7_75t_R _24581_ (.A1(_09052_),
    .A2(_09204_),
    .B(_09205_),
    .Y(_02857_));
 NAND2x1_ASAP7_75t_R _24582_ (.A(_08605_),
    .B(_08657_),
    .Y(_09206_));
 OA211x2_ASAP7_75t_R _24583_ (.A1(_08271_),
    .A2(_08660_),
    .B(_09206_),
    .C(_08597_),
    .Y(_09207_));
 OA21x2_ASAP7_75t_R _24584_ (.A1(_00225_),
    .A2(_09152_),
    .B(_00229_),
    .Y(_09208_));
 OA21x2_ASAP7_75t_R _24585_ (.A1(_00228_),
    .A2(_09208_),
    .B(_00232_),
    .Y(_09209_));
 XNOR2x2_ASAP7_75t_R _24586_ (.A(_00231_),
    .B(_09209_),
    .Y(_09210_));
 NAND2x1_ASAP7_75t_R _24587_ (.A(_08902_),
    .B(_09210_),
    .Y(_09211_));
 OA211x2_ASAP7_75t_R _24588_ (.A1(_08902_),
    .A2(_08649_),
    .B(_09211_),
    .C(_05241_),
    .Y(_09212_));
 AND3x1_ASAP7_75t_R _24589_ (.A(_08348_),
    .B(_09156_),
    .C(_09157_),
    .Y(_09213_));
 AO211x2_ASAP7_75t_R _24590_ (.A1(_18685_),
    .A2(_08352_),
    .B(_08966_),
    .C(_05930_),
    .Y(_09214_));
 OR3x1_ASAP7_75t_R _24591_ (.A(_13452_),
    .B(_08957_),
    .C(_08958_),
    .Y(_09215_));
 AND3x1_ASAP7_75t_R _24592_ (.A(_08357_),
    .B(_09214_),
    .C(_09215_),
    .Y(_09216_));
 NOR3x1_ASAP7_75t_R _24593_ (.A(_08316_),
    .B(_09213_),
    .C(_09216_),
    .Y(_09217_));
 AOI21x1_ASAP7_75t_R _24594_ (.A1(_08316_),
    .A2(_08521_),
    .B(_09217_),
    .Y(_09218_));
 OA222x2_ASAP7_75t_R _24595_ (.A1(_08513_),
    .A2(_08624_),
    .B1(_08723_),
    .B2(_08769_),
    .C1(_09218_),
    .C2(_08457_),
    .Y(_09219_));
 AOI21x1_ASAP7_75t_R _24596_ (.A1(_08456_),
    .A2(_08640_),
    .B(_09165_),
    .Y(_09220_));
 NAND2x1_ASAP7_75t_R _24597_ (.A(_08434_),
    .B(_09220_),
    .Y(_09221_));
 OA211x2_ASAP7_75t_R _24598_ (.A1(_08434_),
    .A2(_09219_),
    .B(_09221_),
    .C(_08437_),
    .Y(_09222_));
 INVx1_ASAP7_75t_R _24599_ (.A(_02319_),
    .Y(_09223_));
 OA222x2_ASAP7_75t_R _24600_ (.A1(_00321_),
    .A2(_08485_),
    .B1(_08815_),
    .B2(_09223_),
    .C1(_08695_),
    .C2(_00320_),
    .Y(_09224_));
 OA21x2_ASAP7_75t_R _24601_ (.A1(_04495_),
    .A2(_08730_),
    .B(_09224_),
    .Y(_09225_));
 NOR2x1_ASAP7_75t_R _24602_ (.A(_08880_),
    .B(_09225_),
    .Y(_09226_));
 OAI21x1_ASAP7_75t_R _24603_ (.A1(_04310_),
    .A2(_08901_),
    .B(_06389_),
    .Y(_09227_));
 OR5x1_ASAP7_75t_R _24604_ (.A(_08593_),
    .B(_09212_),
    .C(_09222_),
    .D(_09226_),
    .E(_09227_),
    .Y(_09228_));
 OA21x2_ASAP7_75t_R _24605_ (.A1(_09024_),
    .A2(_09207_),
    .B(_09228_),
    .Y(_09229_));
 BUFx6f_ASAP7_75t_R _24606_ (.A(_09229_),
    .Y(_09230_));
 AND2x2_ASAP7_75t_R _24607_ (.A(_04281_),
    .B(_09050_),
    .Y(_09231_));
 AO21x1_ASAP7_75t_R _24608_ (.A1(_09052_),
    .A2(_09230_),
    .B(_09231_),
    .Y(_02858_));
 NAND2x1_ASAP7_75t_R _24609_ (.A(_08605_),
    .B(_08708_),
    .Y(_09232_));
 OA211x2_ASAP7_75t_R _24610_ (.A1(_08271_),
    .A2(_08710_),
    .B(_09232_),
    .C(_08597_),
    .Y(_09233_));
 OR3x1_ASAP7_75t_R _24611_ (.A(_00225_),
    .B(_00228_),
    .C(_00231_),
    .Y(_09234_));
 OA21x2_ASAP7_75t_R _24612_ (.A1(_00229_),
    .A2(_00228_),
    .B(_00232_),
    .Y(_09235_));
 OA22x2_ASAP7_75t_R _24613_ (.A1(_09181_),
    .A2(_09234_),
    .B1(_09235_),
    .B2(_00231_),
    .Y(_09236_));
 NAND2x1_ASAP7_75t_R _24614_ (.A(_00235_),
    .B(_09236_),
    .Y(_09237_));
 XNOR2x2_ASAP7_75t_R _24615_ (.A(_00234_),
    .B(_09237_),
    .Y(_09238_));
 NAND2x1_ASAP7_75t_R _24616_ (.A(_09060_),
    .B(_08701_),
    .Y(_09239_));
 OA211x2_ASAP7_75t_R _24617_ (.A1(_09060_),
    .A2(_09238_),
    .B(_09239_),
    .C(_05242_),
    .Y(_09240_));
 AND2x2_ASAP7_75t_R _24618_ (.A(_08833_),
    .B(_08973_),
    .Y(_09241_));
 NOR2x1_ASAP7_75t_R _24619_ (.A(_04480_),
    .B(_09169_),
    .Y(_09242_));
 INVx1_ASAP7_75t_R _24620_ (.A(_02320_),
    .Y(_09243_));
 OA222x2_ASAP7_75t_R _24621_ (.A1(_00323_),
    .A2(_08731_),
    .B1(_08732_),
    .B2(_09243_),
    .C1(_08695_),
    .C2(_00322_),
    .Y(_09244_));
 OAI22x1_ASAP7_75t_R _24622_ (.A1(_04422_),
    .A2(_08901_),
    .B1(_08880_),
    .B2(_09244_),
    .Y(_09245_));
 OAI21x1_ASAP7_75t_R _24623_ (.A1(_08617_),
    .A2(_08680_),
    .B(_08996_),
    .Y(_09246_));
 NAND2x1_ASAP7_75t_R _24624_ (.A(_06410_),
    .B(_09246_),
    .Y(_09247_));
 OR5x1_ASAP7_75t_R _24625_ (.A(_08835_),
    .B(_09241_),
    .C(_09242_),
    .D(_09245_),
    .E(_09247_),
    .Y(_09248_));
 OA22x2_ASAP7_75t_R _24626_ (.A1(_09024_),
    .A2(_09233_),
    .B1(_09240_),
    .B2(_09248_),
    .Y(_09249_));
 BUFx6f_ASAP7_75t_R _24627_ (.A(_09249_),
    .Y(_09250_));
 AND2x2_ASAP7_75t_R _24628_ (.A(_04394_),
    .B(_09050_),
    .Y(_09251_));
 AO21x1_ASAP7_75t_R _24629_ (.A1(_09052_),
    .A2(_09250_),
    .B(_09251_),
    .Y(_02859_));
 AO221x1_ASAP7_75t_R _24630_ (.A1(net61),
    .A2(_08981_),
    .B1(_08982_),
    .B2(net31),
    .C(_08596_),
    .Y(_09252_));
 INVx1_ASAP7_75t_R _24631_ (.A(_01420_),
    .Y(_09253_));
 AO221x1_ASAP7_75t_R _24632_ (.A1(_08791_),
    .A2(_08981_),
    .B1(_08982_),
    .B2(_09253_),
    .C(_08286_),
    .Y(_09254_));
 INVx1_ASAP7_75t_R _24633_ (.A(net69),
    .Y(_09255_));
 OAI22x1_ASAP7_75t_R _24634_ (.A1(_09255_),
    .A2(_08298_),
    .B1(_08799_),
    .B2(_01426_),
    .Y(_09256_));
 AO222x2_ASAP7_75t_R _24635_ (.A1(net75),
    .A2(_08796_),
    .B1(_09252_),
    .B2(_09254_),
    .C1(_09256_),
    .C2(_08987_),
    .Y(_09257_));
 INVx1_ASAP7_75t_R _24636_ (.A(_06599_),
    .Y(_09258_));
 NAND2x1_ASAP7_75t_R _24637_ (.A(_08439_),
    .B(_09220_),
    .Y(_09259_));
 OA211x2_ASAP7_75t_R _24638_ (.A1(_08833_),
    .A2(_09219_),
    .B(_09259_),
    .C(_08437_),
    .Y(_09260_));
 INVx1_ASAP7_75t_R _24639_ (.A(_02298_),
    .Y(_09261_));
 OA222x2_ASAP7_75t_R _24640_ (.A1(_00279_),
    .A2(_08485_),
    .B1(_08815_),
    .B2(_09261_),
    .C1(_05212_),
    .C2(_08484_),
    .Y(_09262_));
 OAI21x1_ASAP7_75t_R _24641_ (.A1(_00278_),
    .A2(_08558_),
    .B(_09262_),
    .Y(_09263_));
 OAI22x1_ASAP7_75t_R _24642_ (.A1(_00120_),
    .A2(_08567_),
    .B1(_08570_),
    .B2(_00114_),
    .Y(_09264_));
 AO21x1_ASAP7_75t_R _24643_ (.A1(_08721_),
    .A2(_09263_),
    .B(_09264_),
    .Y(_09265_));
 OR4x1_ASAP7_75t_R _24644_ (.A(_09258_),
    .B(_08593_),
    .C(_09260_),
    .D(_09265_),
    .Y(_09266_));
 OA21x2_ASAP7_75t_R _24645_ (.A1(_08853_),
    .A2(_09257_),
    .B(_09266_),
    .Y(_09267_));
 BUFx12f_ASAP7_75t_R _24646_ (.A(_09267_),
    .Y(_09268_));
 NOR2x1_ASAP7_75t_R _24647_ (.A(_00536_),
    .B(_08994_),
    .Y(_09269_));
 AO21x1_ASAP7_75t_R _24648_ (.A1(_08956_),
    .A2(_09268_),
    .B(_09269_),
    .Y(_02860_));
 OR4x1_ASAP7_75t_R _24649_ (.A(_00225_),
    .B(_00228_),
    .C(_00231_),
    .D(_00234_),
    .Y(_09270_));
 OA21x2_ASAP7_75t_R _24650_ (.A1(_00232_),
    .A2(_00231_),
    .B(_00235_),
    .Y(_09271_));
 OR4x1_ASAP7_75t_R _24651_ (.A(_00229_),
    .B(_00228_),
    .C(_00231_),
    .D(_00234_),
    .Y(_09272_));
 OA211x2_ASAP7_75t_R _24652_ (.A1(_00234_),
    .A2(_09271_),
    .B(_09272_),
    .C(_00238_),
    .Y(_09273_));
 OA21x2_ASAP7_75t_R _24653_ (.A1(_09152_),
    .A2(_09270_),
    .B(_09273_),
    .Y(_09274_));
 XOR2x2_ASAP7_75t_R _24654_ (.A(_00237_),
    .B(_09274_),
    .Y(_09275_));
 OR2x2_ASAP7_75t_R _24655_ (.A(_08902_),
    .B(_08741_),
    .Y(_09276_));
 OA211x2_ASAP7_75t_R _24656_ (.A1(_09060_),
    .A2(_09275_),
    .B(_09276_),
    .C(_05242_),
    .Y(_09277_));
 AND2x2_ASAP7_75t_R _24657_ (.A(_08311_),
    .B(_08678_),
    .Y(_09278_));
 AO211x2_ASAP7_75t_R _24658_ (.A1(_08555_),
    .A2(_08685_),
    .B(_09278_),
    .C(_08513_),
    .Y(_09279_));
 OA21x2_ASAP7_75t_R _24659_ (.A1(_08688_),
    .A2(_08691_),
    .B(_08311_),
    .Y(_09280_));
 AND2x2_ASAP7_75t_R _24660_ (.A(_18695_),
    .B(_08352_),
    .Y(_09281_));
 AND2x4_ASAP7_75t_R _24661_ (.A(_18567_),
    .B(_08323_),
    .Y(_09282_));
 AO211x2_ASAP7_75t_R _24662_ (.A1(_18572_),
    .A2(_08349_),
    .B(_08964_),
    .C(_13452_),
    .Y(_09283_));
 OA31x2_ASAP7_75t_R _24663_ (.A1(_18555_),
    .A2(_09281_),
    .A3(_09282_),
    .B1(_09283_),
    .Y(_09284_));
 AND3x1_ASAP7_75t_R _24664_ (.A(_08348_),
    .B(_09214_),
    .C(_09215_),
    .Y(_09285_));
 AO211x2_ASAP7_75t_R _24665_ (.A1(_08337_),
    .A2(_09284_),
    .B(_09285_),
    .C(_08528_),
    .Y(_09286_));
 OA211x2_ASAP7_75t_R _24666_ (.A1(_08514_),
    .A2(_09159_),
    .B(_09286_),
    .C(_08367_),
    .Y(_09287_));
 OR3x1_ASAP7_75t_R _24667_ (.A(_08308_),
    .B(_09280_),
    .C(_09287_),
    .Y(_09288_));
 AND3x1_ASAP7_75t_R _24668_ (.A(_08833_),
    .B(_09279_),
    .C(_09288_),
    .Y(_09289_));
 AO21x1_ASAP7_75t_R _24669_ (.A1(_08456_),
    .A2(_08673_),
    .B(_09165_),
    .Y(_09290_));
 AND2x2_ASAP7_75t_R _24670_ (.A(_08511_),
    .B(_09290_),
    .Y(_09291_));
 INVx1_ASAP7_75t_R _24671_ (.A(_02321_),
    .Y(_09292_));
 OA222x2_ASAP7_75t_R _24672_ (.A1(_00325_),
    .A2(_08559_),
    .B1(_08486_),
    .B2(_09292_),
    .C1(_08489_),
    .C2(_00324_),
    .Y(_09293_));
 OA22x2_ASAP7_75t_R _24673_ (.A1(_04558_),
    .A2(_08901_),
    .B1(_08482_),
    .B2(_09293_),
    .Y(_09294_));
 NAND2x1_ASAP7_75t_R _24674_ (.A(_06431_),
    .B(_09294_),
    .Y(_09295_));
 NOR2x1_ASAP7_75t_R _24675_ (.A(_04729_),
    .B(_09169_),
    .Y(_09296_));
 OR5x2_ASAP7_75t_R _24676_ (.A(_08835_),
    .B(_09289_),
    .C(_09291_),
    .D(_09295_),
    .E(_09296_),
    .Y(_09297_));
 NOR2x1_ASAP7_75t_R _24677_ (.A(_08605_),
    .B(_08753_),
    .Y(_09298_));
 AO21x1_ASAP7_75t_R _24678_ (.A1(_08605_),
    .A2(_08750_),
    .B(_09298_),
    .Y(_09299_));
 AO21x2_ASAP7_75t_R _24679_ (.A1(_08597_),
    .A2(_09299_),
    .B(_08922_),
    .Y(_09300_));
 OA21x2_ASAP7_75t_R _24680_ (.A1(_09277_),
    .A2(_09297_),
    .B(_09300_),
    .Y(_09301_));
 BUFx6f_ASAP7_75t_R _24681_ (.A(_09301_),
    .Y(_09302_));
 AND2x2_ASAP7_75t_R _24682_ (.A(_04518_),
    .B(_09050_),
    .Y(_09303_));
 AO21x1_ASAP7_75t_R _24683_ (.A1(_09052_),
    .A2(_09302_),
    .B(_09303_),
    .Y(_02861_));
 AND2x2_ASAP7_75t_R _24684_ (.A(net31),
    .B(_08279_),
    .Y(_09304_));
 AO21x1_ASAP7_75t_R _24685_ (.A1(net61),
    .A2(_08290_),
    .B(_09304_),
    .Y(_09305_));
 OA211x2_ASAP7_75t_R _24686_ (.A1(_09255_),
    .A2(_08290_),
    .B(_08794_),
    .C(_08602_),
    .Y(_09306_));
 INVx1_ASAP7_75t_R _24687_ (.A(_09306_),
    .Y(_09307_));
 OA211x2_ASAP7_75t_R _24688_ (.A1(_08271_),
    .A2(_09305_),
    .B(_09307_),
    .C(_08596_),
    .Y(_09308_));
 AND4x1_ASAP7_75t_R _24689_ (.A(_00235_),
    .B(_00238_),
    .C(_00241_),
    .D(_09236_),
    .Y(_09309_));
 AND3x1_ASAP7_75t_R _24690_ (.A(_00234_),
    .B(_00238_),
    .C(_00241_),
    .Y(_09310_));
 AO21x1_ASAP7_75t_R _24691_ (.A1(_00237_),
    .A2(_00241_),
    .B(_09310_),
    .Y(_09311_));
 NOR2x1_ASAP7_75t_R _24692_ (.A(_09309_),
    .B(_09311_),
    .Y(_09312_));
 XNOR2x2_ASAP7_75t_R _24693_ (.A(_00240_),
    .B(_09312_),
    .Y(_09313_));
 NAND2x1_ASAP7_75t_R _24694_ (.A(_09060_),
    .B(_08780_),
    .Y(_09314_));
 OA211x2_ASAP7_75t_R _24695_ (.A1(_09060_),
    .A2(_09313_),
    .B(_09314_),
    .C(_05242_),
    .Y(_09315_));
 INVx1_ASAP7_75t_R _24696_ (.A(_06453_),
    .Y(_09316_));
 AND2x4_ASAP7_75t_R _24697_ (.A(_08307_),
    .B(_08310_),
    .Y(_09317_));
 OR3x1_ASAP7_75t_R _24698_ (.A(_08448_),
    .B(_09187_),
    .C(_09188_),
    .Y(_09318_));
 AND3x1_ASAP7_75t_R _24699_ (.A(_04666_),
    .B(_04669_),
    .C(_08326_),
    .Y(_09319_));
 AO211x2_ASAP7_75t_R _24700_ (.A1(_18562_),
    .A2(_08323_),
    .B(_09319_),
    .C(_08328_),
    .Y(_09320_));
 OA31x2_ASAP7_75t_R _24701_ (.A1(_08409_),
    .A2(_09281_),
    .A3(_09282_),
    .B1(_09320_),
    .Y(_09321_));
 AND3x1_ASAP7_75t_R _24702_ (.A(_08348_),
    .B(_08965_),
    .C(_08967_),
    .Y(_09322_));
 AO211x2_ASAP7_75t_R _24703_ (.A1(_08337_),
    .A2(_09321_),
    .B(_09322_),
    .C(_08315_),
    .Y(_09323_));
 AO33x2_ASAP7_75t_R _24704_ (.A1(_08633_),
    .A2(_08636_),
    .A3(_08722_),
    .B1(_09318_),
    .B2(_09323_),
    .B3(_08455_),
    .Y(_09324_));
 AO221x1_ASAP7_75t_R _24705_ (.A1(_08725_),
    .A2(_08630_),
    .B1(_08640_),
    .B2(_09317_),
    .C(_09324_),
    .Y(_09325_));
 AND2x2_ASAP7_75t_R _24706_ (.A(_08456_),
    .B(_08622_),
    .Y(_09326_));
 OR3x1_ASAP7_75t_R _24707_ (.A(_08439_),
    .B(_09165_),
    .C(_09326_),
    .Y(_09327_));
 OA211x2_ASAP7_75t_R _24708_ (.A1(_08434_),
    .A2(_09325_),
    .B(_09327_),
    .C(_08437_),
    .Y(_09328_));
 NOR2x1_ASAP7_75t_R _24709_ (.A(_04722_),
    .B(_09169_),
    .Y(_09329_));
 INVx1_ASAP7_75t_R _24710_ (.A(_02322_),
    .Y(_09330_));
 OA222x2_ASAP7_75t_R _24711_ (.A1(_00327_),
    .A2(_08731_),
    .B1(_08732_),
    .B2(_09330_),
    .C1(_08695_),
    .C2(_00326_),
    .Y(_09331_));
 OAI22x1_ASAP7_75t_R _24712_ (.A1(_04670_),
    .A2(_08901_),
    .B1(_08483_),
    .B2(_09331_),
    .Y(_09332_));
 OR5x1_ASAP7_75t_R _24713_ (.A(_09316_),
    .B(_08835_),
    .C(_09328_),
    .D(_09329_),
    .E(_09332_),
    .Y(_09333_));
 OA22x2_ASAP7_75t_R _24714_ (.A1(_09024_),
    .A2(_09308_),
    .B1(_09315_),
    .B2(_09333_),
    .Y(_09334_));
 BUFx6f_ASAP7_75t_R _24715_ (.A(_09334_),
    .Y(_09335_));
 AND2x2_ASAP7_75t_R _24716_ (.A(_04642_),
    .B(_08508_),
    .Y(_09336_));
 AO21x1_ASAP7_75t_R _24717_ (.A1(_09052_),
    .A2(_09335_),
    .B(_09336_),
    .Y(_02862_));
 OR2x2_ASAP7_75t_R _24718_ (.A(_00237_),
    .B(_00240_),
    .Y(_09337_));
 OA21x2_ASAP7_75t_R _24719_ (.A1(_00241_),
    .A2(_00240_),
    .B(_00244_),
    .Y(_09338_));
 OA21x2_ASAP7_75t_R _24720_ (.A1(_09274_),
    .A2(_09337_),
    .B(_09338_),
    .Y(_09339_));
 XNOR2x2_ASAP7_75t_R _24721_ (.A(_00243_),
    .B(_09339_),
    .Y(_09340_));
 NAND2x1_ASAP7_75t_R _24722_ (.A(_08902_),
    .B(_09340_),
    .Y(_09341_));
 OA211x2_ASAP7_75t_R _24723_ (.A1(_08902_),
    .A2(_08811_),
    .B(_09341_),
    .C(_05241_),
    .Y(_09342_));
 AND2x2_ASAP7_75t_R _24724_ (.A(_08307_),
    .B(_08430_),
    .Y(_09343_));
 AO21x1_ASAP7_75t_R _24725_ (.A1(_08513_),
    .A2(_08827_),
    .B(_09343_),
    .Y(_09344_));
 AND3x1_ASAP7_75t_R _24726_ (.A(_04788_),
    .B(_04790_),
    .C(_08371_),
    .Y(_09345_));
 AO21x1_ASAP7_75t_R _24727_ (.A1(_18558_),
    .A2(_08349_),
    .B(_09345_),
    .Y(_09346_));
 AO211x2_ASAP7_75t_R _24728_ (.A1(_18562_),
    .A2(_08349_),
    .B(_09319_),
    .C(_08409_),
    .Y(_09347_));
 OA211x2_ASAP7_75t_R _24729_ (.A1(_18555_),
    .A2(_09346_),
    .B(_09347_),
    .C(_08357_),
    .Y(_09348_));
 AO211x2_ASAP7_75t_R _24730_ (.A1(_08320_),
    .A2(_09284_),
    .B(_09348_),
    .C(_08528_),
    .Y(_09349_));
 OR3x1_ASAP7_75t_R _24731_ (.A(_08347_),
    .B(_09213_),
    .C(_09216_),
    .Y(_09350_));
 AO32x1_ASAP7_75t_R _24732_ (.A1(_08456_),
    .A2(_09349_),
    .A3(_09350_),
    .B1(_08539_),
    .B2(_09317_),
    .Y(_09351_));
 AO221x1_ASAP7_75t_R _24733_ (.A1(_08725_),
    .A2(_08830_),
    .B1(_08530_),
    .B2(_08722_),
    .C(_09351_),
    .Y(_09352_));
 OAI21x1_ASAP7_75t_R _24734_ (.A1(_04791_),
    .A2(_08901_),
    .B(_14388_),
    .Y(_09353_));
 AO221x1_ASAP7_75t_R _24735_ (.A1(_08512_),
    .A2(_09344_),
    .B1(_09352_),
    .B2(_08440_),
    .C(_09353_),
    .Y(_09354_));
 INVx1_ASAP7_75t_R _24736_ (.A(_02323_),
    .Y(_09355_));
 OA222x2_ASAP7_75t_R _24737_ (.A1(_00329_),
    .A2(_08731_),
    .B1(_08732_),
    .B2(_09355_),
    .C1(_08695_),
    .C2(_00328_),
    .Y(_09356_));
 OA21x2_ASAP7_75t_R _24738_ (.A1(_04983_),
    .A2(_08730_),
    .B(_09356_),
    .Y(_09357_));
 NOR2x1_ASAP7_75t_R _24739_ (.A(_08880_),
    .B(_09357_),
    .Y(_09358_));
 OR3x1_ASAP7_75t_R _24740_ (.A(_09342_),
    .B(_09354_),
    .C(_09358_),
    .Y(_09359_));
 AOI21x1_ASAP7_75t_R _24741_ (.A1(_14120_),
    .A2(_06478_),
    .B(_08504_),
    .Y(_09360_));
 NOR2x1_ASAP7_75t_R _24742_ (.A(_08270_),
    .B(_08846_),
    .Y(_09361_));
 AO21x1_ASAP7_75t_R _24743_ (.A1(_08270_),
    .A2(_08844_),
    .B(_09361_),
    .Y(_09362_));
 OA21x2_ASAP7_75t_R _24744_ (.A1(_08286_),
    .A2(_09362_),
    .B(_08912_),
    .Y(_09363_));
 NOR2x1_ASAP7_75t_R _24745_ (.A(_08853_),
    .B(_09363_),
    .Y(_09364_));
 AO21x2_ASAP7_75t_R _24746_ (.A1(_09359_),
    .A2(_09360_),
    .B(_09364_),
    .Y(_09365_));
 BUFx6f_ASAP7_75t_R _24747_ (.A(_09365_),
    .Y(_09366_));
 NAND2x1_ASAP7_75t_R _24748_ (.A(_01356_),
    .B(_08804_),
    .Y(_09367_));
 OA21x2_ASAP7_75t_R _24749_ (.A1(_08804_),
    .A2(_09366_),
    .B(_09367_),
    .Y(_02863_));
 OR3x1_ASAP7_75t_R _24750_ (.A(_08514_),
    .B(_08963_),
    .C(_08968_),
    .Y(_09368_));
 NAND2x1_ASAP7_75t_R _24751_ (.A(_18070_),
    .B(_08352_),
    .Y(_09369_));
 AO21x1_ASAP7_75t_R _24752_ (.A1(_14390_),
    .A2(_14444_),
    .B(_08352_),
    .Y(_09370_));
 AO21x1_ASAP7_75t_R _24753_ (.A1(_09369_),
    .A2(_09370_),
    .B(_18555_),
    .Y(_09371_));
 OA211x2_ASAP7_75t_R _24754_ (.A1(_13453_),
    .A2(_09346_),
    .B(_09371_),
    .C(_08337_),
    .Y(_09372_));
 AO211x2_ASAP7_75t_R _24755_ (.A1(_08320_),
    .A2(_09321_),
    .B(_09372_),
    .C(_08316_),
    .Y(_09373_));
 AND3x1_ASAP7_75t_R _24756_ (.A(_08456_),
    .B(_09368_),
    .C(_09373_),
    .Y(_09374_));
 AOI21x1_ASAP7_75t_R _24757_ (.A1(_08425_),
    .A2(_09317_),
    .B(_09374_),
    .Y(_09375_));
 AOI22x1_ASAP7_75t_R _24758_ (.A1(_08869_),
    .A2(_08725_),
    .B1(_08722_),
    .B2(_08395_),
    .Y(_09376_));
 AO21x1_ASAP7_75t_R _24759_ (.A1(_09375_),
    .A2(_09376_),
    .B(_08434_),
    .Y(_09377_));
 OA21x2_ASAP7_75t_R _24760_ (.A1(_08307_),
    .A2(_08873_),
    .B(_08459_),
    .Y(_09378_));
 INVx1_ASAP7_75t_R _24761_ (.A(_02224_),
    .Y(_09379_));
 OA222x2_ASAP7_75t_R _24762_ (.A1(_00330_),
    .A2(_08485_),
    .B1(_08815_),
    .B2(_09379_),
    .C1(_08489_),
    .C2(_01390_),
    .Y(_09380_));
 OAI22x1_ASAP7_75t_R _24763_ (.A1(_04959_),
    .A2(_08901_),
    .B1(_08483_),
    .B2(_09380_),
    .Y(_09381_));
 AOI21x1_ASAP7_75t_R _24764_ (.A1(_08512_),
    .A2(_09378_),
    .B(_09381_),
    .Y(_09382_));
 AND4x1_ASAP7_75t_R _24765_ (.A(_06502_),
    .B(_08268_),
    .C(_09377_),
    .D(_09382_),
    .Y(_09383_));
 OAI21x1_ASAP7_75t_R _24766_ (.A1(net1952),
    .A2(_09169_),
    .B(_09383_),
    .Y(_09384_));
 OA31x2_ASAP7_75t_R _24767_ (.A1(_00240_),
    .A2(_09309_),
    .A3(_09311_),
    .B1(_00244_),
    .Y(_09385_));
 OA21x2_ASAP7_75t_R _24768_ (.A1(_00243_),
    .A2(_09385_),
    .B(_00247_),
    .Y(_09386_));
 XOR2x2_ASAP7_75t_R _24769_ (.A(_00246_),
    .B(_09386_),
    .Y(_09387_));
 NAND2x1_ASAP7_75t_R _24770_ (.A(_09060_),
    .B(_08886_),
    .Y(_09388_));
 OA211x2_ASAP7_75t_R _24771_ (.A1(_09060_),
    .A2(_09387_),
    .B(_09388_),
    .C(_05242_),
    .Y(_09389_));
 NAND2x1_ASAP7_75t_R _24772_ (.A(_08605_),
    .B(_08864_),
    .Y(_09390_));
 OA211x2_ASAP7_75t_R _24773_ (.A1(_08271_),
    .A2(_08861_),
    .B(_09390_),
    .C(_08597_),
    .Y(_09391_));
 OA22x2_ASAP7_75t_R _24774_ (.A1(_09384_),
    .A2(_09389_),
    .B1(_09391_),
    .B2(_09024_),
    .Y(_09392_));
 BUFx6f_ASAP7_75t_R _24775_ (.A(_09392_),
    .Y(_09393_));
 AND2x2_ASAP7_75t_R _24776_ (.A(_04843_),
    .B(_08508_),
    .Y(_09394_));
 AO21x1_ASAP7_75t_R _24777_ (.A1(_08264_),
    .A2(_09393_),
    .B(_09394_),
    .Y(_02864_));
 NAND2x1_ASAP7_75t_R _24778_ (.A(_08440_),
    .B(_09194_),
    .Y(_09395_));
 INVx1_ASAP7_75t_R _24779_ (.A(_02299_),
    .Y(_09396_));
 OA222x2_ASAP7_75t_R _24780_ (.A1(_00281_),
    .A2(_08731_),
    .B1(_08732_),
    .B2(_09396_),
    .C1(_08695_),
    .C2(_00280_),
    .Y(_09397_));
 NAND2x1_ASAP7_75t_R _24781_ (.A(\alu_adder_result_ex[6] ),
    .B(_08818_),
    .Y(_09398_));
 AO21x1_ASAP7_75t_R _24782_ (.A1(_09397_),
    .A2(_09398_),
    .B(_08483_),
    .Y(_09399_));
 OA22x2_ASAP7_75t_R _24783_ (.A1(_00127_),
    .A2(_08567_),
    .B1(_08570_),
    .B2(_00121_),
    .Y(_09400_));
 AND4x1_ASAP7_75t_R _24784_ (.A(_06623_),
    .B(_09395_),
    .C(_09399_),
    .D(_09400_),
    .Y(_09401_));
 OAI21x1_ASAP7_75t_R _24785_ (.A1(_08438_),
    .A2(_09193_),
    .B(_09401_),
    .Y(_09402_));
 AO221x1_ASAP7_75t_R _24786_ (.A1(net62),
    .A2(_08790_),
    .B1(_08787_),
    .B2(net53),
    .C(_08595_),
    .Y(_09403_));
 INVx1_ASAP7_75t_R _24787_ (.A(_01419_),
    .Y(_09404_));
 AO221x1_ASAP7_75t_R _24788_ (.A1(_08839_),
    .A2(_08790_),
    .B1(_08787_),
    .B2(_09404_),
    .C(_08285_),
    .Y(_09405_));
 AND3x1_ASAP7_75t_R _24789_ (.A(_08289_),
    .B(_09403_),
    .C(_09405_),
    .Y(_09406_));
 OR2x2_ASAP7_75t_R _24790_ (.A(_09102_),
    .B(_09406_),
    .Y(_09407_));
 OAI22x1_ASAP7_75t_R _24791_ (.A1(_08843_),
    .A2(_08298_),
    .B1(_08799_),
    .B2(_01425_),
    .Y(_09408_));
 AO221x1_ASAP7_75t_R _24792_ (.A1(_09403_),
    .A2(_09405_),
    .B1(_09408_),
    .B2(_08290_),
    .C(_08270_),
    .Y(_09409_));
 OA211x2_ASAP7_75t_R _24793_ (.A1(_08287_),
    .A2(_09407_),
    .B(_09409_),
    .C(_08835_),
    .Y(_09410_));
 AO21x2_ASAP7_75t_R _24794_ (.A1(_08853_),
    .A2(_09402_),
    .B(_09410_),
    .Y(_09411_));
 BUFx6f_ASAP7_75t_R _24795_ (.A(_09411_),
    .Y(_09412_));
 NAND2x1_ASAP7_75t_R _24796_ (.A(_08950_),
    .B(_08954_),
    .Y(_09413_));
 BUFx12f_ASAP7_75t_R _24797_ (.A(_09413_),
    .Y(_09414_));
 AND2x2_ASAP7_75t_R _24798_ (.A(_13875_),
    .B(_09414_),
    .Y(_09415_));
 AO21x1_ASAP7_75t_R _24799_ (.A1(_08956_),
    .A2(_09412_),
    .B(_09415_),
    .Y(_02865_));
 NOR2x1_ASAP7_75t_R _24800_ (.A(_01418_),
    .B(_08285_),
    .Y(_09416_));
 AO21x1_ASAP7_75t_R _24801_ (.A1(net54),
    .A2(_08285_),
    .B(_09416_),
    .Y(_09417_));
 AO32x1_ASAP7_75t_R _24802_ (.A1(net63),
    .A2(_08285_),
    .A3(_08981_),
    .B1(_08982_),
    .B2(_09417_),
    .Y(_09418_));
 OA21x2_ASAP7_75t_R _24803_ (.A1(_08275_),
    .A2(_09418_),
    .B(_08299_),
    .Y(_09419_));
 OAI22x1_ASAP7_75t_R _24804_ (.A1(_08863_),
    .A2(_08298_),
    .B1(_08799_),
    .B2(_01424_),
    .Y(_09420_));
 AND3x1_ASAP7_75t_R _24805_ (.A(_08856_),
    .B(_08274_),
    .C(_08595_),
    .Y(_09421_));
 AO21x1_ASAP7_75t_R _24806_ (.A1(_08290_),
    .A2(_09420_),
    .B(_09421_),
    .Y(_09422_));
 OR3x1_ASAP7_75t_R _24807_ (.A(_08605_),
    .B(_09418_),
    .C(_09422_),
    .Y(_09423_));
 OA21x2_ASAP7_75t_R _24808_ (.A1(_08287_),
    .A2(_09419_),
    .B(_09423_),
    .Y(_09424_));
 INVx1_ASAP7_75t_R _24809_ (.A(_06648_),
    .Y(_09425_));
 NAND2x1_ASAP7_75t_R _24810_ (.A(_08439_),
    .B(_09166_),
    .Y(_09426_));
 OA211x2_ASAP7_75t_R _24811_ (.A1(_08833_),
    .A2(_09164_),
    .B(_09426_),
    .C(_08437_),
    .Y(_09427_));
 INVx1_ASAP7_75t_R _24812_ (.A(_02300_),
    .Y(_09428_));
 OA222x2_ASAP7_75t_R _24813_ (.A1(_00283_),
    .A2(_08485_),
    .B1(_08815_),
    .B2(_09428_),
    .C1(_15040_),
    .C2(_08484_),
    .Y(_09429_));
 OAI21x1_ASAP7_75t_R _24814_ (.A1(_00282_),
    .A2(_08558_),
    .B(_09429_),
    .Y(_09430_));
 INVx1_ASAP7_75t_R _24815_ (.A(_02209_),
    .Y(_09431_));
 OAI22x1_ASAP7_75t_R _24816_ (.A1(_09431_),
    .A2(_08567_),
    .B1(_08570_),
    .B2(_00128_),
    .Y(_09432_));
 AO21x1_ASAP7_75t_R _24817_ (.A1(_08721_),
    .A2(_09430_),
    .B(_09432_),
    .Y(_09433_));
 OR4x1_ASAP7_75t_R _24818_ (.A(_09425_),
    .B(_08835_),
    .C(_09427_),
    .D(_09433_),
    .Y(_09434_));
 OA21x2_ASAP7_75t_R _24819_ (.A1(_08853_),
    .A2(_09424_),
    .B(_09434_),
    .Y(_09435_));
 BUFx6f_ASAP7_75t_R _24820_ (.A(_09435_),
    .Y(_09436_));
 NOR2x1_ASAP7_75t_R _24821_ (.A(_00596_),
    .B(_08994_),
    .Y(_09437_));
 AO21x1_ASAP7_75t_R _24822_ (.A1(_08956_),
    .A2(_09436_),
    .B(_09437_),
    .Y(_02866_));
 BUFx6f_ASAP7_75t_R _24823_ (.A(_08506_),
    .Y(_09438_));
 BUFx12f_ASAP7_75t_R _24824_ (.A(_08955_),
    .Y(_09439_));
 NOR2x1_ASAP7_75t_R _24825_ (.A(_00626_),
    .B(_09439_),
    .Y(_09440_));
 AO21x1_ASAP7_75t_R _24826_ (.A1(_09438_),
    .A2(_08994_),
    .B(_09440_),
    .Y(_02867_));
 BUFx12f_ASAP7_75t_R _24827_ (.A(_08615_),
    .Y(_09441_));
 NOR2x1_ASAP7_75t_R _24828_ (.A(_00656_),
    .B(_09439_),
    .Y(_09442_));
 AO21x1_ASAP7_75t_R _24829_ (.A1(_09441_),
    .A2(_08994_),
    .B(_09442_),
    .Y(_02868_));
 BUFx6f_ASAP7_75t_R _24830_ (.A(_08669_),
    .Y(_09443_));
 NOR2x1_ASAP7_75t_R _24831_ (.A(_00686_),
    .B(_09439_),
    .Y(_09444_));
 AO21x1_ASAP7_75t_R _24832_ (.A1(_09443_),
    .A2(_08994_),
    .B(_09444_),
    .Y(_02869_));
 BUFx6f_ASAP7_75t_R _24833_ (.A(_08719_),
    .Y(_09445_));
 NOR2x1_ASAP7_75t_R _24834_ (.A(_00716_),
    .B(_09439_),
    .Y(_09446_));
 AO21x1_ASAP7_75t_R _24835_ (.A1(_09445_),
    .A2(_08994_),
    .B(_09446_),
    .Y(_02870_));
 BUFx6f_ASAP7_75t_R _24836_ (.A(_08757_),
    .Y(_09447_));
 NOR2x1_ASAP7_75t_R _24837_ (.A(_00346_),
    .B(_09439_),
    .Y(_09448_));
 AO21x1_ASAP7_75t_R _24838_ (.A1(_09447_),
    .A2(_08994_),
    .B(_09448_),
    .Y(_02871_));
 BUFx12f_ASAP7_75t_R _24839_ (.A(_08802_),
    .Y(_09449_));
 NOR2x1_ASAP7_75t_R _24840_ (.A(_00784_),
    .B(_09439_),
    .Y(_09450_));
 AO21x1_ASAP7_75t_R _24841_ (.A1(_09449_),
    .A2(_08994_),
    .B(_09450_),
    .Y(_02872_));
 BUFx12f_ASAP7_75t_R _24842_ (.A(_08850_),
    .Y(_09451_));
 AND2x2_ASAP7_75t_R _24843_ (.A(_09451_),
    .B(_08955_),
    .Y(_09452_));
 AOI21x1_ASAP7_75t_R _24844_ (.A1(_00816_),
    .A2(_09414_),
    .B(_09452_),
    .Y(_02873_));
 BUFx6f_ASAP7_75t_R _24845_ (.A(_08892_),
    .Y(_09453_));
 NAND2x1_ASAP7_75t_R _24846_ (.A(_00848_),
    .B(_09414_),
    .Y(_09454_));
 OA21x2_ASAP7_75t_R _24847_ (.A1(_09453_),
    .A2(_09414_),
    .B(_09454_),
    .Y(_02874_));
 BUFx6f_ASAP7_75t_R _24848_ (.A(_08920_),
    .Y(_09455_));
 NOR2x1_ASAP7_75t_R _24849_ (.A(_00880_),
    .B(_09439_),
    .Y(_09456_));
 AO21x1_ASAP7_75t_R _24850_ (.A1(_09455_),
    .A2(_08994_),
    .B(_09456_),
    .Y(_02875_));
 BUFx6f_ASAP7_75t_R _24851_ (.A(_08947_),
    .Y(_09457_));
 AND2x2_ASAP7_75t_R _24852_ (.A(_09457_),
    .B(_08955_),
    .Y(_09458_));
 AOI21x1_ASAP7_75t_R _24853_ (.A1(_00912_),
    .A2(_09414_),
    .B(_09458_),
    .Y(_02876_));
 NOR2x1_ASAP7_75t_R _24854_ (.A(_00944_),
    .B(_09439_),
    .Y(_09459_));
 AO21x1_ASAP7_75t_R _24855_ (.A1(_08956_),
    .A2(_09021_),
    .B(_09459_),
    .Y(_02877_));
 NOR2x1_ASAP7_75t_R _24856_ (.A(_00976_),
    .B(_09439_),
    .Y(_09460_));
 AO21x1_ASAP7_75t_R _24857_ (.A1(_08956_),
    .A2(_09048_),
    .B(_09460_),
    .Y(_02878_));
 NOR2x1_ASAP7_75t_R _24858_ (.A(_01008_),
    .B(_09439_),
    .Y(_09461_));
 AO21x1_ASAP7_75t_R _24859_ (.A1(_08956_),
    .A2(_09074_),
    .B(_09461_),
    .Y(_02879_));
 BUFx12f_ASAP7_75t_R _24860_ (.A(_08955_),
    .Y(_09462_));
 NOR2x1_ASAP7_75t_R _24861_ (.A(_01040_),
    .B(_09462_),
    .Y(_09463_));
 AO21x1_ASAP7_75t_R _24862_ (.A1(_08956_),
    .A2(_09099_),
    .B(_09463_),
    .Y(_02880_));
 BUFx6f_ASAP7_75t_R _24863_ (.A(_08955_),
    .Y(_09464_));
 NOR2x1_ASAP7_75t_R _24864_ (.A(_01072_),
    .B(_09462_),
    .Y(_09465_));
 AO21x1_ASAP7_75t_R _24865_ (.A1(_09464_),
    .A2(_09123_),
    .B(_09465_),
    .Y(_02881_));
 NOR2x1_ASAP7_75t_R _24866_ (.A(_01104_),
    .B(_09462_),
    .Y(_09466_));
 AO21x1_ASAP7_75t_R _24867_ (.A1(_09464_),
    .A2(_09144_),
    .B(_09466_),
    .Y(_02882_));
 NOR2x1_ASAP7_75t_R _24868_ (.A(_01136_),
    .B(_09462_),
    .Y(_09467_));
 AO21x1_ASAP7_75t_R _24869_ (.A1(_09464_),
    .A2(_09176_),
    .B(_09467_),
    .Y(_02883_));
 NOR2x1_ASAP7_75t_R _24870_ (.A(_01168_),
    .B(_09462_),
    .Y(_09468_));
 AO21x1_ASAP7_75t_R _24871_ (.A1(_09464_),
    .A2(_09203_),
    .B(_09468_),
    .Y(_02884_));
 NOR2x1_ASAP7_75t_R _24872_ (.A(_01200_),
    .B(_09462_),
    .Y(_09469_));
 AO21x1_ASAP7_75t_R _24873_ (.A1(_09464_),
    .A2(_09229_),
    .B(_09469_),
    .Y(_02885_));
 NOR2x1_ASAP7_75t_R _24874_ (.A(_01232_),
    .B(_09462_),
    .Y(_09470_));
 AO21x1_ASAP7_75t_R _24875_ (.A1(_09464_),
    .A2(_09249_),
    .B(_09470_),
    .Y(_02886_));
 NOR2x1_ASAP7_75t_R _24876_ (.A(_01264_),
    .B(_09462_),
    .Y(_09471_));
 AO21x1_ASAP7_75t_R _24877_ (.A1(_09464_),
    .A2(_09301_),
    .B(_09471_),
    .Y(_02887_));
 NOR2x1_ASAP7_75t_R _24878_ (.A(_01296_),
    .B(_09462_),
    .Y(_09472_));
 AO21x1_ASAP7_75t_R _24879_ (.A1(_09464_),
    .A2(_09334_),
    .B(_09472_),
    .Y(_02888_));
 NAND2x1_ASAP7_75t_R _24880_ (.A(_01328_),
    .B(_09414_),
    .Y(_09473_));
 OA21x2_ASAP7_75t_R _24881_ (.A1(_09414_),
    .A2(_09365_),
    .B(_09473_),
    .Y(_02889_));
 AND2x2_ASAP7_75t_R _24882_ (.A(_04894_),
    .B(_09413_),
    .Y(_09474_));
 AO21x1_ASAP7_75t_R _24883_ (.A1(_09464_),
    .A2(_09392_),
    .B(_09474_),
    .Y(_02890_));
 NAND2x1_ASAP7_75t_R _24884_ (.A(_08256_),
    .B(_08592_),
    .Y(_09475_));
 AND2x4_ASAP7_75t_R _24885_ (.A(_13685_),
    .B(_13603_),
    .Y(_09476_));
 AND5x2_ASAP7_75t_R _24886_ (.A(_07799_),
    .B(_13455_),
    .C(_13430_),
    .D(_09475_),
    .E(_09476_),
    .Y(_09477_));
 BUFx12f_ASAP7_75t_R _24887_ (.A(_09477_),
    .Y(_09478_));
 BUFx6f_ASAP7_75t_R _24888_ (.A(_09478_),
    .Y(_09479_));
 AO21x1_ASAP7_75t_R _24889_ (.A1(_09375_),
    .A2(_09376_),
    .B(_08438_),
    .Y(_09480_));
 INVx1_ASAP7_75t_R _24890_ (.A(_02293_),
    .Y(_09481_));
 OA22x2_ASAP7_75t_R _24891_ (.A1(_00064_),
    .A2(_08566_),
    .B1(_08569_),
    .B2(_00062_),
    .Y(_09482_));
 OA22x2_ASAP7_75t_R _24892_ (.A1(_16999_),
    .A2(_08468_),
    .B1(_08475_),
    .B2(_00269_),
    .Y(_09483_));
 OA211x2_ASAP7_75t_R _24893_ (.A1(_09481_),
    .A2(_08815_),
    .B(_09482_),
    .C(_09483_),
    .Y(_09484_));
 NAND2x1_ASAP7_75t_R _24894_ (.A(_08439_),
    .B(_09378_),
    .Y(_09485_));
 OA211x2_ASAP7_75t_R _24895_ (.A1(_02292_),
    .A2(_08558_),
    .B(_09484_),
    .C(_09485_),
    .Y(_09486_));
 AO32x2_ASAP7_75t_R _24896_ (.A1(_06857_),
    .A2(_06882_),
    .A3(_06888_),
    .B1(_08471_),
    .B2(_06874_),
    .Y(_09487_));
 NAND3x1_ASAP7_75t_R _24897_ (.A(_09480_),
    .B(_09486_),
    .C(_09487_),
    .Y(_09488_));
 AOI21x1_ASAP7_75t_R _24898_ (.A1(_08880_),
    .A2(_09482_),
    .B(_14120_),
    .Y(_09489_));
 AOI21x1_ASAP7_75t_R _24899_ (.A1(_09488_),
    .A2(_09489_),
    .B(_05805_),
    .Y(_09490_));
 AND3x1_ASAP7_75t_R _24900_ (.A(_01417_),
    .B(_08296_),
    .C(_08298_),
    .Y(_09491_));
 AO21x1_ASAP7_75t_R _24901_ (.A1(_08293_),
    .A2(_08285_),
    .B(_09491_),
    .Y(_09492_));
 NAND2x1_ASAP7_75t_R _24902_ (.A(net64),
    .B(_05738_),
    .Y(_09493_));
 OA211x2_ASAP7_75t_R _24903_ (.A1(_01432_),
    .A2(_08799_),
    .B(_09493_),
    .C(_08289_),
    .Y(_09494_));
 AO21x1_ASAP7_75t_R _24904_ (.A1(_08279_),
    .A2(_09492_),
    .B(_09494_),
    .Y(_09495_));
 AND3x1_ASAP7_75t_R _24905_ (.A(_01439_),
    .B(_08296_),
    .C(_08298_),
    .Y(_09496_));
 AO21x1_ASAP7_75t_R _24906_ (.A1(_08915_),
    .A2(_08285_),
    .B(_09496_),
    .Y(_09497_));
 OA211x2_ASAP7_75t_R _24907_ (.A1(_08609_),
    .A2(_09497_),
    .B(_08916_),
    .C(_08294_),
    .Y(_09498_));
 AO21x1_ASAP7_75t_R _24908_ (.A1(_08287_),
    .A2(_09495_),
    .B(_09498_),
    .Y(_09499_));
 AND2x2_ASAP7_75t_R _24909_ (.A(_08835_),
    .B(_09499_),
    .Y(_09500_));
 AO21x2_ASAP7_75t_R _24910_ (.A1(_08853_),
    .A2(_09490_),
    .B(_09500_),
    .Y(_09501_));
 BUFx12f_ASAP7_75t_R _24911_ (.A(_09501_),
    .Y(_09502_));
 BUFx12f_ASAP7_75t_R _24912_ (.A(_09502_),
    .Y(_09503_));
 NAND2x1_ASAP7_75t_R _24913_ (.A(_13455_),
    .B(_13430_),
    .Y(_09504_));
 AND2x2_ASAP7_75t_R _24914_ (.A(_08256_),
    .B(_08592_),
    .Y(_09505_));
 NAND2x2_ASAP7_75t_R _24915_ (.A(_13685_),
    .B(_13603_),
    .Y(_09506_));
 OR4x1_ASAP7_75t_R _24916_ (.A(_13692_),
    .B(_09504_),
    .C(_09505_),
    .D(_09506_),
    .Y(_09507_));
 BUFx12f_ASAP7_75t_R _24917_ (.A(_09507_),
    .Y(_09508_));
 AND2x2_ASAP7_75t_R _24918_ (.A(_00383_),
    .B(_09508_),
    .Y(_09509_));
 AOI21x1_ASAP7_75t_R _24919_ (.A1(_09479_),
    .A2(_09503_),
    .B(_09509_),
    .Y(_02891_));
 INVx1_ASAP7_75t_R _24920_ (.A(_02294_),
    .Y(_09510_));
 OA222x2_ASAP7_75t_R _24921_ (.A1(_00271_),
    .A2(_08475_),
    .B1(_08478_),
    .B2(_09510_),
    .C1(_18712_),
    .C2(_08468_),
    .Y(_09511_));
 OAI21x1_ASAP7_75t_R _24922_ (.A1(_00270_),
    .A2(_08489_),
    .B(_09511_),
    .Y(_09512_));
 AO21x1_ASAP7_75t_R _24923_ (.A1(_08352_),
    .A2(_09344_),
    .B(_09512_),
    .Y(_09513_));
 AO21x1_ASAP7_75t_R _24924_ (.A1(_08434_),
    .A2(_09352_),
    .B(_09513_),
    .Y(_09514_));
 OA21x2_ASAP7_75t_R _24925_ (.A1(_08437_),
    .A2(_09512_),
    .B(_08721_),
    .Y(_09515_));
 NAND2x1_ASAP7_75t_R _24926_ (.A(_09514_),
    .B(_09515_),
    .Y(_09516_));
 OA22x2_ASAP7_75t_R _24927_ (.A1(_00099_),
    .A2(_08567_),
    .B1(_08570_),
    .B2(_00097_),
    .Y(_09517_));
 AND3x1_ASAP7_75t_R _24928_ (.A(_06231_),
    .B(_09516_),
    .C(_09517_),
    .Y(_09518_));
 AO221x1_ASAP7_75t_R _24929_ (.A1(net56),
    .A2(_08790_),
    .B1(_08787_),
    .B2(net79),
    .C(_08595_),
    .Y(_09519_));
 INVx1_ASAP7_75t_R _24930_ (.A(_01428_),
    .Y(_09520_));
 AO221x1_ASAP7_75t_R _24931_ (.A1(_08600_),
    .A2(_08981_),
    .B1(_08982_),
    .B2(_09520_),
    .C(_08285_),
    .Y(_09521_));
 OAI22x1_ASAP7_75t_R _24932_ (.A1(_08608_),
    .A2(_08298_),
    .B1(_08799_),
    .B2(_01431_),
    .Y(_09522_));
 AO222x2_ASAP7_75t_R _24933_ (.A1(net59),
    .A2(_08796_),
    .B1(_09519_),
    .B2(_09521_),
    .C1(_09522_),
    .C2(_08987_),
    .Y(_09523_));
 NOR2x1_ASAP7_75t_R _24934_ (.A(_08268_),
    .B(_09523_),
    .Y(_09524_));
 AO21x2_ASAP7_75t_R _24935_ (.A1(_08853_),
    .A2(_09518_),
    .B(_09524_),
    .Y(_09525_));
 BUFx12f_ASAP7_75t_R _24936_ (.A(_09525_),
    .Y(_09526_));
 BUFx12f_ASAP7_75t_R _24937_ (.A(_09526_),
    .Y(_09527_));
 AND2x2_ASAP7_75t_R _24938_ (.A(_00416_),
    .B(_09508_),
    .Y(_09528_));
 AOI21x1_ASAP7_75t_R _24939_ (.A1(_09479_),
    .A2(_09527_),
    .B(_09528_),
    .Y(_02892_));
 AO221x1_ASAP7_75t_R _24940_ (.A1(net57),
    .A2(_08981_),
    .B1(_08982_),
    .B2(net28),
    .C(_08596_),
    .Y(_09529_));
 INVx1_ASAP7_75t_R _24941_ (.A(_01423_),
    .Y(_09530_));
 AO221x1_ASAP7_75t_R _24942_ (.A1(_08664_),
    .A2(_08981_),
    .B1(_08982_),
    .B2(_09530_),
    .C(_08285_),
    .Y(_09531_));
 OAI22x1_ASAP7_75t_R _24943_ (.A1(_08655_),
    .A2(_08298_),
    .B1(_08799_),
    .B2(_01430_),
    .Y(_09532_));
 AO222x2_ASAP7_75t_R _24944_ (.A1(net70),
    .A2(_08796_),
    .B1(_09529_),
    .B2(_09531_),
    .C1(_09532_),
    .C2(_08987_),
    .Y(_09533_));
 OR3x1_ASAP7_75t_R _24945_ (.A(_08349_),
    .B(_09165_),
    .C(_09326_),
    .Y(_09534_));
 OA211x2_ASAP7_75t_R _24946_ (.A1(_08439_),
    .A2(_09325_),
    .B(_09534_),
    .C(_08437_),
    .Y(_09535_));
 INVx1_ASAP7_75t_R _24947_ (.A(_02295_),
    .Y(_09536_));
 OA222x2_ASAP7_75t_R _24948_ (.A1(_00273_),
    .A2(_08559_),
    .B1(_08486_),
    .B2(_09536_),
    .C1(_08489_),
    .C2(_00272_),
    .Y(_09537_));
 OAI21x1_ASAP7_75t_R _24949_ (.A1(_05219_),
    .A2(_08484_),
    .B(_09537_),
    .Y(_09538_));
 OAI22x1_ASAP7_75t_R _24950_ (.A1(_00103_),
    .A2(_08567_),
    .B1(_08570_),
    .B2(_00100_),
    .Y(_09539_));
 AO21x1_ASAP7_75t_R _24951_ (.A1(_08721_),
    .A2(_09538_),
    .B(_09539_),
    .Y(_09540_));
 OR4x1_ASAP7_75t_R _24952_ (.A(_05844_),
    .B(_08835_),
    .C(_09535_),
    .D(_09540_),
    .Y(_09541_));
 OAI21x1_ASAP7_75t_R _24953_ (.A1(_08853_),
    .A2(_09533_),
    .B(_09541_),
    .Y(_09542_));
 BUFx6f_ASAP7_75t_R _24954_ (.A(_09542_),
    .Y(_09543_));
 AND2x2_ASAP7_75t_R _24955_ (.A(_09478_),
    .B(_09543_),
    .Y(_09544_));
 AOI21x1_ASAP7_75t_R _24956_ (.A1(_00447_),
    .A2(_09508_),
    .B(_09544_),
    .Y(_02893_));
 AO221x1_ASAP7_75t_R _24957_ (.A1(net58),
    .A2(_08981_),
    .B1(_08982_),
    .B2(net29),
    .C(_08596_),
    .Y(_09545_));
 INVx1_ASAP7_75t_R _24958_ (.A(_01422_),
    .Y(_09546_));
 AO221x1_ASAP7_75t_R _24959_ (.A1(_08714_),
    .A2(_08981_),
    .B1(_08982_),
    .B2(_09546_),
    .C(_08286_),
    .Y(_09547_));
 OAI22x1_ASAP7_75t_R _24960_ (.A1(_08706_),
    .A2(_08298_),
    .B1(_08799_),
    .B2(_01429_),
    .Y(_09548_));
 AO222x2_ASAP7_75t_R _24961_ (.A1(net73),
    .A2(_08796_),
    .B1(_09545_),
    .B2(_09547_),
    .C1(_09548_),
    .C2(_08987_),
    .Y(_09549_));
 INVx1_ASAP7_75t_R _24962_ (.A(_06554_),
    .Y(_09550_));
 INVx1_ASAP7_75t_R _24963_ (.A(_02296_),
    .Y(_09551_));
 OA222x2_ASAP7_75t_R _24964_ (.A1(_00275_),
    .A2(_08559_),
    .B1(_08486_),
    .B2(_09551_),
    .C1(_05214_),
    .C2(_08468_),
    .Y(_09552_));
 OAI21x1_ASAP7_75t_R _24965_ (.A1(_00274_),
    .A2(_08558_),
    .B(_09552_),
    .Y(_09553_));
 AO21x1_ASAP7_75t_R _24966_ (.A1(_08439_),
    .A2(_09290_),
    .B(_09553_),
    .Y(_09554_));
 AND3x1_ASAP7_75t_R _24967_ (.A(_08511_),
    .B(_09279_),
    .C(_09288_),
    .Y(_09555_));
 AO21x1_ASAP7_75t_R _24968_ (.A1(_08721_),
    .A2(_09554_),
    .B(_09555_),
    .Y(_09556_));
 OAI22x1_ASAP7_75t_R _24969_ (.A1(_00108_),
    .A2(_08567_),
    .B1(_08570_),
    .B2(_00104_),
    .Y(_09557_));
 OR4x1_ASAP7_75t_R _24970_ (.A(_09550_),
    .B(_08835_),
    .C(_09556_),
    .D(_09557_),
    .Y(_09558_));
 OA21x2_ASAP7_75t_R _24971_ (.A1(_08853_),
    .A2(_09549_),
    .B(_09558_),
    .Y(_09559_));
 BUFx12f_ASAP7_75t_R _24972_ (.A(_09559_),
    .Y(_09560_));
 BUFx12f_ASAP7_75t_R _24973_ (.A(_09478_),
    .Y(_09561_));
 NOR2x1_ASAP7_75t_R _24974_ (.A(_00477_),
    .B(_09561_),
    .Y(_09562_));
 AO21x1_ASAP7_75t_R _24975_ (.A1(_09479_),
    .A2(_09560_),
    .B(_09562_),
    .Y(_02894_));
 BUFx12f_ASAP7_75t_R _24976_ (.A(_08992_),
    .Y(_09563_));
 NOR2x1_ASAP7_75t_R _24977_ (.A(_00507_),
    .B(_09561_),
    .Y(_09564_));
 AO21x1_ASAP7_75t_R _24978_ (.A1(_09563_),
    .A2(_09479_),
    .B(_09564_),
    .Y(_02895_));
 BUFx12f_ASAP7_75t_R _24979_ (.A(_09267_),
    .Y(_09565_));
 NOR2x1_ASAP7_75t_R _24980_ (.A(_00537_),
    .B(_09561_),
    .Y(_09566_));
 AO21x1_ASAP7_75t_R _24981_ (.A1(_09565_),
    .A2(_09479_),
    .B(_09566_),
    .Y(_02896_));
 BUFx6f_ASAP7_75t_R _24982_ (.A(_09411_),
    .Y(_09567_));
 BUFx12f_ASAP7_75t_R _24983_ (.A(_09478_),
    .Y(_09568_));
 NOR2x1_ASAP7_75t_R _24984_ (.A(_00567_),
    .B(_09568_),
    .Y(_09569_));
 AO21x1_ASAP7_75t_R _24985_ (.A1(_09567_),
    .A2(_09479_),
    .B(_09569_),
    .Y(_02897_));
 BUFx6f_ASAP7_75t_R _24986_ (.A(_09435_),
    .Y(_09570_));
 NOR2x1_ASAP7_75t_R _24987_ (.A(_00597_),
    .B(_09568_),
    .Y(_09571_));
 AO21x1_ASAP7_75t_R _24988_ (.A1(_09570_),
    .A2(_09479_),
    .B(_09571_),
    .Y(_02898_));
 BUFx6f_ASAP7_75t_R _24989_ (.A(_08506_),
    .Y(_09572_));
 NOR2x1_ASAP7_75t_R _24990_ (.A(_00627_),
    .B(_09568_),
    .Y(_09573_));
 AO21x1_ASAP7_75t_R _24991_ (.A1(_09572_),
    .A2(_09479_),
    .B(_09573_),
    .Y(_02899_));
 NOR2x1_ASAP7_75t_R _24992_ (.A(_00657_),
    .B(_09568_),
    .Y(_09574_));
 AO21x1_ASAP7_75t_R _24993_ (.A1(_09441_),
    .A2(_09479_),
    .B(_09574_),
    .Y(_02900_));
 BUFx6f_ASAP7_75t_R _24994_ (.A(_08669_),
    .Y(_09575_));
 NOR2x1_ASAP7_75t_R _24995_ (.A(_00687_),
    .B(_09568_),
    .Y(_09576_));
 AO21x1_ASAP7_75t_R _24996_ (.A1(_09575_),
    .A2(_09479_),
    .B(_09576_),
    .Y(_02901_));
 BUFx6f_ASAP7_75t_R _24997_ (.A(_09478_),
    .Y(_09577_));
 NOR2x1_ASAP7_75t_R _24998_ (.A(_00717_),
    .B(_09568_),
    .Y(_09578_));
 AO21x1_ASAP7_75t_R _24999_ (.A1(_09445_),
    .A2(_09577_),
    .B(_09578_),
    .Y(_02902_));
 BUFx12f_ASAP7_75t_R _25000_ (.A(_08757_),
    .Y(_09579_));
 NOR2x1_ASAP7_75t_R _25001_ (.A(_00347_),
    .B(_09568_),
    .Y(_09580_));
 AO21x1_ASAP7_75t_R _25002_ (.A1(_09579_),
    .A2(_09577_),
    .B(_09580_),
    .Y(_02903_));
 NOR2x1_ASAP7_75t_R _25003_ (.A(_00785_),
    .B(_09568_),
    .Y(_09581_));
 AO21x1_ASAP7_75t_R _25004_ (.A1(_09449_),
    .A2(_09577_),
    .B(_09581_),
    .Y(_02904_));
 AND2x2_ASAP7_75t_R _25005_ (.A(_09451_),
    .B(_09478_),
    .Y(_09582_));
 AOI21x1_ASAP7_75t_R _25006_ (.A1(_00817_),
    .A2(_09508_),
    .B(_09582_),
    .Y(_02905_));
 NAND2x1_ASAP7_75t_R _25007_ (.A(_00849_),
    .B(_09508_),
    .Y(_09583_));
 OA21x2_ASAP7_75t_R _25008_ (.A1(_09453_),
    .A2(_09508_),
    .B(_09583_),
    .Y(_02906_));
 BUFx6f_ASAP7_75t_R _25009_ (.A(_08920_),
    .Y(_09584_));
 NOR2x1_ASAP7_75t_R _25010_ (.A(_00881_),
    .B(_09568_),
    .Y(_09585_));
 AO21x1_ASAP7_75t_R _25011_ (.A1(_09584_),
    .A2(_09577_),
    .B(_09585_),
    .Y(_02907_));
 AND2x2_ASAP7_75t_R _25012_ (.A(_09457_),
    .B(_09478_),
    .Y(_09586_));
 AOI21x1_ASAP7_75t_R _25013_ (.A1(_00913_),
    .A2(_09508_),
    .B(_09586_),
    .Y(_02908_));
 BUFx12f_ASAP7_75t_R _25014_ (.A(_09021_),
    .Y(_09587_));
 NOR2x1_ASAP7_75t_R _25015_ (.A(_00945_),
    .B(_09568_),
    .Y(_09588_));
 AO21x1_ASAP7_75t_R _25016_ (.A1(_09587_),
    .A2(_09577_),
    .B(_09588_),
    .Y(_02909_));
 BUFx12f_ASAP7_75t_R _25017_ (.A(_09048_),
    .Y(_09589_));
 BUFx12f_ASAP7_75t_R _25018_ (.A(_09478_),
    .Y(_09590_));
 NOR2x1_ASAP7_75t_R _25019_ (.A(_00977_),
    .B(_09590_),
    .Y(_09591_));
 AO21x1_ASAP7_75t_R _25020_ (.A1(_09589_),
    .A2(_09577_),
    .B(_09591_),
    .Y(_02910_));
 BUFx6f_ASAP7_75t_R _25021_ (.A(_09074_),
    .Y(_09592_));
 NOR2x1_ASAP7_75t_R _25022_ (.A(_01009_),
    .B(_09590_),
    .Y(_09593_));
 AO21x1_ASAP7_75t_R _25023_ (.A1(_09592_),
    .A2(_09577_),
    .B(_09593_),
    .Y(_02911_));
 BUFx6f_ASAP7_75t_R _25024_ (.A(_09099_),
    .Y(_09594_));
 NOR2x1_ASAP7_75t_R _25025_ (.A(_01041_),
    .B(_09590_),
    .Y(_09595_));
 AO21x1_ASAP7_75t_R _25026_ (.A1(_09594_),
    .A2(_09577_),
    .B(_09595_),
    .Y(_02912_));
 BUFx6f_ASAP7_75t_R _25027_ (.A(_09123_),
    .Y(_09596_));
 NOR2x1_ASAP7_75t_R _25028_ (.A(_01073_),
    .B(_09590_),
    .Y(_09597_));
 AO21x1_ASAP7_75t_R _25029_ (.A1(_09596_),
    .A2(_09577_),
    .B(_09597_),
    .Y(_02913_));
 BUFx6f_ASAP7_75t_R _25030_ (.A(_09144_),
    .Y(_09598_));
 NOR2x1_ASAP7_75t_R _25031_ (.A(_01105_),
    .B(_09590_),
    .Y(_09599_));
 AO21x1_ASAP7_75t_R _25032_ (.A1(_09598_),
    .A2(_09577_),
    .B(_09599_),
    .Y(_02914_));
 BUFx6f_ASAP7_75t_R _25033_ (.A(_09176_),
    .Y(_09600_));
 NOR2x1_ASAP7_75t_R _25034_ (.A(_01137_),
    .B(_09590_),
    .Y(_09601_));
 AO21x1_ASAP7_75t_R _25035_ (.A1(_09600_),
    .A2(_09561_),
    .B(_09601_),
    .Y(_02915_));
 BUFx6f_ASAP7_75t_R _25036_ (.A(_09203_),
    .Y(_09602_));
 NOR2x1_ASAP7_75t_R _25037_ (.A(_01169_),
    .B(_09590_),
    .Y(_09603_));
 AO21x1_ASAP7_75t_R _25038_ (.A1(_09602_),
    .A2(_09561_),
    .B(_09603_),
    .Y(_02916_));
 BUFx6f_ASAP7_75t_R _25039_ (.A(_09229_),
    .Y(_09604_));
 NOR2x1_ASAP7_75t_R _25040_ (.A(_01201_),
    .B(_09590_),
    .Y(_09605_));
 AO21x1_ASAP7_75t_R _25041_ (.A1(_09604_),
    .A2(_09561_),
    .B(_09605_),
    .Y(_02917_));
 BUFx6f_ASAP7_75t_R _25042_ (.A(_09249_),
    .Y(_09606_));
 NOR2x1_ASAP7_75t_R _25043_ (.A(_01233_),
    .B(_09590_),
    .Y(_09607_));
 AO21x1_ASAP7_75t_R _25044_ (.A1(_09606_),
    .A2(_09561_),
    .B(_09607_),
    .Y(_02918_));
 BUFx6f_ASAP7_75t_R _25045_ (.A(_09301_),
    .Y(_09608_));
 NOR2x1_ASAP7_75t_R _25046_ (.A(_01265_),
    .B(_09590_),
    .Y(_09609_));
 AO21x1_ASAP7_75t_R _25047_ (.A1(_09608_),
    .A2(_09561_),
    .B(_09609_),
    .Y(_02919_));
 BUFx6f_ASAP7_75t_R _25048_ (.A(_09334_),
    .Y(_09610_));
 NOR2x1_ASAP7_75t_R _25049_ (.A(_01297_),
    .B(_09478_),
    .Y(_09611_));
 AO21x1_ASAP7_75t_R _25050_ (.A1(_09610_),
    .A2(_09561_),
    .B(_09611_),
    .Y(_02920_));
 BUFx6f_ASAP7_75t_R _25051_ (.A(_09365_),
    .Y(_09612_));
 NAND2x1_ASAP7_75t_R _25052_ (.A(_01329_),
    .B(_09508_),
    .Y(_09613_));
 OA21x2_ASAP7_75t_R _25053_ (.A1(_09612_),
    .A2(_09508_),
    .B(_09613_),
    .Y(_02921_));
 BUFx6f_ASAP7_75t_R _25054_ (.A(_09392_),
    .Y(_09614_));
 NOR2x1_ASAP7_75t_R _25055_ (.A(_01361_),
    .B(_09478_),
    .Y(_09615_));
 AO21x1_ASAP7_75t_R _25056_ (.A1(_09614_),
    .A2(_09561_),
    .B(_09615_),
    .Y(_02922_));
 BUFx12f_ASAP7_75t_R _25057_ (.A(_09476_),
    .Y(_09616_));
 INVx2_ASAP7_75t_R _25058_ (.A(_13430_),
    .Y(_09617_));
 NAND2x1_ASAP7_75t_R _25059_ (.A(_13455_),
    .B(_09617_),
    .Y(_09618_));
 INVx1_ASAP7_75t_R _25060_ (.A(_09618_),
    .Y(_09619_));
 OA211x2_ASAP7_75t_R _25061_ (.A1(_08255_),
    .A2(_08268_),
    .B(_09619_),
    .C(_07799_),
    .Y(_09620_));
 BUFx12f_ASAP7_75t_R _25062_ (.A(_09620_),
    .Y(_09621_));
 AND2x6_ASAP7_75t_R _25063_ (.A(_09616_),
    .B(_09621_),
    .Y(_09622_));
 NAND2x2_ASAP7_75t_R _25064_ (.A(_09616_),
    .B(_09620_),
    .Y(_09623_));
 BUFx12f_ASAP7_75t_R _25065_ (.A(_09623_),
    .Y(_09624_));
 AND2x2_ASAP7_75t_R _25066_ (.A(_00384_),
    .B(_09624_),
    .Y(_09625_));
 AOI21x1_ASAP7_75t_R _25067_ (.A1(_09503_),
    .A2(_09622_),
    .B(_09625_),
    .Y(_02923_));
 AND2x2_ASAP7_75t_R _25068_ (.A(_00417_),
    .B(_09624_),
    .Y(_09626_));
 AOI21x1_ASAP7_75t_R _25069_ (.A1(_09527_),
    .A2(_09622_),
    .B(_09626_),
    .Y(_02924_));
 BUFx12f_ASAP7_75t_R _25070_ (.A(_09623_),
    .Y(_09627_));
 AND2x2_ASAP7_75t_R _25071_ (.A(_09543_),
    .B(_09622_),
    .Y(_09628_));
 AOI21x1_ASAP7_75t_R _25072_ (.A1(_00448_),
    .A2(_09627_),
    .B(_09628_),
    .Y(_02925_));
 BUFx12f_ASAP7_75t_R _25073_ (.A(_09559_),
    .Y(_09629_));
 BUFx12f_ASAP7_75t_R _25074_ (.A(_09623_),
    .Y(_09630_));
 NAND2x1_ASAP7_75t_R _25075_ (.A(_00478_),
    .B(_09630_),
    .Y(_09631_));
 OA21x2_ASAP7_75t_R _25076_ (.A1(_09629_),
    .A2(_09627_),
    .B(_09631_),
    .Y(_02926_));
 NAND2x1_ASAP7_75t_R _25077_ (.A(_00508_),
    .B(_09630_),
    .Y(_09632_));
 OA21x2_ASAP7_75t_R _25078_ (.A1(_09563_),
    .A2(_09627_),
    .B(_09632_),
    .Y(_02927_));
 NAND2x1_ASAP7_75t_R _25079_ (.A(_00538_),
    .B(_09630_),
    .Y(_09633_));
 OA21x2_ASAP7_75t_R _25080_ (.A1(_09565_),
    .A2(_09627_),
    .B(_09633_),
    .Y(_02928_));
 NAND2x1_ASAP7_75t_R _25081_ (.A(_00568_),
    .B(_09630_),
    .Y(_09634_));
 OA21x2_ASAP7_75t_R _25082_ (.A1(_09567_),
    .A2(_09627_),
    .B(_09634_),
    .Y(_02929_));
 NAND2x1_ASAP7_75t_R _25083_ (.A(_00598_),
    .B(_09630_),
    .Y(_09635_));
 OA21x2_ASAP7_75t_R _25084_ (.A1(_09570_),
    .A2(_09627_),
    .B(_09635_),
    .Y(_02930_));
 NAND2x1_ASAP7_75t_R _25085_ (.A(_00628_),
    .B(_09630_),
    .Y(_09636_));
 OA21x2_ASAP7_75t_R _25086_ (.A1(_09438_),
    .A2(_09627_),
    .B(_09636_),
    .Y(_02931_));
 NAND2x1_ASAP7_75t_R _25087_ (.A(_00658_),
    .B(_09630_),
    .Y(_09637_));
 OA21x2_ASAP7_75t_R _25088_ (.A1(_09441_),
    .A2(_09627_),
    .B(_09637_),
    .Y(_02932_));
 BUFx12f_ASAP7_75t_R _25089_ (.A(_09624_),
    .Y(_09638_));
 NAND2x1_ASAP7_75t_R _25090_ (.A(_00688_),
    .B(_09630_),
    .Y(_09639_));
 OA21x2_ASAP7_75t_R _25091_ (.A1(_09443_),
    .A2(_09638_),
    .B(_09639_),
    .Y(_02933_));
 NAND2x1_ASAP7_75t_R _25092_ (.A(_00718_),
    .B(_09630_),
    .Y(_09640_));
 OA21x2_ASAP7_75t_R _25093_ (.A1(_09445_),
    .A2(_09638_),
    .B(_09640_),
    .Y(_02934_));
 NAND2x1_ASAP7_75t_R _25094_ (.A(_00348_),
    .B(_09630_),
    .Y(_09641_));
 OA21x2_ASAP7_75t_R _25095_ (.A1(_09447_),
    .A2(_09638_),
    .B(_09641_),
    .Y(_02935_));
 BUFx12f_ASAP7_75t_R _25096_ (.A(_09623_),
    .Y(_09642_));
 NAND2x1_ASAP7_75t_R _25097_ (.A(_00786_),
    .B(_09642_),
    .Y(_09643_));
 OA21x2_ASAP7_75t_R _25098_ (.A1(_09449_),
    .A2(_09638_),
    .B(_09643_),
    .Y(_02936_));
 AND2x2_ASAP7_75t_R _25099_ (.A(_09451_),
    .B(_09622_),
    .Y(_09644_));
 AOI21x1_ASAP7_75t_R _25100_ (.A1(_00818_),
    .A2(_09627_),
    .B(_09644_),
    .Y(_02937_));
 NAND2x1_ASAP7_75t_R _25101_ (.A(_00850_),
    .B(_09642_),
    .Y(_09645_));
 OA21x2_ASAP7_75t_R _25102_ (.A1(_09453_),
    .A2(_09638_),
    .B(_09645_),
    .Y(_02938_));
 NAND2x1_ASAP7_75t_R _25103_ (.A(_00882_),
    .B(_09642_),
    .Y(_09646_));
 OA21x2_ASAP7_75t_R _25104_ (.A1(_09455_),
    .A2(_09638_),
    .B(_09646_),
    .Y(_02939_));
 AND2x2_ASAP7_75t_R _25105_ (.A(_09457_),
    .B(_09622_),
    .Y(_09647_));
 AOI21x1_ASAP7_75t_R _25106_ (.A1(_00914_),
    .A2(_09627_),
    .B(_09647_),
    .Y(_02940_));
 NAND2x1_ASAP7_75t_R _25107_ (.A(_00946_),
    .B(_09642_),
    .Y(_09648_));
 OA21x2_ASAP7_75t_R _25108_ (.A1(_09587_),
    .A2(_09638_),
    .B(_09648_),
    .Y(_02941_));
 NAND2x1_ASAP7_75t_R _25109_ (.A(_00978_),
    .B(_09642_),
    .Y(_09649_));
 OA21x2_ASAP7_75t_R _25110_ (.A1(_09589_),
    .A2(_09638_),
    .B(_09649_),
    .Y(_02942_));
 NAND2x1_ASAP7_75t_R _25111_ (.A(_01010_),
    .B(_09642_),
    .Y(_09650_));
 OA21x2_ASAP7_75t_R _25112_ (.A1(_09592_),
    .A2(_09638_),
    .B(_09650_),
    .Y(_02943_));
 NAND2x1_ASAP7_75t_R _25113_ (.A(_01042_),
    .B(_09642_),
    .Y(_09651_));
 OA21x2_ASAP7_75t_R _25114_ (.A1(_09594_),
    .A2(_09638_),
    .B(_09651_),
    .Y(_02944_));
 BUFx6f_ASAP7_75t_R _25115_ (.A(_09623_),
    .Y(_09652_));
 NAND2x1_ASAP7_75t_R _25116_ (.A(_01074_),
    .B(_09642_),
    .Y(_09653_));
 OA21x2_ASAP7_75t_R _25117_ (.A1(_09596_),
    .A2(_09652_),
    .B(_09653_),
    .Y(_02945_));
 NAND2x1_ASAP7_75t_R _25118_ (.A(_01106_),
    .B(_09642_),
    .Y(_09654_));
 OA21x2_ASAP7_75t_R _25119_ (.A1(_09598_),
    .A2(_09652_),
    .B(_09654_),
    .Y(_02946_));
 NAND2x1_ASAP7_75t_R _25120_ (.A(_01138_),
    .B(_09642_),
    .Y(_09655_));
 OA21x2_ASAP7_75t_R _25121_ (.A1(_09600_),
    .A2(_09652_),
    .B(_09655_),
    .Y(_02947_));
 NAND2x1_ASAP7_75t_R _25122_ (.A(_01170_),
    .B(_09624_),
    .Y(_09656_));
 OA21x2_ASAP7_75t_R _25123_ (.A1(_09602_),
    .A2(_09652_),
    .B(_09656_),
    .Y(_02948_));
 NAND2x1_ASAP7_75t_R _25124_ (.A(_01202_),
    .B(_09624_),
    .Y(_09657_));
 OA21x2_ASAP7_75t_R _25125_ (.A1(_09604_),
    .A2(_09652_),
    .B(_09657_),
    .Y(_02949_));
 NAND2x1_ASAP7_75t_R _25126_ (.A(_01234_),
    .B(_09624_),
    .Y(_09658_));
 OA21x2_ASAP7_75t_R _25127_ (.A1(_09606_),
    .A2(_09652_),
    .B(_09658_),
    .Y(_02950_));
 NAND2x1_ASAP7_75t_R _25128_ (.A(_01266_),
    .B(_09624_),
    .Y(_09659_));
 OA21x2_ASAP7_75t_R _25129_ (.A1(_09608_),
    .A2(_09652_),
    .B(_09659_),
    .Y(_02951_));
 NAND2x1_ASAP7_75t_R _25130_ (.A(_01298_),
    .B(_09624_),
    .Y(_09660_));
 OA21x2_ASAP7_75t_R _25131_ (.A1(_09610_),
    .A2(_09652_),
    .B(_09660_),
    .Y(_02952_));
 NAND2x1_ASAP7_75t_R _25132_ (.A(_01330_),
    .B(_09624_),
    .Y(_09661_));
 OA21x2_ASAP7_75t_R _25133_ (.A1(_09612_),
    .A2(_09652_),
    .B(_09661_),
    .Y(_02953_));
 NAND2x1_ASAP7_75t_R _25134_ (.A(_01362_),
    .B(_09624_),
    .Y(_09662_));
 OA21x2_ASAP7_75t_R _25135_ (.A1(_09614_),
    .A2(_09652_),
    .B(_09662_),
    .Y(_02954_));
 NAND2x1_ASAP7_75t_R _25136_ (.A(_13456_),
    .B(_13430_),
    .Y(_09663_));
 INVx1_ASAP7_75t_R _25137_ (.A(_09663_),
    .Y(_09664_));
 OA211x2_ASAP7_75t_R _25138_ (.A1(_08255_),
    .A2(_08268_),
    .B(_09664_),
    .C(_00339_),
    .Y(_09665_));
 BUFx12f_ASAP7_75t_R _25139_ (.A(_09665_),
    .Y(_09666_));
 BUFx6f_ASAP7_75t_R _25140_ (.A(_09666_),
    .Y(_09667_));
 AND2x6_ASAP7_75t_R _25141_ (.A(_09616_),
    .B(_09667_),
    .Y(_09668_));
 BUFx6f_ASAP7_75t_R _25142_ (.A(_09668_),
    .Y(_09669_));
 NAND2x2_ASAP7_75t_R _25143_ (.A(_09616_),
    .B(_09666_),
    .Y(_09670_));
 BUFx12f_ASAP7_75t_R _25144_ (.A(_09670_),
    .Y(_09671_));
 AND2x2_ASAP7_75t_R _25145_ (.A(_00385_),
    .B(_09671_),
    .Y(_09672_));
 AOI21x1_ASAP7_75t_R _25146_ (.A1(_09503_),
    .A2(_09669_),
    .B(_09672_),
    .Y(_02955_));
 BUFx6f_ASAP7_75t_R _25147_ (.A(_09670_),
    .Y(_09673_));
 AND2x2_ASAP7_75t_R _25148_ (.A(_00418_),
    .B(_09673_),
    .Y(_09674_));
 AOI21x1_ASAP7_75t_R _25149_ (.A1(_09527_),
    .A2(_09669_),
    .B(_09674_),
    .Y(_02956_));
 BUFx12f_ASAP7_75t_R _25150_ (.A(_09542_),
    .Y(_09675_));
 NOR2x1_ASAP7_75t_R _25151_ (.A(_09675_),
    .B(_09671_),
    .Y(_09676_));
 AO21x1_ASAP7_75t_R _25152_ (.A1(_13556_),
    .A2(_09671_),
    .B(_09676_),
    .Y(_02957_));
 AND2x2_ASAP7_75t_R _25153_ (.A(_13679_),
    .B(_09673_),
    .Y(_09677_));
 AO21x1_ASAP7_75t_R _25154_ (.A1(_09629_),
    .A2(_09669_),
    .B(_09677_),
    .Y(_02958_));
 AND2x2_ASAP7_75t_R _25155_ (.A(_14795_),
    .B(_09673_),
    .Y(_09678_));
 AO21x1_ASAP7_75t_R _25156_ (.A1(_09563_),
    .A2(_09669_),
    .B(_09678_),
    .Y(_02959_));
 BUFx6f_ASAP7_75t_R _25157_ (.A(_09267_),
    .Y(_09679_));
 AND2x2_ASAP7_75t_R _25158_ (.A(_13774_),
    .B(_09673_),
    .Y(_09680_));
 AO21x1_ASAP7_75t_R _25159_ (.A1(_09679_),
    .A2(_09669_),
    .B(_09680_),
    .Y(_02960_));
 AND2x2_ASAP7_75t_R _25160_ (.A(_13901_),
    .B(_09673_),
    .Y(_09681_));
 AO21x1_ASAP7_75t_R _25161_ (.A1(_09567_),
    .A2(_09669_),
    .B(_09681_),
    .Y(_02961_));
 AND2x2_ASAP7_75t_R _25162_ (.A(_13952_),
    .B(_09673_),
    .Y(_09682_));
 AO21x1_ASAP7_75t_R _25163_ (.A1(_09570_),
    .A2(_09669_),
    .B(_09682_),
    .Y(_02962_));
 AND2x2_ASAP7_75t_R _25164_ (.A(_14010_),
    .B(_09673_),
    .Y(_09683_));
 AO21x1_ASAP7_75t_R _25165_ (.A1(_09572_),
    .A2(_09669_),
    .B(_09683_),
    .Y(_02963_));
 AND2x2_ASAP7_75t_R _25166_ (.A(_14032_),
    .B(_09673_),
    .Y(_09684_));
 AO21x1_ASAP7_75t_R _25167_ (.A1(_09441_),
    .A2(_09669_),
    .B(_09684_),
    .Y(_02964_));
 AND2x2_ASAP7_75t_R _25168_ (.A(_14177_),
    .B(_09673_),
    .Y(_09685_));
 AO21x1_ASAP7_75t_R _25169_ (.A1(_09575_),
    .A2(_09669_),
    .B(_09685_),
    .Y(_02965_));
 BUFx12f_ASAP7_75t_R _25170_ (.A(_09668_),
    .Y(_09686_));
 AND2x2_ASAP7_75t_R _25171_ (.A(_14214_),
    .B(_09673_),
    .Y(_09687_));
 AO21x1_ASAP7_75t_R _25172_ (.A1(_09445_),
    .A2(_09686_),
    .B(_09687_),
    .Y(_02966_));
 BUFx6f_ASAP7_75t_R _25173_ (.A(_09670_),
    .Y(_09688_));
 AND2x2_ASAP7_75t_R _25174_ (.A(_13144_),
    .B(_09688_),
    .Y(_09689_));
 AO21x1_ASAP7_75t_R _25175_ (.A1(_09579_),
    .A2(_09686_),
    .B(_09689_),
    .Y(_02967_));
 BUFx12f_ASAP7_75t_R _25176_ (.A(_08802_),
    .Y(_09690_));
 AND2x2_ASAP7_75t_R _25177_ (.A(_15386_),
    .B(_09688_),
    .Y(_09691_));
 AO21x1_ASAP7_75t_R _25178_ (.A1(_09690_),
    .A2(_09686_),
    .B(_09691_),
    .Y(_02968_));
 NOR2x1_ASAP7_75t_R _25179_ (.A(_08851_),
    .B(_09671_),
    .Y(_09692_));
 AO21x1_ASAP7_75t_R _25180_ (.A1(_15539_),
    .A2(_09671_),
    .B(_09692_),
    .Y(_02969_));
 AO21x1_ASAP7_75t_R _25181_ (.A1(_09616_),
    .A2(_09667_),
    .B(_15662_),
    .Y(_09693_));
 OA21x2_ASAP7_75t_R _25182_ (.A1(_09453_),
    .A2(_09671_),
    .B(_09693_),
    .Y(_02970_));
 AND2x2_ASAP7_75t_R _25183_ (.A(_09584_),
    .B(_09668_),
    .Y(_09694_));
 AO21x1_ASAP7_75t_R _25184_ (.A1(_15818_),
    .A2(_09671_),
    .B(_09694_),
    .Y(_02971_));
 BUFx12f_ASAP7_75t_R _25185_ (.A(_08947_),
    .Y(_09695_));
 NOR2x1_ASAP7_75t_R _25186_ (.A(_09695_),
    .B(_09671_),
    .Y(_09696_));
 AO21x1_ASAP7_75t_R _25187_ (.A1(_15900_),
    .A2(_09671_),
    .B(_09696_),
    .Y(_02972_));
 BUFx6f_ASAP7_75t_R _25188_ (.A(_09021_),
    .Y(_09697_));
 AND2x2_ASAP7_75t_R _25189_ (.A(_16065_),
    .B(_09688_),
    .Y(_09698_));
 AO21x1_ASAP7_75t_R _25190_ (.A1(_09697_),
    .A2(_09686_),
    .B(_09698_),
    .Y(_02973_));
 BUFx6f_ASAP7_75t_R _25191_ (.A(_09048_),
    .Y(_09699_));
 AND2x2_ASAP7_75t_R _25192_ (.A(_16147_),
    .B(_09688_),
    .Y(_09700_));
 AO21x1_ASAP7_75t_R _25193_ (.A1(_09699_),
    .A2(_09686_),
    .B(_09700_),
    .Y(_02974_));
 BUFx6f_ASAP7_75t_R _25194_ (.A(_09074_),
    .Y(_09701_));
 AND2x2_ASAP7_75t_R _25195_ (.A(_16282_),
    .B(_09688_),
    .Y(_09702_));
 AO21x1_ASAP7_75t_R _25196_ (.A1(_09701_),
    .A2(_09686_),
    .B(_09702_),
    .Y(_02975_));
 AND2x2_ASAP7_75t_R _25197_ (.A(_16405_),
    .B(_09688_),
    .Y(_09703_));
 AO21x1_ASAP7_75t_R _25198_ (.A1(_09594_),
    .A2(_09686_),
    .B(_09703_),
    .Y(_02976_));
 AND2x2_ASAP7_75t_R _25199_ (.A(_16543_),
    .B(_09688_),
    .Y(_09704_));
 AO21x1_ASAP7_75t_R _25200_ (.A1(_09596_),
    .A2(_09686_),
    .B(_09704_),
    .Y(_02977_));
 AND2x2_ASAP7_75t_R _25201_ (.A(_16653_),
    .B(_09688_),
    .Y(_09705_));
 AO21x1_ASAP7_75t_R _25202_ (.A1(_09598_),
    .A2(_09686_),
    .B(_09705_),
    .Y(_02978_));
 BUFx6f_ASAP7_75t_R _25203_ (.A(_09176_),
    .Y(_09706_));
 AND2x2_ASAP7_75t_R _25204_ (.A(_16776_),
    .B(_09688_),
    .Y(_09707_));
 AO21x1_ASAP7_75t_R _25205_ (.A1(_09706_),
    .A2(_09686_),
    .B(_09707_),
    .Y(_02979_));
 BUFx6f_ASAP7_75t_R _25206_ (.A(_09203_),
    .Y(_09708_));
 AND2x2_ASAP7_75t_R _25207_ (.A(_16918_),
    .B(_09688_),
    .Y(_09709_));
 AO21x1_ASAP7_75t_R _25208_ (.A1(_09708_),
    .A2(_09668_),
    .B(_09709_),
    .Y(_02980_));
 AND2x2_ASAP7_75t_R _25209_ (.A(_04261_),
    .B(_09670_),
    .Y(_09710_));
 AO21x1_ASAP7_75t_R _25210_ (.A1(_09604_),
    .A2(_09668_),
    .B(_09710_),
    .Y(_02981_));
 AND2x2_ASAP7_75t_R _25211_ (.A(_04374_),
    .B(_09670_),
    .Y(_09711_));
 AO21x1_ASAP7_75t_R _25212_ (.A1(_09606_),
    .A2(_09668_),
    .B(_09711_),
    .Y(_02982_));
 AND2x2_ASAP7_75t_R _25213_ (.A(_04541_),
    .B(_09670_),
    .Y(_09712_));
 AO21x1_ASAP7_75t_R _25214_ (.A1(_09608_),
    .A2(_09668_),
    .B(_09712_),
    .Y(_02983_));
 BUFx6f_ASAP7_75t_R _25215_ (.A(_09334_),
    .Y(_09713_));
 AND2x2_ASAP7_75t_R _25216_ (.A(_04622_),
    .B(_09670_),
    .Y(_09714_));
 AO21x1_ASAP7_75t_R _25217_ (.A1(_09713_),
    .A2(_09668_),
    .B(_09714_),
    .Y(_02984_));
 AO21x1_ASAP7_75t_R _25218_ (.A1(_09616_),
    .A2(_09667_),
    .B(_04744_),
    .Y(_09715_));
 OA21x2_ASAP7_75t_R _25219_ (.A1(_09612_),
    .A2(_09671_),
    .B(_09715_),
    .Y(_02985_));
 AND2x2_ASAP7_75t_R _25220_ (.A(_04889_),
    .B(_09670_),
    .Y(_09716_));
 AO21x1_ASAP7_75t_R _25221_ (.A1(_09614_),
    .A2(_09668_),
    .B(_09716_),
    .Y(_02986_));
 AND2x6_ASAP7_75t_R _25222_ (.A(_08954_),
    .B(_09616_),
    .Y(_09717_));
 BUFx6f_ASAP7_75t_R _25223_ (.A(_09717_),
    .Y(_09718_));
 NAND2x2_ASAP7_75t_R _25224_ (.A(_08953_),
    .B(_09616_),
    .Y(_09719_));
 BUFx12f_ASAP7_75t_R _25225_ (.A(_09719_),
    .Y(_09720_));
 AND2x2_ASAP7_75t_R _25226_ (.A(_00386_),
    .B(_09720_),
    .Y(_09721_));
 AOI21x1_ASAP7_75t_R _25227_ (.A1(_09503_),
    .A2(_09718_),
    .B(_09721_),
    .Y(_02987_));
 BUFx6f_ASAP7_75t_R _25228_ (.A(_09719_),
    .Y(_09722_));
 AND2x2_ASAP7_75t_R _25229_ (.A(_00419_),
    .B(_09722_),
    .Y(_09723_));
 AOI21x1_ASAP7_75t_R _25230_ (.A1(_09527_),
    .A2(_09718_),
    .B(_09723_),
    .Y(_02988_));
 NOR2x1_ASAP7_75t_R _25231_ (.A(_09675_),
    .B(_09720_),
    .Y(_09724_));
 AO21x1_ASAP7_75t_R _25232_ (.A1(_13559_),
    .A2(_09720_),
    .B(_09724_),
    .Y(_02989_));
 AND2x2_ASAP7_75t_R _25233_ (.A(_13676_),
    .B(_09722_),
    .Y(_09725_));
 AO21x1_ASAP7_75t_R _25234_ (.A1(_09629_),
    .A2(_09718_),
    .B(_09725_),
    .Y(_02990_));
 BUFx6f_ASAP7_75t_R _25235_ (.A(_08992_),
    .Y(_09726_));
 AND2x2_ASAP7_75t_R _25236_ (.A(_14791_),
    .B(_09722_),
    .Y(_09727_));
 AO21x1_ASAP7_75t_R _25237_ (.A1(_09726_),
    .A2(_09718_),
    .B(_09727_),
    .Y(_02991_));
 AND2x2_ASAP7_75t_R _25238_ (.A(_13770_),
    .B(_09722_),
    .Y(_09728_));
 AO21x1_ASAP7_75t_R _25239_ (.A1(_09679_),
    .A2(_09718_),
    .B(_09728_),
    .Y(_02992_));
 BUFx6f_ASAP7_75t_R _25240_ (.A(_09411_),
    .Y(_09729_));
 AND2x2_ASAP7_75t_R _25241_ (.A(_13897_),
    .B(_09722_),
    .Y(_09730_));
 AO21x1_ASAP7_75t_R _25242_ (.A1(_09729_),
    .A2(_09718_),
    .B(_09730_),
    .Y(_02993_));
 BUFx6f_ASAP7_75t_R _25243_ (.A(_09435_),
    .Y(_09731_));
 AND2x2_ASAP7_75t_R _25244_ (.A(_13959_),
    .B(_09722_),
    .Y(_09732_));
 AO21x1_ASAP7_75t_R _25245_ (.A1(_09731_),
    .A2(_09718_),
    .B(_09732_),
    .Y(_02994_));
 AND2x2_ASAP7_75t_R _25246_ (.A(_14013_),
    .B(_09722_),
    .Y(_09733_));
 AO21x1_ASAP7_75t_R _25247_ (.A1(_09572_),
    .A2(_09718_),
    .B(_09733_),
    .Y(_02995_));
 AND2x2_ASAP7_75t_R _25248_ (.A(_14029_),
    .B(_09722_),
    .Y(_09734_));
 AO21x1_ASAP7_75t_R _25249_ (.A1(_09441_),
    .A2(_09718_),
    .B(_09734_),
    .Y(_02996_));
 AND2x2_ASAP7_75t_R _25250_ (.A(_14174_),
    .B(_09722_),
    .Y(_09735_));
 AO21x1_ASAP7_75t_R _25251_ (.A1(_09575_),
    .A2(_09718_),
    .B(_09735_),
    .Y(_02997_));
 BUFx6f_ASAP7_75t_R _25252_ (.A(_08719_),
    .Y(_09736_));
 BUFx12f_ASAP7_75t_R _25253_ (.A(_09717_),
    .Y(_09737_));
 AND2x2_ASAP7_75t_R _25254_ (.A(_14211_),
    .B(_09722_),
    .Y(_09738_));
 AO21x1_ASAP7_75t_R _25255_ (.A1(_09736_),
    .A2(_09737_),
    .B(_09738_),
    .Y(_02998_));
 BUFx6f_ASAP7_75t_R _25256_ (.A(_09719_),
    .Y(_09739_));
 AND2x2_ASAP7_75t_R _25257_ (.A(_13134_),
    .B(_09739_),
    .Y(_09740_));
 AO21x1_ASAP7_75t_R _25258_ (.A1(_09579_),
    .A2(_09737_),
    .B(_09740_),
    .Y(_02999_));
 AND2x2_ASAP7_75t_R _25259_ (.A(_15383_),
    .B(_09739_),
    .Y(_09741_));
 AO21x1_ASAP7_75t_R _25260_ (.A1(_09690_),
    .A2(_09737_),
    .B(_09741_),
    .Y(_03000_));
 NOR2x1_ASAP7_75t_R _25261_ (.A(_08851_),
    .B(_09720_),
    .Y(_09742_));
 AO21x1_ASAP7_75t_R _25262_ (.A1(_15536_),
    .A2(_09720_),
    .B(_09742_),
    .Y(_03001_));
 AO21x1_ASAP7_75t_R _25263_ (.A1(_08954_),
    .A2(_09616_),
    .B(_15659_),
    .Y(_09743_));
 OA21x2_ASAP7_75t_R _25264_ (.A1(_09453_),
    .A2(_09720_),
    .B(_09743_),
    .Y(_03002_));
 AND2x2_ASAP7_75t_R _25265_ (.A(_09584_),
    .B(_09717_),
    .Y(_09744_));
 AO21x1_ASAP7_75t_R _25266_ (.A1(_15815_),
    .A2(_09720_),
    .B(_09744_),
    .Y(_03003_));
 NOR2x1_ASAP7_75t_R _25267_ (.A(_09695_),
    .B(_09720_),
    .Y(_09745_));
 AO21x1_ASAP7_75t_R _25268_ (.A1(_15897_),
    .A2(_09720_),
    .B(_09745_),
    .Y(_03004_));
 AND2x2_ASAP7_75t_R _25269_ (.A(_16062_),
    .B(_09739_),
    .Y(_09746_));
 AO21x1_ASAP7_75t_R _25270_ (.A1(_09697_),
    .A2(_09737_),
    .B(_09746_),
    .Y(_03005_));
 AND2x2_ASAP7_75t_R _25271_ (.A(_16144_),
    .B(_09739_),
    .Y(_09747_));
 AO21x1_ASAP7_75t_R _25272_ (.A1(_09699_),
    .A2(_09737_),
    .B(_09747_),
    .Y(_03006_));
 AND2x2_ASAP7_75t_R _25273_ (.A(_16279_),
    .B(_09739_),
    .Y(_09748_));
 AO21x1_ASAP7_75t_R _25274_ (.A1(_09701_),
    .A2(_09737_),
    .B(_09748_),
    .Y(_03007_));
 BUFx6f_ASAP7_75t_R _25275_ (.A(_09099_),
    .Y(_09749_));
 AND2x2_ASAP7_75t_R _25276_ (.A(_16402_),
    .B(_09739_),
    .Y(_09750_));
 AO21x1_ASAP7_75t_R _25277_ (.A1(_09749_),
    .A2(_09737_),
    .B(_09750_),
    .Y(_03008_));
 BUFx6f_ASAP7_75t_R _25278_ (.A(_09123_),
    .Y(_09751_));
 AND2x2_ASAP7_75t_R _25279_ (.A(_16540_),
    .B(_09739_),
    .Y(_09752_));
 AO21x1_ASAP7_75t_R _25280_ (.A1(_09751_),
    .A2(_09737_),
    .B(_09752_),
    .Y(_03009_));
 BUFx6f_ASAP7_75t_R _25281_ (.A(_09144_),
    .Y(_09753_));
 AND2x2_ASAP7_75t_R _25282_ (.A(_16650_),
    .B(_09739_),
    .Y(_09754_));
 AO21x1_ASAP7_75t_R _25283_ (.A1(_09753_),
    .A2(_09737_),
    .B(_09754_),
    .Y(_03010_));
 AND2x2_ASAP7_75t_R _25284_ (.A(_16773_),
    .B(_09739_),
    .Y(_09755_));
 AO21x1_ASAP7_75t_R _25285_ (.A1(_09706_),
    .A2(_09737_),
    .B(_09755_),
    .Y(_03011_));
 AND2x2_ASAP7_75t_R _25286_ (.A(_16915_),
    .B(_09739_),
    .Y(_09756_));
 AO21x1_ASAP7_75t_R _25287_ (.A1(_09708_),
    .A2(_09717_),
    .B(_09756_),
    .Y(_03012_));
 BUFx6f_ASAP7_75t_R _25288_ (.A(_09229_),
    .Y(_09757_));
 AND2x2_ASAP7_75t_R _25289_ (.A(_04258_),
    .B(_09719_),
    .Y(_09758_));
 AO21x1_ASAP7_75t_R _25290_ (.A1(_09757_),
    .A2(_09717_),
    .B(_09758_),
    .Y(_03013_));
 BUFx6f_ASAP7_75t_R _25291_ (.A(_09249_),
    .Y(_09759_));
 AND2x2_ASAP7_75t_R _25292_ (.A(_04371_),
    .B(_09719_),
    .Y(_09760_));
 AO21x1_ASAP7_75t_R _25293_ (.A1(_09759_),
    .A2(_09717_),
    .B(_09760_),
    .Y(_03014_));
 BUFx6f_ASAP7_75t_R _25294_ (.A(_09301_),
    .Y(_09761_));
 AND2x2_ASAP7_75t_R _25295_ (.A(_04538_),
    .B(_09719_),
    .Y(_09762_));
 AO21x1_ASAP7_75t_R _25296_ (.A1(_09761_),
    .A2(_09717_),
    .B(_09762_),
    .Y(_03015_));
 AND2x2_ASAP7_75t_R _25297_ (.A(_04619_),
    .B(_09719_),
    .Y(_09763_));
 AO21x1_ASAP7_75t_R _25298_ (.A1(_09713_),
    .A2(_09717_),
    .B(_09763_),
    .Y(_03016_));
 AO21x1_ASAP7_75t_R _25299_ (.A1(_08954_),
    .A2(_09616_),
    .B(_04741_),
    .Y(_09764_));
 OA21x2_ASAP7_75t_R _25300_ (.A1(_09612_),
    .A2(_09720_),
    .B(_09764_),
    .Y(_03017_));
 AND2x2_ASAP7_75t_R _25301_ (.A(_04886_),
    .B(_09719_),
    .Y(_09765_));
 AO21x1_ASAP7_75t_R _25302_ (.A1(_09614_),
    .A2(_09717_),
    .B(_09765_),
    .Y(_03018_));
 AND2x6_ASAP7_75t_R _25303_ (.A(_13686_),
    .B(_13602_),
    .Y(_09766_));
 AND5x2_ASAP7_75t_R _25304_ (.A(_07799_),
    .B(_13455_),
    .C(_13430_),
    .D(_09475_),
    .E(_09766_),
    .Y(_09767_));
 BUFx12f_ASAP7_75t_R _25305_ (.A(_09767_),
    .Y(_09768_));
 BUFx12f_ASAP7_75t_R _25306_ (.A(_09768_),
    .Y(_09769_));
 NAND2x2_ASAP7_75t_R _25307_ (.A(_13686_),
    .B(_13602_),
    .Y(_09770_));
 OR4x1_ASAP7_75t_R _25308_ (.A(_13692_),
    .B(_09504_),
    .C(_09505_),
    .D(_09770_),
    .Y(_09771_));
 BUFx6f_ASAP7_75t_R _25309_ (.A(_09771_),
    .Y(_09772_));
 AND2x2_ASAP7_75t_R _25310_ (.A(_00387_),
    .B(_09772_),
    .Y(_09773_));
 AOI21x1_ASAP7_75t_R _25311_ (.A1(_09503_),
    .A2(_09769_),
    .B(_09773_),
    .Y(_03019_));
 AND2x2_ASAP7_75t_R _25312_ (.A(_00420_),
    .B(_09772_),
    .Y(_09774_));
 AOI21x1_ASAP7_75t_R _25313_ (.A1(_09527_),
    .A2(_09769_),
    .B(_09774_),
    .Y(_03020_));
 AND2x2_ASAP7_75t_R _25314_ (.A(_00451_),
    .B(_09772_),
    .Y(_09775_));
 AOI21x1_ASAP7_75t_R _25315_ (.A1(_09675_),
    .A2(_09769_),
    .B(_09775_),
    .Y(_03021_));
 BUFx12f_ASAP7_75t_R _25316_ (.A(_09768_),
    .Y(_09776_));
 NOR2x1_ASAP7_75t_R _25317_ (.A(_00481_),
    .B(_09776_),
    .Y(_09777_));
 AO21x1_ASAP7_75t_R _25318_ (.A1(_09629_),
    .A2(_09769_),
    .B(_09777_),
    .Y(_03022_));
 NOR2x1_ASAP7_75t_R _25319_ (.A(_00511_),
    .B(_09776_),
    .Y(_09778_));
 AO21x1_ASAP7_75t_R _25320_ (.A1(_09726_),
    .A2(_09769_),
    .B(_09778_),
    .Y(_03023_));
 NOR2x1_ASAP7_75t_R _25321_ (.A(_00541_),
    .B(_09776_),
    .Y(_09779_));
 AO21x1_ASAP7_75t_R _25322_ (.A1(_09679_),
    .A2(_09769_),
    .B(_09779_),
    .Y(_03024_));
 NOR2x1_ASAP7_75t_R _25323_ (.A(_00571_),
    .B(_09776_),
    .Y(_09780_));
 AO21x1_ASAP7_75t_R _25324_ (.A1(_09729_),
    .A2(_09769_),
    .B(_09780_),
    .Y(_03025_));
 NOR2x1_ASAP7_75t_R _25325_ (.A(_00601_),
    .B(_09776_),
    .Y(_09781_));
 AO21x1_ASAP7_75t_R _25326_ (.A1(_09731_),
    .A2(_09769_),
    .B(_09781_),
    .Y(_03026_));
 BUFx12f_ASAP7_75t_R _25327_ (.A(_09768_),
    .Y(_09782_));
 NOR2x1_ASAP7_75t_R _25328_ (.A(_00631_),
    .B(_09776_),
    .Y(_09783_));
 AO21x1_ASAP7_75t_R _25329_ (.A1(_09572_),
    .A2(_09782_),
    .B(_09783_),
    .Y(_03027_));
 BUFx6f_ASAP7_75t_R _25330_ (.A(_08615_),
    .Y(_09784_));
 AND2x2_ASAP7_75t_R _25331_ (.A(_14057_),
    .B(_09772_),
    .Y(_09785_));
 AO21x1_ASAP7_75t_R _25332_ (.A1(_09784_),
    .A2(_09782_),
    .B(_09785_),
    .Y(_03028_));
 NOR2x1_ASAP7_75t_R _25333_ (.A(_00691_),
    .B(_09776_),
    .Y(_09786_));
 AO21x1_ASAP7_75t_R _25334_ (.A1(_09575_),
    .A2(_09782_),
    .B(_09786_),
    .Y(_03029_));
 NOR2x1_ASAP7_75t_R _25335_ (.A(_00721_),
    .B(_09776_),
    .Y(_09787_));
 AO21x1_ASAP7_75t_R _25336_ (.A1(_09736_),
    .A2(_09782_),
    .B(_09787_),
    .Y(_03030_));
 NOR2x1_ASAP7_75t_R _25337_ (.A(_00351_),
    .B(_09776_),
    .Y(_09788_));
 AO21x1_ASAP7_75t_R _25338_ (.A1(_09579_),
    .A2(_09782_),
    .B(_09788_),
    .Y(_03031_));
 NOR2x1_ASAP7_75t_R _25339_ (.A(_00789_),
    .B(_09776_),
    .Y(_09789_));
 AO21x1_ASAP7_75t_R _25340_ (.A1(_09690_),
    .A2(_09782_),
    .B(_09789_),
    .Y(_03032_));
 BUFx12f_ASAP7_75t_R _25341_ (.A(_09451_),
    .Y(_09790_));
 AND2x2_ASAP7_75t_R _25342_ (.A(_00821_),
    .B(_09772_),
    .Y(_09791_));
 AOI21x1_ASAP7_75t_R _25343_ (.A1(_09790_),
    .A2(_09769_),
    .B(_09791_),
    .Y(_03033_));
 NAND2x1_ASAP7_75t_R _25344_ (.A(_00853_),
    .B(_09772_),
    .Y(_09792_));
 OA21x2_ASAP7_75t_R _25345_ (.A1(_09453_),
    .A2(_09772_),
    .B(_09792_),
    .Y(_03034_));
 BUFx12f_ASAP7_75t_R _25346_ (.A(_09768_),
    .Y(_09793_));
 NOR2x1_ASAP7_75t_R _25347_ (.A(_00885_),
    .B(_09793_),
    .Y(_09794_));
 AO21x1_ASAP7_75t_R _25348_ (.A1(_09584_),
    .A2(_09782_),
    .B(_09794_),
    .Y(_03035_));
 AND2x2_ASAP7_75t_R _25349_ (.A(_00917_),
    .B(_09772_),
    .Y(_09795_));
 AOI21x1_ASAP7_75t_R _25350_ (.A1(_08948_),
    .A2(_09769_),
    .B(_09795_),
    .Y(_03036_));
 NOR2x1_ASAP7_75t_R _25351_ (.A(_00949_),
    .B(_09793_),
    .Y(_09796_));
 AO21x1_ASAP7_75t_R _25352_ (.A1(_09697_),
    .A2(_09782_),
    .B(_09796_),
    .Y(_03037_));
 NOR2x1_ASAP7_75t_R _25353_ (.A(_00981_),
    .B(_09793_),
    .Y(_09797_));
 AO21x1_ASAP7_75t_R _25354_ (.A1(_09699_),
    .A2(_09782_),
    .B(_09797_),
    .Y(_03038_));
 NOR2x1_ASAP7_75t_R _25355_ (.A(_01013_),
    .B(_09793_),
    .Y(_09798_));
 AO21x1_ASAP7_75t_R _25356_ (.A1(_09701_),
    .A2(_09782_),
    .B(_09798_),
    .Y(_03039_));
 BUFx6f_ASAP7_75t_R _25357_ (.A(_09768_),
    .Y(_09799_));
 NOR2x1_ASAP7_75t_R _25358_ (.A(_01045_),
    .B(_09793_),
    .Y(_09800_));
 AO21x1_ASAP7_75t_R _25359_ (.A1(_09749_),
    .A2(_09799_),
    .B(_09800_),
    .Y(_03040_));
 NOR2x1_ASAP7_75t_R _25360_ (.A(_01077_),
    .B(_09793_),
    .Y(_09801_));
 AO21x1_ASAP7_75t_R _25361_ (.A1(_09751_),
    .A2(_09799_),
    .B(_09801_),
    .Y(_03041_));
 NOR2x1_ASAP7_75t_R _25362_ (.A(_01109_),
    .B(_09793_),
    .Y(_09802_));
 AO21x1_ASAP7_75t_R _25363_ (.A1(_09753_),
    .A2(_09799_),
    .B(_09802_),
    .Y(_03042_));
 NOR2x1_ASAP7_75t_R _25364_ (.A(_01141_),
    .B(_09793_),
    .Y(_09803_));
 AO21x1_ASAP7_75t_R _25365_ (.A1(_09706_),
    .A2(_09799_),
    .B(_09803_),
    .Y(_03043_));
 NOR2x1_ASAP7_75t_R _25366_ (.A(_01173_),
    .B(_09793_),
    .Y(_09804_));
 AO21x1_ASAP7_75t_R _25367_ (.A1(_09708_),
    .A2(_09799_),
    .B(_09804_),
    .Y(_03044_));
 NOR2x1_ASAP7_75t_R _25368_ (.A(_01205_),
    .B(_09793_),
    .Y(_09805_));
 AO21x1_ASAP7_75t_R _25369_ (.A1(_09757_),
    .A2(_09799_),
    .B(_09805_),
    .Y(_03045_));
 NOR2x1_ASAP7_75t_R _25370_ (.A(_01237_),
    .B(_09768_),
    .Y(_09806_));
 AO21x1_ASAP7_75t_R _25371_ (.A1(_09759_),
    .A2(_09799_),
    .B(_09806_),
    .Y(_03046_));
 NOR2x1_ASAP7_75t_R _25372_ (.A(_01269_),
    .B(_09768_),
    .Y(_09807_));
 AO21x1_ASAP7_75t_R _25373_ (.A1(_09761_),
    .A2(_09799_),
    .B(_09807_),
    .Y(_03047_));
 NOR2x1_ASAP7_75t_R _25374_ (.A(_01301_),
    .B(_09768_),
    .Y(_09808_));
 AO21x1_ASAP7_75t_R _25375_ (.A1(_09713_),
    .A2(_09799_),
    .B(_09808_),
    .Y(_03048_));
 NAND2x1_ASAP7_75t_R _25376_ (.A(_01333_),
    .B(_09772_),
    .Y(_09809_));
 OA21x2_ASAP7_75t_R _25377_ (.A1(_09612_),
    .A2(_09772_),
    .B(_09809_),
    .Y(_03049_));
 BUFx6f_ASAP7_75t_R _25378_ (.A(_09392_),
    .Y(_09810_));
 NOR2x1_ASAP7_75t_R _25379_ (.A(_01365_),
    .B(_09768_),
    .Y(_09811_));
 AO21x1_ASAP7_75t_R _25380_ (.A1(_09810_),
    .A2(_09799_),
    .B(_09811_),
    .Y(_03050_));
 BUFx6f_ASAP7_75t_R _25381_ (.A(_09766_),
    .Y(_09812_));
 AND2x6_ASAP7_75t_R _25382_ (.A(_09621_),
    .B(_09812_),
    .Y(_09813_));
 BUFx6f_ASAP7_75t_R _25383_ (.A(_09813_),
    .Y(_09814_));
 NAND2x2_ASAP7_75t_R _25384_ (.A(_09621_),
    .B(_09812_),
    .Y(_09815_));
 AND2x2_ASAP7_75t_R _25385_ (.A(_00388_),
    .B(_09815_),
    .Y(_09816_));
 AOI21x1_ASAP7_75t_R _25386_ (.A1(_09503_),
    .A2(_09814_),
    .B(_09816_),
    .Y(_03051_));
 AND2x2_ASAP7_75t_R _25387_ (.A(_00421_),
    .B(_09815_),
    .Y(_09817_));
 AOI21x1_ASAP7_75t_R _25388_ (.A1(_09527_),
    .A2(_09814_),
    .B(_09817_),
    .Y(_03052_));
 AO21x1_ASAP7_75t_R _25389_ (.A1(_09621_),
    .A2(_09812_),
    .B(_00452_),
    .Y(_09818_));
 OAI21x1_ASAP7_75t_R _25390_ (.A1(_09675_),
    .A2(_09815_),
    .B(_09818_),
    .Y(_03053_));
 BUFx12f_ASAP7_75t_R _25391_ (.A(_09559_),
    .Y(_09819_));
 AND2x2_ASAP7_75t_R _25392_ (.A(_13642_),
    .B(_09815_),
    .Y(_09820_));
 AO21x1_ASAP7_75t_R _25393_ (.A1(_09819_),
    .A2(_09814_),
    .B(_09820_),
    .Y(_03054_));
 BUFx12f_ASAP7_75t_R _25394_ (.A(_09813_),
    .Y(_09821_));
 NOR2x1_ASAP7_75t_R _25395_ (.A(_00512_),
    .B(_09821_),
    .Y(_09822_));
 AO21x1_ASAP7_75t_R _25396_ (.A1(_09726_),
    .A2(_09814_),
    .B(_09822_),
    .Y(_03055_));
 NOR2x1_ASAP7_75t_R _25397_ (.A(_00542_),
    .B(_09821_),
    .Y(_09823_));
 AO21x1_ASAP7_75t_R _25398_ (.A1(_09679_),
    .A2(_09814_),
    .B(_09823_),
    .Y(_03056_));
 NOR2x1_ASAP7_75t_R _25399_ (.A(_00572_),
    .B(_09821_),
    .Y(_09824_));
 AO21x1_ASAP7_75t_R _25400_ (.A1(_09729_),
    .A2(_09814_),
    .B(_09824_),
    .Y(_03057_));
 BUFx12f_ASAP7_75t_R _25401_ (.A(_09813_),
    .Y(_09825_));
 NOR2x1_ASAP7_75t_R _25402_ (.A(_00602_),
    .B(_09825_),
    .Y(_09826_));
 AO21x1_ASAP7_75t_R _25403_ (.A1(_09731_),
    .A2(_09814_),
    .B(_09826_),
    .Y(_03058_));
 NOR2x1_ASAP7_75t_R _25404_ (.A(_00632_),
    .B(_09825_),
    .Y(_09827_));
 AO21x1_ASAP7_75t_R _25405_ (.A1(_09572_),
    .A2(_09814_),
    .B(_09827_),
    .Y(_03059_));
 NOR2x1_ASAP7_75t_R _25406_ (.A(_00662_),
    .B(_09825_),
    .Y(_09828_));
 AO21x1_ASAP7_75t_R _25407_ (.A1(_09784_),
    .A2(_09814_),
    .B(_09828_),
    .Y(_03060_));
 NOR2x1_ASAP7_75t_R _25408_ (.A(_00692_),
    .B(_09825_),
    .Y(_09829_));
 AO21x1_ASAP7_75t_R _25409_ (.A1(_09575_),
    .A2(_09814_),
    .B(_09829_),
    .Y(_03061_));
 BUFx12f_ASAP7_75t_R _25410_ (.A(_09813_),
    .Y(_09830_));
 NOR2x1_ASAP7_75t_R _25411_ (.A(_00722_),
    .B(_09825_),
    .Y(_09831_));
 AO21x1_ASAP7_75t_R _25412_ (.A1(_09736_),
    .A2(_09830_),
    .B(_09831_),
    .Y(_03062_));
 NOR2x1_ASAP7_75t_R _25413_ (.A(_00352_),
    .B(_09825_),
    .Y(_09832_));
 AO21x1_ASAP7_75t_R _25414_ (.A1(_09579_),
    .A2(_09830_),
    .B(_09832_),
    .Y(_03063_));
 NOR2x1_ASAP7_75t_R _25415_ (.A(_00790_),
    .B(_09825_),
    .Y(_09833_));
 AO21x1_ASAP7_75t_R _25416_ (.A1(_09690_),
    .A2(_09830_),
    .B(_09833_),
    .Y(_03064_));
 AO21x1_ASAP7_75t_R _25417_ (.A1(_09621_),
    .A2(_09812_),
    .B(_00822_),
    .Y(_09834_));
 OAI21x1_ASAP7_75t_R _25418_ (.A1(_09790_),
    .A2(_09815_),
    .B(_09834_),
    .Y(_03065_));
 NAND2x1_ASAP7_75t_R _25419_ (.A(_00854_),
    .B(_09815_),
    .Y(_09835_));
 OA21x2_ASAP7_75t_R _25420_ (.A1(_09453_),
    .A2(_09815_),
    .B(_09835_),
    .Y(_03066_));
 NOR2x1_ASAP7_75t_R _25421_ (.A(_00886_),
    .B(_09825_),
    .Y(_09836_));
 AO21x1_ASAP7_75t_R _25422_ (.A1(_09584_),
    .A2(_09830_),
    .B(_09836_),
    .Y(_03067_));
 AO21x1_ASAP7_75t_R _25423_ (.A1(_09621_),
    .A2(_09812_),
    .B(_00918_),
    .Y(_09837_));
 OAI21x1_ASAP7_75t_R _25424_ (.A1(_08948_),
    .A2(_09815_),
    .B(_09837_),
    .Y(_03068_));
 NOR2x1_ASAP7_75t_R _25425_ (.A(_00950_),
    .B(_09825_),
    .Y(_09838_));
 AO21x1_ASAP7_75t_R _25426_ (.A1(_09697_),
    .A2(_09830_),
    .B(_09838_),
    .Y(_03069_));
 NOR2x1_ASAP7_75t_R _25427_ (.A(_00982_),
    .B(_09825_),
    .Y(_09839_));
 AO21x1_ASAP7_75t_R _25428_ (.A1(_09699_),
    .A2(_09830_),
    .B(_09839_),
    .Y(_03070_));
 BUFx12f_ASAP7_75t_R _25429_ (.A(_09813_),
    .Y(_09840_));
 NOR2x1_ASAP7_75t_R _25430_ (.A(_01014_),
    .B(_09840_),
    .Y(_09841_));
 AO21x1_ASAP7_75t_R _25431_ (.A1(_09701_),
    .A2(_09830_),
    .B(_09841_),
    .Y(_03071_));
 NOR2x1_ASAP7_75t_R _25432_ (.A(_01046_),
    .B(_09840_),
    .Y(_09842_));
 AO21x1_ASAP7_75t_R _25433_ (.A1(_09749_),
    .A2(_09830_),
    .B(_09842_),
    .Y(_03072_));
 NOR2x1_ASAP7_75t_R _25434_ (.A(_01078_),
    .B(_09840_),
    .Y(_09843_));
 AO21x1_ASAP7_75t_R _25435_ (.A1(_09751_),
    .A2(_09830_),
    .B(_09843_),
    .Y(_03073_));
 NOR2x1_ASAP7_75t_R _25436_ (.A(_01110_),
    .B(_09840_),
    .Y(_09844_));
 AO21x1_ASAP7_75t_R _25437_ (.A1(_09753_),
    .A2(_09830_),
    .B(_09844_),
    .Y(_03074_));
 NOR2x1_ASAP7_75t_R _25438_ (.A(_01142_),
    .B(_09840_),
    .Y(_09845_));
 AO21x1_ASAP7_75t_R _25439_ (.A1(_09706_),
    .A2(_09821_),
    .B(_09845_),
    .Y(_03075_));
 NOR2x1_ASAP7_75t_R _25440_ (.A(_01174_),
    .B(_09840_),
    .Y(_09846_));
 AO21x1_ASAP7_75t_R _25441_ (.A1(_09708_),
    .A2(_09821_),
    .B(_09846_),
    .Y(_03076_));
 NOR2x1_ASAP7_75t_R _25442_ (.A(_01206_),
    .B(_09840_),
    .Y(_09847_));
 AO21x1_ASAP7_75t_R _25443_ (.A1(_09757_),
    .A2(_09821_),
    .B(_09847_),
    .Y(_03077_));
 NOR2x1_ASAP7_75t_R _25444_ (.A(_01238_),
    .B(_09840_),
    .Y(_09848_));
 AO21x1_ASAP7_75t_R _25445_ (.A1(_09759_),
    .A2(_09821_),
    .B(_09848_),
    .Y(_03078_));
 NOR2x1_ASAP7_75t_R _25446_ (.A(_01270_),
    .B(_09840_),
    .Y(_09849_));
 AO21x1_ASAP7_75t_R _25447_ (.A1(_09761_),
    .A2(_09821_),
    .B(_09849_),
    .Y(_03079_));
 NOR2x1_ASAP7_75t_R _25448_ (.A(_01302_),
    .B(_09840_),
    .Y(_09850_));
 AO21x1_ASAP7_75t_R _25449_ (.A1(_09713_),
    .A2(_09821_),
    .B(_09850_),
    .Y(_03080_));
 NAND2x1_ASAP7_75t_R _25450_ (.A(_01334_),
    .B(_09815_),
    .Y(_09851_));
 OA21x2_ASAP7_75t_R _25451_ (.A1(_09612_),
    .A2(_09815_),
    .B(_09851_),
    .Y(_03081_));
 NOR2x1_ASAP7_75t_R _25452_ (.A(_01366_),
    .B(_09813_),
    .Y(_09852_));
 AO21x1_ASAP7_75t_R _25453_ (.A1(_09810_),
    .A2(_09821_),
    .B(_09852_),
    .Y(_03082_));
 AND2x6_ASAP7_75t_R _25454_ (.A(_09666_),
    .B(_09766_),
    .Y(_09853_));
 BUFx12f_ASAP7_75t_R _25455_ (.A(_09853_),
    .Y(_09854_));
 NAND2x2_ASAP7_75t_R _25456_ (.A(_09666_),
    .B(_09766_),
    .Y(_09855_));
 BUFx6f_ASAP7_75t_R _25457_ (.A(_09855_),
    .Y(_09856_));
 AND2x2_ASAP7_75t_R _25458_ (.A(_00389_),
    .B(_09856_),
    .Y(_09857_));
 AOI21x1_ASAP7_75t_R _25459_ (.A1(_09503_),
    .A2(_09854_),
    .B(_09857_),
    .Y(_03083_));
 AND2x2_ASAP7_75t_R _25460_ (.A(_00422_),
    .B(_09856_),
    .Y(_09858_));
 AOI21x1_ASAP7_75t_R _25461_ (.A1(_09527_),
    .A2(_09854_),
    .B(_09858_),
    .Y(_03084_));
 NOR2x1_ASAP7_75t_R _25462_ (.A(_09675_),
    .B(_09856_),
    .Y(_09859_));
 AO21x1_ASAP7_75t_R _25463_ (.A1(_14660_),
    .A2(_09856_),
    .B(_09859_),
    .Y(_03085_));
 AND2x2_ASAP7_75t_R _25464_ (.A(_13645_),
    .B(_09856_),
    .Y(_09860_));
 AO21x1_ASAP7_75t_R _25465_ (.A1(_09819_),
    .A2(_09854_),
    .B(_09860_),
    .Y(_03086_));
 BUFx12f_ASAP7_75t_R _25466_ (.A(_09855_),
    .Y(_09861_));
 AND2x2_ASAP7_75t_R _25467_ (.A(_14786_),
    .B(_09861_),
    .Y(_09862_));
 AO21x1_ASAP7_75t_R _25468_ (.A1(_09726_),
    .A2(_09854_),
    .B(_09862_),
    .Y(_03087_));
 AND2x2_ASAP7_75t_R _25469_ (.A(_14848_),
    .B(_09861_),
    .Y(_09863_));
 AO21x1_ASAP7_75t_R _25470_ (.A1(_09679_),
    .A2(_09854_),
    .B(_09863_),
    .Y(_03088_));
 AND2x2_ASAP7_75t_R _25471_ (.A(_14916_),
    .B(_09861_),
    .Y(_09864_));
 AO21x1_ASAP7_75t_R _25472_ (.A1(_09729_),
    .A2(_09854_),
    .B(_09864_),
    .Y(_03089_));
 AND2x2_ASAP7_75t_R _25473_ (.A(_14980_),
    .B(_09861_),
    .Y(_09865_));
 AO21x1_ASAP7_75t_R _25474_ (.A1(_09731_),
    .A2(_09854_),
    .B(_09865_),
    .Y(_03090_));
 AND2x2_ASAP7_75t_R _25475_ (.A(_15056_),
    .B(_09861_),
    .Y(_09866_));
 AO21x1_ASAP7_75t_R _25476_ (.A1(_09572_),
    .A2(_09854_),
    .B(_09866_),
    .Y(_03091_));
 AND2x2_ASAP7_75t_R _25477_ (.A(_15112_),
    .B(_09861_),
    .Y(_09867_));
 AO21x1_ASAP7_75t_R _25478_ (.A1(_09784_),
    .A2(_09854_),
    .B(_09867_),
    .Y(_03092_));
 AND2x4_ASAP7_75t_R _25479_ (.A(_08950_),
    .B(_09621_),
    .Y(_09868_));
 NAND2x2_ASAP7_75t_R _25480_ (.A(_08950_),
    .B(_09620_),
    .Y(_09869_));
 BUFx12f_ASAP7_75t_R _25481_ (.A(_09869_),
    .Y(_09870_));
 AND2x2_ASAP7_75t_R _25482_ (.A(_01796_),
    .B(_09870_),
    .Y(_09871_));
 AOI21x1_ASAP7_75t_R _25483_ (.A1(_09503_),
    .A2(_09868_),
    .B(_09871_),
    .Y(_03093_));
 BUFx12f_ASAP7_75t_R _25484_ (.A(_09853_),
    .Y(_09872_));
 BUFx12f_ASAP7_75t_R _25485_ (.A(_09872_),
    .Y(_09873_));
 AND2x2_ASAP7_75t_R _25486_ (.A(_15186_),
    .B(_09861_),
    .Y(_09874_));
 AO21x1_ASAP7_75t_R _25487_ (.A1(_09575_),
    .A2(_09873_),
    .B(_09874_),
    .Y(_03094_));
 AND2x2_ASAP7_75t_R _25488_ (.A(_14236_),
    .B(_09861_),
    .Y(_09875_));
 AO21x1_ASAP7_75t_R _25489_ (.A1(_09736_),
    .A2(_09873_),
    .B(_09875_),
    .Y(_03095_));
 AND2x2_ASAP7_75t_R _25490_ (.A(_13117_),
    .B(_09861_),
    .Y(_09876_));
 AO21x1_ASAP7_75t_R _25491_ (.A1(_09579_),
    .A2(_09873_),
    .B(_09876_),
    .Y(_03096_));
 AND2x2_ASAP7_75t_R _25492_ (.A(_15378_),
    .B(_09861_),
    .Y(_09877_));
 AO21x1_ASAP7_75t_R _25493_ (.A1(_09690_),
    .A2(_09873_),
    .B(_09877_),
    .Y(_03097_));
 NAND2x1_ASAP7_75t_R _25494_ (.A(_08851_),
    .B(_09872_),
    .Y(_09878_));
 OA21x2_ASAP7_75t_R _25495_ (.A1(_15531_),
    .A2(_09854_),
    .B(_09878_),
    .Y(_03098_));
 AO21x1_ASAP7_75t_R _25496_ (.A1(_09667_),
    .A2(_09812_),
    .B(_15654_),
    .Y(_09879_));
 OA21x2_ASAP7_75t_R _25497_ (.A1(_09453_),
    .A2(_09856_),
    .B(_09879_),
    .Y(_03099_));
 AND2x2_ASAP7_75t_R _25498_ (.A(_09584_),
    .B(_09872_),
    .Y(_09880_));
 AO21x1_ASAP7_75t_R _25499_ (.A1(_15810_),
    .A2(_09856_),
    .B(_09880_),
    .Y(_03100_));
 NOR2x1_ASAP7_75t_R _25500_ (.A(_09695_),
    .B(_09856_),
    .Y(_09881_));
 AO21x1_ASAP7_75t_R _25501_ (.A1(_15892_),
    .A2(_09856_),
    .B(_09881_),
    .Y(_03101_));
 BUFx6f_ASAP7_75t_R _25502_ (.A(_09855_),
    .Y(_09882_));
 AND2x2_ASAP7_75t_R _25503_ (.A(_16057_),
    .B(_09882_),
    .Y(_09883_));
 AO21x1_ASAP7_75t_R _25504_ (.A1(_09697_),
    .A2(_09873_),
    .B(_09883_),
    .Y(_03102_));
 AND2x2_ASAP7_75t_R _25505_ (.A(_16139_),
    .B(_09882_),
    .Y(_09884_));
 AO21x1_ASAP7_75t_R _25506_ (.A1(_09699_),
    .A2(_09873_),
    .B(_09884_),
    .Y(_03103_));
 AND2x2_ASAP7_75t_R _25507_ (.A(_01795_),
    .B(_09870_),
    .Y(_09885_));
 AOI21x1_ASAP7_75t_R _25508_ (.A1(_09527_),
    .A2(_09868_),
    .B(_09885_),
    .Y(_03104_));
 AND2x2_ASAP7_75t_R _25509_ (.A(_16274_),
    .B(_09882_),
    .Y(_09886_));
 AO21x1_ASAP7_75t_R _25510_ (.A1(_09701_),
    .A2(_09873_),
    .B(_09886_),
    .Y(_03105_));
 AND2x2_ASAP7_75t_R _25511_ (.A(_16397_),
    .B(_09882_),
    .Y(_09887_));
 AO21x1_ASAP7_75t_R _25512_ (.A1(_09749_),
    .A2(_09873_),
    .B(_09887_),
    .Y(_03106_));
 AND2x2_ASAP7_75t_R _25513_ (.A(_16535_),
    .B(_09882_),
    .Y(_09888_));
 AO21x1_ASAP7_75t_R _25514_ (.A1(_09751_),
    .A2(_09873_),
    .B(_09888_),
    .Y(_03107_));
 AND2x2_ASAP7_75t_R _25515_ (.A(_16645_),
    .B(_09882_),
    .Y(_09889_));
 AO21x1_ASAP7_75t_R _25516_ (.A1(_09753_),
    .A2(_09873_),
    .B(_09889_),
    .Y(_03108_));
 AND2x2_ASAP7_75t_R _25517_ (.A(_16768_),
    .B(_09882_),
    .Y(_09890_));
 AO21x1_ASAP7_75t_R _25518_ (.A1(_09706_),
    .A2(_09872_),
    .B(_09890_),
    .Y(_03109_));
 AND2x2_ASAP7_75t_R _25519_ (.A(_16910_),
    .B(_09882_),
    .Y(_09891_));
 AO21x1_ASAP7_75t_R _25520_ (.A1(_09708_),
    .A2(_09872_),
    .B(_09891_),
    .Y(_03110_));
 AND2x2_ASAP7_75t_R _25521_ (.A(_04253_),
    .B(_09882_),
    .Y(_09892_));
 AO21x1_ASAP7_75t_R _25522_ (.A1(_09757_),
    .A2(_09872_),
    .B(_09892_),
    .Y(_03111_));
 AND2x2_ASAP7_75t_R _25523_ (.A(_04366_),
    .B(_09882_),
    .Y(_09893_));
 AO21x1_ASAP7_75t_R _25524_ (.A1(_09759_),
    .A2(_09872_),
    .B(_09893_),
    .Y(_03112_));
 AND2x2_ASAP7_75t_R _25525_ (.A(_04533_),
    .B(_09855_),
    .Y(_09894_));
 AO21x1_ASAP7_75t_R _25526_ (.A1(_09761_),
    .A2(_09872_),
    .B(_09894_),
    .Y(_03113_));
 AND2x2_ASAP7_75t_R _25527_ (.A(_04614_),
    .B(_09855_),
    .Y(_09895_));
 AO21x1_ASAP7_75t_R _25528_ (.A1(_09713_),
    .A2(_09872_),
    .B(_09895_),
    .Y(_03114_));
 INVx1_ASAP7_75t_R _25529_ (.A(_01794_),
    .Y(_09896_));
 BUFx12f_ASAP7_75t_R _25530_ (.A(_09869_),
    .Y(_09897_));
 BUFx12f_ASAP7_75t_R _25531_ (.A(_09542_),
    .Y(_09898_));
 NOR2x1_ASAP7_75t_R _25532_ (.A(_09898_),
    .B(_09870_),
    .Y(_09899_));
 AO21x1_ASAP7_75t_R _25533_ (.A1(_09896_),
    .A2(_09897_),
    .B(_09899_),
    .Y(_03115_));
 AO21x1_ASAP7_75t_R _25534_ (.A1(_09667_),
    .A2(_09812_),
    .B(_04736_),
    .Y(_09900_));
 OA21x2_ASAP7_75t_R _25535_ (.A1(_09612_),
    .A2(_09856_),
    .B(_09900_),
    .Y(_03116_));
 AND2x2_ASAP7_75t_R _25536_ (.A(_04920_),
    .B(_09855_),
    .Y(_09901_));
 AO21x1_ASAP7_75t_R _25537_ (.A1(_09810_),
    .A2(_09872_),
    .B(_09901_),
    .Y(_03117_));
 BUFx12f_ASAP7_75t_R _25538_ (.A(_09502_),
    .Y(_09902_));
 AND2x6_ASAP7_75t_R _25539_ (.A(_08954_),
    .B(_09812_),
    .Y(_09903_));
 BUFx6f_ASAP7_75t_R _25540_ (.A(_09903_),
    .Y(_09904_));
 NAND2x2_ASAP7_75t_R _25541_ (.A(_08953_),
    .B(_09766_),
    .Y(_09905_));
 BUFx12f_ASAP7_75t_R _25542_ (.A(_09905_),
    .Y(_09906_));
 AND2x2_ASAP7_75t_R _25543_ (.A(_00390_),
    .B(_09906_),
    .Y(_09907_));
 AOI21x1_ASAP7_75t_R _25544_ (.A1(_09902_),
    .A2(_09904_),
    .B(_09907_),
    .Y(_03118_));
 BUFx12f_ASAP7_75t_R _25545_ (.A(_09526_),
    .Y(_09908_));
 BUFx6f_ASAP7_75t_R _25546_ (.A(_09905_),
    .Y(_09909_));
 AND2x2_ASAP7_75t_R _25547_ (.A(_00423_),
    .B(_09909_),
    .Y(_09910_));
 AOI21x1_ASAP7_75t_R _25548_ (.A1(_09908_),
    .A2(_09904_),
    .B(_09910_),
    .Y(_03119_));
 NOR2x1_ASAP7_75t_R _25549_ (.A(_09898_),
    .B(_09906_),
    .Y(_09911_));
 AO21x1_ASAP7_75t_R _25550_ (.A1(_14657_),
    .A2(_09906_),
    .B(_09911_),
    .Y(_03120_));
 AND2x2_ASAP7_75t_R _25551_ (.A(_14727_),
    .B(_09909_),
    .Y(_09912_));
 AO21x1_ASAP7_75t_R _25552_ (.A1(_09819_),
    .A2(_09904_),
    .B(_09912_),
    .Y(_03121_));
 AND2x2_ASAP7_75t_R _25553_ (.A(_14783_),
    .B(_09909_),
    .Y(_09913_));
 AO21x1_ASAP7_75t_R _25554_ (.A1(_09726_),
    .A2(_09904_),
    .B(_09913_),
    .Y(_03122_));
 AND2x2_ASAP7_75t_R _25555_ (.A(_14845_),
    .B(_09909_),
    .Y(_09914_));
 AO21x1_ASAP7_75t_R _25556_ (.A1(_09679_),
    .A2(_09904_),
    .B(_09914_),
    .Y(_03123_));
 AND2x2_ASAP7_75t_R _25557_ (.A(_14912_),
    .B(_09909_),
    .Y(_09915_));
 AO21x1_ASAP7_75t_R _25558_ (.A1(_09729_),
    .A2(_09904_),
    .B(_09915_),
    .Y(_03124_));
 AND2x2_ASAP7_75t_R _25559_ (.A(_14977_),
    .B(_09909_),
    .Y(_09916_));
 AO21x1_ASAP7_75t_R _25560_ (.A1(_09731_),
    .A2(_09904_),
    .B(_09916_),
    .Y(_03125_));
 BUFx6f_ASAP7_75t_R _25561_ (.A(_09869_),
    .Y(_09917_));
 BUFx12f_ASAP7_75t_R _25562_ (.A(_09869_),
    .Y(_09918_));
 NAND2x1_ASAP7_75t_R _25563_ (.A(_01793_),
    .B(_09918_),
    .Y(_09919_));
 OA21x2_ASAP7_75t_R _25564_ (.A1(_09629_),
    .A2(_09917_),
    .B(_09919_),
    .Y(_03126_));
 AND2x2_ASAP7_75t_R _25565_ (.A(_15053_),
    .B(_09909_),
    .Y(_09920_));
 AO21x1_ASAP7_75t_R _25566_ (.A1(_09572_),
    .A2(_09904_),
    .B(_09920_),
    .Y(_03127_));
 AND2x2_ASAP7_75t_R _25567_ (.A(_15109_),
    .B(_09909_),
    .Y(_09921_));
 AO21x1_ASAP7_75t_R _25568_ (.A1(_09784_),
    .A2(_09904_),
    .B(_09921_),
    .Y(_03128_));
 AND2x2_ASAP7_75t_R _25569_ (.A(_15183_),
    .B(_09909_),
    .Y(_09922_));
 AO21x1_ASAP7_75t_R _25570_ (.A1(_09575_),
    .A2(_09904_),
    .B(_09922_),
    .Y(_03129_));
 BUFx12f_ASAP7_75t_R _25571_ (.A(_09903_),
    .Y(_09923_));
 AND2x2_ASAP7_75t_R _25572_ (.A(_14240_),
    .B(_09909_),
    .Y(_09924_));
 AO21x1_ASAP7_75t_R _25573_ (.A1(_09736_),
    .A2(_09923_),
    .B(_09924_),
    .Y(_03130_));
 BUFx6f_ASAP7_75t_R _25574_ (.A(_09905_),
    .Y(_09925_));
 AND2x2_ASAP7_75t_R _25575_ (.A(_13108_),
    .B(_09925_),
    .Y(_09926_));
 AO21x1_ASAP7_75t_R _25576_ (.A1(_09579_),
    .A2(_09923_),
    .B(_09926_),
    .Y(_03131_));
 AND2x2_ASAP7_75t_R _25577_ (.A(_15375_),
    .B(_09925_),
    .Y(_09927_));
 AO21x1_ASAP7_75t_R _25578_ (.A1(_09690_),
    .A2(_09923_),
    .B(_09927_),
    .Y(_03132_));
 NOR2x1_ASAP7_75t_R _25579_ (.A(_08851_),
    .B(_09906_),
    .Y(_09928_));
 AO21x1_ASAP7_75t_R _25580_ (.A1(_15528_),
    .A2(_09906_),
    .B(_09928_),
    .Y(_03133_));
 AO21x1_ASAP7_75t_R _25581_ (.A1(_08954_),
    .A2(_09812_),
    .B(_15651_),
    .Y(_09929_));
 OA21x2_ASAP7_75t_R _25582_ (.A1(_09453_),
    .A2(_09906_),
    .B(_09929_),
    .Y(_03134_));
 BUFx6f_ASAP7_75t_R _25583_ (.A(_08920_),
    .Y(_09930_));
 AND2x2_ASAP7_75t_R _25584_ (.A(_09930_),
    .B(_09903_),
    .Y(_09931_));
 AO21x1_ASAP7_75t_R _25585_ (.A1(_15807_),
    .A2(_09906_),
    .B(_09931_),
    .Y(_03135_));
 NOR2x1_ASAP7_75t_R _25586_ (.A(_09695_),
    .B(_09906_),
    .Y(_09932_));
 AO21x1_ASAP7_75t_R _25587_ (.A1(_15889_),
    .A2(_09906_),
    .B(_09932_),
    .Y(_03136_));
 NAND2x1_ASAP7_75t_R _25588_ (.A(_01792_),
    .B(_09918_),
    .Y(_09933_));
 OA21x2_ASAP7_75t_R _25589_ (.A1(_09563_),
    .A2(_09917_),
    .B(_09933_),
    .Y(_03137_));
 AND2x2_ASAP7_75t_R _25590_ (.A(_16054_),
    .B(_09925_),
    .Y(_09934_));
 AO21x1_ASAP7_75t_R _25591_ (.A1(_09697_),
    .A2(_09923_),
    .B(_09934_),
    .Y(_03138_));
 AND2x2_ASAP7_75t_R _25592_ (.A(_16136_),
    .B(_09925_),
    .Y(_09935_));
 AO21x1_ASAP7_75t_R _25593_ (.A1(_09699_),
    .A2(_09923_),
    .B(_09935_),
    .Y(_03139_));
 AND2x2_ASAP7_75t_R _25594_ (.A(_16271_),
    .B(_09925_),
    .Y(_09936_));
 AO21x1_ASAP7_75t_R _25595_ (.A1(_09701_),
    .A2(_09923_),
    .B(_09936_),
    .Y(_03140_));
 AND2x2_ASAP7_75t_R _25596_ (.A(_16394_),
    .B(_09925_),
    .Y(_09937_));
 AO21x1_ASAP7_75t_R _25597_ (.A1(_09749_),
    .A2(_09923_),
    .B(_09937_),
    .Y(_03141_));
 AND2x2_ASAP7_75t_R _25598_ (.A(_16532_),
    .B(_09925_),
    .Y(_09938_));
 AO21x1_ASAP7_75t_R _25599_ (.A1(_09751_),
    .A2(_09923_),
    .B(_09938_),
    .Y(_03142_));
 AND2x2_ASAP7_75t_R _25600_ (.A(_16642_),
    .B(_09925_),
    .Y(_09939_));
 AO21x1_ASAP7_75t_R _25601_ (.A1(_09753_),
    .A2(_09923_),
    .B(_09939_),
    .Y(_03143_));
 AND2x2_ASAP7_75t_R _25602_ (.A(_16765_),
    .B(_09925_),
    .Y(_09940_));
 AO21x1_ASAP7_75t_R _25603_ (.A1(_09706_),
    .A2(_09923_),
    .B(_09940_),
    .Y(_03144_));
 AND2x2_ASAP7_75t_R _25604_ (.A(_16907_),
    .B(_09925_),
    .Y(_09941_));
 AO21x1_ASAP7_75t_R _25605_ (.A1(_09708_),
    .A2(_09903_),
    .B(_09941_),
    .Y(_03145_));
 AND2x2_ASAP7_75t_R _25606_ (.A(_04250_),
    .B(_09905_),
    .Y(_09942_));
 AO21x1_ASAP7_75t_R _25607_ (.A1(_09757_),
    .A2(_09903_),
    .B(_09942_),
    .Y(_03146_));
 AND2x2_ASAP7_75t_R _25608_ (.A(_04363_),
    .B(_09905_),
    .Y(_09943_));
 AO21x1_ASAP7_75t_R _25609_ (.A1(_09759_),
    .A2(_09903_),
    .B(_09943_),
    .Y(_03147_));
 NAND2x1_ASAP7_75t_R _25610_ (.A(_01791_),
    .B(_09918_),
    .Y(_09944_));
 OA21x2_ASAP7_75t_R _25611_ (.A1(_09565_),
    .A2(_09917_),
    .B(_09944_),
    .Y(_03148_));
 AND2x2_ASAP7_75t_R _25612_ (.A(_04530_),
    .B(_09905_),
    .Y(_09945_));
 AO21x1_ASAP7_75t_R _25613_ (.A1(_09761_),
    .A2(_09903_),
    .B(_09945_),
    .Y(_03149_));
 AND2x2_ASAP7_75t_R _25614_ (.A(_04611_),
    .B(_09905_),
    .Y(_09946_));
 AO21x1_ASAP7_75t_R _25615_ (.A1(_09713_),
    .A2(_09903_),
    .B(_09946_),
    .Y(_03150_));
 AO21x1_ASAP7_75t_R _25616_ (.A1(_08954_),
    .A2(_09812_),
    .B(_04733_),
    .Y(_09947_));
 OA21x2_ASAP7_75t_R _25617_ (.A1(_09612_),
    .A2(_09906_),
    .B(_09947_),
    .Y(_03151_));
 AND2x2_ASAP7_75t_R _25618_ (.A(_04917_),
    .B(_09905_),
    .Y(_09948_));
 AO21x1_ASAP7_75t_R _25619_ (.A1(_09810_),
    .A2(_09903_),
    .B(_09948_),
    .Y(_03152_));
 NOR2x1_ASAP7_75t_R _25620_ (.A(_13685_),
    .B(_13602_),
    .Y(_09949_));
 AND5x2_ASAP7_75t_R _25621_ (.A(_07799_),
    .B(_13455_),
    .C(_13430_),
    .D(_09949_),
    .E(_09475_),
    .Y(_09950_));
 BUFx12f_ASAP7_75t_R _25622_ (.A(_09950_),
    .Y(_09951_));
 OR4x1_ASAP7_75t_R _25623_ (.A(_13692_),
    .B(_09504_),
    .C(_08254_),
    .D(_09505_),
    .Y(_09952_));
 BUFx12f_ASAP7_75t_R _25624_ (.A(_09952_),
    .Y(_09953_));
 BUFx12f_ASAP7_75t_R _25625_ (.A(_09953_),
    .Y(_09954_));
 AND2x2_ASAP7_75t_R _25626_ (.A(_00391_),
    .B(_09954_),
    .Y(_09955_));
 AOI21x1_ASAP7_75t_R _25627_ (.A1(_09902_),
    .A2(_09951_),
    .B(_09955_),
    .Y(_03153_));
 AND2x2_ASAP7_75t_R _25628_ (.A(_00424_),
    .B(_09954_),
    .Y(_09956_));
 AOI21x1_ASAP7_75t_R _25629_ (.A1(_09908_),
    .A2(_09951_),
    .B(_09956_),
    .Y(_03154_));
 NOR2x1_ASAP7_75t_R _25630_ (.A(_09898_),
    .B(_09954_),
    .Y(_09957_));
 AO21x1_ASAP7_75t_R _25631_ (.A1(_13545_),
    .A2(_09954_),
    .B(_09957_),
    .Y(_03155_));
 AND2x2_ASAP7_75t_R _25632_ (.A(_13633_),
    .B(_09953_),
    .Y(_09958_));
 AO21x1_ASAP7_75t_R _25633_ (.A1(_09819_),
    .A2(_09951_),
    .B(_09958_),
    .Y(_03156_));
 AND2x2_ASAP7_75t_R _25634_ (.A(_13699_),
    .B(_09953_),
    .Y(_09959_));
 AO21x1_ASAP7_75t_R _25635_ (.A1(_09726_),
    .A2(_09951_),
    .B(_09959_),
    .Y(_03157_));
 AND2x2_ASAP7_75t_R _25636_ (.A(_13825_),
    .B(_09953_),
    .Y(_09960_));
 AO21x1_ASAP7_75t_R _25637_ (.A1(_09679_),
    .A2(_09951_),
    .B(_09960_),
    .Y(_03158_));
 NAND2x1_ASAP7_75t_R _25638_ (.A(_01790_),
    .B(_09918_),
    .Y(_09961_));
 OA21x2_ASAP7_75t_R _25639_ (.A1(_09567_),
    .A2(_09917_),
    .B(_09961_),
    .Y(_03159_));
 AND2x2_ASAP7_75t_R _25640_ (.A(_13845_),
    .B(_09953_),
    .Y(_09962_));
 AO21x1_ASAP7_75t_R _25641_ (.A1(_09729_),
    .A2(_09951_),
    .B(_09962_),
    .Y(_03160_));
 AND2x2_ASAP7_75t_R _25642_ (.A(_13914_),
    .B(_09953_),
    .Y(_09963_));
 AO21x1_ASAP7_75t_R _25643_ (.A1(_09731_),
    .A2(_09951_),
    .B(_09963_),
    .Y(_03161_));
 AND2x2_ASAP7_75t_R _25644_ (.A(_14006_),
    .B(_09953_),
    .Y(_09964_));
 AO21x1_ASAP7_75t_R _25645_ (.A1(_09572_),
    .A2(_09951_),
    .B(_09964_),
    .Y(_03162_));
 BUFx12f_ASAP7_75t_R _25646_ (.A(_09950_),
    .Y(_09965_));
 NOR2x1_ASAP7_75t_R _25647_ (.A(_00665_),
    .B(_09965_),
    .Y(_09966_));
 AO21x1_ASAP7_75t_R _25648_ (.A1(_09784_),
    .A2(_09951_),
    .B(_09966_),
    .Y(_03163_));
 BUFx12f_ASAP7_75t_R _25649_ (.A(_09950_),
    .Y(_09967_));
 AND2x2_ASAP7_75t_R _25650_ (.A(_14170_),
    .B(_09953_),
    .Y(_09968_));
 AO21x1_ASAP7_75t_R _25651_ (.A1(_09575_),
    .A2(_09967_),
    .B(_09968_),
    .Y(_03164_));
 AND2x2_ASAP7_75t_R _25652_ (.A(_14233_),
    .B(_09953_),
    .Y(_09969_));
 AO21x1_ASAP7_75t_R _25653_ (.A1(_09736_),
    .A2(_09967_),
    .B(_09969_),
    .Y(_03165_));
 NOR2x1_ASAP7_75t_R _25654_ (.A(_00355_),
    .B(_09965_),
    .Y(_09970_));
 AO21x1_ASAP7_75t_R _25655_ (.A1(_09579_),
    .A2(_09967_),
    .B(_09970_),
    .Y(_03166_));
 BUFx12f_ASAP7_75t_R _25656_ (.A(_09950_),
    .Y(_09971_));
 NOR2x1_ASAP7_75t_R _25657_ (.A(_00793_),
    .B(_09971_),
    .Y(_09972_));
 AO21x1_ASAP7_75t_R _25658_ (.A1(_09690_),
    .A2(_09967_),
    .B(_09972_),
    .Y(_03167_));
 AND2x2_ASAP7_75t_R _25659_ (.A(_00825_),
    .B(_09954_),
    .Y(_09973_));
 AOI21x1_ASAP7_75t_R _25660_ (.A1(_09790_),
    .A2(_09951_),
    .B(_09973_),
    .Y(_03168_));
 NAND2x1_ASAP7_75t_R _25661_ (.A(_00857_),
    .B(_09954_),
    .Y(_09974_));
 OA21x2_ASAP7_75t_R _25662_ (.A1(_09453_),
    .A2(_09954_),
    .B(_09974_),
    .Y(_03169_));
 NAND2x1_ASAP7_75t_R _25663_ (.A(_01789_),
    .B(_09918_),
    .Y(_09975_));
 OA21x2_ASAP7_75t_R _25664_ (.A1(_09570_),
    .A2(_09917_),
    .B(_09975_),
    .Y(_03170_));
 NOR2x1_ASAP7_75t_R _25665_ (.A(_00889_),
    .B(_09971_),
    .Y(_09976_));
 AO21x1_ASAP7_75t_R _25666_ (.A1(_09584_),
    .A2(_09967_),
    .B(_09976_),
    .Y(_03171_));
 AND2x2_ASAP7_75t_R _25667_ (.A(_09457_),
    .B(_09950_),
    .Y(_09977_));
 AOI21x1_ASAP7_75t_R _25668_ (.A1(_00921_),
    .A2(_09954_),
    .B(_09977_),
    .Y(_03172_));
 NOR2x1_ASAP7_75t_R _25669_ (.A(_00953_),
    .B(_09971_),
    .Y(_09978_));
 AO21x1_ASAP7_75t_R _25670_ (.A1(_09697_),
    .A2(_09967_),
    .B(_09978_),
    .Y(_03173_));
 NOR2x1_ASAP7_75t_R _25671_ (.A(_00985_),
    .B(_09971_),
    .Y(_09979_));
 AO21x1_ASAP7_75t_R _25672_ (.A1(_09699_),
    .A2(_09967_),
    .B(_09979_),
    .Y(_03174_));
 NOR2x1_ASAP7_75t_R _25673_ (.A(_01017_),
    .B(_09971_),
    .Y(_09980_));
 AO21x1_ASAP7_75t_R _25674_ (.A1(_09701_),
    .A2(_09967_),
    .B(_09980_),
    .Y(_03175_));
 NOR2x1_ASAP7_75t_R _25675_ (.A(_01049_),
    .B(_09971_),
    .Y(_09981_));
 AO21x1_ASAP7_75t_R _25676_ (.A1(_09749_),
    .A2(_09967_),
    .B(_09981_),
    .Y(_03176_));
 NOR2x1_ASAP7_75t_R _25677_ (.A(_01081_),
    .B(_09971_),
    .Y(_09982_));
 AO21x1_ASAP7_75t_R _25678_ (.A1(_09751_),
    .A2(_09967_),
    .B(_09982_),
    .Y(_03177_));
 NOR2x1_ASAP7_75t_R _25679_ (.A(_01113_),
    .B(_09971_),
    .Y(_09983_));
 AO21x1_ASAP7_75t_R _25680_ (.A1(_09753_),
    .A2(_09965_),
    .B(_09983_),
    .Y(_03178_));
 NOR2x1_ASAP7_75t_R _25681_ (.A(_01145_),
    .B(_09971_),
    .Y(_09984_));
 AO21x1_ASAP7_75t_R _25682_ (.A1(_09706_),
    .A2(_09965_),
    .B(_09984_),
    .Y(_03179_));
 NOR2x1_ASAP7_75t_R _25683_ (.A(_01177_),
    .B(_09971_),
    .Y(_09985_));
 AO21x1_ASAP7_75t_R _25684_ (.A1(_09708_),
    .A2(_09965_),
    .B(_09985_),
    .Y(_03180_));
 NAND2x1_ASAP7_75t_R _25685_ (.A(_01788_),
    .B(_09918_),
    .Y(_09986_));
 OA21x2_ASAP7_75t_R _25686_ (.A1(_09438_),
    .A2(_09917_),
    .B(_09986_),
    .Y(_03181_));
 NOR2x1_ASAP7_75t_R _25687_ (.A(_01209_),
    .B(_09950_),
    .Y(_09987_));
 AO21x1_ASAP7_75t_R _25688_ (.A1(_09757_),
    .A2(_09965_),
    .B(_09987_),
    .Y(_03182_));
 NOR2x1_ASAP7_75t_R _25689_ (.A(_01241_),
    .B(_09950_),
    .Y(_09988_));
 AO21x1_ASAP7_75t_R _25690_ (.A1(_09759_),
    .A2(_09965_),
    .B(_09988_),
    .Y(_03183_));
 NOR2x1_ASAP7_75t_R _25691_ (.A(_01273_),
    .B(_09950_),
    .Y(_09989_));
 AO21x1_ASAP7_75t_R _25692_ (.A1(_09761_),
    .A2(_09965_),
    .B(_09989_),
    .Y(_03184_));
 NOR2x1_ASAP7_75t_R _25693_ (.A(_01305_),
    .B(_09950_),
    .Y(_09990_));
 AO21x1_ASAP7_75t_R _25694_ (.A1(_09713_),
    .A2(_09965_),
    .B(_09990_),
    .Y(_03185_));
 NAND2x1_ASAP7_75t_R _25695_ (.A(_01337_),
    .B(_09954_),
    .Y(_09991_));
 OA21x2_ASAP7_75t_R _25696_ (.A1(_09612_),
    .A2(_09954_),
    .B(_09991_),
    .Y(_03186_));
 AND2x2_ASAP7_75t_R _25697_ (.A(_04871_),
    .B(_09953_),
    .Y(_09992_));
 AO21x1_ASAP7_75t_R _25698_ (.A1(_09810_),
    .A2(_09965_),
    .B(_09992_),
    .Y(_03187_));
 BUFx12f_ASAP7_75t_R _25699_ (.A(_09949_),
    .Y(_09993_));
 AND2x6_ASAP7_75t_R _25700_ (.A(_09993_),
    .B(_09620_),
    .Y(_09994_));
 BUFx12f_ASAP7_75t_R _25701_ (.A(_09994_),
    .Y(_09995_));
 BUFx6f_ASAP7_75t_R _25702_ (.A(_09995_),
    .Y(_09996_));
 NAND2x2_ASAP7_75t_R _25703_ (.A(_09993_),
    .B(_09621_),
    .Y(_09997_));
 BUFx12f_ASAP7_75t_R _25704_ (.A(_09997_),
    .Y(_09998_));
 AND2x2_ASAP7_75t_R _25705_ (.A(_00392_),
    .B(_09998_),
    .Y(_09999_));
 AOI21x1_ASAP7_75t_R _25706_ (.A1(_09902_),
    .A2(_09996_),
    .B(_09999_),
    .Y(_03188_));
 AND2x2_ASAP7_75t_R _25707_ (.A(_00425_),
    .B(_09998_),
    .Y(_10000_));
 AOI21x1_ASAP7_75t_R _25708_ (.A1(_09908_),
    .A2(_09996_),
    .B(_10000_),
    .Y(_03189_));
 NOR2x1_ASAP7_75t_R _25709_ (.A(_09898_),
    .B(_09998_),
    .Y(_10001_));
 AO21x1_ASAP7_75t_R _25710_ (.A1(_13564_),
    .A2(_09998_),
    .B(_10001_),
    .Y(_03190_));
 BUFx12f_ASAP7_75t_R _25711_ (.A(_09994_),
    .Y(_10002_));
 NOR2x1_ASAP7_75t_R _25712_ (.A(_00486_),
    .B(_10002_),
    .Y(_10003_));
 AO21x1_ASAP7_75t_R _25713_ (.A1(_09819_),
    .A2(_09996_),
    .B(_10003_),
    .Y(_03191_));
 NAND2x1_ASAP7_75t_R _25714_ (.A(_01787_),
    .B(_09918_),
    .Y(_10004_));
 OA21x2_ASAP7_75t_R _25715_ (.A1(_09441_),
    .A2(_09917_),
    .B(_10004_),
    .Y(_03192_));
 AND2x2_ASAP7_75t_R _25716_ (.A(_13713_),
    .B(_09997_),
    .Y(_10005_));
 AO21x1_ASAP7_75t_R _25717_ (.A1(_09726_),
    .A2(_09996_),
    .B(_10005_),
    .Y(_03193_));
 AND2x2_ASAP7_75t_R _25718_ (.A(_13800_),
    .B(_09997_),
    .Y(_10006_));
 AO21x1_ASAP7_75t_R _25719_ (.A1(_09679_),
    .A2(_09996_),
    .B(_10006_),
    .Y(_03194_));
 AND2x2_ASAP7_75t_R _25720_ (.A(_13870_),
    .B(_09997_),
    .Y(_10007_));
 AO21x1_ASAP7_75t_R _25721_ (.A1(_09729_),
    .A2(_09996_),
    .B(_10007_),
    .Y(_03195_));
 NOR2x1_ASAP7_75t_R _25722_ (.A(_00606_),
    .B(_10002_),
    .Y(_10008_));
 AO21x1_ASAP7_75t_R _25723_ (.A1(_09731_),
    .A2(_09996_),
    .B(_10008_),
    .Y(_03196_));
 AND2x2_ASAP7_75t_R _25724_ (.A(_13999_),
    .B(_09997_),
    .Y(_10009_));
 AO21x1_ASAP7_75t_R _25725_ (.A1(_09572_),
    .A2(_09996_),
    .B(_10009_),
    .Y(_03197_));
 NOR2x1_ASAP7_75t_R _25726_ (.A(_00666_),
    .B(_10002_),
    .Y(_10010_));
 AO21x1_ASAP7_75t_R _25727_ (.A1(_09784_),
    .A2(_09996_),
    .B(_10010_),
    .Y(_03198_));
 AND2x2_ASAP7_75t_R _25728_ (.A(_14184_),
    .B(_09997_),
    .Y(_10011_));
 AO21x1_ASAP7_75t_R _25729_ (.A1(_09575_),
    .A2(_09996_),
    .B(_10011_),
    .Y(_03199_));
 BUFx12f_ASAP7_75t_R _25730_ (.A(_09995_),
    .Y(_10012_));
 BUFx12f_ASAP7_75t_R _25731_ (.A(_09994_),
    .Y(_10013_));
 NOR2x1_ASAP7_75t_R _25732_ (.A(_00726_),
    .B(_10013_),
    .Y(_10014_));
 AO21x1_ASAP7_75t_R _25733_ (.A1(_09736_),
    .A2(_10012_),
    .B(_10014_),
    .Y(_03200_));
 NOR2x1_ASAP7_75t_R _25734_ (.A(_00356_),
    .B(_10013_),
    .Y(_10015_));
 AO21x1_ASAP7_75t_R _25735_ (.A1(_09579_),
    .A2(_10012_),
    .B(_10015_),
    .Y(_03201_));
 NOR2x1_ASAP7_75t_R _25736_ (.A(_00794_),
    .B(_10013_),
    .Y(_10016_));
 AO21x1_ASAP7_75t_R _25737_ (.A1(_09690_),
    .A2(_10012_),
    .B(_10016_),
    .Y(_03202_));
 NAND2x1_ASAP7_75t_R _25738_ (.A(_01786_),
    .B(_09918_),
    .Y(_10017_));
 OA21x2_ASAP7_75t_R _25739_ (.A1(_09443_),
    .A2(_09917_),
    .B(_10017_),
    .Y(_03203_));
 AND2x2_ASAP7_75t_R _25740_ (.A(_09451_),
    .B(_09995_),
    .Y(_10018_));
 AOI21x1_ASAP7_75t_R _25741_ (.A1(_00826_),
    .A2(_09998_),
    .B(_10018_),
    .Y(_03204_));
 BUFx6f_ASAP7_75t_R _25742_ (.A(_08892_),
    .Y(_10019_));
 NAND2x1_ASAP7_75t_R _25743_ (.A(_00858_),
    .B(_09998_),
    .Y(_10020_));
 OA21x2_ASAP7_75t_R _25744_ (.A1(_10019_),
    .A2(_09998_),
    .B(_10020_),
    .Y(_03205_));
 NOR2x1_ASAP7_75t_R _25745_ (.A(_00890_),
    .B(_10013_),
    .Y(_10021_));
 AO21x1_ASAP7_75t_R _25746_ (.A1(_09584_),
    .A2(_10012_),
    .B(_10021_),
    .Y(_03206_));
 AND2x2_ASAP7_75t_R _25747_ (.A(_09457_),
    .B(_09995_),
    .Y(_10022_));
 AOI21x1_ASAP7_75t_R _25748_ (.A1(_00922_),
    .A2(_09998_),
    .B(_10022_),
    .Y(_03207_));
 NOR2x1_ASAP7_75t_R _25749_ (.A(_00954_),
    .B(_10013_),
    .Y(_10023_));
 AO21x1_ASAP7_75t_R _25750_ (.A1(_09697_),
    .A2(_10012_),
    .B(_10023_),
    .Y(_03208_));
 NOR2x1_ASAP7_75t_R _25751_ (.A(_00986_),
    .B(_10013_),
    .Y(_10024_));
 AO21x1_ASAP7_75t_R _25752_ (.A1(_09699_),
    .A2(_10012_),
    .B(_10024_),
    .Y(_03209_));
 NOR2x1_ASAP7_75t_R _25753_ (.A(_01018_),
    .B(_10013_),
    .Y(_10025_));
 AO21x1_ASAP7_75t_R _25754_ (.A1(_09701_),
    .A2(_10012_),
    .B(_10025_),
    .Y(_03210_));
 NOR2x1_ASAP7_75t_R _25755_ (.A(_01050_),
    .B(_10013_),
    .Y(_10026_));
 AO21x1_ASAP7_75t_R _25756_ (.A1(_09749_),
    .A2(_10012_),
    .B(_10026_),
    .Y(_03211_));
 NOR2x1_ASAP7_75t_R _25757_ (.A(_01082_),
    .B(_10013_),
    .Y(_10027_));
 AO21x1_ASAP7_75t_R _25758_ (.A1(_09751_),
    .A2(_10012_),
    .B(_10027_),
    .Y(_03212_));
 NOR2x1_ASAP7_75t_R _25759_ (.A(_01114_),
    .B(_10013_),
    .Y(_10028_));
 AO21x1_ASAP7_75t_R _25760_ (.A1(_09753_),
    .A2(_10012_),
    .B(_10028_),
    .Y(_03213_));
 BUFx6f_ASAP7_75t_R _25761_ (.A(_09869_),
    .Y(_10029_));
 NAND2x1_ASAP7_75t_R _25762_ (.A(_01785_),
    .B(_09918_),
    .Y(_10030_));
 OA21x2_ASAP7_75t_R _25763_ (.A1(_09445_),
    .A2(_10029_),
    .B(_10030_),
    .Y(_03214_));
 NOR2x1_ASAP7_75t_R _25764_ (.A(_01146_),
    .B(_09995_),
    .Y(_10031_));
 AO21x1_ASAP7_75t_R _25765_ (.A1(_09706_),
    .A2(_10002_),
    .B(_10031_),
    .Y(_03215_));
 NOR2x1_ASAP7_75t_R _25766_ (.A(_01178_),
    .B(_09995_),
    .Y(_10032_));
 AO21x1_ASAP7_75t_R _25767_ (.A1(_09708_),
    .A2(_10002_),
    .B(_10032_),
    .Y(_03216_));
 NOR2x1_ASAP7_75t_R _25768_ (.A(_01210_),
    .B(_09995_),
    .Y(_10033_));
 AO21x1_ASAP7_75t_R _25769_ (.A1(_09757_),
    .A2(_10002_),
    .B(_10033_),
    .Y(_03217_));
 NOR2x1_ASAP7_75t_R _25770_ (.A(_01242_),
    .B(_09995_),
    .Y(_10034_));
 AO21x1_ASAP7_75t_R _25771_ (.A1(_09759_),
    .A2(_10002_),
    .B(_10034_),
    .Y(_03218_));
 NOR2x1_ASAP7_75t_R _25772_ (.A(_01274_),
    .B(_09995_),
    .Y(_10035_));
 AO21x1_ASAP7_75t_R _25773_ (.A1(_09761_),
    .A2(_10002_),
    .B(_10035_),
    .Y(_03219_));
 NOR2x1_ASAP7_75t_R _25774_ (.A(_01306_),
    .B(_09995_),
    .Y(_10036_));
 AO21x1_ASAP7_75t_R _25775_ (.A1(_09713_),
    .A2(_10002_),
    .B(_10036_),
    .Y(_03220_));
 NAND2x1_ASAP7_75t_R _25776_ (.A(_01338_),
    .B(_09998_),
    .Y(_10037_));
 OA21x2_ASAP7_75t_R _25777_ (.A1(_09612_),
    .A2(_09998_),
    .B(_10037_),
    .Y(_03221_));
 AND2x2_ASAP7_75t_R _25778_ (.A(_04874_),
    .B(_09997_),
    .Y(_10038_));
 AO21x1_ASAP7_75t_R _25779_ (.A1(_09810_),
    .A2(_10002_),
    .B(_10038_),
    .Y(_03222_));
 AND2x6_ASAP7_75t_R _25780_ (.A(_09993_),
    .B(_09666_),
    .Y(_10039_));
 BUFx12f_ASAP7_75t_R _25781_ (.A(_10039_),
    .Y(_10040_));
 NAND2x2_ASAP7_75t_R _25782_ (.A(_09993_),
    .B(_09666_),
    .Y(_10041_));
 BUFx12f_ASAP7_75t_R _25783_ (.A(_10041_),
    .Y(_10042_));
 AND2x2_ASAP7_75t_R _25784_ (.A(_00393_),
    .B(_10042_),
    .Y(_10043_));
 AOI21x1_ASAP7_75t_R _25785_ (.A1(_09902_),
    .A2(_10040_),
    .B(_10043_),
    .Y(_03223_));
 AND2x2_ASAP7_75t_R _25786_ (.A(_00426_),
    .B(_10042_),
    .Y(_10044_));
 AOI21x1_ASAP7_75t_R _25787_ (.A1(_09908_),
    .A2(_10040_),
    .B(_10044_),
    .Y(_03224_));
 NAND2x1_ASAP7_75t_R _25788_ (.A(_01784_),
    .B(_09918_),
    .Y(_10045_));
 OA21x2_ASAP7_75t_R _25789_ (.A1(_09447_),
    .A2(_10029_),
    .B(_10045_),
    .Y(_03225_));
 NOR2x1_ASAP7_75t_R _25790_ (.A(_09898_),
    .B(_10042_),
    .Y(_10046_));
 AO21x1_ASAP7_75t_R _25791_ (.A1(_13548_),
    .A2(_10042_),
    .B(_10046_),
    .Y(_03226_));
 BUFx12f_ASAP7_75t_R _25792_ (.A(_10039_),
    .Y(_10047_));
 NOR2x1_ASAP7_75t_R _25793_ (.A(_00487_),
    .B(_10047_),
    .Y(_10048_));
 AO21x1_ASAP7_75t_R _25794_ (.A1(_09819_),
    .A2(_10040_),
    .B(_10048_),
    .Y(_03227_));
 AND2x2_ASAP7_75t_R _25795_ (.A(_13703_),
    .B(_10042_),
    .Y(_10049_));
 AO21x1_ASAP7_75t_R _25796_ (.A1(_09726_),
    .A2(_10040_),
    .B(_10049_),
    .Y(_03228_));
 BUFx12f_ASAP7_75t_R _25797_ (.A(_10041_),
    .Y(_10050_));
 AND2x2_ASAP7_75t_R _25798_ (.A(_13822_),
    .B(_10050_),
    .Y(_10051_));
 AO21x1_ASAP7_75t_R _25799_ (.A1(_09679_),
    .A2(_10040_),
    .B(_10051_),
    .Y(_03229_));
 AND2x2_ASAP7_75t_R _25800_ (.A(_13841_),
    .B(_10050_),
    .Y(_10052_));
 AO21x1_ASAP7_75t_R _25801_ (.A1(_09729_),
    .A2(_10040_),
    .B(_10052_),
    .Y(_03230_));
 AND2x2_ASAP7_75t_R _25802_ (.A(_13911_),
    .B(_10050_),
    .Y(_10053_));
 AO21x1_ASAP7_75t_R _25803_ (.A1(_09731_),
    .A2(_10040_),
    .B(_10053_),
    .Y(_03231_));
 AND2x2_ASAP7_75t_R _25804_ (.A(_14003_),
    .B(_10050_),
    .Y(_10054_));
 AO21x1_ASAP7_75t_R _25805_ (.A1(_09572_),
    .A2(_10040_),
    .B(_10054_),
    .Y(_03232_));
 AND2x2_ASAP7_75t_R _25806_ (.A(_14060_),
    .B(_10050_),
    .Y(_10055_));
 AO21x1_ASAP7_75t_R _25807_ (.A1(_09784_),
    .A2(_10040_),
    .B(_10055_),
    .Y(_03233_));
 BUFx12f_ASAP7_75t_R _25808_ (.A(_10039_),
    .Y(_10056_));
 AND2x2_ASAP7_75t_R _25809_ (.A(_14167_),
    .B(_10050_),
    .Y(_10057_));
 AO21x1_ASAP7_75t_R _25810_ (.A1(_09575_),
    .A2(_10056_),
    .B(_10057_),
    .Y(_03234_));
 AND2x2_ASAP7_75t_R _25811_ (.A(_14332_),
    .B(_10050_),
    .Y(_10058_));
 AO21x1_ASAP7_75t_R _25812_ (.A1(_09736_),
    .A2(_10056_),
    .B(_10058_),
    .Y(_03235_));
 BUFx12f_ASAP7_75t_R _25813_ (.A(_09869_),
    .Y(_10059_));
 NAND2x1_ASAP7_75t_R _25814_ (.A(_01783_),
    .B(_10059_),
    .Y(_10060_));
 OA21x2_ASAP7_75t_R _25815_ (.A1(_09449_),
    .A2(_10029_),
    .B(_10060_),
    .Y(_03236_));
 AND2x2_ASAP7_75t_R _25816_ (.A(_13157_),
    .B(_10050_),
    .Y(_10061_));
 AO21x1_ASAP7_75t_R _25817_ (.A1(_09579_),
    .A2(_10056_),
    .B(_10061_),
    .Y(_03237_));
 AND2x2_ASAP7_75t_R _25818_ (.A(_15393_),
    .B(_10050_),
    .Y(_10062_));
 AO21x1_ASAP7_75t_R _25819_ (.A1(_09690_),
    .A2(_10056_),
    .B(_10062_),
    .Y(_03238_));
 NAND2x1_ASAP7_75t_R _25820_ (.A(_08851_),
    .B(_10047_),
    .Y(_10063_));
 OA21x2_ASAP7_75t_R _25821_ (.A1(_15546_),
    .A2(_10040_),
    .B(_10063_),
    .Y(_03239_));
 AO21x1_ASAP7_75t_R _25822_ (.A1(_09993_),
    .A2(_09667_),
    .B(_15669_),
    .Y(_10064_));
 OA21x2_ASAP7_75t_R _25823_ (.A1(_10019_),
    .A2(_10042_),
    .B(_10064_),
    .Y(_03240_));
 AND2x2_ASAP7_75t_R _25824_ (.A(_09930_),
    .B(_10047_),
    .Y(_10065_));
 AO21x1_ASAP7_75t_R _25825_ (.A1(_15825_),
    .A2(_10042_),
    .B(_10065_),
    .Y(_03241_));
 NOR2x1_ASAP7_75t_R _25826_ (.A(_09695_),
    .B(_10042_),
    .Y(_10066_));
 AO21x1_ASAP7_75t_R _25827_ (.A1(_15907_),
    .A2(_10042_),
    .B(_10066_),
    .Y(_03242_));
 AND2x2_ASAP7_75t_R _25828_ (.A(_16072_),
    .B(_10050_),
    .Y(_10067_));
 AO21x1_ASAP7_75t_R _25829_ (.A1(_09697_),
    .A2(_10056_),
    .B(_10067_),
    .Y(_03243_));
 BUFx6f_ASAP7_75t_R _25830_ (.A(_10041_),
    .Y(_10068_));
 AND2x2_ASAP7_75t_R _25831_ (.A(_16154_),
    .B(_10068_),
    .Y(_10069_));
 AO21x1_ASAP7_75t_R _25832_ (.A1(_09699_),
    .A2(_10056_),
    .B(_10069_),
    .Y(_03244_));
 AND2x2_ASAP7_75t_R _25833_ (.A(_16289_),
    .B(_10068_),
    .Y(_10070_));
 AO21x1_ASAP7_75t_R _25834_ (.A1(_09701_),
    .A2(_10056_),
    .B(_10070_),
    .Y(_03245_));
 AND2x2_ASAP7_75t_R _25835_ (.A(_16412_),
    .B(_10068_),
    .Y(_10071_));
 AO21x1_ASAP7_75t_R _25836_ (.A1(_09749_),
    .A2(_10056_),
    .B(_10071_),
    .Y(_03246_));
 AO21x1_ASAP7_75t_R _25837_ (.A1(_08950_),
    .A2(_09621_),
    .B(_01782_),
    .Y(_10072_));
 OAI21x1_ASAP7_75t_R _25838_ (.A1(_09790_),
    .A2(_09917_),
    .B(_10072_),
    .Y(_03247_));
 AND2x2_ASAP7_75t_R _25839_ (.A(_16550_),
    .B(_10068_),
    .Y(_10073_));
 AO21x1_ASAP7_75t_R _25840_ (.A1(_09751_),
    .A2(_10056_),
    .B(_10073_),
    .Y(_03248_));
 AND2x2_ASAP7_75t_R _25841_ (.A(_16660_),
    .B(_10068_),
    .Y(_10074_));
 AO21x1_ASAP7_75t_R _25842_ (.A1(_09753_),
    .A2(_10056_),
    .B(_10074_),
    .Y(_03249_));
 AND2x2_ASAP7_75t_R _25843_ (.A(_16783_),
    .B(_10068_),
    .Y(_10075_));
 AO21x1_ASAP7_75t_R _25844_ (.A1(_09706_),
    .A2(_10047_),
    .B(_10075_),
    .Y(_03250_));
 AND2x2_ASAP7_75t_R _25845_ (.A(_16925_),
    .B(_10068_),
    .Y(_10076_));
 AO21x1_ASAP7_75t_R _25846_ (.A1(_09708_),
    .A2(_10047_),
    .B(_10076_),
    .Y(_03251_));
 AND2x2_ASAP7_75t_R _25847_ (.A(_04268_),
    .B(_10068_),
    .Y(_10077_));
 AO21x1_ASAP7_75t_R _25848_ (.A1(_09757_),
    .A2(_10047_),
    .B(_10077_),
    .Y(_03252_));
 AND2x2_ASAP7_75t_R _25849_ (.A(_04381_),
    .B(_10068_),
    .Y(_10078_));
 AO21x1_ASAP7_75t_R _25850_ (.A1(_09759_),
    .A2(_10047_),
    .B(_10078_),
    .Y(_03253_));
 AND2x2_ASAP7_75t_R _25851_ (.A(_04548_),
    .B(_10068_),
    .Y(_10079_));
 AO21x1_ASAP7_75t_R _25852_ (.A1(_09761_),
    .A2(_10047_),
    .B(_10079_),
    .Y(_03254_));
 AND2x2_ASAP7_75t_R _25853_ (.A(_04629_),
    .B(_10041_),
    .Y(_10080_));
 AO21x1_ASAP7_75t_R _25854_ (.A1(_09713_),
    .A2(_10047_),
    .B(_10080_),
    .Y(_03255_));
 BUFx6f_ASAP7_75t_R _25855_ (.A(_09365_),
    .Y(_10081_));
 AO21x1_ASAP7_75t_R _25856_ (.A1(_09993_),
    .A2(_09667_),
    .B(_04751_),
    .Y(_10082_));
 OA21x2_ASAP7_75t_R _25857_ (.A1(_10081_),
    .A2(_10042_),
    .B(_10082_),
    .Y(_03256_));
 AND2x2_ASAP7_75t_R _25858_ (.A(_04866_),
    .B(_10041_),
    .Y(_10083_));
 AO21x1_ASAP7_75t_R _25859_ (.A1(_09810_),
    .A2(_10047_),
    .B(_10083_),
    .Y(_03257_));
 NAND2x1_ASAP7_75t_R _25860_ (.A(_01781_),
    .B(_10059_),
    .Y(_10084_));
 OA21x2_ASAP7_75t_R _25861_ (.A1(_10019_),
    .A2(_10029_),
    .B(_10084_),
    .Y(_03258_));
 AND2x6_ASAP7_75t_R _25862_ (.A(_09993_),
    .B(_08953_),
    .Y(_10085_));
 BUFx12f_ASAP7_75t_R _25863_ (.A(_10085_),
    .Y(_10086_));
 NAND2x2_ASAP7_75t_R _25864_ (.A(_09993_),
    .B(_08953_),
    .Y(_10087_));
 BUFx12f_ASAP7_75t_R _25865_ (.A(_10087_),
    .Y(_10088_));
 AND2x2_ASAP7_75t_R _25866_ (.A(_00394_),
    .B(_10088_),
    .Y(_10089_));
 AOI21x1_ASAP7_75t_R _25867_ (.A1(_09902_),
    .A2(_10086_),
    .B(_10089_),
    .Y(_03259_));
 AND2x2_ASAP7_75t_R _25868_ (.A(_00427_),
    .B(_10088_),
    .Y(_10090_));
 AOI21x1_ASAP7_75t_R _25869_ (.A1(_09908_),
    .A2(_10086_),
    .B(_10090_),
    .Y(_03260_));
 NOR2x1_ASAP7_75t_R _25870_ (.A(_09898_),
    .B(_10088_),
    .Y(_10091_));
 AO21x1_ASAP7_75t_R _25871_ (.A1(_13567_),
    .A2(_10088_),
    .B(_10091_),
    .Y(_03261_));
 AND2x2_ASAP7_75t_R _25872_ (.A(_13636_),
    .B(_10088_),
    .Y(_10092_));
 AO21x1_ASAP7_75t_R _25873_ (.A1(_09819_),
    .A2(_10086_),
    .B(_10092_),
    .Y(_03262_));
 BUFx12f_ASAP7_75t_R _25874_ (.A(_10087_),
    .Y(_10093_));
 AND2x2_ASAP7_75t_R _25875_ (.A(_14799_),
    .B(_10093_),
    .Y(_10094_));
 AO21x1_ASAP7_75t_R _25876_ (.A1(_09726_),
    .A2(_10086_),
    .B(_10094_),
    .Y(_03263_));
 AND2x2_ASAP7_75t_R _25877_ (.A(_14862_),
    .B(_10093_),
    .Y(_10095_));
 AO21x1_ASAP7_75t_R _25878_ (.A1(_09679_),
    .A2(_10086_),
    .B(_10095_),
    .Y(_03264_));
 AND2x2_ASAP7_75t_R _25879_ (.A(_13867_),
    .B(_10093_),
    .Y(_10096_));
 AO21x1_ASAP7_75t_R _25880_ (.A1(_09729_),
    .A2(_10086_),
    .B(_10096_),
    .Y(_03265_));
 AND2x2_ASAP7_75t_R _25881_ (.A(_14991_),
    .B(_10093_),
    .Y(_10097_));
 AO21x1_ASAP7_75t_R _25882_ (.A1(_09731_),
    .A2(_10086_),
    .B(_10097_),
    .Y(_03266_));
 BUFx6f_ASAP7_75t_R _25883_ (.A(_08506_),
    .Y(_10098_));
 AND2x2_ASAP7_75t_R _25884_ (.A(_13996_),
    .B(_10093_),
    .Y(_10099_));
 AO21x1_ASAP7_75t_R _25885_ (.A1(_10098_),
    .A2(_10086_),
    .B(_10099_),
    .Y(_03267_));
 AND2x2_ASAP7_75t_R _25886_ (.A(_15125_),
    .B(_10093_),
    .Y(_10100_));
 AO21x1_ASAP7_75t_R _25887_ (.A1(_09784_),
    .A2(_10086_),
    .B(_10100_),
    .Y(_03268_));
 NAND2x1_ASAP7_75t_R _25888_ (.A(_01780_),
    .B(_10059_),
    .Y(_10101_));
 OA21x2_ASAP7_75t_R _25889_ (.A1(_09455_),
    .A2(_10029_),
    .B(_10101_),
    .Y(_03269_));
 BUFx6f_ASAP7_75t_R _25890_ (.A(_08669_),
    .Y(_10102_));
 BUFx12f_ASAP7_75t_R _25891_ (.A(_10085_),
    .Y(_10103_));
 BUFx12f_ASAP7_75t_R _25892_ (.A(_10103_),
    .Y(_10104_));
 AND2x2_ASAP7_75t_R _25893_ (.A(_14181_),
    .B(_10093_),
    .Y(_10105_));
 AO21x1_ASAP7_75t_R _25894_ (.A1(_10102_),
    .A2(_10104_),
    .B(_10105_),
    .Y(_03270_));
 AND2x2_ASAP7_75t_R _25895_ (.A(_14230_),
    .B(_10093_),
    .Y(_10106_));
 AO21x1_ASAP7_75t_R _25896_ (.A1(_09736_),
    .A2(_10104_),
    .B(_10106_),
    .Y(_03271_));
 BUFx6f_ASAP7_75t_R _25897_ (.A(_08757_),
    .Y(_10107_));
 AND2x2_ASAP7_75t_R _25898_ (.A(_13154_),
    .B(_10093_),
    .Y(_10108_));
 AO21x1_ASAP7_75t_R _25899_ (.A1(_10107_),
    .A2(_10104_),
    .B(_10108_),
    .Y(_03272_));
 AND2x2_ASAP7_75t_R _25900_ (.A(_15390_),
    .B(_10093_),
    .Y(_10109_));
 AO21x1_ASAP7_75t_R _25901_ (.A1(_09690_),
    .A2(_10104_),
    .B(_10109_),
    .Y(_03273_));
 NAND2x1_ASAP7_75t_R _25902_ (.A(_08851_),
    .B(_10103_),
    .Y(_10110_));
 OA21x2_ASAP7_75t_R _25903_ (.A1(_15543_),
    .A2(_10086_),
    .B(_10110_),
    .Y(_03274_));
 AO21x1_ASAP7_75t_R _25904_ (.A1(_09993_),
    .A2(_08954_),
    .B(_15666_),
    .Y(_10111_));
 OA21x2_ASAP7_75t_R _25905_ (.A1(_10019_),
    .A2(_10088_),
    .B(_10111_),
    .Y(_03275_));
 AND2x2_ASAP7_75t_R _25906_ (.A(_09930_),
    .B(_10103_),
    .Y(_10112_));
 AO21x1_ASAP7_75t_R _25907_ (.A1(_15822_),
    .A2(_10088_),
    .B(_10112_),
    .Y(_03276_));
 NOR2x1_ASAP7_75t_R _25908_ (.A(_09695_),
    .B(_10088_),
    .Y(_10113_));
 AO21x1_ASAP7_75t_R _25909_ (.A1(_15904_),
    .A2(_10088_),
    .B(_10113_),
    .Y(_03277_));
 BUFx6f_ASAP7_75t_R _25910_ (.A(_10087_),
    .Y(_10114_));
 AND2x2_ASAP7_75t_R _25911_ (.A(_16069_),
    .B(_10114_),
    .Y(_10115_));
 AO21x1_ASAP7_75t_R _25912_ (.A1(_09697_),
    .A2(_10104_),
    .B(_10115_),
    .Y(_03278_));
 AND2x2_ASAP7_75t_R _25913_ (.A(_16151_),
    .B(_10114_),
    .Y(_10116_));
 AO21x1_ASAP7_75t_R _25914_ (.A1(_09699_),
    .A2(_10104_),
    .B(_10116_),
    .Y(_03279_));
 AO21x1_ASAP7_75t_R _25915_ (.A1(_08950_),
    .A2(_09621_),
    .B(_01779_),
    .Y(_10117_));
 OAI21x1_ASAP7_75t_R _25916_ (.A1(_08948_),
    .A2(_09917_),
    .B(_10117_),
    .Y(_03280_));
 AND2x2_ASAP7_75t_R _25917_ (.A(_16286_),
    .B(_10114_),
    .Y(_10118_));
 AO21x1_ASAP7_75t_R _25918_ (.A1(_09701_),
    .A2(_10104_),
    .B(_10118_),
    .Y(_03281_));
 AND2x2_ASAP7_75t_R _25919_ (.A(_16409_),
    .B(_10114_),
    .Y(_10119_));
 AO21x1_ASAP7_75t_R _25920_ (.A1(_09749_),
    .A2(_10104_),
    .B(_10119_),
    .Y(_03282_));
 AND2x2_ASAP7_75t_R _25921_ (.A(_16547_),
    .B(_10114_),
    .Y(_10120_));
 AO21x1_ASAP7_75t_R _25922_ (.A1(_09751_),
    .A2(_10104_),
    .B(_10120_),
    .Y(_03283_));
 AND2x2_ASAP7_75t_R _25923_ (.A(_16657_),
    .B(_10114_),
    .Y(_10121_));
 AO21x1_ASAP7_75t_R _25924_ (.A1(_09753_),
    .A2(_10104_),
    .B(_10121_),
    .Y(_03284_));
 AND2x2_ASAP7_75t_R _25925_ (.A(_16780_),
    .B(_10114_),
    .Y(_10122_));
 AO21x1_ASAP7_75t_R _25926_ (.A1(_09706_),
    .A2(_10103_),
    .B(_10122_),
    .Y(_03285_));
 AND2x2_ASAP7_75t_R _25927_ (.A(_16922_),
    .B(_10114_),
    .Y(_10123_));
 AO21x1_ASAP7_75t_R _25928_ (.A1(_09708_),
    .A2(_10103_),
    .B(_10123_),
    .Y(_03286_));
 AND2x2_ASAP7_75t_R _25929_ (.A(_04265_),
    .B(_10114_),
    .Y(_10124_));
 AO21x1_ASAP7_75t_R _25930_ (.A1(_09757_),
    .A2(_10103_),
    .B(_10124_),
    .Y(_03287_));
 AND2x2_ASAP7_75t_R _25931_ (.A(_04378_),
    .B(_10114_),
    .Y(_10125_));
 AO21x1_ASAP7_75t_R _25932_ (.A1(_09759_),
    .A2(_10103_),
    .B(_10125_),
    .Y(_03288_));
 AND2x2_ASAP7_75t_R _25933_ (.A(_04545_),
    .B(_10087_),
    .Y(_10126_));
 AO21x1_ASAP7_75t_R _25934_ (.A1(_09761_),
    .A2(_10103_),
    .B(_10126_),
    .Y(_03289_));
 AND2x2_ASAP7_75t_R _25935_ (.A(_04626_),
    .B(_10087_),
    .Y(_10127_));
 AO21x1_ASAP7_75t_R _25936_ (.A1(_09713_),
    .A2(_10103_),
    .B(_10127_),
    .Y(_03290_));
 NAND2x1_ASAP7_75t_R _25937_ (.A(_01778_),
    .B(_10059_),
    .Y(_10128_));
 OA21x2_ASAP7_75t_R _25938_ (.A1(_09587_),
    .A2(_10029_),
    .B(_10128_),
    .Y(_03291_));
 AO21x1_ASAP7_75t_R _25939_ (.A1(_09993_),
    .A2(_08954_),
    .B(_04748_),
    .Y(_10129_));
 OA21x2_ASAP7_75t_R _25940_ (.A1(_10081_),
    .A2(_10088_),
    .B(_10129_),
    .Y(_03292_));
 AND2x2_ASAP7_75t_R _25941_ (.A(_04863_),
    .B(_10087_),
    .Y(_10130_));
 AO21x1_ASAP7_75t_R _25942_ (.A1(_09810_),
    .A2(_10103_),
    .B(_10130_),
    .Y(_03293_));
 NAND2x2_ASAP7_75t_R _25943_ (.A(_13685_),
    .B(_13602_),
    .Y(_10131_));
 AO211x2_ASAP7_75t_R _25944_ (.A1(_08256_),
    .A2(_08261_),
    .B(_07799_),
    .C(_09504_),
    .Y(_10132_));
 NOR2x2_ASAP7_75t_R _25945_ (.A(_10131_),
    .B(_10132_),
    .Y(_10133_));
 OR2x6_ASAP7_75t_R _25946_ (.A(_10131_),
    .B(_10132_),
    .Y(_10134_));
 BUFx12f_ASAP7_75t_R _25947_ (.A(_10134_),
    .Y(_10135_));
 AND2x2_ASAP7_75t_R _25948_ (.A(_00395_),
    .B(_10135_),
    .Y(_10136_));
 AOI21x1_ASAP7_75t_R _25949_ (.A1(_09902_),
    .A2(_10133_),
    .B(_10136_),
    .Y(_03294_));
 AND2x2_ASAP7_75t_R _25950_ (.A(_00428_),
    .B(_10135_),
    .Y(_10137_));
 AOI21x1_ASAP7_75t_R _25951_ (.A1(_09908_),
    .A2(_10133_),
    .B(_10137_),
    .Y(_03295_));
 BUFx12f_ASAP7_75t_R _25952_ (.A(_10135_),
    .Y(_10138_));
 AND2x2_ASAP7_75t_R _25953_ (.A(_09543_),
    .B(_10133_),
    .Y(_10139_));
 AOI21x1_ASAP7_75t_R _25954_ (.A1(_00459_),
    .A2(_10138_),
    .B(_10139_),
    .Y(_03296_));
 BUFx12f_ASAP7_75t_R _25955_ (.A(_10134_),
    .Y(_10140_));
 NAND2x1_ASAP7_75t_R _25956_ (.A(_00489_),
    .B(_10140_),
    .Y(_10141_));
 OA21x2_ASAP7_75t_R _25957_ (.A1(_09629_),
    .A2(_10138_),
    .B(_10141_),
    .Y(_03297_));
 BUFx12f_ASAP7_75t_R _25958_ (.A(_10134_),
    .Y(_10142_));
 NAND2x1_ASAP7_75t_R _25959_ (.A(_00519_),
    .B(_10142_),
    .Y(_10143_));
 OA21x2_ASAP7_75t_R _25960_ (.A1(_09563_),
    .A2(_10138_),
    .B(_10143_),
    .Y(_03298_));
 NAND2x1_ASAP7_75t_R _25961_ (.A(_00549_),
    .B(_10142_),
    .Y(_10144_));
 OA21x2_ASAP7_75t_R _25962_ (.A1(_09565_),
    .A2(_10138_),
    .B(_10144_),
    .Y(_03299_));
 NAND2x1_ASAP7_75t_R _25963_ (.A(_00579_),
    .B(_10142_),
    .Y(_10145_));
 OA21x2_ASAP7_75t_R _25964_ (.A1(_09567_),
    .A2(_10138_),
    .B(_10145_),
    .Y(_03300_));
 NAND2x1_ASAP7_75t_R _25965_ (.A(_00609_),
    .B(_10142_),
    .Y(_10146_));
 OA21x2_ASAP7_75t_R _25966_ (.A1(_09570_),
    .A2(_10138_),
    .B(_10146_),
    .Y(_03301_));
 NAND2x1_ASAP7_75t_R _25967_ (.A(_01777_),
    .B(_10059_),
    .Y(_10147_));
 OA21x2_ASAP7_75t_R _25968_ (.A1(_09589_),
    .A2(_10029_),
    .B(_10147_),
    .Y(_03302_));
 NAND2x1_ASAP7_75t_R _25969_ (.A(_00639_),
    .B(_10142_),
    .Y(_10148_));
 OA21x2_ASAP7_75t_R _25970_ (.A1(_09438_),
    .A2(_10138_),
    .B(_10148_),
    .Y(_03303_));
 AND2x2_ASAP7_75t_R _25971_ (.A(_14049_),
    .B(_10135_),
    .Y(_10149_));
 AO21x1_ASAP7_75t_R _25972_ (.A1(_09784_),
    .A2(_10133_),
    .B(_10149_),
    .Y(_03304_));
 NAND2x1_ASAP7_75t_R _25973_ (.A(_00699_),
    .B(_10142_),
    .Y(_10150_));
 OA21x2_ASAP7_75t_R _25974_ (.A1(_09443_),
    .A2(_10138_),
    .B(_10150_),
    .Y(_03305_));
 BUFx6f_ASAP7_75t_R _25975_ (.A(_10135_),
    .Y(_10151_));
 NAND2x1_ASAP7_75t_R _25976_ (.A(_00729_),
    .B(_10142_),
    .Y(_10152_));
 OA21x2_ASAP7_75t_R _25977_ (.A1(_09445_),
    .A2(_10151_),
    .B(_10152_),
    .Y(_03306_));
 NAND2x1_ASAP7_75t_R _25978_ (.A(_00359_),
    .B(_10142_),
    .Y(_10153_));
 OA21x2_ASAP7_75t_R _25979_ (.A1(_09447_),
    .A2(_10151_),
    .B(_10153_),
    .Y(_03307_));
 NAND2x1_ASAP7_75t_R _25980_ (.A(_00797_),
    .B(_10142_),
    .Y(_10154_));
 OA21x2_ASAP7_75t_R _25981_ (.A1(_09449_),
    .A2(_10151_),
    .B(_10154_),
    .Y(_03308_));
 AND2x2_ASAP7_75t_R _25982_ (.A(_09451_),
    .B(_10133_),
    .Y(_10155_));
 AOI21x1_ASAP7_75t_R _25983_ (.A1(_00829_),
    .A2(_10138_),
    .B(_10155_),
    .Y(_03309_));
 NAND2x1_ASAP7_75t_R _25984_ (.A(_00861_),
    .B(_10142_),
    .Y(_10156_));
 OA21x2_ASAP7_75t_R _25985_ (.A1(_10019_),
    .A2(_10151_),
    .B(_10156_),
    .Y(_03310_));
 BUFx12f_ASAP7_75t_R _25986_ (.A(_10134_),
    .Y(_10157_));
 NAND2x1_ASAP7_75t_R _25987_ (.A(_00893_),
    .B(_10157_),
    .Y(_10158_));
 OA21x2_ASAP7_75t_R _25988_ (.A1(_09455_),
    .A2(_10151_),
    .B(_10158_),
    .Y(_03311_));
 AND2x2_ASAP7_75t_R _25989_ (.A(_09457_),
    .B(_10133_),
    .Y(_10159_));
 AOI21x1_ASAP7_75t_R _25990_ (.A1(_00925_),
    .A2(_10138_),
    .B(_10159_),
    .Y(_03312_));
 NAND2x1_ASAP7_75t_R _25991_ (.A(_01776_),
    .B(_10059_),
    .Y(_10160_));
 OA21x2_ASAP7_75t_R _25992_ (.A1(_09592_),
    .A2(_10029_),
    .B(_10160_),
    .Y(_03313_));
 NAND2x1_ASAP7_75t_R _25993_ (.A(_00957_),
    .B(_10157_),
    .Y(_10161_));
 OA21x2_ASAP7_75t_R _25994_ (.A1(_09587_),
    .A2(_10151_),
    .B(_10161_),
    .Y(_03314_));
 NAND2x1_ASAP7_75t_R _25995_ (.A(_00989_),
    .B(_10157_),
    .Y(_10162_));
 OA21x2_ASAP7_75t_R _25996_ (.A1(_09589_),
    .A2(_10151_),
    .B(_10162_),
    .Y(_03315_));
 NAND2x1_ASAP7_75t_R _25997_ (.A(_01021_),
    .B(_10157_),
    .Y(_10163_));
 OA21x2_ASAP7_75t_R _25998_ (.A1(_09592_),
    .A2(_10151_),
    .B(_10163_),
    .Y(_03316_));
 NAND2x1_ASAP7_75t_R _25999_ (.A(_01053_),
    .B(_10157_),
    .Y(_10164_));
 OA21x2_ASAP7_75t_R _26000_ (.A1(_09594_),
    .A2(_10151_),
    .B(_10164_),
    .Y(_03317_));
 NAND2x1_ASAP7_75t_R _26001_ (.A(_01085_),
    .B(_10157_),
    .Y(_10165_));
 OA21x2_ASAP7_75t_R _26002_ (.A1(_09596_),
    .A2(_10151_),
    .B(_10165_),
    .Y(_03318_));
 NAND2x1_ASAP7_75t_R _26003_ (.A(_01117_),
    .B(_10157_),
    .Y(_10166_));
 OA21x2_ASAP7_75t_R _26004_ (.A1(_09598_),
    .A2(_10140_),
    .B(_10166_),
    .Y(_03319_));
 NAND2x1_ASAP7_75t_R _26005_ (.A(_01149_),
    .B(_10157_),
    .Y(_10167_));
 OA21x2_ASAP7_75t_R _26006_ (.A1(_09600_),
    .A2(_10140_),
    .B(_10167_),
    .Y(_03320_));
 NAND2x1_ASAP7_75t_R _26007_ (.A(_01181_),
    .B(_10157_),
    .Y(_10168_));
 OA21x2_ASAP7_75t_R _26008_ (.A1(_09602_),
    .A2(_10140_),
    .B(_10168_),
    .Y(_03321_));
 NAND2x1_ASAP7_75t_R _26009_ (.A(_01213_),
    .B(_10157_),
    .Y(_10169_));
 OA21x2_ASAP7_75t_R _26010_ (.A1(_09604_),
    .A2(_10140_),
    .B(_10169_),
    .Y(_03322_));
 NAND2x1_ASAP7_75t_R _26011_ (.A(_01245_),
    .B(_10135_),
    .Y(_10170_));
 OA21x2_ASAP7_75t_R _26012_ (.A1(_09606_),
    .A2(_10140_),
    .B(_10170_),
    .Y(_03323_));
 NAND2x1_ASAP7_75t_R _26013_ (.A(_01775_),
    .B(_10059_),
    .Y(_10171_));
 OA21x2_ASAP7_75t_R _26014_ (.A1(_09594_),
    .A2(_10029_),
    .B(_10171_),
    .Y(_03324_));
 NAND2x1_ASAP7_75t_R _26015_ (.A(_01277_),
    .B(_10135_),
    .Y(_10172_));
 OA21x2_ASAP7_75t_R _26016_ (.A1(_09608_),
    .A2(_10140_),
    .B(_10172_),
    .Y(_03325_));
 NAND2x1_ASAP7_75t_R _26017_ (.A(_01309_),
    .B(_10135_),
    .Y(_10173_));
 OA21x2_ASAP7_75t_R _26018_ (.A1(_09610_),
    .A2(_10140_),
    .B(_10173_),
    .Y(_03326_));
 NAND2x1_ASAP7_75t_R _26019_ (.A(_01341_),
    .B(_10135_),
    .Y(_10174_));
 OA21x2_ASAP7_75t_R _26020_ (.A1(_10081_),
    .A2(_10140_),
    .B(_10174_),
    .Y(_03327_));
 NAND2x1_ASAP7_75t_R _26021_ (.A(_01373_),
    .B(_10135_),
    .Y(_10175_));
 OA21x2_ASAP7_75t_R _26022_ (.A1(_09614_),
    .A2(_10140_),
    .B(_10175_),
    .Y(_03328_));
 AO211x2_ASAP7_75t_R _26023_ (.A1(_08256_),
    .A2(_08261_),
    .B(_09618_),
    .C(_07799_),
    .Y(_10176_));
 NOR2x2_ASAP7_75t_R _26024_ (.A(_10131_),
    .B(_10176_),
    .Y(_10177_));
 OR2x6_ASAP7_75t_R _26025_ (.A(_10131_),
    .B(_10176_),
    .Y(_10178_));
 BUFx12f_ASAP7_75t_R _26026_ (.A(_10178_),
    .Y(_10179_));
 BUFx12f_ASAP7_75t_R _26027_ (.A(_10179_),
    .Y(_10180_));
 AND2x2_ASAP7_75t_R _26028_ (.A(_00396_),
    .B(_10180_),
    .Y(_10181_));
 AOI21x1_ASAP7_75t_R _26029_ (.A1(_09902_),
    .A2(_10177_),
    .B(_10181_),
    .Y(_03329_));
 AND2x2_ASAP7_75t_R _26030_ (.A(_00429_),
    .B(_10180_),
    .Y(_10182_));
 AOI21x1_ASAP7_75t_R _26031_ (.A1(_09908_),
    .A2(_10177_),
    .B(_10182_),
    .Y(_03330_));
 AND2x2_ASAP7_75t_R _26032_ (.A(_00460_),
    .B(_10180_),
    .Y(_10183_));
 AOI21x1_ASAP7_75t_R _26033_ (.A1(_09675_),
    .A2(_10177_),
    .B(_10183_),
    .Y(_03331_));
 BUFx6f_ASAP7_75t_R _26034_ (.A(_10180_),
    .Y(_10184_));
 BUFx12f_ASAP7_75t_R _26035_ (.A(_10179_),
    .Y(_10185_));
 NAND2x1_ASAP7_75t_R _26036_ (.A(_00490_),
    .B(_10185_),
    .Y(_10186_));
 OA21x2_ASAP7_75t_R _26037_ (.A1(_09629_),
    .A2(_10184_),
    .B(_10186_),
    .Y(_03332_));
 NAND2x1_ASAP7_75t_R _26038_ (.A(_00520_),
    .B(_10185_),
    .Y(_10187_));
 OA21x2_ASAP7_75t_R _26039_ (.A1(_09563_),
    .A2(_10184_),
    .B(_10187_),
    .Y(_03333_));
 NAND2x1_ASAP7_75t_R _26040_ (.A(_00550_),
    .B(_10185_),
    .Y(_10188_));
 OA21x2_ASAP7_75t_R _26041_ (.A1(_09565_),
    .A2(_10184_),
    .B(_10188_),
    .Y(_03334_));
 NAND2x1_ASAP7_75t_R _26042_ (.A(_01774_),
    .B(_10059_),
    .Y(_10189_));
 OA21x2_ASAP7_75t_R _26043_ (.A1(_09596_),
    .A2(_10029_),
    .B(_10189_),
    .Y(_03335_));
 BUFx12f_ASAP7_75t_R _26044_ (.A(_10179_),
    .Y(_10190_));
 NAND2x1_ASAP7_75t_R _26045_ (.A(_00580_),
    .B(_10190_),
    .Y(_10191_));
 OA21x2_ASAP7_75t_R _26046_ (.A1(_09567_),
    .A2(_10184_),
    .B(_10191_),
    .Y(_03336_));
 NAND2x1_ASAP7_75t_R _26047_ (.A(_00610_),
    .B(_10190_),
    .Y(_10192_));
 OA21x2_ASAP7_75t_R _26048_ (.A1(_09570_),
    .A2(_10184_),
    .B(_10192_),
    .Y(_03337_));
 NAND2x1_ASAP7_75t_R _26049_ (.A(_00640_),
    .B(_10190_),
    .Y(_10193_));
 OA21x2_ASAP7_75t_R _26050_ (.A1(_09438_),
    .A2(_10184_),
    .B(_10193_),
    .Y(_03338_));
 NAND2x1_ASAP7_75t_R _26051_ (.A(_00670_),
    .B(_10190_),
    .Y(_10194_));
 OA21x2_ASAP7_75t_R _26052_ (.A1(_09441_),
    .A2(_10184_),
    .B(_10194_),
    .Y(_03339_));
 NAND2x1_ASAP7_75t_R _26053_ (.A(_00700_),
    .B(_10190_),
    .Y(_10195_));
 OA21x2_ASAP7_75t_R _26054_ (.A1(_09443_),
    .A2(_10184_),
    .B(_10195_),
    .Y(_03340_));
 NAND2x1_ASAP7_75t_R _26055_ (.A(_00730_),
    .B(_10190_),
    .Y(_10196_));
 OA21x2_ASAP7_75t_R _26056_ (.A1(_09445_),
    .A2(_10184_),
    .B(_10196_),
    .Y(_03341_));
 NAND2x1_ASAP7_75t_R _26057_ (.A(_00360_),
    .B(_10190_),
    .Y(_10197_));
 OA21x2_ASAP7_75t_R _26058_ (.A1(_09447_),
    .A2(_10184_),
    .B(_10197_),
    .Y(_03342_));
 BUFx6f_ASAP7_75t_R _26059_ (.A(_10179_),
    .Y(_10198_));
 NAND2x1_ASAP7_75t_R _26060_ (.A(_00798_),
    .B(_10190_),
    .Y(_10199_));
 OA21x2_ASAP7_75t_R _26061_ (.A1(_09449_),
    .A2(_10198_),
    .B(_10199_),
    .Y(_03343_));
 AND2x2_ASAP7_75t_R _26062_ (.A(_00830_),
    .B(_10180_),
    .Y(_10200_));
 AOI21x1_ASAP7_75t_R _26063_ (.A1(_09790_),
    .A2(_10177_),
    .B(_10200_),
    .Y(_03344_));
 NAND2x1_ASAP7_75t_R _26064_ (.A(_00862_),
    .B(_10190_),
    .Y(_10201_));
 OA21x2_ASAP7_75t_R _26065_ (.A1(_10019_),
    .A2(_10198_),
    .B(_10201_),
    .Y(_03345_));
 NAND2x1_ASAP7_75t_R _26066_ (.A(_01773_),
    .B(_10059_),
    .Y(_10202_));
 OA21x2_ASAP7_75t_R _26067_ (.A1(_09598_),
    .A2(_09897_),
    .B(_10202_),
    .Y(_03346_));
 NAND2x1_ASAP7_75t_R _26068_ (.A(_00894_),
    .B(_10190_),
    .Y(_10203_));
 OA21x2_ASAP7_75t_R _26069_ (.A1(_09455_),
    .A2(_10198_),
    .B(_10203_),
    .Y(_03347_));
 AND2x2_ASAP7_75t_R _26070_ (.A(_00926_),
    .B(_10180_),
    .Y(_10204_));
 AOI21x1_ASAP7_75t_R _26071_ (.A1(_08948_),
    .A2(_10177_),
    .B(_10204_),
    .Y(_03348_));
 BUFx12f_ASAP7_75t_R _26072_ (.A(_10179_),
    .Y(_10205_));
 NAND2x1_ASAP7_75t_R _26073_ (.A(_00958_),
    .B(_10205_),
    .Y(_10206_));
 OA21x2_ASAP7_75t_R _26074_ (.A1(_09587_),
    .A2(_10198_),
    .B(_10206_),
    .Y(_03349_));
 NAND2x1_ASAP7_75t_R _26075_ (.A(_00990_),
    .B(_10205_),
    .Y(_10207_));
 OA21x2_ASAP7_75t_R _26076_ (.A1(_09589_),
    .A2(_10198_),
    .B(_10207_),
    .Y(_03350_));
 NAND2x1_ASAP7_75t_R _26077_ (.A(_01022_),
    .B(_10205_),
    .Y(_10208_));
 OA21x2_ASAP7_75t_R _26078_ (.A1(_09592_),
    .A2(_10198_),
    .B(_10208_),
    .Y(_03351_));
 NAND2x1_ASAP7_75t_R _26079_ (.A(_01054_),
    .B(_10205_),
    .Y(_10209_));
 OA21x2_ASAP7_75t_R _26080_ (.A1(_09594_),
    .A2(_10198_),
    .B(_10209_),
    .Y(_03352_));
 NAND2x1_ASAP7_75t_R _26081_ (.A(_01086_),
    .B(_10205_),
    .Y(_10210_));
 OA21x2_ASAP7_75t_R _26082_ (.A1(_09596_),
    .A2(_10198_),
    .B(_10210_),
    .Y(_03353_));
 NAND2x1_ASAP7_75t_R _26083_ (.A(_01118_),
    .B(_10205_),
    .Y(_10211_));
 OA21x2_ASAP7_75t_R _26084_ (.A1(_09598_),
    .A2(_10198_),
    .B(_10211_),
    .Y(_03354_));
 NAND2x1_ASAP7_75t_R _26085_ (.A(_01150_),
    .B(_10205_),
    .Y(_10212_));
 OA21x2_ASAP7_75t_R _26086_ (.A1(_09600_),
    .A2(_10198_),
    .B(_10212_),
    .Y(_03355_));
 NAND2x1_ASAP7_75t_R _26087_ (.A(_01182_),
    .B(_10205_),
    .Y(_10213_));
 OA21x2_ASAP7_75t_R _26088_ (.A1(_09602_),
    .A2(_10185_),
    .B(_10213_),
    .Y(_03356_));
 NAND2x1_ASAP7_75t_R _26089_ (.A(_01772_),
    .B(_10059_),
    .Y(_10214_));
 OA21x2_ASAP7_75t_R _26090_ (.A1(_09600_),
    .A2(_09897_),
    .B(_10214_),
    .Y(_03357_));
 NAND2x1_ASAP7_75t_R _26091_ (.A(_01214_),
    .B(_10205_),
    .Y(_10215_));
 OA21x2_ASAP7_75t_R _26092_ (.A1(_09604_),
    .A2(_10185_),
    .B(_10215_),
    .Y(_03358_));
 NAND2x1_ASAP7_75t_R _26093_ (.A(_01246_),
    .B(_10205_),
    .Y(_10216_));
 OA21x2_ASAP7_75t_R _26094_ (.A1(_09606_),
    .A2(_10185_),
    .B(_10216_),
    .Y(_03359_));
 NAND2x1_ASAP7_75t_R _26095_ (.A(_01278_),
    .B(_10180_),
    .Y(_10217_));
 OA21x2_ASAP7_75t_R _26096_ (.A1(_09608_),
    .A2(_10185_),
    .B(_10217_),
    .Y(_03360_));
 NAND2x1_ASAP7_75t_R _26097_ (.A(_01310_),
    .B(_10180_),
    .Y(_10218_));
 OA21x2_ASAP7_75t_R _26098_ (.A1(_09610_),
    .A2(_10185_),
    .B(_10218_),
    .Y(_03361_));
 NAND2x1_ASAP7_75t_R _26099_ (.A(_01342_),
    .B(_10180_),
    .Y(_10219_));
 OA21x2_ASAP7_75t_R _26100_ (.A1(_10081_),
    .A2(_10185_),
    .B(_10219_),
    .Y(_03362_));
 NAND2x1_ASAP7_75t_R _26101_ (.A(_01374_),
    .B(_10180_),
    .Y(_10220_));
 OA21x2_ASAP7_75t_R _26102_ (.A1(_09614_),
    .A2(_10185_),
    .B(_10220_),
    .Y(_03363_));
 AO211x2_ASAP7_75t_R _26103_ (.A1(_08256_),
    .A2(_08261_),
    .B(_09663_),
    .C(_07799_),
    .Y(_10221_));
 NOR2x2_ASAP7_75t_R _26104_ (.A(_10131_),
    .B(_10221_),
    .Y(_10222_));
 BUFx12f_ASAP7_75t_R _26105_ (.A(_10222_),
    .Y(_10223_));
 OR2x6_ASAP7_75t_R _26106_ (.A(_10131_),
    .B(_10221_),
    .Y(_10224_));
 BUFx12f_ASAP7_75t_R _26107_ (.A(_10224_),
    .Y(_10225_));
 BUFx6f_ASAP7_75t_R _26108_ (.A(_10225_),
    .Y(_10226_));
 AND2x2_ASAP7_75t_R _26109_ (.A(_00397_),
    .B(_10226_),
    .Y(_10227_));
 AOI21x1_ASAP7_75t_R _26110_ (.A1(_09902_),
    .A2(_10223_),
    .B(_10227_),
    .Y(_03364_));
 AND2x2_ASAP7_75t_R _26111_ (.A(_00430_),
    .B(_10226_),
    .Y(_10228_));
 AOI21x1_ASAP7_75t_R _26112_ (.A1(_09908_),
    .A2(_10223_),
    .B(_10228_),
    .Y(_03365_));
 BUFx6f_ASAP7_75t_R _26113_ (.A(_10225_),
    .Y(_10229_));
 NOR2x1_ASAP7_75t_R _26114_ (.A(_09898_),
    .B(_10229_),
    .Y(_10230_));
 AO21x1_ASAP7_75t_R _26115_ (.A1(_13581_),
    .A2(_10229_),
    .B(_10230_),
    .Y(_03366_));
 AND2x2_ASAP7_75t_R _26116_ (.A(_13663_),
    .B(_10226_),
    .Y(_10231_));
 AO21x1_ASAP7_75t_R _26117_ (.A1(_09819_),
    .A2(_10223_),
    .B(_10231_),
    .Y(_03367_));
 NAND2x1_ASAP7_75t_R _26118_ (.A(_01771_),
    .B(_09870_),
    .Y(_10232_));
 OA21x2_ASAP7_75t_R _26119_ (.A1(_09602_),
    .A2(_09897_),
    .B(_10232_),
    .Y(_03368_));
 AND2x2_ASAP7_75t_R _26120_ (.A(_13757_),
    .B(_10226_),
    .Y(_10233_));
 AO21x1_ASAP7_75t_R _26121_ (.A1(_09726_),
    .A2(_10223_),
    .B(_10233_),
    .Y(_03369_));
 AND2x2_ASAP7_75t_R _26122_ (.A(_13792_),
    .B(_10226_),
    .Y(_10234_));
 AO21x1_ASAP7_75t_R _26123_ (.A1(_09268_),
    .A2(_10223_),
    .B(_10234_),
    .Y(_03370_));
 AND2x2_ASAP7_75t_R _26124_ (.A(_13881_),
    .B(_10226_),
    .Y(_10235_));
 AO21x1_ASAP7_75t_R _26125_ (.A1(_09729_),
    .A2(_10223_),
    .B(_10235_),
    .Y(_03371_));
 AND2x2_ASAP7_75t_R _26126_ (.A(_13944_),
    .B(_10226_),
    .Y(_10236_));
 AO21x1_ASAP7_75t_R _26127_ (.A1(_09731_),
    .A2(_10223_),
    .B(_10236_),
    .Y(_03372_));
 AND2x2_ASAP7_75t_R _26128_ (.A(_13988_),
    .B(_10226_),
    .Y(_10237_));
 AO21x1_ASAP7_75t_R _26129_ (.A1(_10098_),
    .A2(_10223_),
    .B(_10237_),
    .Y(_03373_));
 AND2x2_ASAP7_75t_R _26130_ (.A(_15151_),
    .B(_10226_),
    .Y(_10238_));
 AO21x1_ASAP7_75t_R _26131_ (.A1(_09784_),
    .A2(_10223_),
    .B(_10238_),
    .Y(_03374_));
 BUFx12f_ASAP7_75t_R _26132_ (.A(_10225_),
    .Y(_10239_));
 AND2x2_ASAP7_75t_R _26133_ (.A(_14196_),
    .B(_10239_),
    .Y(_10240_));
 AO21x1_ASAP7_75t_R _26134_ (.A1(_10102_),
    .A2(_10223_),
    .B(_10240_),
    .Y(_03375_));
 BUFx12f_ASAP7_75t_R _26135_ (.A(_10222_),
    .Y(_10241_));
 AND2x2_ASAP7_75t_R _26136_ (.A(_14225_),
    .B(_10239_),
    .Y(_10242_));
 AO21x1_ASAP7_75t_R _26137_ (.A1(_09736_),
    .A2(_10241_),
    .B(_10242_),
    .Y(_03376_));
 AND2x2_ASAP7_75t_R _26138_ (.A(_13210_),
    .B(_10239_),
    .Y(_10243_));
 AO21x1_ASAP7_75t_R _26139_ (.A1(_10107_),
    .A2(_10241_),
    .B(_10243_),
    .Y(_03377_));
 BUFx6f_ASAP7_75t_R _26140_ (.A(_08802_),
    .Y(_10244_));
 AND2x2_ASAP7_75t_R _26141_ (.A(_15424_),
    .B(_10239_),
    .Y(_10245_));
 AO21x1_ASAP7_75t_R _26142_ (.A1(_10244_),
    .A2(_10241_),
    .B(_10245_),
    .Y(_03378_));
 NAND2x1_ASAP7_75t_R _26143_ (.A(_01770_),
    .B(_09870_),
    .Y(_10246_));
 OA21x2_ASAP7_75t_R _26144_ (.A1(_09604_),
    .A2(_09897_),
    .B(_10246_),
    .Y(_03379_));
 NOR2x1_ASAP7_75t_R _26145_ (.A(_08851_),
    .B(_10229_),
    .Y(_10247_));
 AO21x1_ASAP7_75t_R _26146_ (.A1(_15577_),
    .A2(_10229_),
    .B(_10247_),
    .Y(_03380_));
 NAND2x1_ASAP7_75t_R _26147_ (.A(_00863_),
    .B(_10229_),
    .Y(_10248_));
 OA21x2_ASAP7_75t_R _26148_ (.A1(_10019_),
    .A2(_10229_),
    .B(_10248_),
    .Y(_03381_));
 AND2x2_ASAP7_75t_R _26149_ (.A(_09930_),
    .B(_10222_),
    .Y(_10249_));
 AO21x1_ASAP7_75t_R _26150_ (.A1(_15783_),
    .A2(_10229_),
    .B(_10249_),
    .Y(_03382_));
 NOR2x1_ASAP7_75t_R _26151_ (.A(_09695_),
    .B(_10226_),
    .Y(_10250_));
 AO21x1_ASAP7_75t_R _26152_ (.A1(_15938_),
    .A2(_10229_),
    .B(_10250_),
    .Y(_03383_));
 AND2x2_ASAP7_75t_R _26153_ (.A(_16030_),
    .B(_10239_),
    .Y(_10251_));
 AO21x1_ASAP7_75t_R _26154_ (.A1(_09022_),
    .A2(_10241_),
    .B(_10251_),
    .Y(_03384_));
 AND2x2_ASAP7_75t_R _26155_ (.A(_16185_),
    .B(_10239_),
    .Y(_10252_));
 AO21x1_ASAP7_75t_R _26156_ (.A1(_09049_),
    .A2(_10241_),
    .B(_10252_),
    .Y(_03385_));
 AND2x2_ASAP7_75t_R _26157_ (.A(_16320_),
    .B(_10239_),
    .Y(_10253_));
 AO21x1_ASAP7_75t_R _26158_ (.A1(_09075_),
    .A2(_10241_),
    .B(_10253_),
    .Y(_03386_));
 AND2x2_ASAP7_75t_R _26159_ (.A(_16443_),
    .B(_10239_),
    .Y(_10254_));
 AO21x1_ASAP7_75t_R _26160_ (.A1(_09749_),
    .A2(_10241_),
    .B(_10254_),
    .Y(_03387_));
 AND2x2_ASAP7_75t_R _26161_ (.A(_16581_),
    .B(_10239_),
    .Y(_10255_));
 AO21x1_ASAP7_75t_R _26162_ (.A1(_09751_),
    .A2(_10241_),
    .B(_10255_),
    .Y(_03388_));
 AND2x2_ASAP7_75t_R _26163_ (.A(_16691_),
    .B(_10239_),
    .Y(_10256_));
 AO21x1_ASAP7_75t_R _26164_ (.A1(_09753_),
    .A2(_10241_),
    .B(_10256_),
    .Y(_03389_));
 NAND2x1_ASAP7_75t_R _26165_ (.A(_01769_),
    .B(_09870_),
    .Y(_10257_));
 OA21x2_ASAP7_75t_R _26166_ (.A1(_09606_),
    .A2(_09897_),
    .B(_10257_),
    .Y(_03390_));
 AND2x2_ASAP7_75t_R _26167_ (.A(_16814_),
    .B(_10225_),
    .Y(_10258_));
 AO21x1_ASAP7_75t_R _26168_ (.A1(_09177_),
    .A2(_10241_),
    .B(_10258_),
    .Y(_03391_));
 AND2x2_ASAP7_75t_R _26169_ (.A(_16883_),
    .B(_10225_),
    .Y(_10259_));
 AO21x1_ASAP7_75t_R _26170_ (.A1(_09204_),
    .A2(_10222_),
    .B(_10259_),
    .Y(_03392_));
 AND2x2_ASAP7_75t_R _26171_ (.A(_04299_),
    .B(_10225_),
    .Y(_10260_));
 AO21x1_ASAP7_75t_R _26172_ (.A1(_09757_),
    .A2(_10222_),
    .B(_10260_),
    .Y(_03393_));
 AND2x2_ASAP7_75t_R _26173_ (.A(_04412_),
    .B(_10225_),
    .Y(_10261_));
 AO21x1_ASAP7_75t_R _26174_ (.A1(_09759_),
    .A2(_10222_),
    .B(_10261_),
    .Y(_03394_));
 AND2x2_ASAP7_75t_R _26175_ (.A(_04506_),
    .B(_10225_),
    .Y(_10262_));
 AO21x1_ASAP7_75t_R _26176_ (.A1(_09761_),
    .A2(_10222_),
    .B(_10262_),
    .Y(_03395_));
 AND2x2_ASAP7_75t_R _26177_ (.A(_04660_),
    .B(_10225_),
    .Y(_10263_));
 AO21x1_ASAP7_75t_R _26178_ (.A1(_09335_),
    .A2(_10222_),
    .B(_10263_),
    .Y(_03396_));
 NAND2x1_ASAP7_75t_R _26179_ (.A(_01343_),
    .B(_10229_),
    .Y(_10264_));
 OA21x2_ASAP7_75t_R _26180_ (.A1(_10081_),
    .A2(_10229_),
    .B(_10264_),
    .Y(_03397_));
 AND2x2_ASAP7_75t_R _26181_ (.A(_04859_),
    .B(_10225_),
    .Y(_10265_));
 AO21x1_ASAP7_75t_R _26182_ (.A1(_09810_),
    .A2(_10222_),
    .B(_10265_),
    .Y(_03398_));
 NOR2x2_ASAP7_75t_R _26183_ (.A(_10131_),
    .B(_08263_),
    .Y(_10266_));
 BUFx6f_ASAP7_75t_R _26184_ (.A(_10266_),
    .Y(_10267_));
 OR2x6_ASAP7_75t_R _26185_ (.A(_10131_),
    .B(_08263_),
    .Y(_10268_));
 BUFx12f_ASAP7_75t_R _26186_ (.A(_10268_),
    .Y(_10269_));
 BUFx6f_ASAP7_75t_R _26187_ (.A(_10269_),
    .Y(_10270_));
 AND2x2_ASAP7_75t_R _26188_ (.A(_00398_),
    .B(_10270_),
    .Y(_10271_));
 AOI21x1_ASAP7_75t_R _26189_ (.A1(_09902_),
    .A2(_10267_),
    .B(_10271_),
    .Y(_03399_));
 AND2x2_ASAP7_75t_R _26190_ (.A(_00431_),
    .B(_10270_),
    .Y(_10272_));
 AOI21x1_ASAP7_75t_R _26191_ (.A1(_09908_),
    .A2(_10267_),
    .B(_10272_),
    .Y(_03400_));
 NAND2x1_ASAP7_75t_R _26192_ (.A(_01768_),
    .B(_09870_),
    .Y(_10273_));
 OA21x2_ASAP7_75t_R _26193_ (.A1(_09608_),
    .A2(_09897_),
    .B(_10273_),
    .Y(_03401_));
 BUFx6f_ASAP7_75t_R _26194_ (.A(_10269_),
    .Y(_10274_));
 NOR2x1_ASAP7_75t_R _26195_ (.A(_09898_),
    .B(_10274_),
    .Y(_10275_));
 AO21x1_ASAP7_75t_R _26196_ (.A1(_13578_),
    .A2(_10274_),
    .B(_10275_),
    .Y(_03402_));
 AND2x2_ASAP7_75t_R _26197_ (.A(_13660_),
    .B(_10270_),
    .Y(_10276_));
 AO21x1_ASAP7_75t_R _26198_ (.A1(_09819_),
    .A2(_10267_),
    .B(_10276_),
    .Y(_03403_));
 AND2x2_ASAP7_75t_R _26199_ (.A(_13754_),
    .B(_10270_),
    .Y(_10277_));
 AO21x1_ASAP7_75t_R _26200_ (.A1(_08993_),
    .A2(_10267_),
    .B(_10277_),
    .Y(_03404_));
 AND2x2_ASAP7_75t_R _26201_ (.A(_13789_),
    .B(_10270_),
    .Y(_10278_));
 AO21x1_ASAP7_75t_R _26202_ (.A1(_09268_),
    .A2(_10267_),
    .B(_10278_),
    .Y(_03405_));
 AND2x2_ASAP7_75t_R _26203_ (.A(_13884_),
    .B(_10270_),
    .Y(_10279_));
 AO21x1_ASAP7_75t_R _26204_ (.A1(_09412_),
    .A2(_10267_),
    .B(_10279_),
    .Y(_03406_));
 AND2x2_ASAP7_75t_R _26205_ (.A(_13947_),
    .B(_10270_),
    .Y(_10280_));
 AO21x1_ASAP7_75t_R _26206_ (.A1(_09436_),
    .A2(_10267_),
    .B(_10280_),
    .Y(_03407_));
 AND2x2_ASAP7_75t_R _26207_ (.A(_13985_),
    .B(_10270_),
    .Y(_10281_));
 AO21x1_ASAP7_75t_R _26208_ (.A1(_10098_),
    .A2(_10267_),
    .B(_10281_),
    .Y(_03408_));
 BUFx6f_ASAP7_75t_R _26209_ (.A(_08615_),
    .Y(_10282_));
 AND2x2_ASAP7_75t_R _26210_ (.A(_14052_),
    .B(_10270_),
    .Y(_10283_));
 AO21x1_ASAP7_75t_R _26211_ (.A1(_10282_),
    .A2(_10267_),
    .B(_10283_),
    .Y(_03409_));
 BUFx6f_ASAP7_75t_R _26212_ (.A(_10269_),
    .Y(_10284_));
 AND2x2_ASAP7_75t_R _26213_ (.A(_14193_),
    .B(_10284_),
    .Y(_10285_));
 AO21x1_ASAP7_75t_R _26214_ (.A1(_10102_),
    .A2(_10267_),
    .B(_10285_),
    .Y(_03410_));
 BUFx6f_ASAP7_75t_R _26215_ (.A(_08719_),
    .Y(_10286_));
 BUFx6f_ASAP7_75t_R _26216_ (.A(_10266_),
    .Y(_10287_));
 AND2x2_ASAP7_75t_R _26217_ (.A(_14222_),
    .B(_10284_),
    .Y(_10288_));
 AO21x1_ASAP7_75t_R _26218_ (.A1(_10286_),
    .A2(_10287_),
    .B(_10288_),
    .Y(_03411_));
 NAND2x1_ASAP7_75t_R _26219_ (.A(_01767_),
    .B(_09870_),
    .Y(_10289_));
 OA21x2_ASAP7_75t_R _26220_ (.A1(_09610_),
    .A2(_09897_),
    .B(_10289_),
    .Y(_03412_));
 AND2x2_ASAP7_75t_R _26221_ (.A(_13207_),
    .B(_10284_),
    .Y(_10290_));
 AO21x1_ASAP7_75t_R _26222_ (.A1(_10107_),
    .A2(_10287_),
    .B(_10290_),
    .Y(_03413_));
 AND2x2_ASAP7_75t_R _26223_ (.A(_15421_),
    .B(_10284_),
    .Y(_10291_));
 AO21x1_ASAP7_75t_R _26224_ (.A1(_10244_),
    .A2(_10287_),
    .B(_10291_),
    .Y(_03414_));
 NOR2x1_ASAP7_75t_R _26225_ (.A(_08851_),
    .B(_10274_),
    .Y(_10292_));
 AO21x1_ASAP7_75t_R _26226_ (.A1(_15574_),
    .A2(_10274_),
    .B(_10292_),
    .Y(_03415_));
 NAND2x1_ASAP7_75t_R _26227_ (.A(_00864_),
    .B(_10274_),
    .Y(_10293_));
 OA21x2_ASAP7_75t_R _26228_ (.A1(_10019_),
    .A2(_10274_),
    .B(_10293_),
    .Y(_03416_));
 AND2x2_ASAP7_75t_R _26229_ (.A(_09930_),
    .B(_10266_),
    .Y(_10294_));
 AO21x1_ASAP7_75t_R _26230_ (.A1(_15780_),
    .A2(_10274_),
    .B(_10294_),
    .Y(_03417_));
 NOR2x1_ASAP7_75t_R _26231_ (.A(_09695_),
    .B(_10270_),
    .Y(_10295_));
 AO21x1_ASAP7_75t_R _26232_ (.A1(_15935_),
    .A2(_10274_),
    .B(_10295_),
    .Y(_03418_));
 AND2x2_ASAP7_75t_R _26233_ (.A(_16027_),
    .B(_10284_),
    .Y(_10296_));
 AO21x1_ASAP7_75t_R _26234_ (.A1(_09022_),
    .A2(_10287_),
    .B(_10296_),
    .Y(_03419_));
 AND2x2_ASAP7_75t_R _26235_ (.A(_16182_),
    .B(_10284_),
    .Y(_10297_));
 AO21x1_ASAP7_75t_R _26236_ (.A1(_09049_),
    .A2(_10287_),
    .B(_10297_),
    .Y(_03420_));
 AND2x2_ASAP7_75t_R _26237_ (.A(_16317_),
    .B(_10284_),
    .Y(_10298_));
 AO21x1_ASAP7_75t_R _26238_ (.A1(_09075_),
    .A2(_10287_),
    .B(_10298_),
    .Y(_03421_));
 AND2x2_ASAP7_75t_R _26239_ (.A(_16440_),
    .B(_10284_),
    .Y(_10299_));
 AO21x1_ASAP7_75t_R _26240_ (.A1(_09100_),
    .A2(_10287_),
    .B(_10299_),
    .Y(_03422_));
 NAND2x1_ASAP7_75t_R _26241_ (.A(_01766_),
    .B(_09870_),
    .Y(_10300_));
 OA21x2_ASAP7_75t_R _26242_ (.A1(_10081_),
    .A2(_09897_),
    .B(_10300_),
    .Y(_03423_));
 AND2x2_ASAP7_75t_R _26243_ (.A(_16578_),
    .B(_10284_),
    .Y(_10301_));
 AO21x1_ASAP7_75t_R _26244_ (.A1(_09124_),
    .A2(_10287_),
    .B(_10301_),
    .Y(_03424_));
 AND2x2_ASAP7_75t_R _26245_ (.A(_16688_),
    .B(_10284_),
    .Y(_10302_));
 AO21x1_ASAP7_75t_R _26246_ (.A1(_09145_),
    .A2(_10287_),
    .B(_10302_),
    .Y(_03425_));
 AND2x2_ASAP7_75t_R _26247_ (.A(_16811_),
    .B(_10269_),
    .Y(_10303_));
 AO21x1_ASAP7_75t_R _26248_ (.A1(_09177_),
    .A2(_10287_),
    .B(_10303_),
    .Y(_03426_));
 AND2x2_ASAP7_75t_R _26249_ (.A(_16880_),
    .B(_10269_),
    .Y(_10304_));
 AO21x1_ASAP7_75t_R _26250_ (.A1(_09204_),
    .A2(_10266_),
    .B(_10304_),
    .Y(_03427_));
 AND2x2_ASAP7_75t_R _26251_ (.A(_04296_),
    .B(_10269_),
    .Y(_10305_));
 AO21x1_ASAP7_75t_R _26252_ (.A1(_09230_),
    .A2(_10266_),
    .B(_10305_),
    .Y(_03428_));
 AND2x2_ASAP7_75t_R _26253_ (.A(_04409_),
    .B(_10269_),
    .Y(_10306_));
 AO21x1_ASAP7_75t_R _26254_ (.A1(_09250_),
    .A2(_10266_),
    .B(_10306_),
    .Y(_03429_));
 AND2x2_ASAP7_75t_R _26255_ (.A(_04503_),
    .B(_10269_),
    .Y(_10307_));
 AO21x1_ASAP7_75t_R _26256_ (.A1(_09302_),
    .A2(_10266_),
    .B(_10307_),
    .Y(_03430_));
 AND2x2_ASAP7_75t_R _26257_ (.A(_04657_),
    .B(_10269_),
    .Y(_10308_));
 AO21x1_ASAP7_75t_R _26258_ (.A1(_09335_),
    .A2(_10266_),
    .B(_10308_),
    .Y(_03431_));
 NAND2x1_ASAP7_75t_R _26259_ (.A(_01344_),
    .B(_10274_),
    .Y(_10309_));
 OA21x2_ASAP7_75t_R _26260_ (.A1(_10081_),
    .A2(_10274_),
    .B(_10309_),
    .Y(_03432_));
 AND2x2_ASAP7_75t_R _26261_ (.A(_04856_),
    .B(_10269_),
    .Y(_10310_));
 AO21x1_ASAP7_75t_R _26262_ (.A1(_09810_),
    .A2(_10266_),
    .B(_10310_),
    .Y(_03433_));
 NAND2x1_ASAP7_75t_R _26263_ (.A(_01765_),
    .B(_09870_),
    .Y(_10311_));
 OA21x2_ASAP7_75t_R _26264_ (.A1(_09614_),
    .A2(_09897_),
    .B(_10311_),
    .Y(_03434_));
 NOR2x2_ASAP7_75t_R _26265_ (.A(_09506_),
    .B(_10132_),
    .Y(_10312_));
 BUFx12f_ASAP7_75t_R _26266_ (.A(_10312_),
    .Y(_10313_));
 OR2x6_ASAP7_75t_R _26267_ (.A(_09506_),
    .B(_10132_),
    .Y(_10314_));
 BUFx12f_ASAP7_75t_R _26268_ (.A(_10314_),
    .Y(_10315_));
 AND2x2_ASAP7_75t_R _26269_ (.A(_00399_),
    .B(_10315_),
    .Y(_10316_));
 AOI21x1_ASAP7_75t_R _26270_ (.A1(_09902_),
    .A2(_10313_),
    .B(_10316_),
    .Y(_03435_));
 AND2x2_ASAP7_75t_R _26271_ (.A(_00432_),
    .B(_10315_),
    .Y(_10317_));
 AOI21x1_ASAP7_75t_R _26272_ (.A1(_09908_),
    .A2(_10313_),
    .B(_10317_),
    .Y(_03436_));
 BUFx6f_ASAP7_75t_R _26273_ (.A(_10315_),
    .Y(_10318_));
 AND2x2_ASAP7_75t_R _26274_ (.A(_09543_),
    .B(_10312_),
    .Y(_10319_));
 AOI21x1_ASAP7_75t_R _26275_ (.A1(_00463_),
    .A2(_10318_),
    .B(_10319_),
    .Y(_03437_));
 BUFx12f_ASAP7_75t_R _26276_ (.A(_10312_),
    .Y(_10320_));
 NOR2x1_ASAP7_75t_R _26277_ (.A(_00493_),
    .B(_10320_),
    .Y(_10321_));
 AO21x1_ASAP7_75t_R _26278_ (.A1(_09819_),
    .A2(_10313_),
    .B(_10321_),
    .Y(_03438_));
 BUFx12f_ASAP7_75t_R _26279_ (.A(_10314_),
    .Y(_10322_));
 NAND2x1_ASAP7_75t_R _26280_ (.A(_00523_),
    .B(_10322_),
    .Y(_10323_));
 OA21x2_ASAP7_75t_R _26281_ (.A1(_09563_),
    .A2(_10318_),
    .B(_10323_),
    .Y(_03439_));
 AND2x2_ASAP7_75t_R _26282_ (.A(_13778_),
    .B(_10315_),
    .Y(_10324_));
 AO21x1_ASAP7_75t_R _26283_ (.A1(_09268_),
    .A2(_10313_),
    .B(_10324_),
    .Y(_03440_));
 NAND2x1_ASAP7_75t_R _26284_ (.A(_00583_),
    .B(_10322_),
    .Y(_10325_));
 OA21x2_ASAP7_75t_R _26285_ (.A1(_09567_),
    .A2(_10318_),
    .B(_10325_),
    .Y(_03441_));
 NOR2x1_ASAP7_75t_R _26286_ (.A(_00613_),
    .B(_10320_),
    .Y(_10326_));
 AO21x1_ASAP7_75t_R _26287_ (.A1(_09436_),
    .A2(_10313_),
    .B(_10326_),
    .Y(_03442_));
 NAND2x1_ASAP7_75t_R _26288_ (.A(_00643_),
    .B(_10322_),
    .Y(_10327_));
 OA21x2_ASAP7_75t_R _26289_ (.A1(_09438_),
    .A2(_10318_),
    .B(_10327_),
    .Y(_03443_));
 NAND2x1_ASAP7_75t_R _26290_ (.A(_00673_),
    .B(_10322_),
    .Y(_10328_));
 OA21x2_ASAP7_75t_R _26291_ (.A1(_09441_),
    .A2(_10318_),
    .B(_10328_),
    .Y(_03444_));
 BUFx12f_ASAP7_75t_R _26292_ (.A(_09502_),
    .Y(_10329_));
 AND2x6_ASAP7_75t_R _26293_ (.A(_08950_),
    .B(_09667_),
    .Y(_10330_));
 NAND2x2_ASAP7_75t_R _26294_ (.A(_08950_),
    .B(_09666_),
    .Y(_10331_));
 BUFx12f_ASAP7_75t_R _26295_ (.A(_10331_),
    .Y(_10332_));
 AND2x2_ASAP7_75t_R _26296_ (.A(_00381_),
    .B(_10332_),
    .Y(_10333_));
 AOI21x1_ASAP7_75t_R _26297_ (.A1(_10329_),
    .A2(_10330_),
    .B(_10333_),
    .Y(_03445_));
 BUFx12f_ASAP7_75t_R _26298_ (.A(_10315_),
    .Y(_10334_));
 NAND2x1_ASAP7_75t_R _26299_ (.A(_00703_),
    .B(_10334_),
    .Y(_10335_));
 OA21x2_ASAP7_75t_R _26300_ (.A1(_09443_),
    .A2(_10318_),
    .B(_10335_),
    .Y(_03446_));
 AND2x2_ASAP7_75t_R _26301_ (.A(_14204_),
    .B(_10315_),
    .Y(_10336_));
 AO21x1_ASAP7_75t_R _26302_ (.A1(_10286_),
    .A2(_10313_),
    .B(_10336_),
    .Y(_03447_));
 NAND2x1_ASAP7_75t_R _26303_ (.A(_00363_),
    .B(_10334_),
    .Y(_10337_));
 OA21x2_ASAP7_75t_R _26304_ (.A1(_09447_),
    .A2(_10318_),
    .B(_10337_),
    .Y(_03448_));
 NOR2x1_ASAP7_75t_R _26305_ (.A(_00801_),
    .B(_10320_),
    .Y(_10338_));
 AO21x1_ASAP7_75t_R _26306_ (.A1(_10244_),
    .A2(_10313_),
    .B(_10338_),
    .Y(_03449_));
 AND2x2_ASAP7_75t_R _26307_ (.A(_00833_),
    .B(_10315_),
    .Y(_10339_));
 AOI21x1_ASAP7_75t_R _26308_ (.A1(_09790_),
    .A2(_10313_),
    .B(_10339_),
    .Y(_03450_));
 NAND2x1_ASAP7_75t_R _26309_ (.A(_00865_),
    .B(_10334_),
    .Y(_10340_));
 OA21x2_ASAP7_75t_R _26310_ (.A1(_10019_),
    .A2(_10318_),
    .B(_10340_),
    .Y(_03451_));
 NAND2x1_ASAP7_75t_R _26311_ (.A(_00897_),
    .B(_10334_),
    .Y(_10341_));
 OA21x2_ASAP7_75t_R _26312_ (.A1(_09455_),
    .A2(_10318_),
    .B(_10341_),
    .Y(_03452_));
 AND2x2_ASAP7_75t_R _26313_ (.A(_00929_),
    .B(_10315_),
    .Y(_10342_));
 AOI21x1_ASAP7_75t_R _26314_ (.A1(_08948_),
    .A2(_10313_),
    .B(_10342_),
    .Y(_03453_));
 NAND2x1_ASAP7_75t_R _26315_ (.A(_00961_),
    .B(_10334_),
    .Y(_10343_));
 OA21x2_ASAP7_75t_R _26316_ (.A1(_09587_),
    .A2(_10318_),
    .B(_10343_),
    .Y(_03454_));
 NAND2x1_ASAP7_75t_R _26317_ (.A(_00993_),
    .B(_10334_),
    .Y(_10344_));
 OA21x2_ASAP7_75t_R _26318_ (.A1(_09589_),
    .A2(_10322_),
    .B(_10344_),
    .Y(_03455_));
 BUFx12f_ASAP7_75t_R _26319_ (.A(_09526_),
    .Y(_10345_));
 AND2x2_ASAP7_75t_R _26320_ (.A(_00414_),
    .B(_10332_),
    .Y(_10346_));
 AOI21x1_ASAP7_75t_R _26321_ (.A1(_10345_),
    .A2(_10330_),
    .B(_10346_),
    .Y(_03456_));
 NAND2x1_ASAP7_75t_R _26322_ (.A(_01025_),
    .B(_10334_),
    .Y(_10347_));
 OA21x2_ASAP7_75t_R _26323_ (.A1(_09592_),
    .A2(_10322_),
    .B(_10347_),
    .Y(_03457_));
 NOR2x1_ASAP7_75t_R _26324_ (.A(_01057_),
    .B(_10320_),
    .Y(_10348_));
 AO21x1_ASAP7_75t_R _26325_ (.A1(_09100_),
    .A2(_10313_),
    .B(_10348_),
    .Y(_03458_));
 NOR2x1_ASAP7_75t_R _26326_ (.A(_01089_),
    .B(_10312_),
    .Y(_10349_));
 AO21x1_ASAP7_75t_R _26327_ (.A1(_09124_),
    .A2(_10320_),
    .B(_10349_),
    .Y(_03459_));
 NOR2x1_ASAP7_75t_R _26328_ (.A(_01121_),
    .B(_10312_),
    .Y(_10350_));
 AO21x1_ASAP7_75t_R _26329_ (.A1(_09145_),
    .A2(_10320_),
    .B(_10350_),
    .Y(_03460_));
 NAND2x1_ASAP7_75t_R _26330_ (.A(_01153_),
    .B(_10334_),
    .Y(_10351_));
 OA21x2_ASAP7_75t_R _26331_ (.A1(_09600_),
    .A2(_10322_),
    .B(_10351_),
    .Y(_03461_));
 NAND2x1_ASAP7_75t_R _26332_ (.A(_01185_),
    .B(_10334_),
    .Y(_10352_));
 OA21x2_ASAP7_75t_R _26333_ (.A1(_09602_),
    .A2(_10322_),
    .B(_10352_),
    .Y(_03462_));
 NOR2x1_ASAP7_75t_R _26334_ (.A(_01217_),
    .B(_10312_),
    .Y(_10353_));
 AO21x1_ASAP7_75t_R _26335_ (.A1(_09230_),
    .A2(_10320_),
    .B(_10353_),
    .Y(_03463_));
 NOR2x1_ASAP7_75t_R _26336_ (.A(_01249_),
    .B(_10312_),
    .Y(_10354_));
 AO21x1_ASAP7_75t_R _26337_ (.A1(_09250_),
    .A2(_10320_),
    .B(_10354_),
    .Y(_03464_));
 NOR2x1_ASAP7_75t_R _26338_ (.A(_01281_),
    .B(_10312_),
    .Y(_10355_));
 AO21x1_ASAP7_75t_R _26339_ (.A1(_09302_),
    .A2(_10320_),
    .B(_10355_),
    .Y(_03465_));
 NAND2x1_ASAP7_75t_R _26340_ (.A(_01313_),
    .B(_10334_),
    .Y(_10356_));
 OA21x2_ASAP7_75t_R _26341_ (.A1(_09610_),
    .A2(_10322_),
    .B(_10356_),
    .Y(_03466_));
 BUFx12f_ASAP7_75t_R _26342_ (.A(_10331_),
    .Y(_10357_));
 NOR2x1_ASAP7_75t_R _26343_ (.A(_09898_),
    .B(_10332_),
    .Y(_10358_));
 AO21x1_ASAP7_75t_R _26344_ (.A1(_13554_),
    .A2(_10357_),
    .B(_10358_),
    .Y(_03467_));
 NAND2x1_ASAP7_75t_R _26345_ (.A(_01345_),
    .B(_10315_),
    .Y(_10359_));
 OA21x2_ASAP7_75t_R _26346_ (.A1(_10081_),
    .A2(_10322_),
    .B(_10359_),
    .Y(_03468_));
 AND2x2_ASAP7_75t_R _26347_ (.A(_04851_),
    .B(_10315_),
    .Y(_10360_));
 AO21x1_ASAP7_75t_R _26348_ (.A1(_09393_),
    .A2(_10320_),
    .B(_10360_),
    .Y(_03469_));
 NOR2x2_ASAP7_75t_R _26349_ (.A(_09506_),
    .B(_10176_),
    .Y(_10361_));
 BUFx6f_ASAP7_75t_R _26350_ (.A(_10361_),
    .Y(_10362_));
 OR2x6_ASAP7_75t_R _26351_ (.A(_09506_),
    .B(_10176_),
    .Y(_10363_));
 BUFx12f_ASAP7_75t_R _26352_ (.A(_10363_),
    .Y(_10364_));
 AND2x2_ASAP7_75t_R _26353_ (.A(_00400_),
    .B(_10364_),
    .Y(_10365_));
 AOI21x1_ASAP7_75t_R _26354_ (.A1(_10329_),
    .A2(_10362_),
    .B(_10365_),
    .Y(_03470_));
 AND2x2_ASAP7_75t_R _26355_ (.A(_00433_),
    .B(_10364_),
    .Y(_10366_));
 AOI21x1_ASAP7_75t_R _26356_ (.A1(_10345_),
    .A2(_10362_),
    .B(_10366_),
    .Y(_03471_));
 AND2x2_ASAP7_75t_R _26357_ (.A(_09543_),
    .B(_10361_),
    .Y(_10367_));
 AOI21x1_ASAP7_75t_R _26358_ (.A1(_00464_),
    .A2(_10364_),
    .B(_10367_),
    .Y(_03472_));
 BUFx12f_ASAP7_75t_R _26359_ (.A(_10361_),
    .Y(_10368_));
 NOR2x1_ASAP7_75t_R _26360_ (.A(_00494_),
    .B(_10368_),
    .Y(_10369_));
 AO21x1_ASAP7_75t_R _26361_ (.A1(_09560_),
    .A2(_10362_),
    .B(_10369_),
    .Y(_03473_));
 AND2x2_ASAP7_75t_R _26362_ (.A(_13726_),
    .B(_10364_),
    .Y(_10370_));
 AO21x1_ASAP7_75t_R _26363_ (.A1(_08993_),
    .A2(_10362_),
    .B(_10370_),
    .Y(_03474_));
 NOR2x1_ASAP7_75t_R _26364_ (.A(_00554_),
    .B(_10368_),
    .Y(_10371_));
 AO21x1_ASAP7_75t_R _26365_ (.A1(_09268_),
    .A2(_10362_),
    .B(_10371_),
    .Y(_03475_));
 NOR2x1_ASAP7_75t_R _26366_ (.A(_00584_),
    .B(_10368_),
    .Y(_10372_));
 AO21x1_ASAP7_75t_R _26367_ (.A1(_09412_),
    .A2(_10362_),
    .B(_10372_),
    .Y(_03476_));
 BUFx12f_ASAP7_75t_R _26368_ (.A(_10361_),
    .Y(_10373_));
 NOR2x1_ASAP7_75t_R _26369_ (.A(_00614_),
    .B(_10373_),
    .Y(_10374_));
 AO21x1_ASAP7_75t_R _26370_ (.A1(_09436_),
    .A2(_10362_),
    .B(_10374_),
    .Y(_03477_));
 BUFx6f_ASAP7_75t_R _26371_ (.A(_10332_),
    .Y(_10375_));
 NAND2x1_ASAP7_75t_R _26372_ (.A(_00475_),
    .B(_10357_),
    .Y(_10376_));
 OA21x2_ASAP7_75t_R _26373_ (.A1(_09629_),
    .A2(_10375_),
    .B(_10376_),
    .Y(_03478_));
 NOR2x1_ASAP7_75t_R _26374_ (.A(_00644_),
    .B(_10373_),
    .Y(_10377_));
 AO21x1_ASAP7_75t_R _26375_ (.A1(_10098_),
    .A2(_10362_),
    .B(_10377_),
    .Y(_03479_));
 NOR2x1_ASAP7_75t_R _26376_ (.A(_00674_),
    .B(_10373_),
    .Y(_10378_));
 AO21x1_ASAP7_75t_R _26377_ (.A1(_10282_),
    .A2(_10362_),
    .B(_10378_),
    .Y(_03480_));
 NOR2x1_ASAP7_75t_R _26378_ (.A(_00704_),
    .B(_10373_),
    .Y(_10379_));
 AO21x1_ASAP7_75t_R _26379_ (.A1(_10102_),
    .A2(_10362_),
    .B(_10379_),
    .Y(_03481_));
 BUFx6f_ASAP7_75t_R _26380_ (.A(_10361_),
    .Y(_10380_));
 NOR2x1_ASAP7_75t_R _26381_ (.A(_00734_),
    .B(_10373_),
    .Y(_10381_));
 AO21x1_ASAP7_75t_R _26382_ (.A1(_10286_),
    .A2(_10380_),
    .B(_10381_),
    .Y(_03482_));
 NOR2x1_ASAP7_75t_R _26383_ (.A(_00364_),
    .B(_10373_),
    .Y(_10382_));
 AO21x1_ASAP7_75t_R _26384_ (.A1(_10107_),
    .A2(_10380_),
    .B(_10382_),
    .Y(_03483_));
 NOR2x1_ASAP7_75t_R _26385_ (.A(_00802_),
    .B(_10373_),
    .Y(_10383_));
 AO21x1_ASAP7_75t_R _26386_ (.A1(_10244_),
    .A2(_10380_),
    .B(_10383_),
    .Y(_03484_));
 AND2x2_ASAP7_75t_R _26387_ (.A(_08850_),
    .B(_10361_),
    .Y(_10384_));
 AOI21x1_ASAP7_75t_R _26388_ (.A1(_00834_),
    .A2(_10364_),
    .B(_10384_),
    .Y(_03485_));
 NAND2x1_ASAP7_75t_R _26389_ (.A(_00866_),
    .B(_10364_),
    .Y(_10385_));
 OA21x2_ASAP7_75t_R _26390_ (.A1(_10019_),
    .A2(_10364_),
    .B(_10385_),
    .Y(_03486_));
 NOR2x1_ASAP7_75t_R _26391_ (.A(_00898_),
    .B(_10373_),
    .Y(_10386_));
 AO21x1_ASAP7_75t_R _26392_ (.A1(_09584_),
    .A2(_10380_),
    .B(_10386_),
    .Y(_03487_));
 AND2x2_ASAP7_75t_R _26393_ (.A(_09457_),
    .B(_10361_),
    .Y(_10387_));
 AOI21x1_ASAP7_75t_R _26394_ (.A1(_00930_),
    .A2(_10364_),
    .B(_10387_),
    .Y(_03488_));
 NAND2x1_ASAP7_75t_R _26395_ (.A(_00505_),
    .B(_10357_),
    .Y(_10388_));
 OA21x2_ASAP7_75t_R _26396_ (.A1(_09563_),
    .A2(_10375_),
    .B(_10388_),
    .Y(_03489_));
 NOR2x1_ASAP7_75t_R _26397_ (.A(_00962_),
    .B(_10373_),
    .Y(_10389_));
 AO21x1_ASAP7_75t_R _26398_ (.A1(_09022_),
    .A2(_10380_),
    .B(_10389_),
    .Y(_03490_));
 NOR2x1_ASAP7_75t_R _26399_ (.A(_00994_),
    .B(_10373_),
    .Y(_10390_));
 AO21x1_ASAP7_75t_R _26400_ (.A1(_09049_),
    .A2(_10380_),
    .B(_10390_),
    .Y(_03491_));
 BUFx12f_ASAP7_75t_R _26401_ (.A(_10361_),
    .Y(_10391_));
 NOR2x1_ASAP7_75t_R _26402_ (.A(_01026_),
    .B(_10391_),
    .Y(_10392_));
 AO21x1_ASAP7_75t_R _26403_ (.A1(_09075_),
    .A2(_10380_),
    .B(_10392_),
    .Y(_03492_));
 NOR2x1_ASAP7_75t_R _26404_ (.A(_01058_),
    .B(_10391_),
    .Y(_10393_));
 AO21x1_ASAP7_75t_R _26405_ (.A1(_09100_),
    .A2(_10380_),
    .B(_10393_),
    .Y(_03493_));
 NOR2x1_ASAP7_75t_R _26406_ (.A(_01090_),
    .B(_10391_),
    .Y(_10394_));
 AO21x1_ASAP7_75t_R _26407_ (.A1(_09124_),
    .A2(_10380_),
    .B(_10394_),
    .Y(_03494_));
 NOR2x1_ASAP7_75t_R _26408_ (.A(_01122_),
    .B(_10391_),
    .Y(_10395_));
 AO21x1_ASAP7_75t_R _26409_ (.A1(_09145_),
    .A2(_10380_),
    .B(_10395_),
    .Y(_03495_));
 NOR2x1_ASAP7_75t_R _26410_ (.A(_01154_),
    .B(_10391_),
    .Y(_10396_));
 AO21x1_ASAP7_75t_R _26411_ (.A1(_09177_),
    .A2(_10368_),
    .B(_10396_),
    .Y(_03496_));
 NOR2x1_ASAP7_75t_R _26412_ (.A(_01186_),
    .B(_10391_),
    .Y(_10397_));
 AO21x1_ASAP7_75t_R _26413_ (.A1(_09204_),
    .A2(_10368_),
    .B(_10397_),
    .Y(_03497_));
 NOR2x1_ASAP7_75t_R _26414_ (.A(_01218_),
    .B(_10391_),
    .Y(_10398_));
 AO21x1_ASAP7_75t_R _26415_ (.A1(_09230_),
    .A2(_10368_),
    .B(_10398_),
    .Y(_03498_));
 NOR2x1_ASAP7_75t_R _26416_ (.A(_01250_),
    .B(_10391_),
    .Y(_10399_));
 AO21x1_ASAP7_75t_R _26417_ (.A1(_09250_),
    .A2(_10368_),
    .B(_10399_),
    .Y(_03499_));
 BUFx12f_ASAP7_75t_R _26418_ (.A(_10331_),
    .Y(_10400_));
 NAND2x1_ASAP7_75t_R _26419_ (.A(_00535_),
    .B(_10400_),
    .Y(_10401_));
 OA21x2_ASAP7_75t_R _26420_ (.A1(_09565_),
    .A2(_10375_),
    .B(_10401_),
    .Y(_03500_));
 NOR2x1_ASAP7_75t_R _26421_ (.A(_01282_),
    .B(_10391_),
    .Y(_10402_));
 AO21x1_ASAP7_75t_R _26422_ (.A1(_09302_),
    .A2(_10368_),
    .B(_10402_),
    .Y(_03501_));
 NOR2x1_ASAP7_75t_R _26423_ (.A(_01314_),
    .B(_10391_),
    .Y(_10403_));
 AO21x1_ASAP7_75t_R _26424_ (.A1(_09335_),
    .A2(_10368_),
    .B(_10403_),
    .Y(_03502_));
 NAND2x1_ASAP7_75t_R _26425_ (.A(_01346_),
    .B(_10364_),
    .Y(_10404_));
 OA21x2_ASAP7_75t_R _26426_ (.A1(_10081_),
    .A2(_10364_),
    .B(_10404_),
    .Y(_03503_));
 NOR2x1_ASAP7_75t_R _26427_ (.A(_01378_),
    .B(_10361_),
    .Y(_10405_));
 AO21x1_ASAP7_75t_R _26428_ (.A1(_09393_),
    .A2(_10368_),
    .B(_10405_),
    .Y(_03504_));
 NOR2x2_ASAP7_75t_R _26429_ (.A(_09506_),
    .B(_10221_),
    .Y(_10406_));
 BUFx6f_ASAP7_75t_R _26430_ (.A(_10406_),
    .Y(_10407_));
 OR2x2_ASAP7_75t_R _26431_ (.A(_09506_),
    .B(_10221_),
    .Y(_10408_));
 BUFx6f_ASAP7_75t_R _26432_ (.A(_10408_),
    .Y(_10409_));
 BUFx6f_ASAP7_75t_R _26433_ (.A(_10409_),
    .Y(_10410_));
 AND2x2_ASAP7_75t_R _26434_ (.A(_00401_),
    .B(_10410_),
    .Y(_10411_));
 AOI21x1_ASAP7_75t_R _26435_ (.A1(_10329_),
    .A2(_10407_),
    .B(_10411_),
    .Y(_03505_));
 AND2x2_ASAP7_75t_R _26436_ (.A(_00434_),
    .B(_10410_),
    .Y(_10412_));
 AOI21x1_ASAP7_75t_R _26437_ (.A1(_10345_),
    .A2(_10407_),
    .B(_10412_),
    .Y(_03506_));
 BUFx6f_ASAP7_75t_R _26438_ (.A(_10409_),
    .Y(_10413_));
 NOR2x1_ASAP7_75t_R _26439_ (.A(_09898_),
    .B(_10413_),
    .Y(_10414_));
 AO21x1_ASAP7_75t_R _26440_ (.A1(_13574_),
    .A2(_10413_),
    .B(_10414_),
    .Y(_03507_));
 AND2x2_ASAP7_75t_R _26441_ (.A(_13620_),
    .B(_10410_),
    .Y(_10415_));
 AO21x1_ASAP7_75t_R _26442_ (.A1(_09560_),
    .A2(_10407_),
    .B(_10415_),
    .Y(_03508_));
 AND2x2_ASAP7_75t_R _26443_ (.A(_13729_),
    .B(_10410_),
    .Y(_10416_));
 AO21x1_ASAP7_75t_R _26444_ (.A1(_08993_),
    .A2(_10407_),
    .B(_10416_),
    .Y(_03509_));
 AND2x2_ASAP7_75t_R _26445_ (.A(_14872_),
    .B(_10410_),
    .Y(_10417_));
 AO21x1_ASAP7_75t_R _26446_ (.A1(_09268_),
    .A2(_10407_),
    .B(_10417_),
    .Y(_03510_));
 AND2x2_ASAP7_75t_R _26447_ (.A(_13878_),
    .B(_10332_),
    .Y(_10418_));
 AO21x1_ASAP7_75t_R _26448_ (.A1(_09412_),
    .A2(_10330_),
    .B(_10418_),
    .Y(_03511_));
 AND2x2_ASAP7_75t_R _26449_ (.A(_13892_),
    .B(_10410_),
    .Y(_10419_));
 AO21x1_ASAP7_75t_R _26450_ (.A1(_09412_),
    .A2(_10407_),
    .B(_10419_),
    .Y(_03512_));
 AND2x2_ASAP7_75t_R _26451_ (.A(_13955_),
    .B(_10410_),
    .Y(_10420_));
 AO21x1_ASAP7_75t_R _26452_ (.A1(_09436_),
    .A2(_10407_),
    .B(_10420_),
    .Y(_03513_));
 AND2x2_ASAP7_75t_R _26453_ (.A(_14020_),
    .B(_10410_),
    .Y(_10421_));
 AO21x1_ASAP7_75t_R _26454_ (.A1(_10098_),
    .A2(_10407_),
    .B(_10421_),
    .Y(_03514_));
 AND2x2_ASAP7_75t_R _26455_ (.A(_14039_),
    .B(_10410_),
    .Y(_10422_));
 AO21x1_ASAP7_75t_R _26456_ (.A1(_10282_),
    .A2(_10407_),
    .B(_10422_),
    .Y(_03515_));
 BUFx6f_ASAP7_75t_R _26457_ (.A(_10409_),
    .Y(_10423_));
 AND2x2_ASAP7_75t_R _26458_ (.A(_14155_),
    .B(_10423_),
    .Y(_10424_));
 AO21x1_ASAP7_75t_R _26459_ (.A1(_10102_),
    .A2(_10407_),
    .B(_10424_),
    .Y(_03516_));
 BUFx6f_ASAP7_75t_R _26460_ (.A(_10406_),
    .Y(_10425_));
 AND2x2_ASAP7_75t_R _26461_ (.A(_14343_),
    .B(_10423_),
    .Y(_10426_));
 AO21x1_ASAP7_75t_R _26462_ (.A1(_10286_),
    .A2(_10425_),
    .B(_10426_),
    .Y(_03517_));
 AND2x2_ASAP7_75t_R _26463_ (.A(_13171_),
    .B(_10423_),
    .Y(_10427_));
 AO21x1_ASAP7_75t_R _26464_ (.A1(_10107_),
    .A2(_10425_),
    .B(_10427_),
    .Y(_03518_));
 AND2x2_ASAP7_75t_R _26465_ (.A(_15402_),
    .B(_10423_),
    .Y(_10428_));
 AO21x1_ASAP7_75t_R _26466_ (.A1(_10244_),
    .A2(_10425_),
    .B(_10428_),
    .Y(_03519_));
 NOR2x1_ASAP7_75t_R _26467_ (.A(_08851_),
    .B(_10413_),
    .Y(_10429_));
 AO21x1_ASAP7_75t_R _26468_ (.A1(_15555_),
    .A2(_10413_),
    .B(_10429_),
    .Y(_03520_));
 BUFx6f_ASAP7_75t_R _26469_ (.A(_08892_),
    .Y(_10430_));
 NAND2x1_ASAP7_75t_R _26470_ (.A(_00867_),
    .B(_10413_),
    .Y(_10431_));
 OA21x2_ASAP7_75t_R _26471_ (.A1(_10430_),
    .A2(_10413_),
    .B(_10431_),
    .Y(_03521_));
 NAND2x1_ASAP7_75t_R _26472_ (.A(_00595_),
    .B(_10400_),
    .Y(_10432_));
 OA21x2_ASAP7_75t_R _26473_ (.A1(_09570_),
    .A2(_10375_),
    .B(_10432_),
    .Y(_03522_));
 AND2x2_ASAP7_75t_R _26474_ (.A(_09930_),
    .B(_10406_),
    .Y(_10433_));
 AO21x1_ASAP7_75t_R _26475_ (.A1(_15791_),
    .A2(_10413_),
    .B(_10433_),
    .Y(_03523_));
 NOR2x1_ASAP7_75t_R _26476_ (.A(_09695_),
    .B(_10410_),
    .Y(_10434_));
 AO21x1_ASAP7_75t_R _26477_ (.A1(_15916_),
    .A2(_10413_),
    .B(_10434_),
    .Y(_03524_));
 AND2x2_ASAP7_75t_R _26478_ (.A(_16038_),
    .B(_10423_),
    .Y(_10435_));
 AO21x1_ASAP7_75t_R _26479_ (.A1(_09022_),
    .A2(_10425_),
    .B(_10435_),
    .Y(_03525_));
 AND2x2_ASAP7_75t_R _26480_ (.A(_16163_),
    .B(_10423_),
    .Y(_10436_));
 AO21x1_ASAP7_75t_R _26481_ (.A1(_09049_),
    .A2(_10425_),
    .B(_10436_),
    .Y(_03526_));
 AND2x2_ASAP7_75t_R _26482_ (.A(_16298_),
    .B(_10423_),
    .Y(_10437_));
 AO21x1_ASAP7_75t_R _26483_ (.A1(_09075_),
    .A2(_10425_),
    .B(_10437_),
    .Y(_03527_));
 AND2x2_ASAP7_75t_R _26484_ (.A(_16421_),
    .B(_10423_),
    .Y(_10438_));
 AO21x1_ASAP7_75t_R _26485_ (.A1(_09100_),
    .A2(_10425_),
    .B(_10438_),
    .Y(_03528_));
 AND2x2_ASAP7_75t_R _26486_ (.A(_16559_),
    .B(_10423_),
    .Y(_10439_));
 AO21x1_ASAP7_75t_R _26487_ (.A1(_09124_),
    .A2(_10425_),
    .B(_10439_),
    .Y(_03529_));
 AND2x2_ASAP7_75t_R _26488_ (.A(_16669_),
    .B(_10423_),
    .Y(_10440_));
 AO21x1_ASAP7_75t_R _26489_ (.A1(_09145_),
    .A2(_10425_),
    .B(_10440_),
    .Y(_03530_));
 AND2x2_ASAP7_75t_R _26490_ (.A(_16792_),
    .B(_10409_),
    .Y(_10441_));
 AO21x1_ASAP7_75t_R _26491_ (.A1(_09177_),
    .A2(_10425_),
    .B(_10441_),
    .Y(_03531_));
 AND2x2_ASAP7_75t_R _26492_ (.A(_16891_),
    .B(_10409_),
    .Y(_10442_));
 AO21x1_ASAP7_75t_R _26493_ (.A1(_09204_),
    .A2(_10406_),
    .B(_10442_),
    .Y(_03532_));
 NAND2x1_ASAP7_75t_R _26494_ (.A(_00625_),
    .B(_10400_),
    .Y(_10443_));
 OA21x2_ASAP7_75t_R _26495_ (.A1(_09438_),
    .A2(_10375_),
    .B(_10443_),
    .Y(_03533_));
 AND2x2_ASAP7_75t_R _26496_ (.A(_04277_),
    .B(_10409_),
    .Y(_10444_));
 AO21x1_ASAP7_75t_R _26497_ (.A1(_09230_),
    .A2(_10406_),
    .B(_10444_),
    .Y(_03534_));
 AND2x2_ASAP7_75t_R _26498_ (.A(_04390_),
    .B(_10409_),
    .Y(_10445_));
 AO21x1_ASAP7_75t_R _26499_ (.A1(_09250_),
    .A2(_10406_),
    .B(_10445_),
    .Y(_03535_));
 AND2x2_ASAP7_75t_R _26500_ (.A(_04514_),
    .B(_10409_),
    .Y(_10446_));
 AO21x1_ASAP7_75t_R _26501_ (.A1(_09302_),
    .A2(_10406_),
    .B(_10446_),
    .Y(_03536_));
 AND2x2_ASAP7_75t_R _26502_ (.A(_04638_),
    .B(_10409_),
    .Y(_10447_));
 AO21x1_ASAP7_75t_R _26503_ (.A1(_09335_),
    .A2(_10406_),
    .B(_10447_),
    .Y(_03537_));
 NAND2x1_ASAP7_75t_R _26504_ (.A(_01347_),
    .B(_10413_),
    .Y(_10448_));
 OA21x2_ASAP7_75t_R _26505_ (.A1(_10081_),
    .A2(_10413_),
    .B(_10448_),
    .Y(_03538_));
 INVx1_ASAP7_75t_R _26506_ (.A(_01379_),
    .Y(_10449_));
 AND2x2_ASAP7_75t_R _26507_ (.A(_10449_),
    .B(_10409_),
    .Y(_10450_));
 AO21x1_ASAP7_75t_R _26508_ (.A1(_09393_),
    .A2(_10406_),
    .B(_10450_),
    .Y(_03539_));
 NOR2x2_ASAP7_75t_R _26509_ (.A(_08263_),
    .B(_09506_),
    .Y(_10451_));
 BUFx6f_ASAP7_75t_R _26510_ (.A(_10451_),
    .Y(_10452_));
 OR2x2_ASAP7_75t_R _26511_ (.A(_08263_),
    .B(_09506_),
    .Y(_10453_));
 BUFx6f_ASAP7_75t_R _26512_ (.A(_10453_),
    .Y(_10454_));
 BUFx6f_ASAP7_75t_R _26513_ (.A(_10454_),
    .Y(_10455_));
 AND2x2_ASAP7_75t_R _26514_ (.A(_00402_),
    .B(_10455_),
    .Y(_10456_));
 AOI21x1_ASAP7_75t_R _26515_ (.A1(_10329_),
    .A2(_10452_),
    .B(_10456_),
    .Y(_03540_));
 AND2x2_ASAP7_75t_R _26516_ (.A(_00435_),
    .B(_10455_),
    .Y(_10457_));
 AOI21x1_ASAP7_75t_R _26517_ (.A1(_10345_),
    .A2(_10452_),
    .B(_10457_),
    .Y(_03541_));
 BUFx6f_ASAP7_75t_R _26518_ (.A(_10454_),
    .Y(_10458_));
 NOR2x1_ASAP7_75t_R _26519_ (.A(_09543_),
    .B(_10458_),
    .Y(_10459_));
 AO21x1_ASAP7_75t_R _26520_ (.A1(_13571_),
    .A2(_10458_),
    .B(_10459_),
    .Y(_03542_));
 AND2x2_ASAP7_75t_R _26521_ (.A(_13627_),
    .B(_10455_),
    .Y(_10460_));
 AO21x1_ASAP7_75t_R _26522_ (.A1(_09560_),
    .A2(_10452_),
    .B(_10460_),
    .Y(_03543_));
 NAND2x1_ASAP7_75t_R _26523_ (.A(_00655_),
    .B(_10400_),
    .Y(_10461_));
 OA21x2_ASAP7_75t_R _26524_ (.A1(_09441_),
    .A2(_10375_),
    .B(_10461_),
    .Y(_03544_));
 AND2x2_ASAP7_75t_R _26525_ (.A(_14809_),
    .B(_10455_),
    .Y(_10462_));
 AO21x1_ASAP7_75t_R _26526_ (.A1(_08993_),
    .A2(_10452_),
    .B(_10462_),
    .Y(_03545_));
 AND2x2_ASAP7_75t_R _26527_ (.A(_13781_),
    .B(_10455_),
    .Y(_10463_));
 AO21x1_ASAP7_75t_R _26528_ (.A1(_09268_),
    .A2(_10452_),
    .B(_10463_),
    .Y(_03546_));
 AND2x2_ASAP7_75t_R _26529_ (.A(_14937_),
    .B(_10455_),
    .Y(_10464_));
 AO21x1_ASAP7_75t_R _26530_ (.A1(_09412_),
    .A2(_10452_),
    .B(_10464_),
    .Y(_03547_));
 AND2x2_ASAP7_75t_R _26531_ (.A(_13962_),
    .B(_10455_),
    .Y(_10465_));
 AO21x1_ASAP7_75t_R _26532_ (.A1(_09436_),
    .A2(_10452_),
    .B(_10465_),
    .Y(_03548_));
 AND2x2_ASAP7_75t_R _26533_ (.A(_14017_),
    .B(_10455_),
    .Y(_10466_));
 AO21x1_ASAP7_75t_R _26534_ (.A1(_10098_),
    .A2(_10452_),
    .B(_10466_),
    .Y(_03549_));
 AND2x2_ASAP7_75t_R _26535_ (.A(_14036_),
    .B(_10455_),
    .Y(_10467_));
 AO21x1_ASAP7_75t_R _26536_ (.A1(_10282_),
    .A2(_10452_),
    .B(_10467_),
    .Y(_03550_));
 BUFx6f_ASAP7_75t_R _26537_ (.A(_10454_),
    .Y(_10468_));
 AND2x2_ASAP7_75t_R _26538_ (.A(_14152_),
    .B(_10468_),
    .Y(_10469_));
 AO21x1_ASAP7_75t_R _26539_ (.A1(_10102_),
    .A2(_10452_),
    .B(_10469_),
    .Y(_03551_));
 BUFx6f_ASAP7_75t_R _26540_ (.A(_10451_),
    .Y(_10470_));
 AND2x2_ASAP7_75t_R _26541_ (.A(_14207_),
    .B(_10468_),
    .Y(_10471_));
 AO21x1_ASAP7_75t_R _26542_ (.A1(_10286_),
    .A2(_10470_),
    .B(_10471_),
    .Y(_03552_));
 AND2x2_ASAP7_75t_R _26543_ (.A(_13167_),
    .B(_10468_),
    .Y(_10472_));
 AO21x1_ASAP7_75t_R _26544_ (.A1(_10107_),
    .A2(_10470_),
    .B(_10472_),
    .Y(_03553_));
 AND2x2_ASAP7_75t_R _26545_ (.A(_15399_),
    .B(_10468_),
    .Y(_10473_));
 AO21x1_ASAP7_75t_R _26546_ (.A1(_10244_),
    .A2(_10470_),
    .B(_10473_),
    .Y(_03554_));
 NAND2x1_ASAP7_75t_R _26547_ (.A(_00685_),
    .B(_10400_),
    .Y(_10474_));
 OA21x2_ASAP7_75t_R _26548_ (.A1(_09443_),
    .A2(_10375_),
    .B(_10474_),
    .Y(_03555_));
 NOR2x1_ASAP7_75t_R _26549_ (.A(_09451_),
    .B(_10458_),
    .Y(_10475_));
 AO21x1_ASAP7_75t_R _26550_ (.A1(_15552_),
    .A2(_10458_),
    .B(_10475_),
    .Y(_03556_));
 NAND2x1_ASAP7_75t_R _26551_ (.A(_00868_),
    .B(_10458_),
    .Y(_10476_));
 OA21x2_ASAP7_75t_R _26552_ (.A1(_10430_),
    .A2(_10458_),
    .B(_10476_),
    .Y(_03557_));
 AND2x2_ASAP7_75t_R _26553_ (.A(_09930_),
    .B(_10451_),
    .Y(_10477_));
 AO21x1_ASAP7_75t_R _26554_ (.A1(_15788_),
    .A2(_10458_),
    .B(_10477_),
    .Y(_03558_));
 NOR2x1_ASAP7_75t_R _26555_ (.A(_09695_),
    .B(_10455_),
    .Y(_10478_));
 AO21x1_ASAP7_75t_R _26556_ (.A1(_15913_),
    .A2(_10458_),
    .B(_10478_),
    .Y(_03559_));
 AND2x2_ASAP7_75t_R _26557_ (.A(_16035_),
    .B(_10468_),
    .Y(_10479_));
 AO21x1_ASAP7_75t_R _26558_ (.A1(_09022_),
    .A2(_10470_),
    .B(_10479_),
    .Y(_03560_));
 AND2x2_ASAP7_75t_R _26559_ (.A(_16160_),
    .B(_10468_),
    .Y(_10480_));
 AO21x1_ASAP7_75t_R _26560_ (.A1(_09049_),
    .A2(_10470_),
    .B(_10480_),
    .Y(_03561_));
 AND2x2_ASAP7_75t_R _26561_ (.A(_16295_),
    .B(_10468_),
    .Y(_10481_));
 AO21x1_ASAP7_75t_R _26562_ (.A1(_09075_),
    .A2(_10470_),
    .B(_10481_),
    .Y(_03562_));
 AND2x2_ASAP7_75t_R _26563_ (.A(_16418_),
    .B(_10468_),
    .Y(_10482_));
 AO21x1_ASAP7_75t_R _26564_ (.A1(_09100_),
    .A2(_10470_),
    .B(_10482_),
    .Y(_03563_));
 AND2x2_ASAP7_75t_R _26565_ (.A(_16556_),
    .B(_10468_),
    .Y(_10483_));
 AO21x1_ASAP7_75t_R _26566_ (.A1(_09124_),
    .A2(_10470_),
    .B(_10483_),
    .Y(_03564_));
 AND2x2_ASAP7_75t_R _26567_ (.A(_16666_),
    .B(_10468_),
    .Y(_10484_));
 AO21x1_ASAP7_75t_R _26568_ (.A1(_09145_),
    .A2(_10470_),
    .B(_10484_),
    .Y(_03565_));
 NAND2x1_ASAP7_75t_R _26569_ (.A(_00715_),
    .B(_10400_),
    .Y(_10485_));
 OA21x2_ASAP7_75t_R _26570_ (.A1(_09445_),
    .A2(_10375_),
    .B(_10485_),
    .Y(_03566_));
 AND2x2_ASAP7_75t_R _26571_ (.A(_16789_),
    .B(_10454_),
    .Y(_10486_));
 AO21x1_ASAP7_75t_R _26572_ (.A1(_09177_),
    .A2(_10470_),
    .B(_10486_),
    .Y(_03567_));
 AND2x2_ASAP7_75t_R _26573_ (.A(_16888_),
    .B(_10454_),
    .Y(_10487_));
 AO21x1_ASAP7_75t_R _26574_ (.A1(_09204_),
    .A2(_10451_),
    .B(_10487_),
    .Y(_03568_));
 AND2x2_ASAP7_75t_R _26575_ (.A(_04274_),
    .B(_10454_),
    .Y(_10488_));
 AO21x1_ASAP7_75t_R _26576_ (.A1(_09230_),
    .A2(_10451_),
    .B(_10488_),
    .Y(_03569_));
 AND2x2_ASAP7_75t_R _26577_ (.A(_04387_),
    .B(_10454_),
    .Y(_10489_));
 AO21x1_ASAP7_75t_R _26578_ (.A1(_09250_),
    .A2(_10451_),
    .B(_10489_),
    .Y(_03570_));
 AND2x2_ASAP7_75t_R _26579_ (.A(_04511_),
    .B(_10454_),
    .Y(_10490_));
 AO21x1_ASAP7_75t_R _26580_ (.A1(_09302_),
    .A2(_10451_),
    .B(_10490_),
    .Y(_03571_));
 AND2x2_ASAP7_75t_R _26581_ (.A(_04635_),
    .B(_10454_),
    .Y(_10491_));
 AO21x1_ASAP7_75t_R _26582_ (.A1(_09335_),
    .A2(_10451_),
    .B(_10491_),
    .Y(_03572_));
 NAND2x1_ASAP7_75t_R _26583_ (.A(_01348_),
    .B(_10458_),
    .Y(_10492_));
 OA21x2_ASAP7_75t_R _26584_ (.A1(_09366_),
    .A2(_10458_),
    .B(_10492_),
    .Y(_03573_));
 AND2x2_ASAP7_75t_R _26585_ (.A(_04848_),
    .B(_10454_),
    .Y(_10493_));
 AO21x1_ASAP7_75t_R _26586_ (.A1(_09393_),
    .A2(_10451_),
    .B(_10493_),
    .Y(_03574_));
 NOR2x2_ASAP7_75t_R _26587_ (.A(_09770_),
    .B(_10132_),
    .Y(_10494_));
 BUFx6f_ASAP7_75t_R _26588_ (.A(_10494_),
    .Y(_10495_));
 OR2x6_ASAP7_75t_R _26589_ (.A(_09770_),
    .B(_10132_),
    .Y(_10496_));
 BUFx12f_ASAP7_75t_R _26590_ (.A(_10496_),
    .Y(_10497_));
 AND2x2_ASAP7_75t_R _26591_ (.A(_00403_),
    .B(_10497_),
    .Y(_10498_));
 AOI21x1_ASAP7_75t_R _26592_ (.A1(_10329_),
    .A2(_10495_),
    .B(_10498_),
    .Y(_03575_));
 BUFx6f_ASAP7_75t_R _26593_ (.A(_10496_),
    .Y(_10499_));
 AND2x2_ASAP7_75t_R _26594_ (.A(_00436_),
    .B(_10499_),
    .Y(_10500_));
 AOI21x1_ASAP7_75t_R _26595_ (.A1(_10345_),
    .A2(_10495_),
    .B(_10500_),
    .Y(_03576_));
 BUFx6f_ASAP7_75t_R _26596_ (.A(_10332_),
    .Y(_10501_));
 NAND2x1_ASAP7_75t_R _26597_ (.A(_00345_),
    .B(_10400_),
    .Y(_10502_));
 OA21x2_ASAP7_75t_R _26598_ (.A1(_09447_),
    .A2(_10501_),
    .B(_10502_),
    .Y(_03577_));
 AND2x2_ASAP7_75t_R _26599_ (.A(_00467_),
    .B(_10499_),
    .Y(_10503_));
 AOI21x1_ASAP7_75t_R _26600_ (.A1(_09675_),
    .A2(_10495_),
    .B(_10503_),
    .Y(_03578_));
 AND2x2_ASAP7_75t_R _26601_ (.A(_13653_),
    .B(_10499_),
    .Y(_10504_));
 AO21x1_ASAP7_75t_R _26602_ (.A1(_09560_),
    .A2(_10495_),
    .B(_10504_),
    .Y(_03579_));
 AND2x2_ASAP7_75t_R _26603_ (.A(_13743_),
    .B(_10499_),
    .Y(_10505_));
 AO21x1_ASAP7_75t_R _26604_ (.A1(_08993_),
    .A2(_10495_),
    .B(_10505_),
    .Y(_03580_));
 AND2x2_ASAP7_75t_R _26605_ (.A(_13815_),
    .B(_10499_),
    .Y(_10506_));
 AO21x1_ASAP7_75t_R _26606_ (.A1(_09268_),
    .A2(_10495_),
    .B(_10506_),
    .Y(_03581_));
 BUFx12f_ASAP7_75t_R _26607_ (.A(_10496_),
    .Y(_10507_));
 NAND2x1_ASAP7_75t_R _26608_ (.A(_00587_),
    .B(_10497_),
    .Y(_10508_));
 OA21x2_ASAP7_75t_R _26609_ (.A1(_09567_),
    .A2(_10507_),
    .B(_10508_),
    .Y(_03582_));
 NAND2x1_ASAP7_75t_R _26610_ (.A(_00617_),
    .B(_10497_),
    .Y(_10509_));
 OA21x2_ASAP7_75t_R _26611_ (.A1(_09570_),
    .A2(_10507_),
    .B(_10509_),
    .Y(_03583_));
 NAND2x1_ASAP7_75t_R _26612_ (.A(_00647_),
    .B(_10497_),
    .Y(_10510_));
 OA21x2_ASAP7_75t_R _26613_ (.A1(_09438_),
    .A2(_10507_),
    .B(_10510_),
    .Y(_03584_));
 AND2x2_ASAP7_75t_R _26614_ (.A(_14064_),
    .B(_10499_),
    .Y(_10511_));
 AO21x1_ASAP7_75t_R _26615_ (.A1(_10282_),
    .A2(_10495_),
    .B(_10511_),
    .Y(_03585_));
 NAND2x1_ASAP7_75t_R _26616_ (.A(_00707_),
    .B(_10497_),
    .Y(_10512_));
 OA21x2_ASAP7_75t_R _26617_ (.A1(_09443_),
    .A2(_10507_),
    .B(_10512_),
    .Y(_03586_));
 AND2x2_ASAP7_75t_R _26618_ (.A(_14355_),
    .B(_10499_),
    .Y(_10513_));
 AO21x1_ASAP7_75t_R _26619_ (.A1(_10286_),
    .A2(_10495_),
    .B(_10513_),
    .Y(_03587_));
 NAND2x1_ASAP7_75t_R _26620_ (.A(_00783_),
    .B(_10400_),
    .Y(_10514_));
 OA21x2_ASAP7_75t_R _26621_ (.A1(_09449_),
    .A2(_10501_),
    .B(_10514_),
    .Y(_03588_));
 AND2x2_ASAP7_75t_R _26622_ (.A(_13191_),
    .B(_10499_),
    .Y(_10515_));
 AO21x1_ASAP7_75t_R _26623_ (.A1(_10107_),
    .A2(_10495_),
    .B(_10515_),
    .Y(_03589_));
 AND2x2_ASAP7_75t_R _26624_ (.A(_15414_),
    .B(_10499_),
    .Y(_10516_));
 AO21x1_ASAP7_75t_R _26625_ (.A1(_10244_),
    .A2(_10495_),
    .B(_10516_),
    .Y(_03590_));
 NOR2x1_ASAP7_75t_R _26626_ (.A(_09451_),
    .B(_10497_),
    .Y(_10517_));
 AO21x1_ASAP7_75t_R _26627_ (.A1(_15567_),
    .A2(_10507_),
    .B(_10517_),
    .Y(_03591_));
 NAND2x1_ASAP7_75t_R _26628_ (.A(_00869_),
    .B(_10497_),
    .Y(_10518_));
 OA21x2_ASAP7_75t_R _26629_ (.A1(_10430_),
    .A2(_10507_),
    .B(_10518_),
    .Y(_03592_));
 AND2x2_ASAP7_75t_R _26630_ (.A(_09930_),
    .B(_10494_),
    .Y(_10519_));
 AO21x1_ASAP7_75t_R _26631_ (.A1(_15773_),
    .A2(_10507_),
    .B(_10519_),
    .Y(_03593_));
 NOR2x1_ASAP7_75t_R _26632_ (.A(_09457_),
    .B(_10497_),
    .Y(_10520_));
 AO21x1_ASAP7_75t_R _26633_ (.A1(_15928_),
    .A2(_10507_),
    .B(_10520_),
    .Y(_03594_));
 BUFx6f_ASAP7_75t_R _26634_ (.A(_10494_),
    .Y(_10521_));
 AND2x2_ASAP7_75t_R _26635_ (.A(_16020_),
    .B(_10499_),
    .Y(_10522_));
 AO21x1_ASAP7_75t_R _26636_ (.A1(_09022_),
    .A2(_10521_),
    .B(_10522_),
    .Y(_03595_));
 BUFx6f_ASAP7_75t_R _26637_ (.A(_10496_),
    .Y(_10523_));
 AND2x2_ASAP7_75t_R _26638_ (.A(_16175_),
    .B(_10523_),
    .Y(_10524_));
 AO21x1_ASAP7_75t_R _26639_ (.A1(_09049_),
    .A2(_10521_),
    .B(_10524_),
    .Y(_03596_));
 AND2x2_ASAP7_75t_R _26640_ (.A(_16310_),
    .B(_10523_),
    .Y(_10525_));
 AO21x1_ASAP7_75t_R _26641_ (.A1(_09075_),
    .A2(_10521_),
    .B(_10525_),
    .Y(_03597_));
 AND2x2_ASAP7_75t_R _26642_ (.A(_16433_),
    .B(_10523_),
    .Y(_10526_));
 AO21x1_ASAP7_75t_R _26643_ (.A1(_09100_),
    .A2(_10521_),
    .B(_10526_),
    .Y(_03598_));
 AO21x1_ASAP7_75t_R _26644_ (.A1(_08950_),
    .A2(_09667_),
    .B(_00815_),
    .Y(_10527_));
 OAI21x1_ASAP7_75t_R _26645_ (.A1(_09790_),
    .A2(_10375_),
    .B(_10527_),
    .Y(_03599_));
 AND2x2_ASAP7_75t_R _26646_ (.A(_16571_),
    .B(_10523_),
    .Y(_10528_));
 AO21x1_ASAP7_75t_R _26647_ (.A1(_09124_),
    .A2(_10521_),
    .B(_10528_),
    .Y(_03600_));
 AND2x2_ASAP7_75t_R _26648_ (.A(_16681_),
    .B(_10523_),
    .Y(_10529_));
 AO21x1_ASAP7_75t_R _26649_ (.A1(_09145_),
    .A2(_10521_),
    .B(_10529_),
    .Y(_03601_));
 AND2x2_ASAP7_75t_R _26650_ (.A(_16804_),
    .B(_10523_),
    .Y(_10530_));
 AO21x1_ASAP7_75t_R _26651_ (.A1(_09177_),
    .A2(_10521_),
    .B(_10530_),
    .Y(_03602_));
 AND2x2_ASAP7_75t_R _26652_ (.A(_16873_),
    .B(_10523_),
    .Y(_10531_));
 AO21x1_ASAP7_75t_R _26653_ (.A1(_09204_),
    .A2(_10521_),
    .B(_10531_),
    .Y(_03603_));
 AND2x2_ASAP7_75t_R _26654_ (.A(_04289_),
    .B(_10523_),
    .Y(_10532_));
 AO21x1_ASAP7_75t_R _26655_ (.A1(_09230_),
    .A2(_10521_),
    .B(_10532_),
    .Y(_03604_));
 AND2x2_ASAP7_75t_R _26656_ (.A(_04402_),
    .B(_10523_),
    .Y(_10533_));
 AO21x1_ASAP7_75t_R _26657_ (.A1(_09250_),
    .A2(_10521_),
    .B(_10533_),
    .Y(_03605_));
 AND2x2_ASAP7_75t_R _26658_ (.A(_04496_),
    .B(_10523_),
    .Y(_10534_));
 AO21x1_ASAP7_75t_R _26659_ (.A1(_09302_),
    .A2(_10494_),
    .B(_10534_),
    .Y(_03606_));
 AND2x2_ASAP7_75t_R _26660_ (.A(_04650_),
    .B(_10496_),
    .Y(_10535_));
 AO21x1_ASAP7_75t_R _26661_ (.A1(_09335_),
    .A2(_10494_),
    .B(_10535_),
    .Y(_03607_));
 NAND2x1_ASAP7_75t_R _26662_ (.A(_01349_),
    .B(_10497_),
    .Y(_10536_));
 OA21x2_ASAP7_75t_R _26663_ (.A1(_09366_),
    .A2(_10507_),
    .B(_10536_),
    .Y(_03608_));
 NAND2x1_ASAP7_75t_R _26664_ (.A(_01381_),
    .B(_10497_),
    .Y(_10537_));
 OA21x2_ASAP7_75t_R _26665_ (.A1(_09614_),
    .A2(_10507_),
    .B(_10537_),
    .Y(_03609_));
 NAND2x1_ASAP7_75t_R _26666_ (.A(_00847_),
    .B(_10400_),
    .Y(_10538_));
 OA21x2_ASAP7_75t_R _26667_ (.A1(_10430_),
    .A2(_10501_),
    .B(_10538_),
    .Y(_03610_));
 NOR2x2_ASAP7_75t_R _26668_ (.A(_09770_),
    .B(_10176_),
    .Y(_10539_));
 OR2x6_ASAP7_75t_R _26669_ (.A(_09770_),
    .B(_10176_),
    .Y(_10540_));
 BUFx12f_ASAP7_75t_R _26670_ (.A(_10540_),
    .Y(_10541_));
 AND2x2_ASAP7_75t_R _26671_ (.A(_00404_),
    .B(_10541_),
    .Y(_10542_));
 AOI21x1_ASAP7_75t_R _26672_ (.A1(_10329_),
    .A2(_10539_),
    .B(_10542_),
    .Y(_03611_));
 AND2x2_ASAP7_75t_R _26673_ (.A(_00437_),
    .B(_10541_),
    .Y(_10543_));
 AOI21x1_ASAP7_75t_R _26674_ (.A1(_10345_),
    .A2(_10539_),
    .B(_10543_),
    .Y(_03612_));
 AND2x2_ASAP7_75t_R _26675_ (.A(_00468_),
    .B(_10541_),
    .Y(_10544_));
 AOI21x1_ASAP7_75t_R _26676_ (.A1(_09675_),
    .A2(_10539_),
    .B(_10544_),
    .Y(_03613_));
 BUFx6f_ASAP7_75t_R _26677_ (.A(_10541_),
    .Y(_10545_));
 BUFx12f_ASAP7_75t_R _26678_ (.A(_10540_),
    .Y(_10546_));
 NAND2x1_ASAP7_75t_R _26679_ (.A(_00498_),
    .B(_10546_),
    .Y(_10547_));
 OA21x2_ASAP7_75t_R _26680_ (.A1(_09629_),
    .A2(_10545_),
    .B(_10547_),
    .Y(_03614_));
 NAND2x1_ASAP7_75t_R _26681_ (.A(_00528_),
    .B(_10546_),
    .Y(_10548_));
 OA21x2_ASAP7_75t_R _26682_ (.A1(_09563_),
    .A2(_10545_),
    .B(_10548_),
    .Y(_03615_));
 NAND2x1_ASAP7_75t_R _26683_ (.A(_00558_),
    .B(_10546_),
    .Y(_10549_));
 OA21x2_ASAP7_75t_R _26684_ (.A1(_09565_),
    .A2(_10545_),
    .B(_10549_),
    .Y(_03616_));
 NAND2x1_ASAP7_75t_R _26685_ (.A(_00588_),
    .B(_10546_),
    .Y(_10550_));
 OA21x2_ASAP7_75t_R _26686_ (.A1(_09567_),
    .A2(_10545_),
    .B(_10550_),
    .Y(_03617_));
 BUFx12f_ASAP7_75t_R _26687_ (.A(_10540_),
    .Y(_10551_));
 NAND2x1_ASAP7_75t_R _26688_ (.A(_00618_),
    .B(_10551_),
    .Y(_10552_));
 OA21x2_ASAP7_75t_R _26689_ (.A1(_09570_),
    .A2(_10545_),
    .B(_10552_),
    .Y(_03618_));
 NAND2x1_ASAP7_75t_R _26690_ (.A(_00648_),
    .B(_10551_),
    .Y(_10553_));
 OA21x2_ASAP7_75t_R _26691_ (.A1(_09438_),
    .A2(_10545_),
    .B(_10553_),
    .Y(_03619_));
 AND2x2_ASAP7_75t_R _26692_ (.A(_14075_),
    .B(_10541_),
    .Y(_10554_));
 AO21x1_ASAP7_75t_R _26693_ (.A1(_10282_),
    .A2(_10539_),
    .B(_10554_),
    .Y(_03620_));
 NAND2x1_ASAP7_75t_R _26694_ (.A(_00879_),
    .B(_10400_),
    .Y(_10555_));
 OA21x2_ASAP7_75t_R _26695_ (.A1(_09455_),
    .A2(_10501_),
    .B(_10555_),
    .Y(_03621_));
 NAND2x1_ASAP7_75t_R _26696_ (.A(_00708_),
    .B(_10551_),
    .Y(_10556_));
 OA21x2_ASAP7_75t_R _26697_ (.A1(_09443_),
    .A2(_10545_),
    .B(_10556_),
    .Y(_03622_));
 NAND2x1_ASAP7_75t_R _26698_ (.A(_00738_),
    .B(_10551_),
    .Y(_10557_));
 OA21x2_ASAP7_75t_R _26699_ (.A1(_09445_),
    .A2(_10545_),
    .B(_10557_),
    .Y(_03623_));
 NAND2x1_ASAP7_75t_R _26700_ (.A(_00368_),
    .B(_10551_),
    .Y(_10558_));
 OA21x2_ASAP7_75t_R _26701_ (.A1(_09447_),
    .A2(_10545_),
    .B(_10558_),
    .Y(_03624_));
 NAND2x1_ASAP7_75t_R _26702_ (.A(_00806_),
    .B(_10551_),
    .Y(_10559_));
 OA21x2_ASAP7_75t_R _26703_ (.A1(_09449_),
    .A2(_10545_),
    .B(_10559_),
    .Y(_03625_));
 AND2x2_ASAP7_75t_R _26704_ (.A(_00838_),
    .B(_10541_),
    .Y(_10560_));
 AOI21x1_ASAP7_75t_R _26705_ (.A1(_09790_),
    .A2(_10539_),
    .B(_10560_),
    .Y(_03626_));
 BUFx6f_ASAP7_75t_R _26706_ (.A(_10541_),
    .Y(_10561_));
 NAND2x1_ASAP7_75t_R _26707_ (.A(_00870_),
    .B(_10551_),
    .Y(_10562_));
 OA21x2_ASAP7_75t_R _26708_ (.A1(_10430_),
    .A2(_10561_),
    .B(_10562_),
    .Y(_03627_));
 NAND2x1_ASAP7_75t_R _26709_ (.A(_00902_),
    .B(_10551_),
    .Y(_10563_));
 OA21x2_ASAP7_75t_R _26710_ (.A1(_09455_),
    .A2(_10561_),
    .B(_10563_),
    .Y(_03628_));
 AND2x2_ASAP7_75t_R _26711_ (.A(_00934_),
    .B(_10541_),
    .Y(_10564_));
 AOI21x1_ASAP7_75t_R _26712_ (.A1(_08948_),
    .A2(_10539_),
    .B(_10564_),
    .Y(_03629_));
 NAND2x1_ASAP7_75t_R _26713_ (.A(_00966_),
    .B(_10551_),
    .Y(_10565_));
 OA21x2_ASAP7_75t_R _26714_ (.A1(_09587_),
    .A2(_10561_),
    .B(_10565_),
    .Y(_03630_));
 NAND2x1_ASAP7_75t_R _26715_ (.A(_00998_),
    .B(_10551_),
    .Y(_10566_));
 OA21x2_ASAP7_75t_R _26716_ (.A1(_09589_),
    .A2(_10561_),
    .B(_10566_),
    .Y(_03631_));
 AO21x1_ASAP7_75t_R _26717_ (.A1(_08950_),
    .A2(_09667_),
    .B(_00911_),
    .Y(_10567_));
 OAI21x1_ASAP7_75t_R _26718_ (.A1(_08948_),
    .A2(_10375_),
    .B(_10567_),
    .Y(_03632_));
 BUFx12f_ASAP7_75t_R _26719_ (.A(_10540_),
    .Y(_10568_));
 NAND2x1_ASAP7_75t_R _26720_ (.A(_01030_),
    .B(_10568_),
    .Y(_10569_));
 OA21x2_ASAP7_75t_R _26721_ (.A1(_09592_),
    .A2(_10561_),
    .B(_10569_),
    .Y(_03633_));
 NAND2x1_ASAP7_75t_R _26722_ (.A(_01062_),
    .B(_10568_),
    .Y(_10570_));
 OA21x2_ASAP7_75t_R _26723_ (.A1(_09594_),
    .A2(_10561_),
    .B(_10570_),
    .Y(_03634_));
 NAND2x1_ASAP7_75t_R _26724_ (.A(_01094_),
    .B(_10568_),
    .Y(_10571_));
 OA21x2_ASAP7_75t_R _26725_ (.A1(_09596_),
    .A2(_10561_),
    .B(_10571_),
    .Y(_03635_));
 NAND2x1_ASAP7_75t_R _26726_ (.A(_01126_),
    .B(_10568_),
    .Y(_10572_));
 OA21x2_ASAP7_75t_R _26727_ (.A1(_09598_),
    .A2(_10561_),
    .B(_10572_),
    .Y(_03636_));
 NAND2x1_ASAP7_75t_R _26728_ (.A(_01158_),
    .B(_10568_),
    .Y(_10573_));
 OA21x2_ASAP7_75t_R _26729_ (.A1(_09600_),
    .A2(_10561_),
    .B(_10573_),
    .Y(_03637_));
 NAND2x1_ASAP7_75t_R _26730_ (.A(_01190_),
    .B(_10568_),
    .Y(_10574_));
 OA21x2_ASAP7_75t_R _26731_ (.A1(_09602_),
    .A2(_10561_),
    .B(_10574_),
    .Y(_03638_));
 NAND2x1_ASAP7_75t_R _26732_ (.A(_01222_),
    .B(_10568_),
    .Y(_10575_));
 OA21x2_ASAP7_75t_R _26733_ (.A1(_09604_),
    .A2(_10546_),
    .B(_10575_),
    .Y(_03639_));
 NAND2x1_ASAP7_75t_R _26734_ (.A(_01254_),
    .B(_10568_),
    .Y(_10576_));
 OA21x2_ASAP7_75t_R _26735_ (.A1(_09606_),
    .A2(_10546_),
    .B(_10576_),
    .Y(_03640_));
 NAND2x1_ASAP7_75t_R _26736_ (.A(_01286_),
    .B(_10568_),
    .Y(_10577_));
 OA21x2_ASAP7_75t_R _26737_ (.A1(_09608_),
    .A2(_10546_),
    .B(_10577_),
    .Y(_03641_));
 NAND2x1_ASAP7_75t_R _26738_ (.A(_01318_),
    .B(_10568_),
    .Y(_10578_));
 OA21x2_ASAP7_75t_R _26739_ (.A1(_09610_),
    .A2(_10546_),
    .B(_10578_),
    .Y(_03642_));
 BUFx12f_ASAP7_75t_R _26740_ (.A(_10331_),
    .Y(_10579_));
 NAND2x1_ASAP7_75t_R _26741_ (.A(_00943_),
    .B(_10579_),
    .Y(_10580_));
 OA21x2_ASAP7_75t_R _26742_ (.A1(_09587_),
    .A2(_10501_),
    .B(_10580_),
    .Y(_03643_));
 NAND2x1_ASAP7_75t_R _26743_ (.A(_01350_),
    .B(_10541_),
    .Y(_10581_));
 OA21x2_ASAP7_75t_R _26744_ (.A1(_09366_),
    .A2(_10546_),
    .B(_10581_),
    .Y(_03644_));
 NAND2x1_ASAP7_75t_R _26745_ (.A(_01382_),
    .B(_10541_),
    .Y(_10582_));
 OA21x2_ASAP7_75t_R _26746_ (.A1(_09614_),
    .A2(_10546_),
    .B(_10582_),
    .Y(_03645_));
 NOR2x2_ASAP7_75t_R _26747_ (.A(_09770_),
    .B(_10221_),
    .Y(_10583_));
 BUFx6f_ASAP7_75t_R _26748_ (.A(_10583_),
    .Y(_10584_));
 OR2x2_ASAP7_75t_R _26749_ (.A(_09770_),
    .B(_10221_),
    .Y(_10585_));
 BUFx6f_ASAP7_75t_R _26750_ (.A(_10585_),
    .Y(_10586_));
 BUFx6f_ASAP7_75t_R _26751_ (.A(_10586_),
    .Y(_10587_));
 AND2x2_ASAP7_75t_R _26752_ (.A(_00405_),
    .B(_10587_),
    .Y(_10588_));
 AOI21x1_ASAP7_75t_R _26753_ (.A1(_10329_),
    .A2(_10584_),
    .B(_10588_),
    .Y(_03646_));
 AND2x2_ASAP7_75t_R _26754_ (.A(_00438_),
    .B(_10587_),
    .Y(_10589_));
 AOI21x1_ASAP7_75t_R _26755_ (.A1(_10345_),
    .A2(_10584_),
    .B(_10589_),
    .Y(_03647_));
 BUFx12f_ASAP7_75t_R _26756_ (.A(_10586_),
    .Y(_10590_));
 NOR2x1_ASAP7_75t_R _26757_ (.A(_09543_),
    .B(_10587_),
    .Y(_10591_));
 AO21x1_ASAP7_75t_R _26758_ (.A1(_13592_),
    .A2(_10590_),
    .B(_10591_),
    .Y(_03648_));
 NOR2x1_ASAP7_75t_R _26759_ (.A(_00499_),
    .B(_10583_),
    .Y(_10592_));
 AO21x1_ASAP7_75t_R _26760_ (.A1(_09560_),
    .A2(_10584_),
    .B(_10592_),
    .Y(_03649_));
 NOR2x1_ASAP7_75t_R _26761_ (.A(_00529_),
    .B(_10583_),
    .Y(_10593_));
 AO21x1_ASAP7_75t_R _26762_ (.A1(_08993_),
    .A2(_10584_),
    .B(_10593_),
    .Y(_03650_));
 BUFx6f_ASAP7_75t_R _26763_ (.A(_10586_),
    .Y(_10594_));
 NAND2x1_ASAP7_75t_R _26764_ (.A(_00559_),
    .B(_10590_),
    .Y(_10595_));
 OA21x2_ASAP7_75t_R _26765_ (.A1(_09565_),
    .A2(_10594_),
    .B(_10595_),
    .Y(_03651_));
 AND2x2_ASAP7_75t_R _26766_ (.A(_14959_),
    .B(_10587_),
    .Y(_10596_));
 AO21x1_ASAP7_75t_R _26767_ (.A1(_09412_),
    .A2(_10584_),
    .B(_10596_),
    .Y(_03652_));
 AND2x2_ASAP7_75t_R _26768_ (.A(_15018_),
    .B(_10587_),
    .Y(_10597_));
 AO21x1_ASAP7_75t_R _26769_ (.A1(_09436_),
    .A2(_10584_),
    .B(_10597_),
    .Y(_03653_));
 NAND2x1_ASAP7_75t_R _26770_ (.A(_00975_),
    .B(_10579_),
    .Y(_10598_));
 OA21x2_ASAP7_75t_R _26771_ (.A1(_09589_),
    .A2(_10501_),
    .B(_10598_),
    .Y(_03654_));
 AND2x2_ASAP7_75t_R _26772_ (.A(_13977_),
    .B(_10587_),
    .Y(_10599_));
 AO21x1_ASAP7_75t_R _26773_ (.A1(_10098_),
    .A2(_10584_),
    .B(_10599_),
    .Y(_03655_));
 NAND2x1_ASAP7_75t_R _26774_ (.A(_00679_),
    .B(_10590_),
    .Y(_10600_));
 OA21x2_ASAP7_75t_R _26775_ (.A1(_09441_),
    .A2(_10594_),
    .B(_10600_),
    .Y(_03656_));
 AND2x2_ASAP7_75t_R _26776_ (.A(_14148_),
    .B(_10587_),
    .Y(_10601_));
 AO21x1_ASAP7_75t_R _26777_ (.A1(_10102_),
    .A2(_10584_),
    .B(_10601_),
    .Y(_03657_));
 NAND2x1_ASAP7_75t_R _26778_ (.A(_00739_),
    .B(_10590_),
    .Y(_10602_));
 OA21x2_ASAP7_75t_R _26779_ (.A1(_09445_),
    .A2(_10594_),
    .B(_10602_),
    .Y(_03658_));
 NAND2x1_ASAP7_75t_R _26780_ (.A(_00369_),
    .B(_10590_),
    .Y(_10603_));
 OA21x2_ASAP7_75t_R _26781_ (.A1(_09447_),
    .A2(_10594_),
    .B(_10603_),
    .Y(_03659_));
 NAND2x1_ASAP7_75t_R _26782_ (.A(_00807_),
    .B(_10590_),
    .Y(_10604_));
 OA21x2_ASAP7_75t_R _26783_ (.A1(_09449_),
    .A2(_10594_),
    .B(_10604_),
    .Y(_03660_));
 AND2x2_ASAP7_75t_R _26784_ (.A(_00839_),
    .B(_10587_),
    .Y(_10605_));
 AOI21x1_ASAP7_75t_R _26785_ (.A1(_09790_),
    .A2(_10584_),
    .B(_10605_),
    .Y(_03661_));
 NAND2x1_ASAP7_75t_R _26786_ (.A(_00871_),
    .B(_10590_),
    .Y(_10606_));
 OA21x2_ASAP7_75t_R _26787_ (.A1(_10430_),
    .A2(_10594_),
    .B(_10606_),
    .Y(_03662_));
 NAND2x1_ASAP7_75t_R _26788_ (.A(_00903_),
    .B(_10590_),
    .Y(_10607_));
 OA21x2_ASAP7_75t_R _26789_ (.A1(_09455_),
    .A2(_10594_),
    .B(_10607_),
    .Y(_03663_));
 AND2x2_ASAP7_75t_R _26790_ (.A(_00935_),
    .B(_10587_),
    .Y(_10608_));
 AOI21x1_ASAP7_75t_R _26791_ (.A1(_08948_),
    .A2(_10584_),
    .B(_10608_),
    .Y(_03664_));
 NAND2x1_ASAP7_75t_R _26792_ (.A(_01007_),
    .B(_10579_),
    .Y(_10609_));
 OA21x2_ASAP7_75t_R _26793_ (.A1(_09592_),
    .A2(_10501_),
    .B(_10609_),
    .Y(_03665_));
 NAND2x1_ASAP7_75t_R _26794_ (.A(_00967_),
    .B(_10590_),
    .Y(_10610_));
 OA21x2_ASAP7_75t_R _26795_ (.A1(_09587_),
    .A2(_10594_),
    .B(_10610_),
    .Y(_03666_));
 NAND2x1_ASAP7_75t_R _26796_ (.A(_00999_),
    .B(_10590_),
    .Y(_10611_));
 OA21x2_ASAP7_75t_R _26797_ (.A1(_09589_),
    .A2(_10594_),
    .B(_10611_),
    .Y(_03667_));
 BUFx12f_ASAP7_75t_R _26798_ (.A(_10586_),
    .Y(_10612_));
 NAND2x1_ASAP7_75t_R _26799_ (.A(_01031_),
    .B(_10612_),
    .Y(_10613_));
 OA21x2_ASAP7_75t_R _26800_ (.A1(_09592_),
    .A2(_10594_),
    .B(_10613_),
    .Y(_03668_));
 BUFx6f_ASAP7_75t_R _26801_ (.A(_10586_),
    .Y(_10614_));
 NAND2x1_ASAP7_75t_R _26802_ (.A(_01063_),
    .B(_10612_),
    .Y(_10615_));
 OA21x2_ASAP7_75t_R _26803_ (.A1(_09594_),
    .A2(_10614_),
    .B(_10615_),
    .Y(_03669_));
 NAND2x1_ASAP7_75t_R _26804_ (.A(_01095_),
    .B(_10612_),
    .Y(_10616_));
 OA21x2_ASAP7_75t_R _26805_ (.A1(_09596_),
    .A2(_10614_),
    .B(_10616_),
    .Y(_03670_));
 NAND2x1_ASAP7_75t_R _26806_ (.A(_01127_),
    .B(_10612_),
    .Y(_10617_));
 OA21x2_ASAP7_75t_R _26807_ (.A1(_09598_),
    .A2(_10614_),
    .B(_10617_),
    .Y(_03671_));
 NAND2x1_ASAP7_75t_R _26808_ (.A(_01159_),
    .B(_10612_),
    .Y(_10618_));
 OA21x2_ASAP7_75t_R _26809_ (.A1(_09600_),
    .A2(_10614_),
    .B(_10618_),
    .Y(_03672_));
 NAND2x1_ASAP7_75t_R _26810_ (.A(_01191_),
    .B(_10612_),
    .Y(_10619_));
 OA21x2_ASAP7_75t_R _26811_ (.A1(_09602_),
    .A2(_10614_),
    .B(_10619_),
    .Y(_03673_));
 NAND2x1_ASAP7_75t_R _26812_ (.A(_01223_),
    .B(_10612_),
    .Y(_10620_));
 OA21x2_ASAP7_75t_R _26813_ (.A1(_09604_),
    .A2(_10614_),
    .B(_10620_),
    .Y(_03674_));
 NAND2x1_ASAP7_75t_R _26814_ (.A(_01255_),
    .B(_10612_),
    .Y(_10621_));
 OA21x2_ASAP7_75t_R _26815_ (.A1(_09606_),
    .A2(_10614_),
    .B(_10621_),
    .Y(_03675_));
 NAND2x1_ASAP7_75t_R _26816_ (.A(_01039_),
    .B(_10579_),
    .Y(_10622_));
 OA21x2_ASAP7_75t_R _26817_ (.A1(_09594_),
    .A2(_10501_),
    .B(_10622_),
    .Y(_03676_));
 NAND2x1_ASAP7_75t_R _26818_ (.A(_01287_),
    .B(_10612_),
    .Y(_10623_));
 OA21x2_ASAP7_75t_R _26819_ (.A1(_09608_),
    .A2(_10614_),
    .B(_10623_),
    .Y(_03677_));
 NAND2x1_ASAP7_75t_R _26820_ (.A(_01319_),
    .B(_10612_),
    .Y(_10624_));
 OA21x2_ASAP7_75t_R _26821_ (.A1(_09610_),
    .A2(_10614_),
    .B(_10624_),
    .Y(_03678_));
 NAND2x1_ASAP7_75t_R _26822_ (.A(_01351_),
    .B(_10587_),
    .Y(_10625_));
 OA21x2_ASAP7_75t_R _26823_ (.A1(_09366_),
    .A2(_10614_),
    .B(_10625_),
    .Y(_03679_));
 AND2x2_ASAP7_75t_R _26824_ (.A(_04878_),
    .B(_10586_),
    .Y(_10626_));
 AO21x1_ASAP7_75t_R _26825_ (.A1(_09393_),
    .A2(_10583_),
    .B(_10626_),
    .Y(_03680_));
 NOR2x2_ASAP7_75t_R _26826_ (.A(_08263_),
    .B(_09770_),
    .Y(_10627_));
 BUFx6f_ASAP7_75t_R _26827_ (.A(_10627_),
    .Y(_10628_));
 OR2x2_ASAP7_75t_R _26828_ (.A(_08263_),
    .B(_09770_),
    .Y(_10629_));
 BUFx6f_ASAP7_75t_R _26829_ (.A(_10629_),
    .Y(_10630_));
 BUFx6f_ASAP7_75t_R _26830_ (.A(_10630_),
    .Y(_10631_));
 AND2x2_ASAP7_75t_R _26831_ (.A(_00406_),
    .B(_10631_),
    .Y(_10632_));
 AOI21x1_ASAP7_75t_R _26832_ (.A1(_10329_),
    .A2(_10628_),
    .B(_10632_),
    .Y(_03681_));
 AND2x2_ASAP7_75t_R _26833_ (.A(_00439_),
    .B(_10631_),
    .Y(_10633_));
 AOI21x1_ASAP7_75t_R _26834_ (.A1(_10345_),
    .A2(_10628_),
    .B(_10633_),
    .Y(_03682_));
 BUFx6f_ASAP7_75t_R _26835_ (.A(_10630_),
    .Y(_10634_));
 NOR2x1_ASAP7_75t_R _26836_ (.A(_09543_),
    .B(_10634_),
    .Y(_10635_));
 AO21x1_ASAP7_75t_R _26837_ (.A1(_13595_),
    .A2(_10634_),
    .B(_10635_),
    .Y(_03683_));
 AND2x2_ASAP7_75t_R _26838_ (.A(_13656_),
    .B(_10631_),
    .Y(_10636_));
 AO21x1_ASAP7_75t_R _26839_ (.A1(_09560_),
    .A2(_10628_),
    .B(_10636_),
    .Y(_03684_));
 AND2x2_ASAP7_75t_R _26840_ (.A(_13747_),
    .B(_10631_),
    .Y(_10637_));
 AO21x1_ASAP7_75t_R _26841_ (.A1(_08993_),
    .A2(_10628_),
    .B(_10637_),
    .Y(_03685_));
 AND2x2_ASAP7_75t_R _26842_ (.A(_14887_),
    .B(_10631_),
    .Y(_10638_));
 AO21x1_ASAP7_75t_R _26843_ (.A1(_09268_),
    .A2(_10628_),
    .B(_10638_),
    .Y(_03686_));
 NAND2x1_ASAP7_75t_R _26844_ (.A(_01071_),
    .B(_10579_),
    .Y(_10639_));
 OA21x2_ASAP7_75t_R _26845_ (.A1(_09596_),
    .A2(_10501_),
    .B(_10639_),
    .Y(_03687_));
 AND2x2_ASAP7_75t_R _26846_ (.A(_14956_),
    .B(_10631_),
    .Y(_10640_));
 AO21x1_ASAP7_75t_R _26847_ (.A1(_09412_),
    .A2(_10628_),
    .B(_10640_),
    .Y(_03688_));
 AND2x2_ASAP7_75t_R _26848_ (.A(_15015_),
    .B(_10631_),
    .Y(_10641_));
 AO21x1_ASAP7_75t_R _26849_ (.A1(_09436_),
    .A2(_10628_),
    .B(_10641_),
    .Y(_03689_));
 AND2x2_ASAP7_75t_R _26850_ (.A(_13971_),
    .B(_10631_),
    .Y(_10642_));
 AO21x1_ASAP7_75t_R _26851_ (.A1(_10098_),
    .A2(_10628_),
    .B(_10642_),
    .Y(_03690_));
 AND2x2_ASAP7_75t_R _26852_ (.A(_14082_),
    .B(_10631_),
    .Y(_10643_));
 AO21x1_ASAP7_75t_R _26853_ (.A1(_10282_),
    .A2(_10628_),
    .B(_10643_),
    .Y(_03691_));
 BUFx6f_ASAP7_75t_R _26854_ (.A(_10630_),
    .Y(_10644_));
 AND2x2_ASAP7_75t_R _26855_ (.A(_14145_),
    .B(_10644_),
    .Y(_10645_));
 AO21x1_ASAP7_75t_R _26856_ (.A1(_10102_),
    .A2(_10628_),
    .B(_10645_),
    .Y(_03692_));
 BUFx6f_ASAP7_75t_R _26857_ (.A(_10627_),
    .Y(_10646_));
 AND2x2_ASAP7_75t_R _26858_ (.A(_14359_),
    .B(_10644_),
    .Y(_10647_));
 AO21x1_ASAP7_75t_R _26859_ (.A1(_10286_),
    .A2(_10646_),
    .B(_10647_),
    .Y(_03693_));
 AND2x2_ASAP7_75t_R _26860_ (.A(_13198_),
    .B(_10644_),
    .Y(_10648_));
 AO21x1_ASAP7_75t_R _26861_ (.A1(_10107_),
    .A2(_10646_),
    .B(_10648_),
    .Y(_03694_));
 AND2x2_ASAP7_75t_R _26862_ (.A(_15417_),
    .B(_10644_),
    .Y(_10649_));
 AO21x1_ASAP7_75t_R _26863_ (.A1(_10244_),
    .A2(_10646_),
    .B(_10649_),
    .Y(_03695_));
 NOR2x1_ASAP7_75t_R _26864_ (.A(_09451_),
    .B(_10634_),
    .Y(_10650_));
 AO21x1_ASAP7_75t_R _26865_ (.A1(_15570_),
    .A2(_10634_),
    .B(_10650_),
    .Y(_03696_));
 NAND2x1_ASAP7_75t_R _26866_ (.A(_00872_),
    .B(_10634_),
    .Y(_10651_));
 OA21x2_ASAP7_75t_R _26867_ (.A1(_10430_),
    .A2(_10634_),
    .B(_10651_),
    .Y(_03697_));
 NAND2x1_ASAP7_75t_R _26868_ (.A(_01103_),
    .B(_10579_),
    .Y(_10652_));
 OA21x2_ASAP7_75t_R _26869_ (.A1(_09598_),
    .A2(_10501_),
    .B(_10652_),
    .Y(_03698_));
 AND2x2_ASAP7_75t_R _26870_ (.A(_09930_),
    .B(_10627_),
    .Y(_10653_));
 AO21x1_ASAP7_75t_R _26871_ (.A1(_15776_),
    .A2(_10634_),
    .B(_10653_),
    .Y(_03699_));
 NOR2x1_ASAP7_75t_R _26872_ (.A(_09457_),
    .B(_10631_),
    .Y(_10654_));
 AO21x1_ASAP7_75t_R _26873_ (.A1(_15931_),
    .A2(_10634_),
    .B(_10654_),
    .Y(_03700_));
 AND2x2_ASAP7_75t_R _26874_ (.A(_16023_),
    .B(_10644_),
    .Y(_10655_));
 AO21x1_ASAP7_75t_R _26875_ (.A1(_09022_),
    .A2(_10646_),
    .B(_10655_),
    .Y(_03701_));
 AND2x2_ASAP7_75t_R _26876_ (.A(_16178_),
    .B(_10644_),
    .Y(_10656_));
 AO21x1_ASAP7_75t_R _26877_ (.A1(_09049_),
    .A2(_10646_),
    .B(_10656_),
    .Y(_03702_));
 AND2x2_ASAP7_75t_R _26878_ (.A(_16313_),
    .B(_10644_),
    .Y(_10657_));
 AO21x1_ASAP7_75t_R _26879_ (.A1(_09075_),
    .A2(_10646_),
    .B(_10657_),
    .Y(_03703_));
 AND2x2_ASAP7_75t_R _26880_ (.A(_16436_),
    .B(_10644_),
    .Y(_10658_));
 AO21x1_ASAP7_75t_R _26881_ (.A1(_09100_),
    .A2(_10646_),
    .B(_10658_),
    .Y(_03704_));
 AND2x2_ASAP7_75t_R _26882_ (.A(_16574_),
    .B(_10644_),
    .Y(_10659_));
 AO21x1_ASAP7_75t_R _26883_ (.A1(_09124_),
    .A2(_10646_),
    .B(_10659_),
    .Y(_03705_));
 AND2x2_ASAP7_75t_R _26884_ (.A(_16684_),
    .B(_10644_),
    .Y(_10660_));
 AO21x1_ASAP7_75t_R _26885_ (.A1(_09145_),
    .A2(_10646_),
    .B(_10660_),
    .Y(_03706_));
 AND2x2_ASAP7_75t_R _26886_ (.A(_16807_),
    .B(_10630_),
    .Y(_10661_));
 AO21x1_ASAP7_75t_R _26887_ (.A1(_09177_),
    .A2(_10646_),
    .B(_10661_),
    .Y(_03707_));
 AND2x2_ASAP7_75t_R _26888_ (.A(_16876_),
    .B(_10630_),
    .Y(_10662_));
 AO21x1_ASAP7_75t_R _26889_ (.A1(_09204_),
    .A2(_10627_),
    .B(_10662_),
    .Y(_03708_));
 NAND2x1_ASAP7_75t_R _26890_ (.A(_01135_),
    .B(_10579_),
    .Y(_10663_));
 OA21x2_ASAP7_75t_R _26891_ (.A1(_09600_),
    .A2(_10357_),
    .B(_10663_),
    .Y(_03709_));
 AND2x2_ASAP7_75t_R _26892_ (.A(_04292_),
    .B(_10630_),
    .Y(_10664_));
 AO21x1_ASAP7_75t_R _26893_ (.A1(_09230_),
    .A2(_10627_),
    .B(_10664_),
    .Y(_03710_));
 AND2x2_ASAP7_75t_R _26894_ (.A(_04405_),
    .B(_10630_),
    .Y(_10665_));
 AO21x1_ASAP7_75t_R _26895_ (.A1(_09250_),
    .A2(_10627_),
    .B(_10665_),
    .Y(_03711_));
 AND2x2_ASAP7_75t_R _26896_ (.A(_04499_),
    .B(_10630_),
    .Y(_10666_));
 AO21x1_ASAP7_75t_R _26897_ (.A1(_09302_),
    .A2(_10627_),
    .B(_10666_),
    .Y(_03712_));
 AND2x2_ASAP7_75t_R _26898_ (.A(_04653_),
    .B(_10630_),
    .Y(_10667_));
 AO21x1_ASAP7_75t_R _26899_ (.A1(_09335_),
    .A2(_10627_),
    .B(_10667_),
    .Y(_03713_));
 NAND2x1_ASAP7_75t_R _26900_ (.A(_01352_),
    .B(_10634_),
    .Y(_10668_));
 OA21x2_ASAP7_75t_R _26901_ (.A1(_09366_),
    .A2(_10634_),
    .B(_10668_),
    .Y(_03714_));
 AND2x2_ASAP7_75t_R _26902_ (.A(_04881_),
    .B(_10630_),
    .Y(_10669_));
 AO21x1_ASAP7_75t_R _26903_ (.A1(_09393_),
    .A2(_10627_),
    .B(_10669_),
    .Y(_03715_));
 NOR2x2_ASAP7_75t_R _26904_ (.A(_08254_),
    .B(_10132_),
    .Y(_10670_));
 BUFx12f_ASAP7_75t_R _26905_ (.A(_10670_),
    .Y(_10671_));
 BUFx6f_ASAP7_75t_R _26906_ (.A(_10671_),
    .Y(_10672_));
 OR2x6_ASAP7_75t_R _26907_ (.A(_08254_),
    .B(_10132_),
    .Y(_10673_));
 BUFx6f_ASAP7_75t_R _26908_ (.A(_10673_),
    .Y(_10674_));
 AND2x2_ASAP7_75t_R _26909_ (.A(_00407_),
    .B(_10674_),
    .Y(_10675_));
 AOI21x1_ASAP7_75t_R _26910_ (.A1(_10329_),
    .A2(_10672_),
    .B(_10675_),
    .Y(_03716_));
 AND2x2_ASAP7_75t_R _26911_ (.A(_00440_),
    .B(_10673_),
    .Y(_10676_));
 AOI21x1_ASAP7_75t_R _26912_ (.A1(_10345_),
    .A2(_10672_),
    .B(_10676_),
    .Y(_03717_));
 AND2x2_ASAP7_75t_R _26913_ (.A(_09543_),
    .B(_10671_),
    .Y(_10677_));
 AOI21x1_ASAP7_75t_R _26914_ (.A1(_00471_),
    .A2(_10674_),
    .B(_10677_),
    .Y(_03718_));
 BUFx12f_ASAP7_75t_R _26915_ (.A(_10670_),
    .Y(_10678_));
 NOR2x1_ASAP7_75t_R _26916_ (.A(_00501_),
    .B(_10678_),
    .Y(_10679_));
 AO21x1_ASAP7_75t_R _26917_ (.A1(_09560_),
    .A2(_10672_),
    .B(_10679_),
    .Y(_03719_));
 NAND2x1_ASAP7_75t_R _26918_ (.A(_01167_),
    .B(_10579_),
    .Y(_10680_));
 OA21x2_ASAP7_75t_R _26919_ (.A1(_09602_),
    .A2(_10357_),
    .B(_10680_),
    .Y(_03720_));
 AND2x2_ASAP7_75t_R _26920_ (.A(_13733_),
    .B(_10673_),
    .Y(_10681_));
 AO21x1_ASAP7_75t_R _26921_ (.A1(_08993_),
    .A2(_10672_),
    .B(_10681_),
    .Y(_03721_));
 NAND2x1_ASAP7_75t_R _26922_ (.A(_00561_),
    .B(_10674_),
    .Y(_10682_));
 OA21x2_ASAP7_75t_R _26923_ (.A1(_09565_),
    .A2(_10674_),
    .B(_10682_),
    .Y(_03722_));
 AND2x2_ASAP7_75t_R _26924_ (.A(_13852_),
    .B(_10673_),
    .Y(_10683_));
 AO21x1_ASAP7_75t_R _26925_ (.A1(_09412_),
    .A2(_10672_),
    .B(_10683_),
    .Y(_03723_));
 AND2x2_ASAP7_75t_R _26926_ (.A(_13921_),
    .B(_10673_),
    .Y(_10684_));
 AO21x1_ASAP7_75t_R _26927_ (.A1(_09436_),
    .A2(_10672_),
    .B(_10684_),
    .Y(_03724_));
 AND2x2_ASAP7_75t_R _26928_ (.A(_13974_),
    .B(_10673_),
    .Y(_10685_));
 AO21x1_ASAP7_75t_R _26929_ (.A1(_10098_),
    .A2(_10672_),
    .B(_10685_),
    .Y(_03725_));
 NOR2x1_ASAP7_75t_R _26930_ (.A(_00681_),
    .B(_10678_),
    .Y(_10686_));
 AO21x1_ASAP7_75t_R _26931_ (.A1(_10282_),
    .A2(_10672_),
    .B(_10686_),
    .Y(_03726_));
 NOR2x1_ASAP7_75t_R _26932_ (.A(_00711_),
    .B(_10678_),
    .Y(_10687_));
 AO21x1_ASAP7_75t_R _26933_ (.A1(_10102_),
    .A2(_10672_),
    .B(_10687_),
    .Y(_03727_));
 AND2x2_ASAP7_75t_R _26934_ (.A(_14247_),
    .B(_10673_),
    .Y(_10688_));
 AO21x1_ASAP7_75t_R _26935_ (.A1(_10286_),
    .A2(_10672_),
    .B(_10688_),
    .Y(_03728_));
 BUFx6f_ASAP7_75t_R _26936_ (.A(_10671_),
    .Y(_10689_));
 NOR2x1_ASAP7_75t_R _26937_ (.A(_00371_),
    .B(_10678_),
    .Y(_10690_));
 AO21x1_ASAP7_75t_R _26938_ (.A1(_10107_),
    .A2(_10689_),
    .B(_10690_),
    .Y(_03729_));
 BUFx12f_ASAP7_75t_R _26939_ (.A(_10670_),
    .Y(_10691_));
 NOR2x1_ASAP7_75t_R _26940_ (.A(_00809_),
    .B(_10691_),
    .Y(_10692_));
 AO21x1_ASAP7_75t_R _26941_ (.A1(_10244_),
    .A2(_10689_),
    .B(_10692_),
    .Y(_03730_));
 NAND2x1_ASAP7_75t_R _26942_ (.A(_01199_),
    .B(_10579_),
    .Y(_10693_));
 OA21x2_ASAP7_75t_R _26943_ (.A1(_09604_),
    .A2(_10357_),
    .B(_10693_),
    .Y(_03731_));
 AND2x2_ASAP7_75t_R _26944_ (.A(_08850_),
    .B(_10671_),
    .Y(_10694_));
 AOI21x1_ASAP7_75t_R _26945_ (.A1(_00841_),
    .A2(_10674_),
    .B(_10694_),
    .Y(_03732_));
 NAND2x1_ASAP7_75t_R _26946_ (.A(_00873_),
    .B(_10674_),
    .Y(_10695_));
 OA21x2_ASAP7_75t_R _26947_ (.A1(_10430_),
    .A2(_10674_),
    .B(_10695_),
    .Y(_03733_));
 NOR2x1_ASAP7_75t_R _26948_ (.A(_00905_),
    .B(_10691_),
    .Y(_10696_));
 AO21x1_ASAP7_75t_R _26949_ (.A1(_09584_),
    .A2(_10689_),
    .B(_10696_),
    .Y(_03734_));
 AND2x2_ASAP7_75t_R _26950_ (.A(_08947_),
    .B(_10671_),
    .Y(_10697_));
 AOI21x1_ASAP7_75t_R _26951_ (.A1(_00937_),
    .A2(_10674_),
    .B(_10697_),
    .Y(_03735_));
 NOR2x1_ASAP7_75t_R _26952_ (.A(_00969_),
    .B(_10691_),
    .Y(_10698_));
 AO21x1_ASAP7_75t_R _26953_ (.A1(_09022_),
    .A2(_10689_),
    .B(_10698_),
    .Y(_03736_));
 NOR2x1_ASAP7_75t_R _26954_ (.A(_01001_),
    .B(_10691_),
    .Y(_10699_));
 AO21x1_ASAP7_75t_R _26955_ (.A1(_09049_),
    .A2(_10689_),
    .B(_10699_),
    .Y(_03737_));
 NOR2x1_ASAP7_75t_R _26956_ (.A(_01033_),
    .B(_10691_),
    .Y(_10700_));
 AO21x1_ASAP7_75t_R _26957_ (.A1(_09075_),
    .A2(_10689_),
    .B(_10700_),
    .Y(_03738_));
 NOR2x1_ASAP7_75t_R _26958_ (.A(_01065_),
    .B(_10691_),
    .Y(_10701_));
 AO21x1_ASAP7_75t_R _26959_ (.A1(_09100_),
    .A2(_10689_),
    .B(_10701_),
    .Y(_03739_));
 NOR2x1_ASAP7_75t_R _26960_ (.A(_01097_),
    .B(_10691_),
    .Y(_10702_));
 AO21x1_ASAP7_75t_R _26961_ (.A1(_09124_),
    .A2(_10689_),
    .B(_10702_),
    .Y(_03740_));
 NOR2x1_ASAP7_75t_R _26962_ (.A(_01129_),
    .B(_10691_),
    .Y(_10703_));
 AO21x1_ASAP7_75t_R _26963_ (.A1(_09145_),
    .A2(_10689_),
    .B(_10703_),
    .Y(_03741_));
 NAND2x1_ASAP7_75t_R _26964_ (.A(_01231_),
    .B(_10579_),
    .Y(_10704_));
 OA21x2_ASAP7_75t_R _26965_ (.A1(_09606_),
    .A2(_10357_),
    .B(_10704_),
    .Y(_03742_));
 NOR2x1_ASAP7_75t_R _26966_ (.A(_01161_),
    .B(_10691_),
    .Y(_10705_));
 AO21x1_ASAP7_75t_R _26967_ (.A1(_09177_),
    .A2(_10689_),
    .B(_10705_),
    .Y(_03743_));
 NOR2x1_ASAP7_75t_R _26968_ (.A(_01193_),
    .B(_10691_),
    .Y(_10706_));
 AO21x1_ASAP7_75t_R _26969_ (.A1(_09204_),
    .A2(_10678_),
    .B(_10706_),
    .Y(_03744_));
 NOR2x1_ASAP7_75t_R _26970_ (.A(_01225_),
    .B(_10671_),
    .Y(_10707_));
 AO21x1_ASAP7_75t_R _26971_ (.A1(_09230_),
    .A2(_10678_),
    .B(_10707_),
    .Y(_03745_));
 NOR2x1_ASAP7_75t_R _26972_ (.A(_01257_),
    .B(_10671_),
    .Y(_10708_));
 AO21x1_ASAP7_75t_R _26973_ (.A1(_09250_),
    .A2(_10678_),
    .B(_10708_),
    .Y(_03746_));
 NOR2x1_ASAP7_75t_R _26974_ (.A(_01289_),
    .B(_10671_),
    .Y(_10709_));
 AO21x1_ASAP7_75t_R _26975_ (.A1(_09302_),
    .A2(_10678_),
    .B(_10709_),
    .Y(_03747_));
 NOR2x1_ASAP7_75t_R _26976_ (.A(_01321_),
    .B(_10671_),
    .Y(_10710_));
 AO21x1_ASAP7_75t_R _26977_ (.A1(_09335_),
    .A2(_10678_),
    .B(_10710_),
    .Y(_03748_));
 NAND2x1_ASAP7_75t_R _26978_ (.A(_01353_),
    .B(_10674_),
    .Y(_10711_));
 OA21x2_ASAP7_75t_R _26979_ (.A1(_09366_),
    .A2(_10674_),
    .B(_10711_),
    .Y(_03749_));
 NOR2x1_ASAP7_75t_R _26980_ (.A(_01385_),
    .B(_10671_),
    .Y(_10712_));
 AO21x1_ASAP7_75t_R _26981_ (.A1(_09393_),
    .A2(_10678_),
    .B(_10712_),
    .Y(_03750_));
 NOR2x2_ASAP7_75t_R _26982_ (.A(_08254_),
    .B(_10176_),
    .Y(_10713_));
 OR2x6_ASAP7_75t_R _26983_ (.A(_08254_),
    .B(_10176_),
    .Y(_10714_));
 BUFx6f_ASAP7_75t_R _26984_ (.A(_10714_),
    .Y(_10715_));
 AND2x2_ASAP7_75t_R _26985_ (.A(_00408_),
    .B(_10715_),
    .Y(_10716_));
 AOI21x1_ASAP7_75t_R _26986_ (.A1(_10329_),
    .A2(_10713_),
    .B(_10716_),
    .Y(_03751_));
 AND2x2_ASAP7_75t_R _26987_ (.A(_00441_),
    .B(_10715_),
    .Y(_10717_));
 AOI21x1_ASAP7_75t_R _26988_ (.A1(_10345_),
    .A2(_10713_),
    .B(_10717_),
    .Y(_03752_));
 NAND2x1_ASAP7_75t_R _26989_ (.A(_01263_),
    .B(_10332_),
    .Y(_10718_));
 OA21x2_ASAP7_75t_R _26990_ (.A1(_09608_),
    .A2(_10357_),
    .B(_10718_),
    .Y(_03753_));
 AND2x2_ASAP7_75t_R _26991_ (.A(_00472_),
    .B(_10715_),
    .Y(_10719_));
 AOI21x1_ASAP7_75t_R _26992_ (.A1(_09675_),
    .A2(_10713_),
    .B(_10719_),
    .Y(_03754_));
 BUFx6f_ASAP7_75t_R _26993_ (.A(_10715_),
    .Y(_10720_));
 BUFx12f_ASAP7_75t_R _26994_ (.A(_10714_),
    .Y(_10721_));
 NAND2x1_ASAP7_75t_R _26995_ (.A(_00502_),
    .B(_10721_),
    .Y(_10722_));
 OA21x2_ASAP7_75t_R _26996_ (.A1(_09629_),
    .A2(_10720_),
    .B(_10722_),
    .Y(_03755_));
 NAND2x1_ASAP7_75t_R _26997_ (.A(_00532_),
    .B(_10721_),
    .Y(_10723_));
 OA21x2_ASAP7_75t_R _26998_ (.A1(_09563_),
    .A2(_10720_),
    .B(_10723_),
    .Y(_03756_));
 NAND2x1_ASAP7_75t_R _26999_ (.A(_00562_),
    .B(_10721_),
    .Y(_10724_));
 OA21x2_ASAP7_75t_R _27000_ (.A1(_09565_),
    .A2(_10720_),
    .B(_10724_),
    .Y(_03757_));
 NAND2x1_ASAP7_75t_R _27001_ (.A(_00592_),
    .B(_10721_),
    .Y(_10725_));
 OA21x2_ASAP7_75t_R _27002_ (.A1(_09567_),
    .A2(_10720_),
    .B(_10725_),
    .Y(_03758_));
 NAND2x1_ASAP7_75t_R _27003_ (.A(_00622_),
    .B(_10721_),
    .Y(_10726_));
 OA21x2_ASAP7_75t_R _27004_ (.A1(_09570_),
    .A2(_10720_),
    .B(_10726_),
    .Y(_03759_));
 BUFx12f_ASAP7_75t_R _27005_ (.A(_10715_),
    .Y(_10727_));
 NAND2x1_ASAP7_75t_R _27006_ (.A(_00652_),
    .B(_10727_),
    .Y(_10728_));
 OA21x2_ASAP7_75t_R _27007_ (.A1(_09438_),
    .A2(_10720_),
    .B(_10728_),
    .Y(_03760_));
 AND2x2_ASAP7_75t_R _27008_ (.A(_14072_),
    .B(_10715_),
    .Y(_10729_));
 AO21x1_ASAP7_75t_R _27009_ (.A1(_10282_),
    .A2(_10713_),
    .B(_10729_),
    .Y(_03761_));
 NAND2x1_ASAP7_75t_R _27010_ (.A(_00712_),
    .B(_10727_),
    .Y(_10730_));
 OA21x2_ASAP7_75t_R _27011_ (.A1(_09443_),
    .A2(_10720_),
    .B(_10730_),
    .Y(_03762_));
 AND2x2_ASAP7_75t_R _27012_ (.A(_14254_),
    .B(_10715_),
    .Y(_10731_));
 AO21x1_ASAP7_75t_R _27013_ (.A1(_10286_),
    .A2(_10713_),
    .B(_10731_),
    .Y(_03763_));
 NAND2x1_ASAP7_75t_R _27014_ (.A(_01295_),
    .B(_10332_),
    .Y(_10732_));
 OA21x2_ASAP7_75t_R _27015_ (.A1(_09610_),
    .A2(_10357_),
    .B(_10732_),
    .Y(_03764_));
 NAND2x1_ASAP7_75t_R _27016_ (.A(_00372_),
    .B(_10727_),
    .Y(_10733_));
 OA21x2_ASAP7_75t_R _27017_ (.A1(_09447_),
    .A2(_10720_),
    .B(_10733_),
    .Y(_03765_));
 NAND2x1_ASAP7_75t_R _27018_ (.A(_00810_),
    .B(_10727_),
    .Y(_10734_));
 OA21x2_ASAP7_75t_R _27019_ (.A1(_09449_),
    .A2(_10720_),
    .B(_10734_),
    .Y(_03766_));
 AND2x2_ASAP7_75t_R _27020_ (.A(_00842_),
    .B(_10715_),
    .Y(_10735_));
 AOI21x1_ASAP7_75t_R _27021_ (.A1(_09790_),
    .A2(_10713_),
    .B(_10735_),
    .Y(_03767_));
 NAND2x1_ASAP7_75t_R _27022_ (.A(_00874_),
    .B(_10727_),
    .Y(_10736_));
 OA21x2_ASAP7_75t_R _27023_ (.A1(_10430_),
    .A2(_10720_),
    .B(_10736_),
    .Y(_03768_));
 BUFx6f_ASAP7_75t_R _27024_ (.A(_10715_),
    .Y(_10737_));
 NAND2x1_ASAP7_75t_R _27025_ (.A(_00906_),
    .B(_10727_),
    .Y(_10738_));
 OA21x2_ASAP7_75t_R _27026_ (.A1(_09455_),
    .A2(_10737_),
    .B(_10738_),
    .Y(_03769_));
 AND2x2_ASAP7_75t_R _27027_ (.A(_00938_),
    .B(_10715_),
    .Y(_10739_));
 AOI21x1_ASAP7_75t_R _27028_ (.A1(_08948_),
    .A2(_10713_),
    .B(_10739_),
    .Y(_03770_));
 NAND2x1_ASAP7_75t_R _27029_ (.A(_00970_),
    .B(_10727_),
    .Y(_10740_));
 OA21x2_ASAP7_75t_R _27030_ (.A1(_09587_),
    .A2(_10737_),
    .B(_10740_),
    .Y(_03771_));
 NAND2x1_ASAP7_75t_R _27031_ (.A(_01002_),
    .B(_10727_),
    .Y(_10741_));
 OA21x2_ASAP7_75t_R _27032_ (.A1(_09589_),
    .A2(_10737_),
    .B(_10741_),
    .Y(_03772_));
 NAND2x1_ASAP7_75t_R _27033_ (.A(_01034_),
    .B(_10727_),
    .Y(_10742_));
 OA21x2_ASAP7_75t_R _27034_ (.A1(_09592_),
    .A2(_10737_),
    .B(_10742_),
    .Y(_03773_));
 NAND2x1_ASAP7_75t_R _27035_ (.A(_01066_),
    .B(_10727_),
    .Y(_10743_));
 OA21x2_ASAP7_75t_R _27036_ (.A1(_09594_),
    .A2(_10737_),
    .B(_10743_),
    .Y(_03774_));
 NAND2x1_ASAP7_75t_R _27037_ (.A(_01327_),
    .B(_10332_),
    .Y(_10744_));
 OA21x2_ASAP7_75t_R _27038_ (.A1(_09366_),
    .A2(_10357_),
    .B(_10744_),
    .Y(_03775_));
 BUFx12f_ASAP7_75t_R _27039_ (.A(_10714_),
    .Y(_10745_));
 NAND2x1_ASAP7_75t_R _27040_ (.A(_01098_),
    .B(_10745_),
    .Y(_10746_));
 OA21x2_ASAP7_75t_R _27041_ (.A1(_09596_),
    .A2(_10737_),
    .B(_10746_),
    .Y(_03776_));
 NAND2x1_ASAP7_75t_R _27042_ (.A(_01130_),
    .B(_10745_),
    .Y(_10747_));
 OA21x2_ASAP7_75t_R _27043_ (.A1(_09598_),
    .A2(_10737_),
    .B(_10747_),
    .Y(_03777_));
 NAND2x1_ASAP7_75t_R _27044_ (.A(_01162_),
    .B(_10745_),
    .Y(_10748_));
 OA21x2_ASAP7_75t_R _27045_ (.A1(_09600_),
    .A2(_10737_),
    .B(_10748_),
    .Y(_03778_));
 NAND2x1_ASAP7_75t_R _27046_ (.A(_01194_),
    .B(_10745_),
    .Y(_10749_));
 OA21x2_ASAP7_75t_R _27047_ (.A1(_09602_),
    .A2(_10737_),
    .B(_10749_),
    .Y(_03779_));
 NAND2x1_ASAP7_75t_R _27048_ (.A(_01226_),
    .B(_10745_),
    .Y(_10750_));
 OA21x2_ASAP7_75t_R _27049_ (.A1(_09604_),
    .A2(_10737_),
    .B(_10750_),
    .Y(_03780_));
 NAND2x1_ASAP7_75t_R _27050_ (.A(_01258_),
    .B(_10745_),
    .Y(_10751_));
 OA21x2_ASAP7_75t_R _27051_ (.A1(_09606_),
    .A2(_10721_),
    .B(_10751_),
    .Y(_03781_));
 NAND2x1_ASAP7_75t_R _27052_ (.A(_01290_),
    .B(_10745_),
    .Y(_10752_));
 OA21x2_ASAP7_75t_R _27053_ (.A1(_09608_),
    .A2(_10721_),
    .B(_10752_),
    .Y(_03782_));
 NAND2x1_ASAP7_75t_R _27054_ (.A(_01322_),
    .B(_10745_),
    .Y(_10753_));
 OA21x2_ASAP7_75t_R _27055_ (.A1(_09610_),
    .A2(_10721_),
    .B(_10753_),
    .Y(_03783_));
 NAND2x1_ASAP7_75t_R _27056_ (.A(_01354_),
    .B(_10745_),
    .Y(_10754_));
 OA21x2_ASAP7_75t_R _27057_ (.A1(_09366_),
    .A2(_10721_),
    .B(_10754_),
    .Y(_03784_));
 NAND2x1_ASAP7_75t_R _27058_ (.A(_01386_),
    .B(_10745_),
    .Y(_10755_));
 OA21x2_ASAP7_75t_R _27059_ (.A1(_09614_),
    .A2(_10721_),
    .B(_10755_),
    .Y(_03785_));
 AND2x2_ASAP7_75t_R _27060_ (.A(_04893_),
    .B(_10332_),
    .Y(_10756_));
 AO21x1_ASAP7_75t_R _27061_ (.A1(_09393_),
    .A2(_10330_),
    .B(_10756_),
    .Y(_03786_));
 NOR2x2_ASAP7_75t_R _27062_ (.A(_08254_),
    .B(_10221_),
    .Y(_10757_));
 BUFx6f_ASAP7_75t_R _27063_ (.A(_10757_),
    .Y(_10758_));
 OR2x6_ASAP7_75t_R _27064_ (.A(_08254_),
    .B(_10221_),
    .Y(_10759_));
 BUFx12f_ASAP7_75t_R _27065_ (.A(_10759_),
    .Y(_10760_));
 BUFx6f_ASAP7_75t_R _27066_ (.A(_10760_),
    .Y(_10761_));
 AND2x2_ASAP7_75t_R _27067_ (.A(_00409_),
    .B(_10761_),
    .Y(_10762_));
 AOI21x1_ASAP7_75t_R _27068_ (.A1(_09502_),
    .A2(_10758_),
    .B(_10762_),
    .Y(_03787_));
 AND2x2_ASAP7_75t_R _27069_ (.A(_00442_),
    .B(_10761_),
    .Y(_10763_));
 AOI21x1_ASAP7_75t_R _27070_ (.A1(_09526_),
    .A2(_10758_),
    .B(_10763_),
    .Y(_03788_));
 BUFx6f_ASAP7_75t_R _27071_ (.A(_10760_),
    .Y(_10764_));
 NOR2x1_ASAP7_75t_R _27072_ (.A(_09543_),
    .B(_10764_),
    .Y(_10765_));
 AO21x1_ASAP7_75t_R _27073_ (.A1(_13585_),
    .A2(_10764_),
    .B(_10765_),
    .Y(_03789_));
 AND2x2_ASAP7_75t_R _27074_ (.A(_13617_),
    .B(_10761_),
    .Y(_10766_));
 AO21x1_ASAP7_75t_R _27075_ (.A1(_09560_),
    .A2(_10758_),
    .B(_10766_),
    .Y(_03790_));
 AND2x2_ASAP7_75t_R _27076_ (.A(_14818_),
    .B(_10761_),
    .Y(_10767_));
 AO21x1_ASAP7_75t_R _27077_ (.A1(_08993_),
    .A2(_10758_),
    .B(_10767_),
    .Y(_03791_));
 AND2x2_ASAP7_75t_R _27078_ (.A(_13818_),
    .B(_10761_),
    .Y(_10768_));
 AO21x1_ASAP7_75t_R _27079_ (.A1(_09268_),
    .A2(_10758_),
    .B(_10768_),
    .Y(_03792_));
 AND2x2_ASAP7_75t_R _27080_ (.A(_13849_),
    .B(_10761_),
    .Y(_10769_));
 AO21x1_ASAP7_75t_R _27081_ (.A1(_09412_),
    .A2(_10758_),
    .B(_10769_),
    .Y(_03793_));
 AND2x2_ASAP7_75t_R _27082_ (.A(_13918_),
    .B(_10761_),
    .Y(_10770_));
 AO21x1_ASAP7_75t_R _27083_ (.A1(_09436_),
    .A2(_10758_),
    .B(_10770_),
    .Y(_03794_));
 AND2x2_ASAP7_75t_R _27084_ (.A(_15081_),
    .B(_10761_),
    .Y(_10771_));
 AO21x1_ASAP7_75t_R _27085_ (.A1(_10098_),
    .A2(_10758_),
    .B(_10771_),
    .Y(_03795_));
 AND2x2_ASAP7_75t_R _27086_ (.A(_14067_),
    .B(_10761_),
    .Y(_10772_));
 AO21x1_ASAP7_75t_R _27087_ (.A1(_10282_),
    .A2(_10758_),
    .B(_10772_),
    .Y(_03796_));
 AND2x2_ASAP7_75t_R _27088_ (.A(_00382_),
    .B(_09414_),
    .Y(_10773_));
 AOI21x1_ASAP7_75t_R _27089_ (.A1(_08956_),
    .A2(_09503_),
    .B(_10773_),
    .Y(_03797_));
 BUFx6f_ASAP7_75t_R _27090_ (.A(_10760_),
    .Y(_10774_));
 AND2x2_ASAP7_75t_R _27091_ (.A(_14163_),
    .B(_10774_),
    .Y(_10775_));
 AO21x1_ASAP7_75t_R _27092_ (.A1(_10102_),
    .A2(_10758_),
    .B(_10775_),
    .Y(_03798_));
 BUFx6f_ASAP7_75t_R _27093_ (.A(_10757_),
    .Y(_10776_));
 AND2x2_ASAP7_75t_R _27094_ (.A(_14244_),
    .B(_10774_),
    .Y(_10777_));
 AO21x1_ASAP7_75t_R _27095_ (.A1(_10286_),
    .A2(_10776_),
    .B(_10777_),
    .Y(_03799_));
 AND2x2_ASAP7_75t_R _27096_ (.A(_13180_),
    .B(_10774_),
    .Y(_10778_));
 AO21x1_ASAP7_75t_R _27097_ (.A1(_10107_),
    .A2(_10776_),
    .B(_10778_),
    .Y(_03800_));
 AND2x2_ASAP7_75t_R _27098_ (.A(_15409_),
    .B(_10774_),
    .Y(_10779_));
 AO21x1_ASAP7_75t_R _27099_ (.A1(_10244_),
    .A2(_10776_),
    .B(_10779_),
    .Y(_03801_));
 NOR2x1_ASAP7_75t_R _27100_ (.A(_09451_),
    .B(_10764_),
    .Y(_10780_));
 AO21x1_ASAP7_75t_R _27101_ (.A1(_15562_),
    .A2(_10764_),
    .B(_10780_),
    .Y(_03802_));
 NAND2x1_ASAP7_75t_R _27102_ (.A(_00875_),
    .B(_10764_),
    .Y(_10781_));
 OA21x2_ASAP7_75t_R _27103_ (.A1(_10430_),
    .A2(_10764_),
    .B(_10781_),
    .Y(_03803_));
 AND2x2_ASAP7_75t_R _27104_ (.A(_09930_),
    .B(_10757_),
    .Y(_10782_));
 AO21x1_ASAP7_75t_R _27105_ (.A1(_15798_),
    .A2(_10764_),
    .B(_10782_),
    .Y(_03804_));
 NOR2x1_ASAP7_75t_R _27106_ (.A(_09457_),
    .B(_10761_),
    .Y(_10783_));
 AO21x1_ASAP7_75t_R _27107_ (.A1(_15923_),
    .A2(_10764_),
    .B(_10783_),
    .Y(_03805_));
 AND2x2_ASAP7_75t_R _27108_ (.A(_16045_),
    .B(_10774_),
    .Y(_10784_));
 AO21x1_ASAP7_75t_R _27109_ (.A1(_09022_),
    .A2(_10776_),
    .B(_10784_),
    .Y(_03806_));
 AND2x2_ASAP7_75t_R _27110_ (.A(_16170_),
    .B(_10774_),
    .Y(_10785_));
 AO21x1_ASAP7_75t_R _27111_ (.A1(_09049_),
    .A2(_10776_),
    .B(_10785_),
    .Y(_03807_));
 AND2x2_ASAP7_75t_R _27112_ (.A(_00415_),
    .B(_09414_),
    .Y(_10786_));
 AOI21x1_ASAP7_75t_R _27113_ (.A1(_08956_),
    .A2(_09527_),
    .B(_10786_),
    .Y(_03808_));
 AND2x2_ASAP7_75t_R _27114_ (.A(_16305_),
    .B(_10774_),
    .Y(_10787_));
 AO21x1_ASAP7_75t_R _27115_ (.A1(_09075_),
    .A2(_10776_),
    .B(_10787_),
    .Y(_03809_));
 AND2x2_ASAP7_75t_R _27116_ (.A(_16428_),
    .B(_10774_),
    .Y(_10788_));
 AO21x1_ASAP7_75t_R _27117_ (.A1(_09100_),
    .A2(_10776_),
    .B(_10788_),
    .Y(_03810_));
 AND2x2_ASAP7_75t_R _27118_ (.A(_16566_),
    .B(_10774_),
    .Y(_10789_));
 AO21x1_ASAP7_75t_R _27119_ (.A1(_09124_),
    .A2(_10776_),
    .B(_10789_),
    .Y(_03811_));
 AND2x2_ASAP7_75t_R _27120_ (.A(_16676_),
    .B(_10774_),
    .Y(_10790_));
 AO21x1_ASAP7_75t_R _27121_ (.A1(_09145_),
    .A2(_10776_),
    .B(_10790_),
    .Y(_03812_));
 AND2x2_ASAP7_75t_R _27122_ (.A(_16799_),
    .B(_10760_),
    .Y(_10791_));
 AO21x1_ASAP7_75t_R _27123_ (.A1(_09177_),
    .A2(_10776_),
    .B(_10791_),
    .Y(_03813_));
 AND2x2_ASAP7_75t_R _27124_ (.A(_16898_),
    .B(_10760_),
    .Y(_10792_));
 AO21x1_ASAP7_75t_R _27125_ (.A1(_09204_),
    .A2(_10757_),
    .B(_10792_),
    .Y(_03814_));
 AND2x2_ASAP7_75t_R _27126_ (.A(_04284_),
    .B(_10760_),
    .Y(_10793_));
 AO21x1_ASAP7_75t_R _27127_ (.A1(_09230_),
    .A2(_10757_),
    .B(_10793_),
    .Y(_03815_));
 AND2x2_ASAP7_75t_R _27128_ (.A(_04397_),
    .B(_10760_),
    .Y(_10794_));
 AO21x1_ASAP7_75t_R _27129_ (.A1(_09250_),
    .A2(_10757_),
    .B(_10794_),
    .Y(_03816_));
 AND2x2_ASAP7_75t_R _27130_ (.A(_04521_),
    .B(_10760_),
    .Y(_10795_));
 AO21x1_ASAP7_75t_R _27131_ (.A1(_09302_),
    .A2(_10757_),
    .B(_10795_),
    .Y(_03817_));
 AND2x2_ASAP7_75t_R _27132_ (.A(_04645_),
    .B(_10760_),
    .Y(_10796_));
 AO21x1_ASAP7_75t_R _27133_ (.A1(_09335_),
    .A2(_10757_),
    .B(_10796_),
    .Y(_03818_));
 AND2x2_ASAP7_75t_R _27134_ (.A(_08955_),
    .B(_09542_),
    .Y(_10797_));
 AOI21x1_ASAP7_75t_R _27135_ (.A1(_00446_),
    .A2(_09414_),
    .B(_10797_),
    .Y(_03819_));
 NAND2x1_ASAP7_75t_R _27136_ (.A(_01355_),
    .B(_10764_),
    .Y(_10798_));
 OA21x2_ASAP7_75t_R _27137_ (.A1(_09366_),
    .A2(_10764_),
    .B(_10798_),
    .Y(_03820_));
 AND2x2_ASAP7_75t_R _27138_ (.A(_04840_),
    .B(_10760_),
    .Y(_10799_));
 AO21x1_ASAP7_75t_R _27139_ (.A1(_09393_),
    .A2(_10757_),
    .B(_10799_),
    .Y(_03821_));
 AND2x2_ASAP7_75t_R _27140_ (.A(_00410_),
    .B(_08509_),
    .Y(_10800_));
 AOI21x1_ASAP7_75t_R _27141_ (.A1(_08265_),
    .A2(_09503_),
    .B(_10800_),
    .Y(_03822_));
 AND2x2_ASAP7_75t_R _27142_ (.A(_00443_),
    .B(_08509_),
    .Y(_10801_));
 AOI21x1_ASAP7_75t_R _27143_ (.A1(_08265_),
    .A2(_09527_),
    .B(_10801_),
    .Y(_03823_));
 NOR2x1_ASAP7_75t_R _27144_ (.A(_08509_),
    .B(_09675_),
    .Y(_10802_));
 AO21x1_ASAP7_75t_R _27145_ (.A1(_13588_),
    .A2(_08804_),
    .B(_10802_),
    .Y(_03824_));
 AND2x2_ASAP7_75t_R _27146_ (.A(_13624_),
    .B(_08508_),
    .Y(_10803_));
 AO21x1_ASAP7_75t_R _27147_ (.A1(_08264_),
    .A2(_09560_),
    .B(_10803_),
    .Y(_03825_));
 AND2x2_ASAP7_75t_R _27148_ (.A(_13739_),
    .B(_08508_),
    .Y(_10804_));
 AO21x1_ASAP7_75t_R _27149_ (.A1(_08264_),
    .A2(_08992_),
    .B(_10804_),
    .Y(_03826_));
 AND2x2_ASAP7_75t_R _27150_ (.A(_13804_),
    .B(_08508_),
    .Y(_10805_));
 AO21x1_ASAP7_75t_R _27151_ (.A1(_08264_),
    .A2(_09267_),
    .B(_10805_),
    .Y(_03827_));
 AND2x2_ASAP7_75t_R _27152_ (.A(_14944_),
    .B(_08508_),
    .Y(_10806_));
 AO21x1_ASAP7_75t_R _27153_ (.A1(_08264_),
    .A2(_09411_),
    .B(_10806_),
    .Y(_03828_));
 AND2x2_ASAP7_75t_R _27154_ (.A(_13928_),
    .B(_08508_),
    .Y(_10807_));
 AO21x1_ASAP7_75t_R _27155_ (.A1(_08264_),
    .A2(_09435_),
    .B(_10807_),
    .Y(_03829_));
 NOR2x1_ASAP7_75t_R _27156_ (.A(_00476_),
    .B(_09462_),
    .Y(_10808_));
 AO21x1_ASAP7_75t_R _27157_ (.A1(_09464_),
    .A2(_09559_),
    .B(_10808_),
    .Y(_03830_));
 NOR2x2_ASAP7_75t_R _27158_ (.A(_06885_),
    .B(_06899_),
    .Y(_10809_));
 AND2x4_ASAP7_75t_R _27159_ (.A(_05449_),
    .B(_05451_),
    .Y(_10810_));
 NOR2x1_ASAP7_75t_R _27160_ (.A(_13233_),
    .B(_01398_),
    .Y(_10811_));
 OA21x2_ASAP7_75t_R _27161_ (.A1(net81),
    .A2(_10811_),
    .B(_04991_),
    .Y(_10812_));
 OR3x2_ASAP7_75t_R _27162_ (.A(_05153_),
    .B(_05173_),
    .C(_10812_),
    .Y(_10813_));
 OR3x1_ASAP7_75t_R _27163_ (.A(_10809_),
    .B(_10810_),
    .C(_10813_),
    .Y(_10814_));
 AO21x1_ASAP7_75t_R _27164_ (.A1(_05404_),
    .A2(_10814_),
    .B(_05402_),
    .Y(_10815_));
 OA21x2_ASAP7_75t_R _27165_ (.A1(_14109_),
    .A2(_14110_),
    .B(_05164_),
    .Y(_10816_));
 AND3x1_ASAP7_75t_R _27166_ (.A(_13724_),
    .B(_02226_),
    .C(_13470_),
    .Y(_10817_));
 INVx1_ASAP7_75t_R _27167_ (.A(_02226_),
    .Y(_10818_));
 AND4x1_ASAP7_75t_R _27168_ (.A(_02228_),
    .B(_10818_),
    .C(_13310_),
    .D(_14105_),
    .Y(_10819_));
 AO21x1_ASAP7_75t_R _27169_ (.A1(_14106_),
    .A2(_10817_),
    .B(_10819_),
    .Y(_10820_));
 AND4x1_ASAP7_75t_R _27170_ (.A(_14107_),
    .B(_05702_),
    .C(_05191_),
    .D(_10820_),
    .Y(_10821_));
 OR3x2_ASAP7_75t_R _27171_ (.A(_06908_),
    .B(_10816_),
    .C(_10821_),
    .Y(_10822_));
 NOR2x1_ASAP7_75t_R _27172_ (.A(\id_stage_i.controller_i.exc_req_d ),
    .B(_10822_),
    .Y(_10823_));
 OR2x6_ASAP7_75t_R _27173_ (.A(_06885_),
    .B(_06899_),
    .Y(_10824_));
 BUFx6f_ASAP7_75t_R _27174_ (.A(_10824_),
    .Y(_10825_));
 OAI21x1_ASAP7_75t_R _27175_ (.A1(net81),
    .A2(_10811_),
    .B(_04991_),
    .Y(_10826_));
 BUFx12f_ASAP7_75t_R _27176_ (.A(_05190_),
    .Y(_10827_));
 BUFx12f_ASAP7_75t_R _27177_ (.A(_10827_),
    .Y(_10828_));
 OA21x2_ASAP7_75t_R _27178_ (.A1(_10825_),
    .A2(_10826_),
    .B(_10828_),
    .Y(_10829_));
 OR3x1_ASAP7_75t_R _27179_ (.A(_05172_),
    .B(_05704_),
    .C(_05154_),
    .Y(_10830_));
 NAND2x1_ASAP7_75t_R _27180_ (.A(_10813_),
    .B(_10830_),
    .Y(_10831_));
 AO21x1_ASAP7_75t_R _27181_ (.A1(_05171_),
    .A2(_05704_),
    .B(_05706_),
    .Y(_10832_));
 OA21x2_ASAP7_75t_R _27182_ (.A1(_05415_),
    .A2(_07269_),
    .B(_10812_),
    .Y(_10833_));
 NOR2x1_ASAP7_75t_R _27183_ (.A(_05174_),
    .B(_10833_),
    .Y(_10834_));
 OA21x2_ASAP7_75t_R _27184_ (.A1(_05166_),
    .A2(_05409_),
    .B(_10834_),
    .Y(_10835_));
 AO221x1_ASAP7_75t_R _27185_ (.A1(_05404_),
    .A2(_10831_),
    .B1(_10832_),
    .B2(_05172_),
    .C(_10835_),
    .Y(_10836_));
 AO21x1_ASAP7_75t_R _27186_ (.A1(_10823_),
    .A2(_10829_),
    .B(_10836_),
    .Y(_10837_));
 AND3x1_ASAP7_75t_R _27187_ (.A(_04991_),
    .B(_07273_),
    .C(_05547_),
    .Y(_10838_));
 AND3x1_ASAP7_75t_R _27188_ (.A(_05404_),
    .B(_05172_),
    .C(_05153_),
    .Y(_10839_));
 AND3x1_ASAP7_75t_R _27189_ (.A(_05173_),
    .B(_10838_),
    .C(_10839_),
    .Y(_10840_));
 AO21x1_ASAP7_75t_R _27190_ (.A1(_10815_),
    .A2(_10837_),
    .B(_10840_),
    .Y(_03831_));
 AO21x1_ASAP7_75t_R _27191_ (.A1(_10809_),
    .A2(_10810_),
    .B(_05153_),
    .Y(_10841_));
 AND4x1_ASAP7_75t_R _27192_ (.A(_05155_),
    .B(_05704_),
    .C(_10810_),
    .D(_10826_),
    .Y(_10842_));
 AO21x1_ASAP7_75t_R _27193_ (.A1(_05172_),
    .A2(_05153_),
    .B(_10842_),
    .Y(_10843_));
 AO21x1_ASAP7_75t_R _27194_ (.A1(_05706_),
    .A2(_10843_),
    .B(_10840_),
    .Y(_10844_));
 INVx1_ASAP7_75t_R _27195_ (.A(_05409_),
    .Y(_10845_));
 AO32x1_ASAP7_75t_R _27196_ (.A1(_05449_),
    .A2(_05451_),
    .A3(_10821_),
    .B1(_05164_),
    .B2(_14110_),
    .Y(_10846_));
 AND3x1_ASAP7_75t_R _27197_ (.A(_10845_),
    .B(_10834_),
    .C(_10846_),
    .Y(_10847_));
 NAND2x2_ASAP7_75t_R _27198_ (.A(_10828_),
    .B(_10822_),
    .Y(_10848_));
 NAND2x1_ASAP7_75t_R _27199_ (.A(_13234_),
    .B(_10828_),
    .Y(_10849_));
 AO21x2_ASAP7_75t_R _27200_ (.A1(_05149_),
    .A2(_05176_),
    .B(_10849_),
    .Y(_10850_));
 NAND2x1_ASAP7_75t_R _27201_ (.A(_10848_),
    .B(_10850_),
    .Y(_10851_));
 OR3x1_ASAP7_75t_R _27202_ (.A(_10844_),
    .B(_10847_),
    .C(_10851_),
    .Y(_10852_));
 AO21x1_ASAP7_75t_R _27203_ (.A1(_10829_),
    .A2(_10841_),
    .B(_10852_),
    .Y(_03832_));
 INVx1_ASAP7_75t_R _27204_ (.A(_10840_),
    .Y(_10853_));
 BUFx6f_ASAP7_75t_R _27205_ (.A(_10824_),
    .Y(_10854_));
 OR4x1_ASAP7_75t_R _27206_ (.A(\id_stage_i.controller_i.exc_req_d ),
    .B(_10854_),
    .C(_10826_),
    .D(_10822_),
    .Y(_10855_));
 OAI22x1_ASAP7_75t_R _27207_ (.A1(_05704_),
    .A2(_05154_),
    .B1(_10813_),
    .B2(_05172_),
    .Y(_10856_));
 AO21x1_ASAP7_75t_R _27208_ (.A1(_05171_),
    .A2(_05704_),
    .B(_05472_),
    .Y(_10857_));
 AO222x2_ASAP7_75t_R _27209_ (.A1(_05404_),
    .A2(_10856_),
    .B1(_10857_),
    .B2(_05172_),
    .C1(_05417_),
    .C2(_10835_),
    .Y(_10858_));
 AO21x1_ASAP7_75t_R _27210_ (.A1(_10828_),
    .A2(_10855_),
    .B(_10858_),
    .Y(_10859_));
 OA211x2_ASAP7_75t_R _27211_ (.A1(_05404_),
    .A2(_05402_),
    .B(_10853_),
    .C(_10859_),
    .Y(_03833_));
 INVx1_ASAP7_75t_R _27212_ (.A(_10855_),
    .Y(_10860_));
 INVx1_ASAP7_75t_R _27213_ (.A(_05417_),
    .Y(_10861_));
 OR3x1_ASAP7_75t_R _27214_ (.A(_05704_),
    .B(_10861_),
    .C(_10833_),
    .Y(_10862_));
 OA211x2_ASAP7_75t_R _27215_ (.A1(_05153_),
    .A2(_10812_),
    .B(_05189_),
    .C(_05154_),
    .Y(_10863_));
 AO22x1_ASAP7_75t_R _27216_ (.A1(_10828_),
    .A2(_10860_),
    .B1(_10862_),
    .B2(_10863_),
    .Y(_03834_));
 AO21x1_ASAP7_75t_R _27217_ (.A1(_05154_),
    .A2(_07273_),
    .B(_07272_),
    .Y(_10864_));
 AND4x1_ASAP7_75t_R _27218_ (.A(_05406_),
    .B(_05167_),
    .C(_05407_),
    .D(_05409_),
    .Y(_10865_));
 AOI21x1_ASAP7_75t_R _27219_ (.A1(_04991_),
    .A2(_10864_),
    .B(_10865_),
    .Y(_03835_));
 AO21x1_ASAP7_75t_R _27220_ (.A1(net166),
    .A2(_07268_),
    .B(_07639_),
    .Y(_10866_));
 AND2x2_ASAP7_75t_R _27221_ (.A(_07266_),
    .B(_10866_),
    .Y(_03836_));
 AND4x1_ASAP7_75t_R _27222_ (.A(_14135_),
    .B(_05394_),
    .C(_06891_),
    .D(_07156_),
    .Y(_10867_));
 OAI21x1_ASAP7_75t_R _27223_ (.A1(_05159_),
    .A2(_06892_),
    .B(_13294_),
    .Y(_10868_));
 OAI21x1_ASAP7_75t_R _27224_ (.A1(_06883_),
    .A2(_10867_),
    .B(_10868_),
    .Y(_03837_));
 AND3x1_ASAP7_75t_R _27225_ (.A(_14624_),
    .B(_04963_),
    .C(_05390_),
    .Y(_10869_));
 BUFx6f_ASAP7_75t_R _27226_ (.A(_10869_),
    .Y(_10870_));
 BUFx6f_ASAP7_75t_R _27227_ (.A(_10870_),
    .Y(_10871_));
 INVx2_ASAP7_75t_R _27228_ (.A(_13420_),
    .Y(_10872_));
 BUFx6f_ASAP7_75t_R _27229_ (.A(_05391_),
    .Y(_10873_));
 NOR2x1_ASAP7_75t_R _27230_ (.A(_10872_),
    .B(_10873_),
    .Y(_10874_));
 AO21x1_ASAP7_75t_R _27231_ (.A1(_05255_),
    .A2(_10871_),
    .B(_10874_),
    .Y(_10875_));
 AO21x1_ASAP7_75t_R _27232_ (.A1(_05724_),
    .A2(_08171_),
    .B(_14638_),
    .Y(_10876_));
 OA21x2_ASAP7_75t_R _27233_ (.A1(_05202_),
    .A2(_10875_),
    .B(_10876_),
    .Y(_03838_));
 NAND3x2_ASAP7_75t_R _27234_ (.B(_04963_),
    .C(_05390_),
    .Y(_10877_),
    .A(_14624_));
 BUFx6f_ASAP7_75t_R _27235_ (.A(_10877_),
    .Y(_10878_));
 AOI22x1_ASAP7_75t_R _27236_ (.A1(_15248_),
    .A2(_10873_),
    .B1(_10878_),
    .B2(_05002_),
    .Y(_10879_));
 BUFx6f_ASAP7_75t_R _27237_ (.A(_05201_),
    .Y(_10880_));
 NAND2x1_ASAP7_75t_R _27238_ (.A(_01755_),
    .B(_10880_),
    .Y(_10881_));
 OA21x2_ASAP7_75t_R _27239_ (.A1(_05202_),
    .A2(_10879_),
    .B(_10881_),
    .Y(_03839_));
 AND2x2_ASAP7_75t_R _27240_ (.A(_14260_),
    .B(_10878_),
    .Y(_10882_));
 AO21x1_ASAP7_75t_R _27241_ (.A1(\alu_adder_result_ex[11] ),
    .A2(_10871_),
    .B(_10882_),
    .Y(_10883_));
 AO21x1_ASAP7_75t_R _27242_ (.A1(_05724_),
    .A2(_08171_),
    .B(_05614_),
    .Y(_10884_));
 OA21x2_ASAP7_75t_R _27243_ (.A1(_05202_),
    .A2(_10883_),
    .B(_10884_),
    .Y(_03840_));
 NOR2x1_ASAP7_75t_R _27244_ (.A(_15363_),
    .B(_10873_),
    .Y(_10885_));
 AO21x1_ASAP7_75t_R _27245_ (.A1(\alu_adder_result_ex[12] ),
    .A2(_10871_),
    .B(_10885_),
    .Y(_10886_));
 NAND2x1_ASAP7_75t_R _27246_ (.A(_01753_),
    .B(_10880_),
    .Y(_10887_));
 OA21x2_ASAP7_75t_R _27247_ (.A1(_05202_),
    .A2(_10886_),
    .B(_10887_),
    .Y(_03841_));
 AND3x1_ASAP7_75t_R _27248_ (.A(_15465_),
    .B(_15501_),
    .C(_10878_),
    .Y(_10888_));
 AO21x1_ASAP7_75t_R _27249_ (.A1(\alu_adder_result_ex[13] ),
    .A2(_10871_),
    .B(_10888_),
    .Y(_10889_));
 NAND2x1_ASAP7_75t_R _27250_ (.A(_01752_),
    .B(_10880_),
    .Y(_10890_));
 OA21x2_ASAP7_75t_R _27251_ (.A1(_05202_),
    .A2(_10889_),
    .B(_10890_),
    .Y(_03842_));
 BUFx6f_ASAP7_75t_R _27252_ (.A(_10870_),
    .Y(_10891_));
 NOR2x1_ASAP7_75t_R _27253_ (.A(_15646_),
    .B(_10891_),
    .Y(_10892_));
 AO21x1_ASAP7_75t_R _27254_ (.A1(\alu_adder_result_ex[14] ),
    .A2(_10871_),
    .B(_10892_),
    .Y(_10893_));
 NAND2x1_ASAP7_75t_R _27255_ (.A(_01751_),
    .B(_10880_),
    .Y(_10894_));
 OA21x2_ASAP7_75t_R _27256_ (.A1(_05202_),
    .A2(_10893_),
    .B(_10894_),
    .Y(_03843_));
 NOR2x1_ASAP7_75t_R _27257_ (.A(_15759_),
    .B(_10891_),
    .Y(_10895_));
 AO21x1_ASAP7_75t_R _27258_ (.A1(\alu_adder_result_ex[15] ),
    .A2(_10871_),
    .B(_10895_),
    .Y(_10896_));
 INVx1_ASAP7_75t_R _27259_ (.A(_01750_),
    .Y(_10897_));
 AO21x1_ASAP7_75t_R _27260_ (.A1(_05724_),
    .A2(_08171_),
    .B(_10897_),
    .Y(_10898_));
 OA21x2_ASAP7_75t_R _27261_ (.A1(_05202_),
    .A2(_10896_),
    .B(_10898_),
    .Y(_03844_));
 NOR2x1_ASAP7_75t_R _27262_ (.A(_15884_),
    .B(_10891_),
    .Y(_10899_));
 AO21x1_ASAP7_75t_R _27263_ (.A1(\alu_adder_result_ex[16] ),
    .A2(_10871_),
    .B(_10899_),
    .Y(_10900_));
 AO21x1_ASAP7_75t_R _27264_ (.A1(_05724_),
    .A2(_08171_),
    .B(_05637_),
    .Y(_10901_));
 OA21x2_ASAP7_75t_R _27265_ (.A1(_05202_),
    .A2(_10900_),
    .B(_10901_),
    .Y(_03845_));
 NOR2x1_ASAP7_75t_R _27266_ (.A(_15995_),
    .B(_10870_),
    .Y(_10902_));
 AO21x1_ASAP7_75t_R _27267_ (.A1(\alu_adder_result_ex[17] ),
    .A2(_10871_),
    .B(_10902_),
    .Y(_10903_));
 NAND2x1_ASAP7_75t_R _27268_ (.A(_01748_),
    .B(_10880_),
    .Y(_10904_));
 OA21x2_ASAP7_75t_R _27269_ (.A1(_05202_),
    .A2(_10903_),
    .B(_10904_),
    .Y(_03846_));
 BUFx12f_ASAP7_75t_R _27270_ (.A(_05201_),
    .Y(_10905_));
 BUFx6f_ASAP7_75t_R _27271_ (.A(_10905_),
    .Y(_10906_));
 NOR2x1_ASAP7_75t_R _27272_ (.A(_16131_),
    .B(_10870_),
    .Y(_10907_));
 AO21x1_ASAP7_75t_R _27273_ (.A1(\alu_adder_result_ex[18] ),
    .A2(_10871_),
    .B(_10907_),
    .Y(_10908_));
 NAND2x1_ASAP7_75t_R _27274_ (.A(_01747_),
    .B(_10880_),
    .Y(_10909_));
 OA21x2_ASAP7_75t_R _27275_ (.A1(_10906_),
    .A2(_10908_),
    .B(_10909_),
    .Y(_03847_));
 AND3x1_ASAP7_75t_R _27276_ (.A(_16217_),
    .B(_16241_),
    .C(_10878_),
    .Y(_10910_));
 AO21x1_ASAP7_75t_R _27277_ (.A1(\alu_adder_result_ex[19] ),
    .A2(_10871_),
    .B(_10910_),
    .Y(_10911_));
 NAND2x1_ASAP7_75t_R _27278_ (.A(_01746_),
    .B(_10880_),
    .Y(_10912_));
 OA21x2_ASAP7_75t_R _27279_ (.A1(_10906_),
    .A2(_10911_),
    .B(_10912_),
    .Y(_03848_));
 BUFx6f_ASAP7_75t_R _27280_ (.A(_10870_),
    .Y(_10913_));
 NOR2x1_ASAP7_75t_R _27281_ (.A(_05556_),
    .B(_10873_),
    .Y(_10914_));
 AO21x1_ASAP7_75t_R _27282_ (.A1(\alu_adder_result_ex[1] ),
    .A2(_10913_),
    .B(_10914_),
    .Y(_10915_));
 NAND2x1_ASAP7_75t_R _27283_ (.A(_01745_),
    .B(_10905_),
    .Y(_10916_));
 OA21x2_ASAP7_75t_R _27284_ (.A1(_10906_),
    .A2(_10915_),
    .B(_10916_),
    .Y(_03849_));
 AND2x2_ASAP7_75t_R _27285_ (.A(_16384_),
    .B(_10878_),
    .Y(_10917_));
 AO21x1_ASAP7_75t_R _27286_ (.A1(\alu_adder_result_ex[20] ),
    .A2(_10913_),
    .B(_10917_),
    .Y(_10918_));
 AO21x1_ASAP7_75t_R _27287_ (.A1(_05724_),
    .A2(_08171_),
    .B(_05655_),
    .Y(_10919_));
 OA21x2_ASAP7_75t_R _27288_ (.A1(_10906_),
    .A2(_10918_),
    .B(_10919_),
    .Y(_03850_));
 AND2x2_ASAP7_75t_R _27289_ (.A(_16498_),
    .B(_10878_),
    .Y(_10920_));
 AO21x1_ASAP7_75t_R _27290_ (.A1(\alu_adder_result_ex[21] ),
    .A2(_10913_),
    .B(_10920_),
    .Y(_10921_));
 BUFx6f_ASAP7_75t_R _27291_ (.A(_05196_),
    .Y(_10922_));
 AO21x1_ASAP7_75t_R _27292_ (.A1(_05724_),
    .A2(_10922_),
    .B(_05660_),
    .Y(_10923_));
 OA21x2_ASAP7_75t_R _27293_ (.A1(_10906_),
    .A2(_10921_),
    .B(_10923_),
    .Y(_03851_));
 NOR2x1_ASAP7_75t_R _27294_ (.A(_16637_),
    .B(_10870_),
    .Y(_10924_));
 AO21x1_ASAP7_75t_R _27295_ (.A1(\alu_adder_result_ex[22] ),
    .A2(_10913_),
    .B(_10924_),
    .Y(_10925_));
 NAND2x1_ASAP7_75t_R _27296_ (.A(_01742_),
    .B(_10905_),
    .Y(_10926_));
 OA21x2_ASAP7_75t_R _27297_ (.A1(_10906_),
    .A2(_10925_),
    .B(_10926_),
    .Y(_03852_));
 AND3x1_ASAP7_75t_R _27298_ (.A(_16723_),
    .B(_16746_),
    .C(_10877_),
    .Y(_10927_));
 AO21x1_ASAP7_75t_R _27299_ (.A1(\alu_adder_result_ex[23] ),
    .A2(_10913_),
    .B(_10927_),
    .Y(_10928_));
 NAND2x1_ASAP7_75t_R _27300_ (.A(_01741_),
    .B(_10905_),
    .Y(_10929_));
 OA21x2_ASAP7_75t_R _27301_ (.A1(_10906_),
    .A2(_10928_),
    .B(_10929_),
    .Y(_03853_));
 AND2x2_ASAP7_75t_R _27302_ (.A(_16870_),
    .B(_10878_),
    .Y(_10930_));
 AO21x1_ASAP7_75t_R _27303_ (.A1(\alu_adder_result_ex[24] ),
    .A2(_10913_),
    .B(_10930_),
    .Y(_10931_));
 AO21x1_ASAP7_75t_R _27304_ (.A1(_05724_),
    .A2(_10922_),
    .B(_05673_),
    .Y(_10932_));
 OA21x2_ASAP7_75t_R _27305_ (.A1(_10906_),
    .A2(_10931_),
    .B(_10932_),
    .Y(_03854_));
 AND3x1_ASAP7_75t_R _27306_ (.A(_16959_),
    .B(_16982_),
    .C(_10877_),
    .Y(_10933_));
 AO21x1_ASAP7_75t_R _27307_ (.A1(\alu_adder_result_ex[25] ),
    .A2(_10913_),
    .B(_10933_),
    .Y(_10934_));
 AO21x1_ASAP7_75t_R _27308_ (.A1(_05724_),
    .A2(_10922_),
    .B(_05677_),
    .Y(_10935_));
 OA21x2_ASAP7_75t_R _27309_ (.A1(_10906_),
    .A2(_10934_),
    .B(_10935_),
    .Y(_03855_));
 AND3x1_ASAP7_75t_R _27310_ (.A(_04333_),
    .B(_04356_),
    .C(_10877_),
    .Y(_10936_));
 AO21x1_ASAP7_75t_R _27311_ (.A1(\alu_adder_result_ex[26] ),
    .A2(_10913_),
    .B(_10936_),
    .Y(_10937_));
 AO21x1_ASAP7_75t_R _27312_ (.A1(_05724_),
    .A2(_10922_),
    .B(_05681_),
    .Y(_10938_));
 OA21x2_ASAP7_75t_R _27313_ (.A1(_10906_),
    .A2(_10937_),
    .B(_10938_),
    .Y(_03856_));
 BUFx6f_ASAP7_75t_R _27314_ (.A(_05201_),
    .Y(_10939_));
 INVx3_ASAP7_75t_R _27315_ (.A(_05391_),
    .Y(_10940_));
 AND3x1_ASAP7_75t_R _27316_ (.A(_04444_),
    .B(_04467_),
    .C(_10940_),
    .Y(_10941_));
 AO21x1_ASAP7_75t_R _27317_ (.A1(\alu_adder_result_ex[27] ),
    .A2(_10913_),
    .B(_10941_),
    .Y(_10942_));
 NAND2x1_ASAP7_75t_R _27318_ (.A(_01737_),
    .B(_10905_),
    .Y(_10943_));
 OA21x2_ASAP7_75t_R _27319_ (.A1(_10939_),
    .A2(_10942_),
    .B(_10943_),
    .Y(_03857_));
 AND3x1_ASAP7_75t_R _27320_ (.A(_04581_),
    .B(_04604_),
    .C(_10877_),
    .Y(_10944_));
 AO21x1_ASAP7_75t_R _27321_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_10913_),
    .B(_10944_),
    .Y(_10945_));
 AO21x1_ASAP7_75t_R _27322_ (.A1(_05200_),
    .A2(_10922_),
    .B(_05689_),
    .Y(_10946_));
 OA21x2_ASAP7_75t_R _27323_ (.A1(_10939_),
    .A2(_10945_),
    .B(_10946_),
    .Y(_03858_));
 AND3x1_ASAP7_75t_R _27324_ (.A(_04693_),
    .B(_04716_),
    .C(_10877_),
    .Y(_10947_));
 AO21x1_ASAP7_75t_R _27325_ (.A1(\alu_adder_result_ex[29] ),
    .A2(_10891_),
    .B(_10947_),
    .Y(_10948_));
 AO21x1_ASAP7_75t_R _27326_ (.A1(_05200_),
    .A2(_10922_),
    .B(_05693_),
    .Y(_10949_));
 OA21x2_ASAP7_75t_R _27327_ (.A1(_10939_),
    .A2(_10948_),
    .B(_10949_),
    .Y(_03859_));
 AND2x2_ASAP7_75t_R _27328_ (.A(_13601_),
    .B(_10878_),
    .Y(_10950_));
 AO21x1_ASAP7_75t_R _27329_ (.A1(\alu_adder_result_ex[2] ),
    .A2(_10891_),
    .B(_10950_),
    .Y(_10951_));
 AO21x1_ASAP7_75t_R _27330_ (.A1(_05200_),
    .A2(_10922_),
    .B(_05568_),
    .Y(_10952_));
 OA21x2_ASAP7_75t_R _27331_ (.A1(_10939_),
    .A2(_10951_),
    .B(_10952_),
    .Y(_03860_));
 AND3x1_ASAP7_75t_R _27332_ (.A(_04813_),
    .B(_04836_),
    .C(_10877_),
    .Y(_10953_));
 AO21x1_ASAP7_75t_R _27333_ (.A1(\alu_adder_result_ex[30] ),
    .A2(_10891_),
    .B(_10953_),
    .Y(_10954_));
 NAND2x1_ASAP7_75t_R _27334_ (.A(_01733_),
    .B(_10905_),
    .Y(_10955_));
 OA21x2_ASAP7_75t_R _27335_ (.A1(_10939_),
    .A2(_10954_),
    .B(_10955_),
    .Y(_03861_));
 NAND2x1_ASAP7_75t_R _27336_ (.A(_15236_),
    .B(_05390_),
    .Y(_10956_));
 OA21x2_ASAP7_75t_R _27337_ (.A1(net1961),
    .A2(_10956_),
    .B(_04963_),
    .Y(_10957_));
 AO21x1_ASAP7_75t_R _27338_ (.A1(_05200_),
    .A2(_10922_),
    .B(_08207_),
    .Y(_10958_));
 OA21x2_ASAP7_75t_R _27339_ (.A1(_10939_),
    .A2(_10957_),
    .B(_10958_),
    .Y(_03862_));
 BUFx6f_ASAP7_75t_R _27340_ (.A(_02198_),
    .Y(_10959_));
 BUFx6f_ASAP7_75t_R _27341_ (.A(_10959_),
    .Y(_10960_));
 NAND2x1_ASAP7_75t_R _27342_ (.A(_05720_),
    .B(_08060_),
    .Y(_10961_));
 BUFx6f_ASAP7_75t_R _27343_ (.A(_10961_),
    .Y(_10962_));
 BUFx6f_ASAP7_75t_R _27344_ (.A(_08208_),
    .Y(_10963_));
 NOR2x1_ASAP7_75t_R _27345_ (.A(_05255_),
    .B(_08223_),
    .Y(_10964_));
 AO21x1_ASAP7_75t_R _27346_ (.A1(_00062_),
    .A2(_10963_),
    .B(_10964_),
    .Y(_10965_));
 AND3x4_ASAP7_75t_R _27347_ (.A(_13262_),
    .B(_15234_),
    .C(_08060_),
    .Y(_10966_));
 BUFx6f_ASAP7_75t_R _27348_ (.A(_10966_),
    .Y(_10967_));
 OA211x2_ASAP7_75t_R _27349_ (.A1(_08078_),
    .A2(_08210_),
    .B(_10967_),
    .C(_00028_),
    .Y(_10968_));
 AO21x1_ASAP7_75t_R _27350_ (.A1(_10962_),
    .A2(_10965_),
    .B(_10968_),
    .Y(_10969_));
 OR3x2_ASAP7_75t_R _27351_ (.A(_14639_),
    .B(_05200_),
    .C(_14641_),
    .Y(_10970_));
 BUFx6f_ASAP7_75t_R _27352_ (.A(_10970_),
    .Y(_10971_));
 BUFx6f_ASAP7_75t_R _27353_ (.A(_10971_),
    .Y(_10972_));
 NAND2x1_ASAP7_75t_R _27354_ (.A(_05559_),
    .B(_05255_),
    .Y(_10973_));
 OA211x2_ASAP7_75t_R _27355_ (.A1(_00095_),
    .A2(_02193_),
    .B(_10972_),
    .C(_10973_),
    .Y(_10974_));
 XOR2x2_ASAP7_75t_R _27356_ (.A(_05186_),
    .B(_02238_),
    .Y(_10975_));
 BUFx6f_ASAP7_75t_R _27357_ (.A(_08068_),
    .Y(_10976_));
 BUFx6f_ASAP7_75t_R _27358_ (.A(_02237_),
    .Y(_10977_));
 NAND2x1_ASAP7_75t_R _27359_ (.A(_10977_),
    .B(_00080_),
    .Y(_10978_));
 OA211x2_ASAP7_75t_R _27360_ (.A1(_10976_),
    .A2(_08106_),
    .B(_10978_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_10979_));
 NAND2x1_ASAP7_75t_R _27361_ (.A(_10977_),
    .B(_00079_),
    .Y(_10980_));
 OA211x2_ASAP7_75t_R _27362_ (.A1(_10976_),
    .A2(_08110_),
    .B(_10980_),
    .C(_05254_),
    .Y(_10981_));
 OR3x1_ASAP7_75t_R _27363_ (.A(_08075_),
    .B(_10979_),
    .C(_10981_),
    .Y(_10982_));
 XNOR2x2_ASAP7_75t_R _27364_ (.A(_05187_),
    .B(_08074_),
    .Y(_10983_));
 NAND2x1_ASAP7_75t_R _27365_ (.A(_10977_),
    .B(_00072_),
    .Y(_10984_));
 OA211x2_ASAP7_75t_R _27366_ (.A1(_10976_),
    .A2(_08187_),
    .B(_10984_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_10985_));
 NAND2x1_ASAP7_75t_R _27367_ (.A(_10977_),
    .B(_00071_),
    .Y(_10986_));
 OA211x2_ASAP7_75t_R _27368_ (.A1(_10976_),
    .A2(_08191_),
    .B(_10986_),
    .C(_05254_),
    .Y(_10987_));
 OR3x1_ASAP7_75t_R _27369_ (.A(_10983_),
    .B(_10985_),
    .C(_10987_),
    .Y(_10988_));
 AND3x1_ASAP7_75t_R _27370_ (.A(_10975_),
    .B(_10982_),
    .C(_10988_),
    .Y(_10989_));
 NAND2x1_ASAP7_75t_R _27371_ (.A(_10977_),
    .B(_00076_),
    .Y(_10990_));
 OA211x2_ASAP7_75t_R _27372_ (.A1(_10976_),
    .A2(_08201_),
    .B(_10990_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_10991_));
 NAND2x1_ASAP7_75t_R _27373_ (.A(_10977_),
    .B(_00075_),
    .Y(_10992_));
 OA211x2_ASAP7_75t_R _27374_ (.A1(_10976_),
    .A2(_08205_),
    .B(_10992_),
    .C(_05254_),
    .Y(_10993_));
 OR3x1_ASAP7_75t_R _27375_ (.A(_08075_),
    .B(_10991_),
    .C(_10993_),
    .Y(_10994_));
 NAND2x1_ASAP7_75t_R _27376_ (.A(_00068_),
    .B(_10976_),
    .Y(_10995_));
 OA211x2_ASAP7_75t_R _27377_ (.A1(_08093_),
    .A2(_10976_),
    .B(_10995_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_10996_));
 NAND2x1_ASAP7_75t_R _27378_ (.A(_00067_),
    .B(_10976_),
    .Y(_10997_));
 OA211x2_ASAP7_75t_R _27379_ (.A1(_08134_),
    .A2(_10976_),
    .B(_10997_),
    .C(_05254_),
    .Y(_10998_));
 OR3x1_ASAP7_75t_R _27380_ (.A(_10983_),
    .B(_10996_),
    .C(_10998_),
    .Y(_10999_));
 AND3x1_ASAP7_75t_R _27381_ (.A(_08071_),
    .B(_10994_),
    .C(_10999_),
    .Y(_11000_));
 XNOR2x2_ASAP7_75t_R _27382_ (.A(_08081_),
    .B(_08082_),
    .Y(_11001_));
 OAI21x1_ASAP7_75t_R _27383_ (.A1(_10989_),
    .A2(_11000_),
    .B(_11001_),
    .Y(_11002_));
 AND2x2_ASAP7_75t_R _27384_ (.A(_08068_),
    .B(_00096_),
    .Y(_11003_));
 AO21x1_ASAP7_75t_R _27385_ (.A1(_08069_),
    .A2(_00094_),
    .B(_11003_),
    .Y(_11004_));
 NAND2x1_ASAP7_75t_R _27386_ (.A(_08068_),
    .B(_00095_),
    .Y(_11005_));
 OA211x2_ASAP7_75t_R _27387_ (.A1(_10977_),
    .A2(_08172_),
    .B(_11005_),
    .C(_18083_),
    .Y(_11006_));
 INVx1_ASAP7_75t_R _27388_ (.A(_11006_),
    .Y(_11007_));
 OA211x2_ASAP7_75t_R _27389_ (.A1(_05254_),
    .A2(_11004_),
    .B(_11007_),
    .C(_10983_),
    .Y(_11008_));
 AND2x2_ASAP7_75t_R _27390_ (.A(_08068_),
    .B(_00088_),
    .Y(_11009_));
 AO21x1_ASAP7_75t_R _27391_ (.A1(_08069_),
    .A2(_00086_),
    .B(_11009_),
    .Y(_11010_));
 NAND2x1_ASAP7_75t_R _27392_ (.A(_08068_),
    .B(_00087_),
    .Y(_11011_));
 OA211x2_ASAP7_75t_R _27393_ (.A1(_10977_),
    .A2(_08142_),
    .B(_11011_),
    .C(_18083_),
    .Y(_11012_));
 INVx1_ASAP7_75t_R _27394_ (.A(_11012_),
    .Y(_11013_));
 OA211x2_ASAP7_75t_R _27395_ (.A1(_05254_),
    .A2(_11010_),
    .B(_11013_),
    .C(_08075_),
    .Y(_11014_));
 OR3x1_ASAP7_75t_R _27396_ (.A(_08071_),
    .B(_11008_),
    .C(_11014_),
    .Y(_11015_));
 AND2x2_ASAP7_75t_R _27397_ (.A(_08068_),
    .B(_00092_),
    .Y(_11016_));
 AO21x1_ASAP7_75t_R _27398_ (.A1(_08069_),
    .A2(_00090_),
    .B(_11016_),
    .Y(_11017_));
 NAND2x1_ASAP7_75t_R _27399_ (.A(_08068_),
    .B(_00091_),
    .Y(_11018_));
 OA211x2_ASAP7_75t_R _27400_ (.A1(_10977_),
    .A2(_08157_),
    .B(_11018_),
    .C(_18083_),
    .Y(_11019_));
 INVx1_ASAP7_75t_R _27401_ (.A(_11019_),
    .Y(_11020_));
 OA211x2_ASAP7_75t_R _27402_ (.A1(_05254_),
    .A2(_11017_),
    .B(_11020_),
    .C(_10983_),
    .Y(_11021_));
 AND2x2_ASAP7_75t_R _27403_ (.A(_08068_),
    .B(_00084_),
    .Y(_11022_));
 AO21x1_ASAP7_75t_R _27404_ (.A1(_08069_),
    .A2(_00082_),
    .B(_11022_),
    .Y(_11023_));
 NAND2x1_ASAP7_75t_R _27405_ (.A(_08068_),
    .B(_00083_),
    .Y(_11024_));
 OA211x2_ASAP7_75t_R _27406_ (.A1(_10977_),
    .A2(_08123_),
    .B(_11024_),
    .C(_18083_),
    .Y(_11025_));
 INVx1_ASAP7_75t_R _27407_ (.A(_11025_),
    .Y(_11026_));
 OA211x2_ASAP7_75t_R _27408_ (.A1(_05254_),
    .A2(_11023_),
    .B(_11026_),
    .C(_08075_),
    .Y(_11027_));
 OR3x1_ASAP7_75t_R _27409_ (.A(_10975_),
    .B(_11021_),
    .C(_11027_),
    .Y(_11028_));
 AO21x1_ASAP7_75t_R _27410_ (.A1(_11015_),
    .A2(_11028_),
    .B(_11001_),
    .Y(_11029_));
 AO21x1_ASAP7_75t_R _27411_ (.A1(_11002_),
    .A2(_11029_),
    .B(_08219_),
    .Y(_11030_));
 OA211x2_ASAP7_75t_R _27412_ (.A1(_10960_),
    .A2(_10969_),
    .B(_10974_),
    .C(_11030_),
    .Y(_11031_));
 OR2x2_ASAP7_75t_R _27413_ (.A(_10966_),
    .B(_10970_),
    .Y(_11032_));
 BUFx6f_ASAP7_75t_R _27414_ (.A(_11032_),
    .Y(_11033_));
 BUFx6f_ASAP7_75t_R _27415_ (.A(_11033_),
    .Y(_11034_));
 AND3x4_ASAP7_75t_R _27416_ (.A(_00753_),
    .B(_02193_),
    .C(_14628_),
    .Y(_11035_));
 AND3x1_ASAP7_75t_R _27417_ (.A(_13262_),
    .B(_02192_),
    .C(_11035_),
    .Y(_11036_));
 AND3x1_ASAP7_75t_R _27418_ (.A(_08086_),
    .B(_05391_),
    .C(_10966_),
    .Y(_11037_));
 AO21x1_ASAP7_75t_R _27419_ (.A1(_05350_),
    .A2(_10940_),
    .B(_11037_),
    .Y(_11038_));
 OR3x1_ASAP7_75t_R _27420_ (.A(_14533_),
    .B(_14636_),
    .C(_08568_),
    .Y(_11039_));
 AOI221x1_ASAP7_75t_R _27421_ (.A1(_05350_),
    .A2(_10961_),
    .B1(_11038_),
    .B2(_01799_),
    .C(_11039_),
    .Y(_11040_));
 OR4x1_ASAP7_75t_R _27422_ (.A(_08568_),
    .B(_06905_),
    .C(_11036_),
    .D(_11040_),
    .Y(_11041_));
 BUFx12f_ASAP7_75t_R _27423_ (.A(_11041_),
    .Y(_11042_));
 NOR2x1_ASAP7_75t_R _27424_ (.A(_09037_),
    .B(_11042_),
    .Y(_11043_));
 BUFx6f_ASAP7_75t_R _27425_ (.A(_11043_),
    .Y(_11044_));
 OAI21x1_ASAP7_75t_R _27426_ (.A1(_14635_),
    .A2(_11034_),
    .B(_11044_),
    .Y(_11045_));
 OR2x6_ASAP7_75t_R _27427_ (.A(_09059_),
    .B(_11042_),
    .Y(_11046_));
 BUFx6f_ASAP7_75t_R _27428_ (.A(_11046_),
    .Y(_11047_));
 NAND2x1_ASAP7_75t_R _27429_ (.A(_14534_),
    .B(_15235_),
    .Y(_11048_));
 BUFx6f_ASAP7_75t_R _27430_ (.A(_11048_),
    .Y(_11049_));
 NOR2x2_ASAP7_75t_R _27431_ (.A(_09060_),
    .B(_11042_),
    .Y(_11050_));
 OA21x2_ASAP7_75t_R _27432_ (.A1(_00064_),
    .A2(_11049_),
    .B(_11050_),
    .Y(_11051_));
 AO21x1_ASAP7_75t_R _27433_ (.A1(_00062_),
    .A2(_11047_),
    .B(_11051_),
    .Y(_11052_));
 OAI21x1_ASAP7_75t_R _27434_ (.A1(_11031_),
    .A2(_11045_),
    .B(_11052_),
    .Y(_03863_));
 NOR2x1_ASAP7_75t_R _27435_ (.A(_10967_),
    .B(_10971_),
    .Y(_11053_));
 NOR2x1_ASAP7_75t_R _27436_ (.A(\alu_adder_result_ex[1] ),
    .B(_08223_),
    .Y(_11054_));
 AO21x1_ASAP7_75t_R _27437_ (.A1(_00097_),
    .A2(_10963_),
    .B(_11054_),
    .Y(_11055_));
 AND2x2_ASAP7_75t_R _27438_ (.A(_00030_),
    .B(_08061_),
    .Y(_11056_));
 AO221x1_ASAP7_75t_R _27439_ (.A1(_10961_),
    .A2(_11055_),
    .B1(_11056_),
    .B2(_08243_),
    .C(_10959_),
    .Y(_11057_));
 OA21x2_ASAP7_75t_R _27440_ (.A1(_14636_),
    .A2(_18712_),
    .B(_10970_),
    .Y(_11058_));
 OA21x2_ASAP7_75t_R _27441_ (.A1(_05197_),
    .A2(_10965_),
    .B(_11058_),
    .Y(_11059_));
 AO221x1_ASAP7_75t_R _27442_ (.A1(_14528_),
    .A2(_11053_),
    .B1(_11057_),
    .B2(_11059_),
    .C(_09037_),
    .Y(_11060_));
 OA211x2_ASAP7_75t_R _27443_ (.A1(_00099_),
    .A2(_11049_),
    .B(_11050_),
    .C(_11060_),
    .Y(_11061_));
 AOI21x1_ASAP7_75t_R _27444_ (.A1(_00097_),
    .A2(_11047_),
    .B(_11061_),
    .Y(_03864_));
 BUFx6f_ASAP7_75t_R _27445_ (.A(_10962_),
    .Y(_11062_));
 BUFx6f_ASAP7_75t_R _27446_ (.A(_08223_),
    .Y(_11063_));
 BUFx6f_ASAP7_75t_R _27447_ (.A(_11063_),
    .Y(_11064_));
 NOR2x1_ASAP7_75t_R _27448_ (.A(\alu_adder_result_ex[2] ),
    .B(_11064_),
    .Y(_11065_));
 AO21x1_ASAP7_75t_R _27449_ (.A1(_00100_),
    .A2(_11064_),
    .B(_11065_),
    .Y(_11066_));
 BUFx3_ASAP7_75t_R _27450_ (.A(_10966_),
    .Y(_11067_));
 BUFx6f_ASAP7_75t_R _27451_ (.A(_11067_),
    .Y(_11068_));
 OA211x2_ASAP7_75t_R _27452_ (.A1(_08078_),
    .A2(_08218_),
    .B(_11068_),
    .C(_00031_),
    .Y(_11069_));
 AO21x1_ASAP7_75t_R _27453_ (.A1(_11062_),
    .A2(_11066_),
    .B(_11069_),
    .Y(_11070_));
 OA21x2_ASAP7_75t_R _27454_ (.A1(_05252_),
    .A2(_05219_),
    .B(_10972_),
    .Y(_11071_));
 OA21x2_ASAP7_75t_R _27455_ (.A1(_05198_),
    .A2(_11055_),
    .B(_11071_),
    .Y(_11072_));
 OAI21x1_ASAP7_75t_R _27456_ (.A1(_10960_),
    .A2(_11070_),
    .B(_11072_),
    .Y(_11073_));
 OA21x2_ASAP7_75t_R _27457_ (.A1(_14703_),
    .A2(_11034_),
    .B(_11044_),
    .Y(_11074_));
 BUFx6f_ASAP7_75t_R _27458_ (.A(_11050_),
    .Y(_11075_));
 OR3x1_ASAP7_75t_R _27459_ (.A(_00103_),
    .B(_11049_),
    .C(_11047_),
    .Y(_11076_));
 OAI21x1_ASAP7_75t_R _27460_ (.A1(_00100_),
    .A2(_11075_),
    .B(_11076_),
    .Y(_11077_));
 AO21x1_ASAP7_75t_R _27461_ (.A1(_11073_),
    .A2(_11074_),
    .B(_11077_),
    .Y(_03865_));
 NOR2x1_ASAP7_75t_R _27462_ (.A(\alu_adder_result_ex[3] ),
    .B(_11064_),
    .Y(_11078_));
 AO21x1_ASAP7_75t_R _27463_ (.A1(_00104_),
    .A2(_11064_),
    .B(_11078_),
    .Y(_11079_));
 OA211x2_ASAP7_75t_R _27464_ (.A1(_08078_),
    .A2(_08225_),
    .B(_11068_),
    .C(_00033_),
    .Y(_11080_));
 AO21x1_ASAP7_75t_R _27465_ (.A1(_11062_),
    .A2(_11079_),
    .B(_11080_),
    .Y(_11081_));
 OA21x2_ASAP7_75t_R _27466_ (.A1(_05252_),
    .A2(_05214_),
    .B(_10972_),
    .Y(_11082_));
 OA21x2_ASAP7_75t_R _27467_ (.A1(_05198_),
    .A2(_11066_),
    .B(_11082_),
    .Y(_11083_));
 OAI21x1_ASAP7_75t_R _27468_ (.A1(_10960_),
    .A2(_11081_),
    .B(_11083_),
    .Y(_11084_));
 OA21x2_ASAP7_75t_R _27469_ (.A1(_14770_),
    .A2(_11034_),
    .B(_11044_),
    .Y(_11085_));
 OR3x1_ASAP7_75t_R _27470_ (.A(_00108_),
    .B(_11049_),
    .C(_11047_),
    .Y(_11086_));
 OAI21x1_ASAP7_75t_R _27471_ (.A1(_00104_),
    .A2(_11075_),
    .B(_11086_),
    .Y(_11087_));
 AO21x1_ASAP7_75t_R _27472_ (.A1(_11084_),
    .A2(_11085_),
    .B(_11087_),
    .Y(_03866_));
 NOR2x1_ASAP7_75t_R _27473_ (.A(\alu_adder_result_ex[4] ),
    .B(_11064_),
    .Y(_11088_));
 AO21x1_ASAP7_75t_R _27474_ (.A1(_00109_),
    .A2(_11064_),
    .B(_11088_),
    .Y(_11089_));
 OA211x2_ASAP7_75t_R _27475_ (.A1(_08210_),
    .A2(_08246_),
    .B(_00034_),
    .C(_11068_),
    .Y(_11090_));
 AO21x1_ASAP7_75t_R _27476_ (.A1(_11062_),
    .A2(_11089_),
    .B(_11090_),
    .Y(_11091_));
 OA21x2_ASAP7_75t_R _27477_ (.A1(_05252_),
    .A2(_05226_),
    .B(_10972_),
    .Y(_11092_));
 OA21x2_ASAP7_75t_R _27478_ (.A1(_05198_),
    .A2(_11079_),
    .B(_11092_),
    .Y(_11093_));
 OAI21x1_ASAP7_75t_R _27479_ (.A1(_10960_),
    .A2(_11091_),
    .B(_11093_),
    .Y(_11094_));
 OA21x2_ASAP7_75t_R _27480_ (.A1(_14835_),
    .A2(_11034_),
    .B(_11044_),
    .Y(_11095_));
 OR3x1_ASAP7_75t_R _27481_ (.A(_00113_),
    .B(_11049_),
    .C(_11047_),
    .Y(_11096_));
 OAI21x1_ASAP7_75t_R _27482_ (.A1(_00109_),
    .A2(_11075_),
    .B(_11096_),
    .Y(_11097_));
 AO21x1_ASAP7_75t_R _27483_ (.A1(_11094_),
    .A2(_11095_),
    .B(_11097_),
    .Y(_03867_));
 NOR2x1_ASAP7_75t_R _27484_ (.A(\alu_adder_result_ex[5] ),
    .B(_11064_),
    .Y(_11098_));
 AO21x1_ASAP7_75t_R _27485_ (.A1(_00114_),
    .A2(_11064_),
    .B(_11098_),
    .Y(_11099_));
 OA211x2_ASAP7_75t_R _27486_ (.A1(_08230_),
    .A2(_08246_),
    .B(_00035_),
    .C(_11068_),
    .Y(_11100_));
 AO21x1_ASAP7_75t_R _27487_ (.A1(_11062_),
    .A2(_11099_),
    .B(_11100_),
    .Y(_11101_));
 OA21x2_ASAP7_75t_R _27488_ (.A1(_05252_),
    .A2(_05212_),
    .B(_10972_),
    .Y(_11102_));
 OA21x2_ASAP7_75t_R _27489_ (.A1(_05198_),
    .A2(_11089_),
    .B(_11102_),
    .Y(_11103_));
 OAI21x1_ASAP7_75t_R _27490_ (.A1(_10960_),
    .A2(_11101_),
    .B(_11103_),
    .Y(_11104_));
 OA21x2_ASAP7_75t_R _27491_ (.A1(_05583_),
    .A2(_11034_),
    .B(_11044_),
    .Y(_11105_));
 OR3x1_ASAP7_75t_R _27492_ (.A(_00120_),
    .B(_11049_),
    .C(_11047_),
    .Y(_11106_));
 OAI21x1_ASAP7_75t_R _27493_ (.A1(_00114_),
    .A2(_11075_),
    .B(_11106_),
    .Y(_11107_));
 AO21x1_ASAP7_75t_R _27494_ (.A1(_11104_),
    .A2(_11105_),
    .B(_11107_),
    .Y(_03868_));
 OR2x2_ASAP7_75t_R _27495_ (.A(_13684_),
    .B(_10873_),
    .Y(_11108_));
 OA21x2_ASAP7_75t_R _27496_ (.A1(\alu_adder_result_ex[3] ),
    .A2(_10940_),
    .B(_11108_),
    .Y(_11109_));
 NAND2x1_ASAP7_75t_R _27497_ (.A(_01731_),
    .B(_10905_),
    .Y(_11110_));
 OA21x2_ASAP7_75t_R _27498_ (.A1(_10939_),
    .A2(_11109_),
    .B(_11110_),
    .Y(_03869_));
 BUFx6f_ASAP7_75t_R _27499_ (.A(_08223_),
    .Y(_11111_));
 NOR2x1_ASAP7_75t_R _27500_ (.A(\alu_adder_result_ex[6] ),
    .B(_11111_),
    .Y(_11112_));
 AO21x1_ASAP7_75t_R _27501_ (.A1(_00121_),
    .A2(_11064_),
    .B(_11112_),
    .Y(_11113_));
 OA211x2_ASAP7_75t_R _27502_ (.A1(_08218_),
    .A2(_08246_),
    .B(_00036_),
    .C(_11068_),
    .Y(_11114_));
 AO21x1_ASAP7_75t_R _27503_ (.A1(_11062_),
    .A2(_11113_),
    .B(_11114_),
    .Y(_11115_));
 OA21x2_ASAP7_75t_R _27504_ (.A1(_05252_),
    .A2(_05207_),
    .B(_10972_),
    .Y(_11116_));
 OA21x2_ASAP7_75t_R _27505_ (.A1(_05198_),
    .A2(_11099_),
    .B(_11116_),
    .Y(_11117_));
 OAI21x1_ASAP7_75t_R _27506_ (.A1(_10960_),
    .A2(_11115_),
    .B(_11117_),
    .Y(_11118_));
 OA21x2_ASAP7_75t_R _27507_ (.A1(_05303_),
    .A2(_11034_),
    .B(_11044_),
    .Y(_11119_));
 OR3x1_ASAP7_75t_R _27508_ (.A(_00127_),
    .B(_11048_),
    .C(_11047_),
    .Y(_11120_));
 OAI21x1_ASAP7_75t_R _27509_ (.A1(_00121_),
    .A2(_11075_),
    .B(_11120_),
    .Y(_11121_));
 AO21x1_ASAP7_75t_R _27510_ (.A1(_11118_),
    .A2(_11119_),
    .B(_11121_),
    .Y(_03870_));
 BUFx6f_ASAP7_75t_R _27511_ (.A(_08223_),
    .Y(_11122_));
 NOR2x1_ASAP7_75t_R _27512_ (.A(\alu_adder_result_ex[7] ),
    .B(_11063_),
    .Y(_11123_));
 AO21x1_ASAP7_75t_R _27513_ (.A1(_00128_),
    .A2(_11122_),
    .B(_11123_),
    .Y(_11124_));
 OA211x2_ASAP7_75t_R _27514_ (.A1(_08225_),
    .A2(_08246_),
    .B(_00037_),
    .C(_11068_),
    .Y(_11125_));
 AO21x1_ASAP7_75t_R _27515_ (.A1(_11062_),
    .A2(_11124_),
    .B(_11125_),
    .Y(_11126_));
 OA21x2_ASAP7_75t_R _27516_ (.A1(_05252_),
    .A2(_15040_),
    .B(_10972_),
    .Y(_11127_));
 OA21x2_ASAP7_75t_R _27517_ (.A1(_05198_),
    .A2(_11113_),
    .B(_11127_),
    .Y(_11128_));
 OAI21x1_ASAP7_75t_R _27518_ (.A1(_10960_),
    .A2(_11126_),
    .B(_11128_),
    .Y(_11129_));
 OA21x2_ASAP7_75t_R _27519_ (.A1(_05595_),
    .A2(_11034_),
    .B(_11044_),
    .Y(_11130_));
 AND3x1_ASAP7_75t_R _27520_ (.A(_02209_),
    .B(_05242_),
    .C(_11050_),
    .Y(_11131_));
 AO21x1_ASAP7_75t_R _27521_ (.A1(_15027_),
    .A2(_11047_),
    .B(_11131_),
    .Y(_11132_));
 AO21x1_ASAP7_75t_R _27522_ (.A1(_11129_),
    .A2(_11130_),
    .B(_11132_),
    .Y(_03871_));
 BUFx6f_ASAP7_75t_R _27523_ (.A(_11042_),
    .Y(_11133_));
 INVx1_ASAP7_75t_R _27524_ (.A(_08500_),
    .Y(_11134_));
 NOR2x1_ASAP7_75t_R _27525_ (.A(\alu_adder_result_ex[8] ),
    .B(_11063_),
    .Y(_11135_));
 AO21x1_ASAP7_75t_R _27526_ (.A1(_00135_),
    .A2(_11111_),
    .B(_11135_),
    .Y(_11136_));
 OA211x2_ASAP7_75t_R _27527_ (.A1(_08210_),
    .A2(_08220_),
    .B(_00038_),
    .C(_11067_),
    .Y(_11137_));
 AO21x1_ASAP7_75t_R _27528_ (.A1(_10962_),
    .A2(_11136_),
    .B(_11137_),
    .Y(_11138_));
 OA211x2_ASAP7_75t_R _27529_ (.A1(_14636_),
    .A2(_15179_),
    .B(_10970_),
    .C(_14541_),
    .Y(_11139_));
 OA21x2_ASAP7_75t_R _27530_ (.A1(_05197_),
    .A2(_11124_),
    .B(_11139_),
    .Y(_11140_));
 OAI21x1_ASAP7_75t_R _27531_ (.A1(_10959_),
    .A2(_11138_),
    .B(_11140_),
    .Y(_11141_));
 OR3x1_ASAP7_75t_R _27532_ (.A(_14534_),
    .B(_15098_),
    .C(_11033_),
    .Y(_11142_));
 AND4x1_ASAP7_75t_R _27533_ (.A(_15236_),
    .B(_11134_),
    .C(_11141_),
    .D(_11142_),
    .Y(_11143_));
 BUFx6f_ASAP7_75t_R _27534_ (.A(_11042_),
    .Y(_11144_));
 NAND2x1_ASAP7_75t_R _27535_ (.A(_00135_),
    .B(_11144_),
    .Y(_11145_));
 OA21x2_ASAP7_75t_R _27536_ (.A1(_11133_),
    .A2(_11143_),
    .B(_11145_),
    .Y(_03872_));
 NOR2x1_ASAP7_75t_R _27537_ (.A(\alu_adder_result_ex[9] ),
    .B(_08223_),
    .Y(_11146_));
 AO21x1_ASAP7_75t_R _27538_ (.A1(_00144_),
    .A2(_11063_),
    .B(_11146_),
    .Y(_11147_));
 OA211x2_ASAP7_75t_R _27539_ (.A1(_08220_),
    .A2(_08230_),
    .B(_00039_),
    .C(_10967_),
    .Y(_11148_));
 AO21x1_ASAP7_75t_R _27540_ (.A1(_11062_),
    .A2(_11147_),
    .B(_11148_),
    .Y(_11149_));
 OA21x2_ASAP7_75t_R _27541_ (.A1(_05252_),
    .A2(_15166_),
    .B(_10972_),
    .Y(_11150_));
 OA21x2_ASAP7_75t_R _27542_ (.A1(_05198_),
    .A2(_11136_),
    .B(_11150_),
    .Y(_11151_));
 OAI21x1_ASAP7_75t_R _27543_ (.A1(_10960_),
    .A2(_11149_),
    .B(_11151_),
    .Y(_11152_));
 OA21x2_ASAP7_75t_R _27544_ (.A1(_05605_),
    .A2(_11034_),
    .B(_11044_),
    .Y(_11153_));
 OR3x1_ASAP7_75t_R _27545_ (.A(_11049_),
    .B(_08565_),
    .C(_11047_),
    .Y(_11154_));
 OAI21x1_ASAP7_75t_R _27546_ (.A1(_00144_),
    .A2(_11075_),
    .B(_11154_),
    .Y(_11155_));
 AO21x1_ASAP7_75t_R _27547_ (.A1(_11152_),
    .A2(_11153_),
    .B(_11155_),
    .Y(_03873_));
 NOR2x1_ASAP7_75t_R _27548_ (.A(_00152_),
    .B(_11075_),
    .Y(_11156_));
 AND3x1_ASAP7_75t_R _27549_ (.A(_05242_),
    .B(_08649_),
    .C(_11050_),
    .Y(_11157_));
 BUFx6f_ASAP7_75t_R _27550_ (.A(_11033_),
    .Y(_11158_));
 BUFx6f_ASAP7_75t_R _27551_ (.A(_08223_),
    .Y(_11159_));
 NOR2x1_ASAP7_75t_R _27552_ (.A(\alu_adder_result_ex[10] ),
    .B(_10963_),
    .Y(_11160_));
 AO21x1_ASAP7_75t_R _27553_ (.A1(_00152_),
    .A2(_11159_),
    .B(_11160_),
    .Y(_11161_));
 OA211x2_ASAP7_75t_R _27554_ (.A1(_08218_),
    .A2(_08220_),
    .B(_00040_),
    .C(_10966_),
    .Y(_11162_));
 AO21x1_ASAP7_75t_R _27555_ (.A1(_10962_),
    .A2(_11161_),
    .B(_11162_),
    .Y(_11163_));
 OA21x2_ASAP7_75t_R _27556_ (.A1(_14636_),
    .A2(_15248_),
    .B(_10970_),
    .Y(_11164_));
 OA21x2_ASAP7_75t_R _27557_ (.A1(_05197_),
    .A2(_11147_),
    .B(_11164_),
    .Y(_11165_));
 OAI21x1_ASAP7_75t_R _27558_ (.A1(_10959_),
    .A2(_11163_),
    .B(_11165_),
    .Y(_11166_));
 OA211x2_ASAP7_75t_R _27559_ (.A1(_05324_),
    .A2(_11158_),
    .B(_11043_),
    .C(_11166_),
    .Y(_11167_));
 OR3x1_ASAP7_75t_R _27560_ (.A(_11156_),
    .B(_11157_),
    .C(_11167_),
    .Y(_03874_));
 NOR2x1_ASAP7_75t_R _27561_ (.A(\alu_adder_result_ex[11] ),
    .B(_11111_),
    .Y(_11168_));
 AO21x1_ASAP7_75t_R _27562_ (.A1(_00160_),
    .A2(_11064_),
    .B(_11168_),
    .Y(_11169_));
 OA211x2_ASAP7_75t_R _27563_ (.A1(_08220_),
    .A2(_08225_),
    .B(_00041_),
    .C(_10967_),
    .Y(_11170_));
 AO21x1_ASAP7_75t_R _27564_ (.A1(_11062_),
    .A2(_11169_),
    .B(_11170_),
    .Y(_11171_));
 OA21x2_ASAP7_75t_R _27565_ (.A1(_05252_),
    .A2(_15240_),
    .B(_10972_),
    .Y(_11172_));
 OA21x2_ASAP7_75t_R _27566_ (.A1(_08219_),
    .A2(_11161_),
    .B(_11172_),
    .Y(_11173_));
 OAI21x1_ASAP7_75t_R _27567_ (.A1(_10960_),
    .A2(_11171_),
    .B(_11173_),
    .Y(_11174_));
 OA21x2_ASAP7_75t_R _27568_ (.A1(_05328_),
    .A2(_11034_),
    .B(_11044_),
    .Y(_11175_));
 OR3x1_ASAP7_75t_R _27569_ (.A(_11049_),
    .B(_08701_),
    .C(_11046_),
    .Y(_11176_));
 OAI21x1_ASAP7_75t_R _27570_ (.A1(_00160_),
    .A2(_11075_),
    .B(_11176_),
    .Y(_11177_));
 AO21x1_ASAP7_75t_R _27571_ (.A1(_11174_),
    .A2(_11175_),
    .B(_11177_),
    .Y(_03875_));
 NOR2x1_ASAP7_75t_R _27572_ (.A(\alu_adder_result_ex[12] ),
    .B(_11122_),
    .Y(_11178_));
 AO21x1_ASAP7_75t_R _27573_ (.A1(_00168_),
    .A2(_11111_),
    .B(_11178_),
    .Y(_11179_));
 OA211x2_ASAP7_75t_R _27574_ (.A1(_08210_),
    .A2(_08227_),
    .B(_00042_),
    .C(_10967_),
    .Y(_11180_));
 AO21x1_ASAP7_75t_R _27575_ (.A1(_11062_),
    .A2(_11179_),
    .B(_11180_),
    .Y(_11181_));
 OA21x2_ASAP7_75t_R _27576_ (.A1(_05252_),
    .A2(_15524_),
    .B(_10972_),
    .Y(_11182_));
 OA21x2_ASAP7_75t_R _27577_ (.A1(_08219_),
    .A2(_11169_),
    .B(_11182_),
    .Y(_11183_));
 OA21x2_ASAP7_75t_R _27578_ (.A1(_10960_),
    .A2(_11181_),
    .B(_11183_),
    .Y(_11184_));
 INVx1_ASAP7_75t_R _27579_ (.A(_11043_),
    .Y(_11185_));
 AO21x1_ASAP7_75t_R _27580_ (.A1(_05618_),
    .A2(_11053_),
    .B(_11185_),
    .Y(_11186_));
 OA21x2_ASAP7_75t_R _27581_ (.A1(_11049_),
    .A2(_08742_),
    .B(_11050_),
    .Y(_11187_));
 AO21x1_ASAP7_75t_R _27582_ (.A1(_00168_),
    .A2(_11047_),
    .B(_11187_),
    .Y(_11188_));
 OAI21x1_ASAP7_75t_R _27583_ (.A1(_11184_),
    .A2(_11186_),
    .B(_11188_),
    .Y(_03876_));
 NOR2x1_ASAP7_75t_R _27584_ (.A(\alu_adder_result_ex[13] ),
    .B(_11063_),
    .Y(_11189_));
 AO21x1_ASAP7_75t_R _27585_ (.A1(_00175_),
    .A2(_11122_),
    .B(_11189_),
    .Y(_11190_));
 OA211x2_ASAP7_75t_R _27586_ (.A1(_08227_),
    .A2(_08230_),
    .B(_00043_),
    .C(_10966_),
    .Y(_11191_));
 AO21x1_ASAP7_75t_R _27587_ (.A1(_10962_),
    .A2(_11190_),
    .B(_11191_),
    .Y(_11192_));
 OR2x2_ASAP7_75t_R _27588_ (.A(_10959_),
    .B(_11192_),
    .Y(_11193_));
 OA21x2_ASAP7_75t_R _27589_ (.A1(_05566_),
    .A2(_15518_),
    .B(_10971_),
    .Y(_11194_));
 OA21x2_ASAP7_75t_R _27590_ (.A1(_05197_),
    .A2(_11179_),
    .B(_11194_),
    .Y(_11195_));
 NOR2x1_ASAP7_75t_R _27591_ (.A(_05624_),
    .B(_11033_),
    .Y(_11196_));
 OA21x2_ASAP7_75t_R _27592_ (.A1(_11195_),
    .A2(_11196_),
    .B(_05722_),
    .Y(_11197_));
 AOI21x1_ASAP7_75t_R _27593_ (.A1(_11193_),
    .A2(_11197_),
    .B(_08783_),
    .Y(_11198_));
 NAND2x1_ASAP7_75t_R _27594_ (.A(_00175_),
    .B(_11144_),
    .Y(_11199_));
 OA21x2_ASAP7_75t_R _27595_ (.A1(_11133_),
    .A2(_11198_),
    .B(_11199_),
    .Y(_03877_));
 OA211x2_ASAP7_75t_R _27596_ (.A1(_08218_),
    .A2(_08227_),
    .B(_00044_),
    .C(_10967_),
    .Y(_11200_));
 NAND2x1_ASAP7_75t_R _27597_ (.A(_00180_),
    .B(_11122_),
    .Y(_11201_));
 OA21x2_ASAP7_75t_R _27598_ (.A1(\alu_adder_result_ex[14] ),
    .A2(_11111_),
    .B(_11201_),
    .Y(_11202_));
 NOR2x1_ASAP7_75t_R _27599_ (.A(_11068_),
    .B(_11202_),
    .Y(_11203_));
 OR3x1_ASAP7_75t_R _27600_ (.A(_10959_),
    .B(_11200_),
    .C(_11203_),
    .Y(_11204_));
 OA211x2_ASAP7_75t_R _27601_ (.A1(_05635_),
    .A2(_15772_),
    .B(_08813_),
    .C(_10971_),
    .Y(_11205_));
 OA21x2_ASAP7_75t_R _27602_ (.A1(_08219_),
    .A2(_11190_),
    .B(_11205_),
    .Y(_11206_));
 AO21x1_ASAP7_75t_R _27603_ (.A1(_15583_),
    .A2(_11053_),
    .B(_14534_),
    .Y(_11207_));
 AOI221x1_ASAP7_75t_R _27604_ (.A1(_11204_),
    .A2(_11206_),
    .B1(_11207_),
    .B2(_08813_),
    .C(_08568_),
    .Y(_11208_));
 NAND2x1_ASAP7_75t_R _27605_ (.A(_00180_),
    .B(_11144_),
    .Y(_11209_));
 OA21x2_ASAP7_75t_R _27606_ (.A1(_11133_),
    .A2(_11208_),
    .B(_11209_),
    .Y(_03878_));
 NOR2x1_ASAP7_75t_R _27607_ (.A(\alu_adder_result_ex[15] ),
    .B(_11159_),
    .Y(_11210_));
 AO21x1_ASAP7_75t_R _27608_ (.A1(_00187_),
    .A2(_11111_),
    .B(_11210_),
    .Y(_11211_));
 OA211x2_ASAP7_75t_R _27609_ (.A1(_08225_),
    .A2(_08227_),
    .B(_00045_),
    .C(_10967_),
    .Y(_11212_));
 AOI21x1_ASAP7_75t_R _27610_ (.A1(_11062_),
    .A2(_11211_),
    .B(_11212_),
    .Y(_11213_));
 BUFx6f_ASAP7_75t_R _27611_ (.A(_11035_),
    .Y(_11214_));
 AO221x1_ASAP7_75t_R _27612_ (.A1(_05559_),
    .A2(\alu_adder_result_ex[15] ),
    .B1(_11202_),
    .B2(_05249_),
    .C(_11214_),
    .Y(_11215_));
 AO21x1_ASAP7_75t_R _27613_ (.A1(_05247_),
    .A2(_11213_),
    .B(_11215_),
    .Y(_11216_));
 OA21x2_ASAP7_75t_R _27614_ (.A1(_15707_),
    .A2(_11034_),
    .B(_11044_),
    .Y(_11217_));
 OR3x1_ASAP7_75t_R _27615_ (.A(_11049_),
    .B(_08886_),
    .C(_11046_),
    .Y(_11218_));
 OAI21x1_ASAP7_75t_R _27616_ (.A1(_00187_),
    .A2(_11075_),
    .B(_11218_),
    .Y(_11219_));
 AO21x1_ASAP7_75t_R _27617_ (.A1(_11216_),
    .A2(_11217_),
    .B(_11219_),
    .Y(_03879_));
 NOR2x1_ASAP7_75t_R _27618_ (.A(_05578_),
    .B(_10873_),
    .Y(_11220_));
 AO21x1_ASAP7_75t_R _27619_ (.A1(\alu_adder_result_ex[4] ),
    .A2(_10873_),
    .B(_11220_),
    .Y(_11221_));
 NAND2x1_ASAP7_75t_R _27620_ (.A(_01730_),
    .B(_10905_),
    .Y(_11222_));
 OA21x2_ASAP7_75t_R _27621_ (.A1(_10939_),
    .A2(_11221_),
    .B(_11222_),
    .Y(_03880_));
 NOR2x1_ASAP7_75t_R _27622_ (.A(\alu_adder_result_ex[16] ),
    .B(_11122_),
    .Y(_11223_));
 AO21x1_ASAP7_75t_R _27623_ (.A1(_15836_),
    .A2(_11111_),
    .B(_11223_),
    .Y(_11224_));
 OA211x2_ASAP7_75t_R _27624_ (.A1(_08078_),
    .A2(_08232_),
    .B(_11067_),
    .C(_00046_),
    .Y(_11225_));
 AO21x1_ASAP7_75t_R _27625_ (.A1(_10962_),
    .A2(_11224_),
    .B(_11225_),
    .Y(_11226_));
 OA211x2_ASAP7_75t_R _27626_ (.A1(_14636_),
    .A2(_16019_),
    .B(_05721_),
    .C(_10971_),
    .Y(_11227_));
 OA21x2_ASAP7_75t_R _27627_ (.A1(_05197_),
    .A2(_11211_),
    .B(_11227_),
    .Y(_11228_));
 OAI21x1_ASAP7_75t_R _27628_ (.A1(_10959_),
    .A2(_11226_),
    .B(_11228_),
    .Y(_11229_));
 OR3x1_ASAP7_75t_R _27629_ (.A(_15831_),
    .B(_09037_),
    .C(_11033_),
    .Y(_11230_));
 AND3x1_ASAP7_75t_R _27630_ (.A(_08909_),
    .B(_11229_),
    .C(_11230_),
    .Y(_11231_));
 NAND2x1_ASAP7_75t_R _27631_ (.A(_15836_),
    .B(_11144_),
    .Y(_11232_));
 OA21x2_ASAP7_75t_R _27632_ (.A1(_11133_),
    .A2(_11231_),
    .B(_11232_),
    .Y(_03881_));
 NOR2x1_ASAP7_75t_R _27633_ (.A(\alu_adder_result_ex[17] ),
    .B(_11063_),
    .Y(_11233_));
 AO21x1_ASAP7_75t_R _27634_ (.A1(_15947_),
    .A2(_11122_),
    .B(_11233_),
    .Y(_11234_));
 OA211x2_ASAP7_75t_R _27635_ (.A1(_08078_),
    .A2(_08235_),
    .B(_11067_),
    .C(_00047_),
    .Y(_11235_));
 AO21x1_ASAP7_75t_R _27636_ (.A1(_10962_),
    .A2(_11234_),
    .B(_11235_),
    .Y(_11236_));
 OR2x2_ASAP7_75t_R _27637_ (.A(_10959_),
    .B(_11236_),
    .Y(_11237_));
 OA21x2_ASAP7_75t_R _27638_ (.A1(_05566_),
    .A2(_16004_),
    .B(_10971_),
    .Y(_11238_));
 OA21x2_ASAP7_75t_R _27639_ (.A1(_05197_),
    .A2(_11224_),
    .B(_11238_),
    .Y(_11239_));
 NOR2x1_ASAP7_75t_R _27640_ (.A(_05281_),
    .B(_11033_),
    .Y(_11240_));
 OA21x2_ASAP7_75t_R _27641_ (.A1(_11239_),
    .A2(_11240_),
    .B(_05722_),
    .Y(_11241_));
 AOI21x1_ASAP7_75t_R _27642_ (.A1(_11237_),
    .A2(_11241_),
    .B(_08942_),
    .Y(_11242_));
 NAND2x1_ASAP7_75t_R _27643_ (.A(_15947_),
    .B(_11144_),
    .Y(_11243_));
 OA21x2_ASAP7_75t_R _27644_ (.A1(_11133_),
    .A2(_11242_),
    .B(_11243_),
    .Y(_03882_));
 NOR2x1_ASAP7_75t_R _27645_ (.A(\alu_adder_result_ex[18] ),
    .B(_11159_),
    .Y(_11244_));
 AO21x1_ASAP7_75t_R _27646_ (.A1(_16083_),
    .A2(_11111_),
    .B(_11244_),
    .Y(_11245_));
 OA211x2_ASAP7_75t_R _27647_ (.A1(_08078_),
    .A2(_08238_),
    .B(_10967_),
    .C(_00048_),
    .Y(_11246_));
 AOI211x1_ASAP7_75t_R _27648_ (.A1(_08063_),
    .A2(_11245_),
    .B(_11246_),
    .C(_10959_),
    .Y(_11247_));
 OA211x2_ASAP7_75t_R _27649_ (.A1(_05635_),
    .A2(_16267_),
    .B(_05194_),
    .C(_10971_),
    .Y(_11248_));
 OAI21x1_ASAP7_75t_R _27650_ (.A1(_05198_),
    .A2(_11234_),
    .B(_11248_),
    .Y(_11249_));
 NOR3x1_ASAP7_75t_R _27651_ (.A(_16078_),
    .B(_09037_),
    .C(_11033_),
    .Y(_11250_));
 NOR2x1_ASAP7_75t_R _27652_ (.A(_09012_),
    .B(_11250_),
    .Y(_11251_));
 OA21x2_ASAP7_75t_R _27653_ (.A1(_11247_),
    .A2(_11249_),
    .B(_11251_),
    .Y(_11252_));
 NAND2x1_ASAP7_75t_R _27654_ (.A(_16083_),
    .B(_11144_),
    .Y(_11253_));
 OA21x2_ASAP7_75t_R _27655_ (.A1(_11133_),
    .A2(_11252_),
    .B(_11253_),
    .Y(_03883_));
 NOR2x1_ASAP7_75t_R _27656_ (.A(\alu_adder_result_ex[19] ),
    .B(_11159_),
    .Y(_11254_));
 AO21x1_ASAP7_75t_R _27657_ (.A1(_16195_),
    .A2(_11111_),
    .B(_11254_),
    .Y(_11255_));
 OA211x2_ASAP7_75t_R _27658_ (.A1(_08078_),
    .A2(_08241_),
    .B(_11067_),
    .C(_00049_),
    .Y(_11256_));
 AOI21x1_ASAP7_75t_R _27659_ (.A1(_10962_),
    .A2(_11255_),
    .B(_11256_),
    .Y(_11257_));
 OA21x2_ASAP7_75t_R _27660_ (.A1(_05566_),
    .A2(_16253_),
    .B(_10971_),
    .Y(_11258_));
 OAI21x1_ASAP7_75t_R _27661_ (.A1(_08219_),
    .A2(_11245_),
    .B(_11258_),
    .Y(_11259_));
 AO21x1_ASAP7_75t_R _27662_ (.A1(_05247_),
    .A2(_11257_),
    .B(_11259_),
    .Y(_11260_));
 AO21x1_ASAP7_75t_R _27663_ (.A1(_16159_),
    .A2(_16190_),
    .B(_11033_),
    .Y(_11261_));
 AO32x1_ASAP7_75t_R _27664_ (.A1(_05194_),
    .A2(_11260_),
    .A3(_11261_),
    .B1(_05242_),
    .B2(_09044_),
    .Y(_11262_));
 NAND2x1_ASAP7_75t_R _27665_ (.A(_16195_),
    .B(_11144_),
    .Y(_11263_));
 OA21x2_ASAP7_75t_R _27666_ (.A1(_11133_),
    .A2(_11262_),
    .B(_11263_),
    .Y(_03884_));
 OA211x2_ASAP7_75t_R _27667_ (.A1(_08232_),
    .A2(_08246_),
    .B(_00050_),
    .C(_08061_),
    .Y(_11264_));
 INVx1_ASAP7_75t_R _27668_ (.A(_11264_),
    .Y(_11265_));
 NAND2x1_ASAP7_75t_R _27669_ (.A(_16329_),
    .B(_11159_),
    .Y(_11266_));
 OA21x2_ASAP7_75t_R _27670_ (.A1(\alu_adder_result_ex[20] ),
    .A2(_11122_),
    .B(_11266_),
    .Y(_11267_));
 OA21x2_ASAP7_75t_R _27671_ (.A1(_08062_),
    .A2(_11267_),
    .B(_05247_),
    .Y(_11268_));
 OA21x2_ASAP7_75t_R _27672_ (.A1(_05566_),
    .A2(_16528_),
    .B(_10971_),
    .Y(_11269_));
 OAI21x1_ASAP7_75t_R _27673_ (.A1(_08219_),
    .A2(_11255_),
    .B(_11269_),
    .Y(_11270_));
 AO21x1_ASAP7_75t_R _27674_ (.A1(_11265_),
    .A2(_11268_),
    .B(_11270_),
    .Y(_11271_));
 OA21x2_ASAP7_75t_R _27675_ (.A1(_05654_),
    .A2(_11158_),
    .B(_05722_),
    .Y(_11272_));
 AO21x1_ASAP7_75t_R _27676_ (.A1(_11271_),
    .A2(_11272_),
    .B(_09065_),
    .Y(_11273_));
 NAND2x1_ASAP7_75t_R _27677_ (.A(_16329_),
    .B(_11144_),
    .Y(_11274_));
 OA21x2_ASAP7_75t_R _27678_ (.A1(_11133_),
    .A2(_11273_),
    .B(_11274_),
    .Y(_03885_));
 OA211x2_ASAP7_75t_R _27679_ (.A1(_08235_),
    .A2(_08246_),
    .B(_00051_),
    .C(_11067_),
    .Y(_11275_));
 INVx1_ASAP7_75t_R _27680_ (.A(_11275_),
    .Y(_11276_));
 NAND2x1_ASAP7_75t_R _27681_ (.A(_00115_),
    .B(_10963_),
    .Y(_11277_));
 OA21x2_ASAP7_75t_R _27682_ (.A1(\alu_adder_result_ex[21] ),
    .A2(_11063_),
    .B(_11277_),
    .Y(_11278_));
 OA21x2_ASAP7_75t_R _27683_ (.A1(_08062_),
    .A2(_11278_),
    .B(_05246_),
    .Y(_11279_));
 AO21x1_ASAP7_75t_R _27684_ (.A1(_05559_),
    .A2(\alu_adder_result_ex[21] ),
    .B(_11214_),
    .Y(_11280_));
 AO221x1_ASAP7_75t_R _27685_ (.A1(_05249_),
    .A2(_11267_),
    .B1(_11276_),
    .B2(_11279_),
    .C(_11280_),
    .Y(_11281_));
 OA21x2_ASAP7_75t_R _27686_ (.A1(_05295_),
    .A2(_11158_),
    .B(_05722_),
    .Y(_11282_));
 AO21x1_ASAP7_75t_R _27687_ (.A1(_11281_),
    .A2(_11282_),
    .B(_09097_),
    .Y(_11283_));
 NAND2x1_ASAP7_75t_R _27688_ (.A(_00115_),
    .B(_11144_),
    .Y(_11284_));
 OA21x2_ASAP7_75t_R _27689_ (.A1(_11133_),
    .A2(_11283_),
    .B(_11284_),
    .Y(_03886_));
 BUFx6f_ASAP7_75t_R _27690_ (.A(_11042_),
    .Y(_11285_));
 OA211x2_ASAP7_75t_R _27691_ (.A1(_08238_),
    .A2(_08246_),
    .B(_00052_),
    .C(_08061_),
    .Y(_11286_));
 INVx1_ASAP7_75t_R _27692_ (.A(_11286_),
    .Y(_11287_));
 NAND2x1_ASAP7_75t_R _27693_ (.A(_16591_),
    .B(_11063_),
    .Y(_11288_));
 OA21x2_ASAP7_75t_R _27694_ (.A1(\alu_adder_result_ex[22] ),
    .A2(_11122_),
    .B(_11288_),
    .Y(_11289_));
 OA21x2_ASAP7_75t_R _27695_ (.A1(_08062_),
    .A2(_11289_),
    .B(_05247_),
    .Y(_11290_));
 AO221x1_ASAP7_75t_R _27696_ (.A1(_05559_),
    .A2(\alu_adder_result_ex[22] ),
    .B1(_11278_),
    .B2(_05249_),
    .C(_11214_),
    .Y(_11291_));
 AO21x1_ASAP7_75t_R _27697_ (.A1(_11287_),
    .A2(_11290_),
    .B(_11291_),
    .Y(_11292_));
 OA21x2_ASAP7_75t_R _27698_ (.A1(_16587_),
    .A2(_11158_),
    .B(_05722_),
    .Y(_11293_));
 AO21x1_ASAP7_75t_R _27699_ (.A1(_11292_),
    .A2(_11293_),
    .B(_09114_),
    .Y(_11294_));
 NAND2x1_ASAP7_75t_R _27700_ (.A(_16591_),
    .B(_11144_),
    .Y(_11295_));
 OA21x2_ASAP7_75t_R _27701_ (.A1(_11285_),
    .A2(_11294_),
    .B(_11295_),
    .Y(_03887_));
 OA211x2_ASAP7_75t_R _27702_ (.A1(_08241_),
    .A2(_08246_),
    .B(_00053_),
    .C(_11067_),
    .Y(_11296_));
 INVx1_ASAP7_75t_R _27703_ (.A(_11296_),
    .Y(_11297_));
 NAND2x1_ASAP7_75t_R _27704_ (.A(_16701_),
    .B(_10963_),
    .Y(_11298_));
 OA21x2_ASAP7_75t_R _27705_ (.A1(\alu_adder_result_ex[23] ),
    .A2(_11159_),
    .B(_11298_),
    .Y(_11299_));
 OA21x2_ASAP7_75t_R _27706_ (.A1(_08062_),
    .A2(_11299_),
    .B(_05246_),
    .Y(_11300_));
 AO21x1_ASAP7_75t_R _27707_ (.A1(_05559_),
    .A2(\alu_adder_result_ex[23] ),
    .B(_11214_),
    .Y(_11301_));
 AO221x1_ASAP7_75t_R _27708_ (.A1(_05249_),
    .A2(_11289_),
    .B1(_11297_),
    .B2(_11300_),
    .C(_11301_),
    .Y(_11302_));
 OA21x2_ASAP7_75t_R _27709_ (.A1(_05308_),
    .A2(_11158_),
    .B(_05722_),
    .Y(_11303_));
 AOI211x1_ASAP7_75t_R _27710_ (.A1(_11302_),
    .A2(_11303_),
    .B(_09135_),
    .C(_11285_),
    .Y(_11304_));
 AOI21x1_ASAP7_75t_R _27711_ (.A1(_16701_),
    .A2(_11133_),
    .B(_11304_),
    .Y(_03888_));
 OA211x2_ASAP7_75t_R _27712_ (.A1(_08220_),
    .A2(_08232_),
    .B(_00054_),
    .C(_10967_),
    .Y(_11305_));
 INVx1_ASAP7_75t_R _27713_ (.A(_11305_),
    .Y(_11306_));
 NAND2x1_ASAP7_75t_R _27714_ (.A(_16823_),
    .B(_11063_),
    .Y(_11307_));
 OA21x2_ASAP7_75t_R _27715_ (.A1(\alu_adder_result_ex[24] ),
    .A2(_11122_),
    .B(_11307_),
    .Y(_11308_));
 OA21x2_ASAP7_75t_R _27716_ (.A1(_08062_),
    .A2(_11308_),
    .B(_05247_),
    .Y(_11309_));
 AO221x1_ASAP7_75t_R _27717_ (.A1(_05559_),
    .A2(\alu_adder_result_ex[24] ),
    .B1(_11299_),
    .B2(_05249_),
    .C(_11214_),
    .Y(_11310_));
 AO21x1_ASAP7_75t_R _27718_ (.A1(_11306_),
    .A2(_11309_),
    .B(_11310_),
    .Y(_11311_));
 OA21x2_ASAP7_75t_R _27719_ (.A1(_05672_),
    .A2(_11158_),
    .B(_05721_),
    .Y(_11312_));
 AO21x1_ASAP7_75t_R _27720_ (.A1(_11311_),
    .A2(_11312_),
    .B(_09155_),
    .Y(_11313_));
 BUFx6f_ASAP7_75t_R _27721_ (.A(_11042_),
    .Y(_11314_));
 NAND2x1_ASAP7_75t_R _27722_ (.A(_16823_),
    .B(_11314_),
    .Y(_11315_));
 OA21x2_ASAP7_75t_R _27723_ (.A1(_11285_),
    .A2(_11313_),
    .B(_11315_),
    .Y(_03889_));
 OA211x2_ASAP7_75t_R _27724_ (.A1(_08220_),
    .A2(_08235_),
    .B(_00055_),
    .C(_11067_),
    .Y(_11316_));
 INVx1_ASAP7_75t_R _27725_ (.A(_11316_),
    .Y(_11317_));
 NAND2x1_ASAP7_75t_R _27726_ (.A(_16935_),
    .B(_10963_),
    .Y(_11318_));
 OA21x2_ASAP7_75t_R _27727_ (.A1(\alu_adder_result_ex[25] ),
    .A2(_11063_),
    .B(_11318_),
    .Y(_11319_));
 OA21x2_ASAP7_75t_R _27728_ (.A1(_08061_),
    .A2(_11319_),
    .B(_05246_),
    .Y(_11320_));
 AO21x1_ASAP7_75t_R _27729_ (.A1(_05559_),
    .A2(\alu_adder_result_ex[25] ),
    .B(_11214_),
    .Y(_11321_));
 AO221x1_ASAP7_75t_R _27730_ (.A1(_05249_),
    .A2(_11308_),
    .B1(_11317_),
    .B2(_11320_),
    .C(_11321_),
    .Y(_11322_));
 OA21x2_ASAP7_75t_R _27731_ (.A1(_16931_),
    .A2(_11158_),
    .B(_05721_),
    .Y(_11323_));
 AO21x1_ASAP7_75t_R _27732_ (.A1(_11322_),
    .A2(_11323_),
    .B(_09185_),
    .Y(_11324_));
 NAND2x1_ASAP7_75t_R _27733_ (.A(_16935_),
    .B(_11314_),
    .Y(_11325_));
 OA21x2_ASAP7_75t_R _27734_ (.A1(_11285_),
    .A2(_11324_),
    .B(_11325_),
    .Y(_03890_));
 AND2x2_ASAP7_75t_R _27735_ (.A(_13830_),
    .B(_10878_),
    .Y(_11326_));
 AO21x1_ASAP7_75t_R _27736_ (.A1(\alu_adder_result_ex[5] ),
    .A2(_10891_),
    .B(_11326_),
    .Y(_11327_));
 AO21x1_ASAP7_75t_R _27737_ (.A1(_05200_),
    .A2(_10922_),
    .B(_05584_),
    .Y(_11328_));
 OA21x2_ASAP7_75t_R _27738_ (.A1(_10939_),
    .A2(_11327_),
    .B(_11328_),
    .Y(_03891_));
 OA211x2_ASAP7_75t_R _27739_ (.A1(_08220_),
    .A2(_08238_),
    .B(_00056_),
    .C(_10967_),
    .Y(_11329_));
 INVx1_ASAP7_75t_R _27740_ (.A(_11329_),
    .Y(_11330_));
 NAND2x1_ASAP7_75t_R _27741_ (.A(_04310_),
    .B(_10963_),
    .Y(_11331_));
 OA21x2_ASAP7_75t_R _27742_ (.A1(\alu_adder_result_ex[26] ),
    .A2(_11159_),
    .B(_11331_),
    .Y(_11332_));
 OA21x2_ASAP7_75t_R _27743_ (.A1(_08062_),
    .A2(_11332_),
    .B(_05247_),
    .Y(_11333_));
 AO221x1_ASAP7_75t_R _27744_ (.A1(_05622_),
    .A2(\alu_adder_result_ex[26] ),
    .B1(_11319_),
    .B2(_05249_),
    .C(_11214_),
    .Y(_11334_));
 AO21x1_ASAP7_75t_R _27745_ (.A1(_11330_),
    .A2(_11333_),
    .B(_11334_),
    .Y(_11335_));
 OA21x2_ASAP7_75t_R _27746_ (.A1(_04305_),
    .A2(_11158_),
    .B(_05721_),
    .Y(_11336_));
 AO21x1_ASAP7_75t_R _27747_ (.A1(_11335_),
    .A2(_11336_),
    .B(_09212_),
    .Y(_11337_));
 NAND2x1_ASAP7_75t_R _27748_ (.A(_04310_),
    .B(_11314_),
    .Y(_11338_));
 OA21x2_ASAP7_75t_R _27749_ (.A1(_11285_),
    .A2(_11337_),
    .B(_11338_),
    .Y(_03892_));
 OA21x2_ASAP7_75t_R _27750_ (.A1(_08220_),
    .A2(_08241_),
    .B(_00057_),
    .Y(_11339_));
 NAND2x1_ASAP7_75t_R _27751_ (.A(_11068_),
    .B(_11339_),
    .Y(_11340_));
 NAND2x1_ASAP7_75t_R _27752_ (.A(_04422_),
    .B(_10963_),
    .Y(_11341_));
 OA21x2_ASAP7_75t_R _27753_ (.A1(\alu_adder_result_ex[27] ),
    .A2(_11159_),
    .B(_11341_),
    .Y(_11342_));
 OA21x2_ASAP7_75t_R _27754_ (.A1(_08062_),
    .A2(_11342_),
    .B(_05247_),
    .Y(_11343_));
 AO221x1_ASAP7_75t_R _27755_ (.A1(_05622_),
    .A2(\alu_adder_result_ex[27] ),
    .B1(_11332_),
    .B2(_05249_),
    .C(_11214_),
    .Y(_11344_));
 AO21x1_ASAP7_75t_R _27756_ (.A1(_11340_),
    .A2(_11343_),
    .B(_11344_),
    .Y(_11345_));
 AOI21x1_ASAP7_75t_R _27757_ (.A1(_05685_),
    .A2(_11053_),
    .B(_09037_),
    .Y(_11346_));
 AO21x1_ASAP7_75t_R _27758_ (.A1(_11345_),
    .A2(_11346_),
    .B(_09240_),
    .Y(_11347_));
 NAND2x1_ASAP7_75t_R _27759_ (.A(_04422_),
    .B(_11314_),
    .Y(_11348_));
 OA21x2_ASAP7_75t_R _27760_ (.A1(_11285_),
    .A2(_11347_),
    .B(_11348_),
    .Y(_03893_));
 OA211x2_ASAP7_75t_R _27761_ (.A1(_08227_),
    .A2(_08232_),
    .B(_00058_),
    .C(_08061_),
    .Y(_11349_));
 INVx1_ASAP7_75t_R _27762_ (.A(_11349_),
    .Y(_11350_));
 NAND2x1_ASAP7_75t_R _27763_ (.A(_04558_),
    .B(_10963_),
    .Y(_11351_));
 OA21x2_ASAP7_75t_R _27764_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_11159_),
    .B(_11351_),
    .Y(_11352_));
 OA21x2_ASAP7_75t_R _27765_ (.A1(_08062_),
    .A2(_11352_),
    .B(_05246_),
    .Y(_11353_));
 AO221x1_ASAP7_75t_R _27766_ (.A1(_05622_),
    .A2(\alu_adder_result_ex[28] ),
    .B1(_11342_),
    .B2(_05248_),
    .C(_11035_),
    .Y(_11354_));
 AO21x1_ASAP7_75t_R _27767_ (.A1(_11350_),
    .A2(_11353_),
    .B(_11354_),
    .Y(_11355_));
 OA21x2_ASAP7_75t_R _27768_ (.A1(_04554_),
    .A2(_11158_),
    .B(_05721_),
    .Y(_11356_));
 AO21x1_ASAP7_75t_R _27769_ (.A1(_11355_),
    .A2(_11356_),
    .B(_09277_),
    .Y(_11357_));
 NAND2x1_ASAP7_75t_R _27770_ (.A(_04558_),
    .B(_11314_),
    .Y(_11358_));
 OA21x2_ASAP7_75t_R _27771_ (.A1(_11285_),
    .A2(_11357_),
    .B(_11358_),
    .Y(_03894_));
 OA211x2_ASAP7_75t_R _27772_ (.A1(_08227_),
    .A2(_08235_),
    .B(_00059_),
    .C(_08061_),
    .Y(_11359_));
 INVx1_ASAP7_75t_R _27773_ (.A(_11359_),
    .Y(_11360_));
 NAND2x1_ASAP7_75t_R _27774_ (.A(_04670_),
    .B(_10963_),
    .Y(_11361_));
 OA21x2_ASAP7_75t_R _27775_ (.A1(\alu_adder_result_ex[29] ),
    .A2(_11159_),
    .B(_11361_),
    .Y(_11362_));
 OA21x2_ASAP7_75t_R _27776_ (.A1(_08062_),
    .A2(_11362_),
    .B(_05246_),
    .Y(_11363_));
 AO221x1_ASAP7_75t_R _27777_ (.A1(_05622_),
    .A2(\alu_adder_result_ex[29] ),
    .B1(_11352_),
    .B2(_05248_),
    .C(_11035_),
    .Y(_11364_));
 AO21x1_ASAP7_75t_R _27778_ (.A1(_11360_),
    .A2(_11363_),
    .B(_11364_),
    .Y(_11365_));
 OA21x2_ASAP7_75t_R _27779_ (.A1(_05343_),
    .A2(_11158_),
    .B(_05721_),
    .Y(_11366_));
 AO21x1_ASAP7_75t_R _27780_ (.A1(_11365_),
    .A2(_11366_),
    .B(_09315_),
    .Y(_11367_));
 NAND2x1_ASAP7_75t_R _27781_ (.A(_04670_),
    .B(_11314_),
    .Y(_11368_));
 OA21x2_ASAP7_75t_R _27782_ (.A1(_11285_),
    .A2(_11367_),
    .B(_11368_),
    .Y(_03895_));
 NOR2x1_ASAP7_75t_R _27783_ (.A(\alu_adder_result_ex[30] ),
    .B(_11122_),
    .Y(_11369_));
 AO21x1_ASAP7_75t_R _27784_ (.A1(_04791_),
    .A2(_11111_),
    .B(_11369_),
    .Y(_11370_));
 OA211x2_ASAP7_75t_R _27785_ (.A1(_08227_),
    .A2(_08238_),
    .B(_00060_),
    .C(_11067_),
    .Y(_11371_));
 AOI21x1_ASAP7_75t_R _27786_ (.A1(_10962_),
    .A2(_11370_),
    .B(_11371_),
    .Y(_11372_));
 AO221x1_ASAP7_75t_R _27787_ (.A1(_05622_),
    .A2(\alu_adder_result_ex[30] ),
    .B1(_11362_),
    .B2(_05248_),
    .C(_11035_),
    .Y(_11373_));
 AO21x1_ASAP7_75t_R _27788_ (.A1(_05247_),
    .A2(_11372_),
    .B(_11373_),
    .Y(_11374_));
 OA21x2_ASAP7_75t_R _27789_ (.A1(_05358_),
    .A2(_11033_),
    .B(_05721_),
    .Y(_11375_));
 AO21x1_ASAP7_75t_R _27790_ (.A1(_11374_),
    .A2(_11375_),
    .B(_09342_),
    .Y(_11376_));
 NAND2x1_ASAP7_75t_R _27791_ (.A(_04791_),
    .B(_11314_),
    .Y(_11377_));
 OA21x2_ASAP7_75t_R _27792_ (.A1(_11285_),
    .A2(_11376_),
    .B(_11377_),
    .Y(_03896_));
 NAND2x1_ASAP7_75t_R _27793_ (.A(_04960_),
    .B(net1961),
    .Y(_11378_));
 OA211x2_ASAP7_75t_R _27794_ (.A1(_08227_),
    .A2(_08241_),
    .B(_00061_),
    .C(_11067_),
    .Y(_11379_));
 AO21x1_ASAP7_75t_R _27795_ (.A1(_10962_),
    .A2(_11378_),
    .B(_11379_),
    .Y(_11380_));
 OA21x2_ASAP7_75t_R _27796_ (.A1(_05566_),
    .A2(_04971_),
    .B(_10971_),
    .Y(_11381_));
 OA21x2_ASAP7_75t_R _27797_ (.A1(_08219_),
    .A2(_11370_),
    .B(_11381_),
    .Y(_11382_));
 OAI21x1_ASAP7_75t_R _27798_ (.A1(_10959_),
    .A2(_11380_),
    .B(_11382_),
    .Y(_11383_));
 OA21x2_ASAP7_75t_R _27799_ (.A1(_04962_),
    .A2(_11033_),
    .B(_05721_),
    .Y(_11384_));
 OA211x2_ASAP7_75t_R _27800_ (.A1(_09060_),
    .A2(_09387_),
    .B(_09388_),
    .C(_09037_),
    .Y(_11385_));
 AO21x1_ASAP7_75t_R _27801_ (.A1(_11383_),
    .A2(_11384_),
    .B(_11385_),
    .Y(_11386_));
 NAND2x1_ASAP7_75t_R _27802_ (.A(_04959_),
    .B(_11314_),
    .Y(_11387_));
 OA21x2_ASAP7_75t_R _27803_ (.A1(_11285_),
    .A2(_11386_),
    .B(_11387_),
    .Y(_03897_));
 OA21x2_ASAP7_75t_R _27804_ (.A1(_00243_),
    .A2(_09339_),
    .B(_00247_),
    .Y(_11388_));
 OA21x2_ASAP7_75t_R _27805_ (.A1(_00246_),
    .A2(_11388_),
    .B(_00253_),
    .Y(_11389_));
 XOR2x2_ASAP7_75t_R _27806_ (.A(_00252_),
    .B(_11389_),
    .Y(_11390_));
 AND3x1_ASAP7_75t_R _27807_ (.A(_09037_),
    .B(_08902_),
    .C(_11390_),
    .Y(_11391_));
 AO32x1_ASAP7_75t_R _27808_ (.A1(_04960_),
    .A2(_05249_),
    .A3(net1961),
    .B1(_11068_),
    .B2(_11214_),
    .Y(_11392_));
 AO21x1_ASAP7_75t_R _27809_ (.A1(_05722_),
    .A2(_11392_),
    .B(_11042_),
    .Y(_11393_));
 NAND2x1_ASAP7_75t_R _27810_ (.A(_01728_),
    .B(_11314_),
    .Y(_11394_));
 OA21x2_ASAP7_75t_R _27811_ (.A1(_11391_),
    .A2(_11393_),
    .B(_11394_),
    .Y(_03898_));
 AO21x1_ASAP7_75t_R _27812_ (.A1(_11068_),
    .A2(_11214_),
    .B(_11042_),
    .Y(_11395_));
 NAND2x1_ASAP7_75t_R _27813_ (.A(_00205_),
    .B(_11314_),
    .Y(_11396_));
 OA21x2_ASAP7_75t_R _27814_ (.A1(_00246_),
    .A2(_09386_),
    .B(_00253_),
    .Y(_11397_));
 OA21x2_ASAP7_75t_R _27815_ (.A1(_00252_),
    .A2(_11397_),
    .B(_00259_),
    .Y(_11398_));
 XOR2x2_ASAP7_75t_R _27816_ (.A(_00255_),
    .B(_17973_),
    .Y(_11399_));
 XNOR2x2_ASAP7_75t_R _27817_ (.A(net32),
    .B(_17937_),
    .Y(_11400_));
 XNOR2x2_ASAP7_75t_R _27818_ (.A(_11399_),
    .B(_11400_),
    .Y(_11401_));
 XNOR2x2_ASAP7_75t_R _27819_ (.A(_00258_),
    .B(_02290_),
    .Y(_11402_));
 XNOR2x2_ASAP7_75t_R _27820_ (.A(_00249_),
    .B(_00257_),
    .Y(_11403_));
 XNOR2x2_ASAP7_75t_R _27821_ (.A(_11402_),
    .B(_11403_),
    .Y(_11404_));
 XNOR2x2_ASAP7_75t_R _27822_ (.A(_11401_),
    .B(_11404_),
    .Y(_11405_));
 XOR2x2_ASAP7_75t_R _27823_ (.A(_02214_),
    .B(_02215_),
    .Y(_11406_));
 XNOR2x2_ASAP7_75t_R _27824_ (.A(_00254_),
    .B(net1962),
    .Y(_11407_));
 XNOR2x2_ASAP7_75t_R _27825_ (.A(_11406_),
    .B(_11407_),
    .Y(_11408_));
 XOR2x2_ASAP7_75t_R _27826_ (.A(_02218_),
    .B(_02219_),
    .Y(_11409_));
 XNOR2x2_ASAP7_75t_R _27827_ (.A(_02216_),
    .B(_11409_),
    .Y(_11410_));
 XNOR2x2_ASAP7_75t_R _27828_ (.A(_11408_),
    .B(_11410_),
    .Y(_11411_));
 XNOR2x2_ASAP7_75t_R _27829_ (.A(_11405_),
    .B(_11411_),
    .Y(_11412_));
 OA21x2_ASAP7_75t_R _27830_ (.A1(_00205_),
    .A2(_05244_),
    .B(_05376_),
    .Y(_11413_));
 XNOR2x2_ASAP7_75t_R _27831_ (.A(_11412_),
    .B(_11413_),
    .Y(_11414_));
 XNOR2x2_ASAP7_75t_R _27832_ (.A(_17365_),
    .B(_11414_),
    .Y(_11415_));
 XNOR2x2_ASAP7_75t_R _27833_ (.A(_17421_),
    .B(_11415_),
    .Y(_11416_));
 XNOR2x2_ASAP7_75t_R _27834_ (.A(_11398_),
    .B(_11416_),
    .Y(_11417_));
 AND3x1_ASAP7_75t_R _27835_ (.A(_05235_),
    .B(_11075_),
    .C(_11417_),
    .Y(_11418_));
 AO21x1_ASAP7_75t_R _27836_ (.A1(_11395_),
    .A2(_11396_),
    .B(_11418_),
    .Y(_03899_));
 NOR2x1_ASAP7_75t_R _27837_ (.A(_05033_),
    .B(_10873_),
    .Y(_11419_));
 AO21x1_ASAP7_75t_R _27838_ (.A1(\alu_adder_result_ex[6] ),
    .A2(_10891_),
    .B(_11419_),
    .Y(_11420_));
 AO21x1_ASAP7_75t_R _27839_ (.A1(_05200_),
    .A2(_10922_),
    .B(_05590_),
    .Y(_11421_));
 OA21x2_ASAP7_75t_R _27840_ (.A1(_10939_),
    .A2(_11420_),
    .B(_11421_),
    .Y(_03900_));
 AND2x2_ASAP7_75t_R _27841_ (.A(_13968_),
    .B(_10878_),
    .Y(_11422_));
 AO21x1_ASAP7_75t_R _27842_ (.A1(\alu_adder_result_ex[7] ),
    .A2(_10891_),
    .B(_11422_),
    .Y(_11423_));
 AO21x1_ASAP7_75t_R _27843_ (.A1(_05200_),
    .A2(_05196_),
    .B(_05594_),
    .Y(_11424_));
 OA21x2_ASAP7_75t_R _27844_ (.A1(_10880_),
    .A2(_11423_),
    .B(_11424_),
    .Y(_03901_));
 NOR2x1_ASAP7_75t_R _27845_ (.A(_04996_),
    .B(_10873_),
    .Y(_11425_));
 AO21x1_ASAP7_75t_R _27846_ (.A1(\alu_adder_result_ex[8] ),
    .A2(_10891_),
    .B(_11425_),
    .Y(_11426_));
 NAND2x1_ASAP7_75t_R _27847_ (.A(_01725_),
    .B(_10905_),
    .Y(_11427_));
 OA21x2_ASAP7_75t_R _27848_ (.A1(_10880_),
    .A2(_11426_),
    .B(_11427_),
    .Y(_03902_));
 OR2x2_ASAP7_75t_R _27849_ (.A(_14089_),
    .B(_10873_),
    .Y(_11428_));
 OA21x2_ASAP7_75t_R _27850_ (.A1(\alu_adder_result_ex[9] ),
    .A2(_10940_),
    .B(_11428_),
    .Y(_11429_));
 NAND2x1_ASAP7_75t_R _27851_ (.A(_02201_),
    .B(_10905_),
    .Y(_11430_));
 OA21x2_ASAP7_75t_R _27852_ (.A1(_10880_),
    .A2(_11429_),
    .B(_11430_),
    .Y(_03903_));
 NAND2x1_ASAP7_75t_R _27853_ (.A(_01723_),
    .B(_05456_),
    .Y(_11431_));
 NAND3x2_ASAP7_75t_R _27854_ (.B(_05474_),
    .C(_05475_),
    .Y(_11432_),
    .A(_05470_));
 AND2x6_ASAP7_75t_R _27855_ (.A(_05462_),
    .B(_11432_),
    .Y(_11433_));
 OA222x2_ASAP7_75t_R _27856_ (.A1(_15040_),
    .A2(_05158_),
    .B1(_05470_),
    .B2(_02029_),
    .C1(_01927_),
    .C2(_05502_),
    .Y(_11434_));
 AOI22x1_ASAP7_75t_R _27857_ (.A1(_01696_),
    .A2(_05456_),
    .B1(_11433_),
    .B2(_11434_),
    .Y(_11435_));
 INVx2_ASAP7_75t_R _27858_ (.A(_02331_),
    .Y(_11436_));
 OAI22x1_ASAP7_75t_R _27859_ (.A1(_01400_),
    .A2(_05471_),
    .B1(_05502_),
    .B2(_01930_),
    .Y(_11437_));
 AO21x1_ASAP7_75t_R _27860_ (.A1(_07268_),
    .A2(_07535_),
    .B(_11437_),
    .Y(_11438_));
 OA211x2_ASAP7_75t_R _27861_ (.A1(_15029_),
    .A2(_05221_),
    .B(_05225_),
    .C(_10827_),
    .Y(_11439_));
 OA21x2_ASAP7_75t_R _27862_ (.A1(_11438_),
    .A2(_11439_),
    .B(_11433_),
    .Y(_11440_));
 NOR2x1_ASAP7_75t_R _27863_ (.A(_01699_),
    .B(_05463_),
    .Y(_11441_));
 OA222x2_ASAP7_75t_R _27864_ (.A1(_01401_),
    .A2(_05470_),
    .B1(_05501_),
    .B2(_01929_),
    .C1(_05158_),
    .C2(_05212_),
    .Y(_11442_));
 AND3x4_ASAP7_75t_R _27865_ (.A(_05463_),
    .B(_07548_),
    .C(_11442_),
    .Y(_11443_));
 AOI21x1_ASAP7_75t_R _27866_ (.A1(_01698_),
    .A2(_05456_),
    .B(_11443_),
    .Y(_11444_));
 OA21x2_ASAP7_75t_R _27867_ (.A1(_11440_),
    .A2(_11441_),
    .B(_11444_),
    .Y(_11445_));
 OR2x2_ASAP7_75t_R _27868_ (.A(_01402_),
    .B(_05470_),
    .Y(_11446_));
 OA211x2_ASAP7_75t_R _27869_ (.A1(_01928_),
    .A2(_05502_),
    .B(_07555_),
    .C(_11446_),
    .Y(_11447_));
 INVx1_ASAP7_75t_R _27870_ (.A(_11447_),
    .Y(_11448_));
 AO21x1_ASAP7_75t_R _27871_ (.A1(\alu_adder_result_ex[6] ),
    .A2(_10827_),
    .B(_11448_),
    .Y(_11449_));
 NOR2x1_ASAP7_75t_R _27872_ (.A(_01697_),
    .B(_05463_),
    .Y(_11450_));
 AO21x2_ASAP7_75t_R _27873_ (.A1(_11433_),
    .A2(_11449_),
    .B(_11450_),
    .Y(_11451_));
 AND3x4_ASAP7_75t_R _27874_ (.A(_11436_),
    .B(_11445_),
    .C(_11451_),
    .Y(_11452_));
 NAND2x1_ASAP7_75t_R _27875_ (.A(_11435_),
    .B(_11452_),
    .Y(_11453_));
 OA21x2_ASAP7_75t_R _27876_ (.A1(_07274_),
    .A2(_05407_),
    .B(_05154_),
    .Y(_11454_));
 OR3x2_ASAP7_75t_R _27877_ (.A(_05704_),
    .B(_05156_),
    .C(_11454_),
    .Y(_11455_));
 OA222x2_ASAP7_75t_R _27878_ (.A1(_02027_),
    .A2(_05470_),
    .B1(_05501_),
    .B2(_01925_),
    .C1(_01404_),
    .C2(_11455_),
    .Y(_11456_));
 OA21x2_ASAP7_75t_R _27879_ (.A1(_08058_),
    .A2(_11432_),
    .B(_11456_),
    .Y(_11457_));
 OA211x2_ASAP7_75t_R _27880_ (.A1(_15166_),
    .A2(_05158_),
    .B(_05462_),
    .C(_11457_),
    .Y(_11458_));
 AOI21x1_ASAP7_75t_R _27881_ (.A1(_01694_),
    .A2(_05456_),
    .B(_11458_),
    .Y(_11459_));
 OA222x2_ASAP7_75t_R _27882_ (.A1(_02028_),
    .A2(_05470_),
    .B1(_05502_),
    .B2(_01926_),
    .C1(_01403_),
    .C2(_11455_),
    .Y(_11460_));
 OAI21x1_ASAP7_75t_R _27883_ (.A1(_08056_),
    .A2(_11432_),
    .B(_11460_),
    .Y(_11461_));
 AO31x2_ASAP7_75t_R _27884_ (.A1(_15177_),
    .A2(_15178_),
    .A3(_10827_),
    .B(_11461_),
    .Y(_11462_));
 NOR2x1_ASAP7_75t_R _27885_ (.A(_01695_),
    .B(_05463_),
    .Y(_11463_));
 AO21x2_ASAP7_75t_R _27886_ (.A1(_05463_),
    .A2(_11462_),
    .B(_11463_),
    .Y(_11464_));
 NAND2x1_ASAP7_75t_R _27887_ (.A(_11459_),
    .B(_11464_),
    .Y(_11465_));
 OR2x2_ASAP7_75t_R _27888_ (.A(_11453_),
    .B(_11465_),
    .Y(_11466_));
 OA222x2_ASAP7_75t_R _27889_ (.A1(_02052_),
    .A2(_05470_),
    .B1(_05501_),
    .B2(_01955_),
    .C1(_01405_),
    .C2(_11455_),
    .Y(_11467_));
 OA211x2_ASAP7_75t_R _27890_ (.A1(_08003_),
    .A2(_11432_),
    .B(_11467_),
    .C(_05463_),
    .Y(_11468_));
 OAI21x1_ASAP7_75t_R _27891_ (.A1(_15248_),
    .A2(_05158_),
    .B(_11468_),
    .Y(_11469_));
 XNOR2x2_ASAP7_75t_R _27892_ (.A(_11466_),
    .B(_11469_),
    .Y(_11470_));
 INVx1_ASAP7_75t_R _27893_ (.A(_01723_),
    .Y(_11471_));
 BUFx6f_ASAP7_75t_R _27894_ (.A(_05716_),
    .Y(_11472_));
 OR3x1_ASAP7_75t_R _27895_ (.A(_11471_),
    .B(_11472_),
    .C(_11466_),
    .Y(_11473_));
 OAI21x1_ASAP7_75t_R _27896_ (.A1(_01723_),
    .A2(_18717_),
    .B(_11473_),
    .Y(_11474_));
 BUFx6f_ASAP7_75t_R _27897_ (.A(_05459_),
    .Y(_11475_));
 AO22x1_ASAP7_75t_R _27898_ (.A1(_11431_),
    .A2(_11470_),
    .B1(_11474_),
    .B2(_11475_),
    .Y(_03904_));
 NAND2x2_ASAP7_75t_R _27899_ (.A(_05458_),
    .B(_05716_),
    .Y(_11476_));
 BUFx6f_ASAP7_75t_R _27900_ (.A(_11476_),
    .Y(_11477_));
 AOI211x1_ASAP7_75t_R _27901_ (.A1(_05189_),
    .A2(_05452_),
    .B(_05473_),
    .C(_07270_),
    .Y(_11478_));
 OA21x2_ASAP7_75t_R _27902_ (.A1(_04991_),
    .A2(_05509_),
    .B(_07272_),
    .Y(_11479_));
 AND2x2_ASAP7_75t_R _27903_ (.A(_00746_),
    .B(_11479_),
    .Y(_11480_));
 OA222x2_ASAP7_75t_R _27904_ (.A1(_02051_),
    .A2(_05470_),
    .B1(_11478_),
    .B2(_11480_),
    .C1(_05501_),
    .C2(_01954_),
    .Y(_11481_));
 OA21x2_ASAP7_75t_R _27905_ (.A1(_08011_),
    .A2(_11432_),
    .B(_11481_),
    .Y(_11482_));
 OA211x2_ASAP7_75t_R _27906_ (.A1(_15240_),
    .A2(_05158_),
    .B(_05462_),
    .C(_11482_),
    .Y(_11483_));
 AOI21x1_ASAP7_75t_R _27907_ (.A1(_01722_),
    .A2(_05456_),
    .B(_11483_),
    .Y(_11484_));
 AND4x1_ASAP7_75t_R _27908_ (.A(_18718_),
    .B(_18719_),
    .C(_11445_),
    .D(_11451_),
    .Y(_11485_));
 AND2x2_ASAP7_75t_R _27909_ (.A(_11431_),
    .B(_11469_),
    .Y(_11486_));
 AND4x1_ASAP7_75t_R _27910_ (.A(_11435_),
    .B(_11459_),
    .C(_11464_),
    .D(_11486_),
    .Y(_11487_));
 NAND2x1_ASAP7_75t_R _27911_ (.A(_11485_),
    .B(_11487_),
    .Y(_11488_));
 XNOR2x2_ASAP7_75t_R _27912_ (.A(_11484_),
    .B(_11488_),
    .Y(_11489_));
 BUFx6f_ASAP7_75t_R _27913_ (.A(_11476_),
    .Y(_11490_));
 NOR2x1_ASAP7_75t_R _27914_ (.A(_01722_),
    .B(_11490_),
    .Y(_11491_));
 AO21x1_ASAP7_75t_R _27915_ (.A1(_11477_),
    .A2(_11489_),
    .B(_11491_),
    .Y(_03905_));
 OA222x2_ASAP7_75t_R _27916_ (.A1(_02050_),
    .A2(_05471_),
    .B1(_05502_),
    .B2(_01953_),
    .C1(_00745_),
    .C2(_11455_),
    .Y(_11492_));
 OA21x2_ASAP7_75t_R _27917_ (.A1(_08013_),
    .A2(_11432_),
    .B(_11492_),
    .Y(_11493_));
 NAND2x1_ASAP7_75t_R _27918_ (.A(_05463_),
    .B(_11493_),
    .Y(_11494_));
 AO21x2_ASAP7_75t_R _27919_ (.A1(\alu_adder_result_ex[12] ),
    .A2(_10827_),
    .B(_11494_),
    .Y(_11495_));
 NAND2x1_ASAP7_75t_R _27920_ (.A(_01721_),
    .B(_05457_),
    .Y(_11496_));
 AND2x4_ASAP7_75t_R _27921_ (.A(_11495_),
    .B(_11496_),
    .Y(_11497_));
 AND3x1_ASAP7_75t_R _27922_ (.A(_11452_),
    .B(_11484_),
    .C(_11487_),
    .Y(_11498_));
 XOR2x2_ASAP7_75t_R _27923_ (.A(_11497_),
    .B(_11498_),
    .Y(_11499_));
 BUFx12f_ASAP7_75t_R _27924_ (.A(_11476_),
    .Y(_11500_));
 NOR2x1_ASAP7_75t_R _27925_ (.A(_01721_),
    .B(_11500_),
    .Y(_11501_));
 AO21x1_ASAP7_75t_R _27926_ (.A1(_11477_),
    .A2(_11499_),
    .B(_11501_),
    .Y(_03906_));
 NOR2x1_ASAP7_75t_R _27927_ (.A(_01720_),
    .B(_05464_),
    .Y(_11502_));
 AND5x1_ASAP7_75t_R _27928_ (.A(_11431_),
    .B(_11435_),
    .C(_11459_),
    .D(_11469_),
    .E(_11484_),
    .Y(_11503_));
 AND4x1_ASAP7_75t_R _27929_ (.A(_11464_),
    .B(_11495_),
    .C(_11496_),
    .D(_11503_),
    .Y(_11504_));
 NAND2x1_ASAP7_75t_R _27930_ (.A(_11485_),
    .B(_11504_),
    .Y(_11505_));
 OA222x2_ASAP7_75t_R _27931_ (.A1(_02049_),
    .A2(_05471_),
    .B1(_05502_),
    .B2(_01952_),
    .C1(_01406_),
    .C2(_11455_),
    .Y(_11506_));
 INVx1_ASAP7_75t_R _27932_ (.A(_11506_),
    .Y(_11507_));
 AO221x1_ASAP7_75t_R _27933_ (.A1(\alu_adder_result_ex[13] ),
    .A2(_10827_),
    .B1(_05476_),
    .B2(net4),
    .C(_11507_),
    .Y(_11508_));
 AND2x6_ASAP7_75t_R _27934_ (.A(_05463_),
    .B(_11508_),
    .Y(_11509_));
 XNOR2x2_ASAP7_75t_R _27935_ (.A(_11505_),
    .B(_11509_),
    .Y(_11510_));
 NAND2x1_ASAP7_75t_R _27936_ (.A(_01720_),
    .B(_11472_),
    .Y(_11511_));
 OR3x1_ASAP7_75t_R _27937_ (.A(_01720_),
    .B(_11472_),
    .C(_11505_),
    .Y(_11512_));
 AO21x1_ASAP7_75t_R _27938_ (.A1(_11511_),
    .A2(_11512_),
    .B(_05467_),
    .Y(_11513_));
 OA21x2_ASAP7_75t_R _27939_ (.A1(_11502_),
    .A2(_11510_),
    .B(_11513_),
    .Y(_03907_));
 NOR2x1_ASAP7_75t_R _27940_ (.A(_01719_),
    .B(_05464_),
    .Y(_11514_));
 INVx1_ASAP7_75t_R _27941_ (.A(_11514_),
    .Y(_11515_));
 OA22x2_ASAP7_75t_R _27942_ (.A1(_02048_),
    .A2(_05471_),
    .B1(_11455_),
    .B2(_01407_),
    .Y(_11516_));
 OAI21x1_ASAP7_75t_R _27943_ (.A1(_01951_),
    .A2(_05503_),
    .B(_11516_),
    .Y(_11517_));
 AO21x2_ASAP7_75t_R _27944_ (.A1(net5),
    .A2(_05476_),
    .B(_11517_),
    .Y(_11518_));
 OA21x2_ASAP7_75t_R _27945_ (.A1(_15770_),
    .A2(_15771_),
    .B(_10827_),
    .Y(_11519_));
 OAI21x1_ASAP7_75t_R _27946_ (.A1(_11518_),
    .A2(_11519_),
    .B(_05466_),
    .Y(_11520_));
 NOR2x1_ASAP7_75t_R _27947_ (.A(_11502_),
    .B(_11509_),
    .Y(_11521_));
 NAND2x1_ASAP7_75t_R _27948_ (.A(_11452_),
    .B(_11504_),
    .Y(_11522_));
 OR2x6_ASAP7_75t_R _27949_ (.A(_11521_),
    .B(_11522_),
    .Y(_11523_));
 AO21x1_ASAP7_75t_R _27950_ (.A1(_11515_),
    .A2(_11520_),
    .B(_11523_),
    .Y(_11524_));
 AND2x6_ASAP7_75t_R _27951_ (.A(_05459_),
    .B(_05716_),
    .Y(_11525_));
 AOI21x1_ASAP7_75t_R _27952_ (.A1(_11523_),
    .A2(_11520_),
    .B(_11525_),
    .Y(_11526_));
 OA21x2_ASAP7_75t_R _27953_ (.A1(_11472_),
    .A2(_11523_),
    .B(_11514_),
    .Y(_11527_));
 AO21x1_ASAP7_75t_R _27954_ (.A1(_11524_),
    .A2(_11526_),
    .B(_11527_),
    .Y(_03908_));
 OA22x2_ASAP7_75t_R _27955_ (.A1(_02047_),
    .A2(_05471_),
    .B1(_11455_),
    .B2(_01408_),
    .Y(_11528_));
 OAI21x1_ASAP7_75t_R _27956_ (.A1(_01950_),
    .A2(_05503_),
    .B(_11528_),
    .Y(_11529_));
 AO221x1_ASAP7_75t_R _27957_ (.A1(\alu_adder_result_ex[15] ),
    .A2(_10827_),
    .B1(_05476_),
    .B2(net6),
    .C(_11529_),
    .Y(_11530_));
 AND2x4_ASAP7_75t_R _27958_ (.A(_05464_),
    .B(_11530_),
    .Y(_11531_));
 NOR2x1_ASAP7_75t_R _27959_ (.A(_01718_),
    .B(_05464_),
    .Y(_11532_));
 NOR2x1_ASAP7_75t_R _27960_ (.A(_11531_),
    .B(_11532_),
    .Y(_11533_));
 AND2x2_ASAP7_75t_R _27961_ (.A(_11515_),
    .B(_11520_),
    .Y(_11534_));
 OR3x1_ASAP7_75t_R _27962_ (.A(_11505_),
    .B(_11521_),
    .C(_11534_),
    .Y(_11535_));
 AND2x2_ASAP7_75t_R _27963_ (.A(_11533_),
    .B(_11535_),
    .Y(_11536_));
 OA21x2_ASAP7_75t_R _27964_ (.A1(_11518_),
    .A2(_11519_),
    .B(_05464_),
    .Y(_11537_));
 OA222x2_ASAP7_75t_R _27965_ (.A1(_11502_),
    .A2(_11509_),
    .B1(_11514_),
    .B2(_11537_),
    .C1(_11531_),
    .C2(_11532_),
    .Y(_11538_));
 AND3x4_ASAP7_75t_R _27966_ (.A(_11485_),
    .B(_11504_),
    .C(_11538_),
    .Y(_11539_));
 OR3x1_ASAP7_75t_R _27967_ (.A(_11525_),
    .B(_11536_),
    .C(_11539_),
    .Y(_11540_));
 OAI21x1_ASAP7_75t_R _27968_ (.A1(_01718_),
    .A2(_11477_),
    .B(_11540_),
    .Y(_03909_));
 BUFx6f_ASAP7_75t_R _27969_ (.A(_05467_),
    .Y(_11541_));
 INVx1_ASAP7_75t_R _27970_ (.A(_01717_),
    .Y(_11542_));
 OR4x1_ASAP7_75t_R _27971_ (.A(_11521_),
    .B(_11522_),
    .C(_11534_),
    .D(_11533_),
    .Y(_11543_));
 OR3x1_ASAP7_75t_R _27972_ (.A(_01717_),
    .B(_05716_),
    .C(_11543_),
    .Y(_11544_));
 OA21x2_ASAP7_75t_R _27973_ (.A1(_11542_),
    .A2(_18717_),
    .B(_11544_),
    .Y(_11545_));
 AND2x2_ASAP7_75t_R _27974_ (.A(_01409_),
    .B(_11479_),
    .Y(_11546_));
 OA222x2_ASAP7_75t_R _27975_ (.A1(_02046_),
    .A2(_05471_),
    .B1(_11478_),
    .B2(_11546_),
    .C1(_05502_),
    .C2(_01949_),
    .Y(_11547_));
 OA21x2_ASAP7_75t_R _27976_ (.A1(_08021_),
    .A2(_11432_),
    .B(_11547_),
    .Y(_11548_));
 AO31x2_ASAP7_75t_R _27977_ (.A1(_16007_),
    .A2(_16014_),
    .A3(_16018_),
    .B(_05158_),
    .Y(_11549_));
 AO21x1_ASAP7_75t_R _27978_ (.A1(_11548_),
    .A2(_11549_),
    .B(_05456_),
    .Y(_11550_));
 BUFx6f_ASAP7_75t_R _27979_ (.A(_11550_),
    .Y(_11551_));
 XOR2x2_ASAP7_75t_R _27980_ (.A(_11543_),
    .B(_11551_),
    .Y(_11552_));
 AO21x1_ASAP7_75t_R _27981_ (.A1(_11542_),
    .A2(_11475_),
    .B(_11552_),
    .Y(_11553_));
 OA21x2_ASAP7_75t_R _27982_ (.A1(_11541_),
    .A2(_11545_),
    .B(_11553_),
    .Y(_03910_));
 NOR2x1_ASAP7_75t_R _27983_ (.A(_01716_),
    .B(_05466_),
    .Y(_11554_));
 OAI21x1_ASAP7_75t_R _27984_ (.A1(_01717_),
    .A2(_05466_),
    .B(_11551_),
    .Y(_11555_));
 AND2x2_ASAP7_75t_R _27985_ (.A(_11539_),
    .B(_11555_),
    .Y(_11556_));
 NAND2x1_ASAP7_75t_R _27986_ (.A(_18717_),
    .B(_11556_),
    .Y(_11557_));
 OA222x2_ASAP7_75t_R _27987_ (.A1(_02045_),
    .A2(_05471_),
    .B1(_05502_),
    .B2(_01948_),
    .C1(_01410_),
    .C2(_11455_),
    .Y(_11558_));
 OA21x2_ASAP7_75t_R _27988_ (.A1(_08023_),
    .A2(_11432_),
    .B(_11558_),
    .Y(_11559_));
 NAND2x1_ASAP7_75t_R _27989_ (.A(\alu_adder_result_ex[17] ),
    .B(_10827_),
    .Y(_11560_));
 AOI21x1_ASAP7_75t_R _27990_ (.A1(_11559_),
    .A2(_11560_),
    .B(_05458_),
    .Y(_11561_));
 AO21x2_ASAP7_75t_R _27991_ (.A1(_11559_),
    .A2(_11560_),
    .B(_05456_),
    .Y(_11562_));
 OA21x2_ASAP7_75t_R _27992_ (.A1(_11551_),
    .A2(_11562_),
    .B(_05464_),
    .Y(_11563_));
 AOI221x1_ASAP7_75t_R _27993_ (.A1(_01717_),
    .A2(_11551_),
    .B1(_11562_),
    .B2(_01716_),
    .C(_11563_),
    .Y(_11564_));
 NAND2x1_ASAP7_75t_R _27994_ (.A(_11539_),
    .B(_11564_),
    .Y(_11565_));
 OA211x2_ASAP7_75t_R _27995_ (.A1(_11556_),
    .A2(_11561_),
    .B(_11565_),
    .C(_11476_),
    .Y(_11566_));
 AO21x1_ASAP7_75t_R _27996_ (.A1(_11554_),
    .A2(_11557_),
    .B(_11566_),
    .Y(_03911_));
 INVx1_ASAP7_75t_R _27997_ (.A(_01715_),
    .Y(_11567_));
 BUFx6f_ASAP7_75t_R _27998_ (.A(_11432_),
    .Y(_11568_));
 BUFx6f_ASAP7_75t_R _27999_ (.A(_11455_),
    .Y(_11569_));
 OA222x2_ASAP7_75t_R _28000_ (.A1(_02044_),
    .A2(_05499_),
    .B1(_05503_),
    .B2(_01947_),
    .C1(_01411_),
    .C2(_11569_),
    .Y(_11570_));
 OA211x2_ASAP7_75t_R _28001_ (.A1(_08025_),
    .A2(_11568_),
    .B(_11570_),
    .C(_05464_),
    .Y(_11571_));
 OAI21x1_ASAP7_75t_R _28002_ (.A1(_16267_),
    .A2(_05477_),
    .B(_11571_),
    .Y(_11572_));
 OA21x2_ASAP7_75t_R _28003_ (.A1(_11567_),
    .A2(_05465_),
    .B(_11572_),
    .Y(_11573_));
 AND4x1_ASAP7_75t_R _28004_ (.A(_11452_),
    .B(_11504_),
    .C(_11538_),
    .D(_11564_),
    .Y(_11574_));
 XNOR2x2_ASAP7_75t_R _28005_ (.A(_11573_),
    .B(_11574_),
    .Y(_11575_));
 NAND2x1_ASAP7_75t_R _28006_ (.A(_11490_),
    .B(_11575_),
    .Y(_11576_));
 OA21x2_ASAP7_75t_R _28007_ (.A1(_11567_),
    .A2(_11477_),
    .B(_11576_),
    .Y(_03912_));
 AND3x4_ASAP7_75t_R _28008_ (.A(_11539_),
    .B(_11564_),
    .C(_11573_),
    .Y(_11577_));
 OA222x2_ASAP7_75t_R _28009_ (.A1(_02043_),
    .A2(_05499_),
    .B1(_05503_),
    .B2(_01946_),
    .C1(_01412_),
    .C2(_11569_),
    .Y(_11578_));
 OA21x2_ASAP7_75t_R _28010_ (.A1(_08027_),
    .A2(_11568_),
    .B(_11578_),
    .Y(_11579_));
 OAI21x1_ASAP7_75t_R _28011_ (.A1(_16253_),
    .A2(_05477_),
    .B(_11579_),
    .Y(_11580_));
 NAND2x1_ASAP7_75t_R _28012_ (.A(_01714_),
    .B(_05457_),
    .Y(_11581_));
 OA21x2_ASAP7_75t_R _28013_ (.A1(_05457_),
    .A2(_11580_),
    .B(_11581_),
    .Y(_11582_));
 XOR2x2_ASAP7_75t_R _28014_ (.A(_11577_),
    .B(_11582_),
    .Y(_11583_));
 NOR2x1_ASAP7_75t_R _28015_ (.A(_01714_),
    .B(_11500_),
    .Y(_11584_));
 AO21x1_ASAP7_75t_R _28016_ (.A1(_11477_),
    .A2(_11583_),
    .B(_11584_),
    .Y(_03913_));
 NOR2x1_ASAP7_75t_R _28017_ (.A(_01713_),
    .B(_05464_),
    .Y(_11585_));
 AND2x2_ASAP7_75t_R _28018_ (.A(_01413_),
    .B(_11479_),
    .Y(_11586_));
 OA222x2_ASAP7_75t_R _28019_ (.A1(_02042_),
    .A2(_05499_),
    .B1(_11478_),
    .B2(_11586_),
    .C1(_05503_),
    .C2(_01944_),
    .Y(_11587_));
 OA21x2_ASAP7_75t_R _28020_ (.A1(_08030_),
    .A2(_11568_),
    .B(_11587_),
    .Y(_11588_));
 NAND2x1_ASAP7_75t_R _28021_ (.A(\alu_adder_result_ex[20] ),
    .B(_10827_),
    .Y(_11589_));
 AOI21x1_ASAP7_75t_R _28022_ (.A1(_11588_),
    .A2(_11589_),
    .B(_05457_),
    .Y(_11590_));
 AND5x2_ASAP7_75t_R _28023_ (.A(_11452_),
    .B(_11504_),
    .C(_11538_),
    .D(_11564_),
    .E(_11573_),
    .Y(_11591_));
 OA211x2_ASAP7_75t_R _28024_ (.A1(_11585_),
    .A2(_11590_),
    .B(_11591_),
    .C(_11582_),
    .Y(_11592_));
 NAND2x1_ASAP7_75t_R _28025_ (.A(_11582_),
    .B(_11591_),
    .Y(_11593_));
 INVx1_ASAP7_75t_R _28026_ (.A(_11590_),
    .Y(_11594_));
 AO21x1_ASAP7_75t_R _28027_ (.A1(_11593_),
    .A2(_11594_),
    .B(_11525_),
    .Y(_11595_));
 OAI21x1_ASAP7_75t_R _28028_ (.A1(_11472_),
    .A2(_11593_),
    .B(_11585_),
    .Y(_11596_));
 OAI21x1_ASAP7_75t_R _28029_ (.A1(_11592_),
    .A2(_11595_),
    .B(_11596_),
    .Y(_03914_));
 AND2x4_ASAP7_75t_R _28030_ (.A(_01712_),
    .B(_05458_),
    .Y(_11597_));
 OA211x2_ASAP7_75t_R _28031_ (.A1(_11585_),
    .A2(_11590_),
    .B(_11577_),
    .C(_11582_),
    .Y(_11598_));
 NAND2x1_ASAP7_75t_R _28032_ (.A(_18717_),
    .B(_11598_),
    .Y(_11599_));
 OA222x2_ASAP7_75t_R _28033_ (.A1(_02041_),
    .A2(_05471_),
    .B1(_05503_),
    .B2(_01943_),
    .C1(_01414_),
    .C2(_11569_),
    .Y(_11600_));
 OA21x2_ASAP7_75t_R _28034_ (.A1(_08034_),
    .A2(_11568_),
    .B(_11600_),
    .Y(_11601_));
 OA211x2_ASAP7_75t_R _28035_ (.A1(_16515_),
    .A2(_05477_),
    .B(_05464_),
    .C(_11601_),
    .Y(_11602_));
 OAI21x1_ASAP7_75t_R _28036_ (.A1(_11597_),
    .A2(_11602_),
    .B(_11598_),
    .Y(_11603_));
 OA211x2_ASAP7_75t_R _28037_ (.A1(_11598_),
    .A2(_11602_),
    .B(_11603_),
    .C(_11476_),
    .Y(_11604_));
 AOI21x1_ASAP7_75t_R _28038_ (.A1(_11597_),
    .A2(_11599_),
    .B(_11604_),
    .Y(_03915_));
 NOR2x1_ASAP7_75t_R _28039_ (.A(_01711_),
    .B(_05465_),
    .Y(_11605_));
 AOI21x1_ASAP7_75t_R _28040_ (.A1(_01712_),
    .A2(_05457_),
    .B(_11602_),
    .Y(_11606_));
 OA211x2_ASAP7_75t_R _28041_ (.A1(_11585_),
    .A2(_11590_),
    .B(_11606_),
    .C(_11582_),
    .Y(_11607_));
 AND2x4_ASAP7_75t_R _28042_ (.A(_11591_),
    .B(_11607_),
    .Y(_11608_));
 NAND2x1_ASAP7_75t_R _28043_ (.A(_18717_),
    .B(_11608_),
    .Y(_11609_));
 OA222x2_ASAP7_75t_R _28044_ (.A1(_02040_),
    .A2(_05499_),
    .B1(_05503_),
    .B2(_01942_),
    .C1(_01415_),
    .C2(_11569_),
    .Y(_11610_));
 OA21x2_ASAP7_75t_R _28045_ (.A1(_08036_),
    .A2(_11568_),
    .B(_11610_),
    .Y(_11611_));
 OA21x2_ASAP7_75t_R _28046_ (.A1(_16761_),
    .A2(_05477_),
    .B(_11611_),
    .Y(_11612_));
 NOR2x2_ASAP7_75t_R _28047_ (.A(_05457_),
    .B(_11612_),
    .Y(_11613_));
 OAI21x1_ASAP7_75t_R _28048_ (.A1(_11605_),
    .A2(_11613_),
    .B(_11608_),
    .Y(_11614_));
 OA211x2_ASAP7_75t_R _28049_ (.A1(_11608_),
    .A2(_11613_),
    .B(_11614_),
    .C(_11476_),
    .Y(_11615_));
 AO21x1_ASAP7_75t_R _28050_ (.A1(_11605_),
    .A2(_11609_),
    .B(_11615_),
    .Y(_03916_));
 OA222x2_ASAP7_75t_R _28051_ (.A1(_02039_),
    .A2(_05499_),
    .B1(_05503_),
    .B2(_01941_),
    .C1(_00007_),
    .C2(_11569_),
    .Y(_11616_));
 OA21x2_ASAP7_75t_R _28052_ (.A1(_08038_),
    .A2(_11568_),
    .B(_11616_),
    .Y(_11617_));
 OA211x2_ASAP7_75t_R _28053_ (.A1(_16753_),
    .A2(_05477_),
    .B(_05465_),
    .C(_11617_),
    .Y(_11618_));
 AOI21x1_ASAP7_75t_R _28054_ (.A1(_01710_),
    .A2(_05458_),
    .B(_11618_),
    .Y(_11619_));
 OA211x2_ASAP7_75t_R _28055_ (.A1(_11605_),
    .A2(_11613_),
    .B(_11607_),
    .C(_11577_),
    .Y(_11620_));
 XOR2x2_ASAP7_75t_R _28056_ (.A(_11619_),
    .B(_11620_),
    .Y(_11621_));
 NOR2x1_ASAP7_75t_R _28057_ (.A(_01710_),
    .B(_11500_),
    .Y(_11622_));
 AO21x1_ASAP7_75t_R _28058_ (.A1(_11477_),
    .A2(_11621_),
    .B(_11622_),
    .Y(_03917_));
 INVx1_ASAP7_75t_R _28059_ (.A(_01709_),
    .Y(_11623_));
 NAND2x1_ASAP7_75t_R _28060_ (.A(_11623_),
    .B(_05458_),
    .Y(_11624_));
 OA222x2_ASAP7_75t_R _28061_ (.A1(_02038_),
    .A2(_05500_),
    .B1(_05504_),
    .B2(_01940_),
    .C1(_00008_),
    .C2(_11569_),
    .Y(_11625_));
 INVx1_ASAP7_75t_R _28062_ (.A(_11625_),
    .Y(_11626_));
 AO221x1_ASAP7_75t_R _28063_ (.A1(\alu_adder_result_ex[24] ),
    .A2(_10828_),
    .B1(_05476_),
    .B2(net15),
    .C(_11626_),
    .Y(_11627_));
 NAND2x2_ASAP7_75t_R _28064_ (.A(_05465_),
    .B(_11627_),
    .Y(_11628_));
 OA211x2_ASAP7_75t_R _28065_ (.A1(_11605_),
    .A2(_11613_),
    .B(_11619_),
    .C(_11607_),
    .Y(_11629_));
 NAND2x1_ASAP7_75t_R _28066_ (.A(_11591_),
    .B(_11629_),
    .Y(_11630_));
 AO21x1_ASAP7_75t_R _28067_ (.A1(_11624_),
    .A2(_11628_),
    .B(_11630_),
    .Y(_11631_));
 AOI21x1_ASAP7_75t_R _28068_ (.A1(_11630_),
    .A2(_11628_),
    .B(_11525_),
    .Y(_11632_));
 OA211x2_ASAP7_75t_R _28069_ (.A1(_11472_),
    .A2(_11630_),
    .B(_11623_),
    .C(_05459_),
    .Y(_11633_));
 AO21x1_ASAP7_75t_R _28070_ (.A1(_11631_),
    .A2(_11632_),
    .B(_11633_),
    .Y(_03918_));
 AND2x2_ASAP7_75t_R _28071_ (.A(_00009_),
    .B(_11479_),
    .Y(_11634_));
 OA222x2_ASAP7_75t_R _28072_ (.A1(_02037_),
    .A2(_05500_),
    .B1(_11478_),
    .B2(_11634_),
    .C1(_05504_),
    .C2(_01939_),
    .Y(_11635_));
 OA21x2_ASAP7_75t_R _28073_ (.A1(_08042_),
    .A2(_11568_),
    .B(_11635_),
    .Y(_11636_));
 OA211x2_ASAP7_75t_R _28074_ (.A1(_16995_),
    .A2(_05477_),
    .B(_05465_),
    .C(_11636_),
    .Y(_11637_));
 AOI21x1_ASAP7_75t_R _28075_ (.A1(_01708_),
    .A2(_05458_),
    .B(_11637_),
    .Y(_11638_));
 NAND2x1_ASAP7_75t_R _28076_ (.A(_11624_),
    .B(_11628_),
    .Y(_11639_));
 AND3x4_ASAP7_75t_R _28077_ (.A(_11577_),
    .B(_11629_),
    .C(_11639_),
    .Y(_11640_));
 XOR2x2_ASAP7_75t_R _28078_ (.A(_11638_),
    .B(_11640_),
    .Y(_11641_));
 NOR2x1_ASAP7_75t_R _28079_ (.A(_01708_),
    .B(_11500_),
    .Y(_11642_));
 AO21x1_ASAP7_75t_R _28080_ (.A1(_11477_),
    .A2(_11641_),
    .B(_11642_),
    .Y(_03919_));
 OA222x2_ASAP7_75t_R _28081_ (.A1(_02036_),
    .A2(_05499_),
    .B1(_05504_),
    .B2(_01938_),
    .C1(_00010_),
    .C2(_11569_),
    .Y(_11643_));
 INVx1_ASAP7_75t_R _28082_ (.A(_11643_),
    .Y(_11644_));
 AO221x1_ASAP7_75t_R _28083_ (.A1(\alu_adder_result_ex[26] ),
    .A2(_10828_),
    .B1(_05476_),
    .B2(net17),
    .C(_11644_),
    .Y(_11645_));
 AND2x6_ASAP7_75t_R _28084_ (.A(_05465_),
    .B(_11645_),
    .Y(_11646_));
 INVx1_ASAP7_75t_R _28085_ (.A(_01707_),
    .Y(_11647_));
 AND2x4_ASAP7_75t_R _28086_ (.A(_11647_),
    .B(_05457_),
    .Y(_11648_));
 NOR2x1_ASAP7_75t_R _28087_ (.A(_11646_),
    .B(_11648_),
    .Y(_11649_));
 AND4x1_ASAP7_75t_R _28088_ (.A(_11591_),
    .B(_11629_),
    .C(_11638_),
    .D(_11639_),
    .Y(_11650_));
 XNOR2x2_ASAP7_75t_R _28089_ (.A(_11649_),
    .B(_11650_),
    .Y(_11651_));
 AND3x1_ASAP7_75t_R _28090_ (.A(_11647_),
    .B(_05459_),
    .C(_11472_),
    .Y(_11652_));
 AO21x1_ASAP7_75t_R _28091_ (.A1(_11477_),
    .A2(_11651_),
    .B(_11652_),
    .Y(_03920_));
 INVx1_ASAP7_75t_R _28092_ (.A(_11649_),
    .Y(_11653_));
 AND3x1_ASAP7_75t_R _28093_ (.A(_11638_),
    .B(_11640_),
    .C(_11653_),
    .Y(_11654_));
 AND2x2_ASAP7_75t_R _28094_ (.A(_00011_),
    .B(_11479_),
    .Y(_11655_));
 OA222x2_ASAP7_75t_R _28095_ (.A1(_02035_),
    .A2(_05499_),
    .B1(_11478_),
    .B2(_11655_),
    .C1(_05504_),
    .C2(_01937_),
    .Y(_11656_));
 OA21x2_ASAP7_75t_R _28096_ (.A1(_08046_),
    .A2(_11568_),
    .B(_11656_),
    .Y(_11657_));
 NAND2x1_ASAP7_75t_R _28097_ (.A(\alu_adder_result_ex[27] ),
    .B(_10828_),
    .Y(_11658_));
 AO21x2_ASAP7_75t_R _28098_ (.A1(_11657_),
    .A2(_11658_),
    .B(_05457_),
    .Y(_11659_));
 OAI21x1_ASAP7_75t_R _28099_ (.A1(_01706_),
    .A2(_05465_),
    .B(_11659_),
    .Y(_11660_));
 XOR2x2_ASAP7_75t_R _28100_ (.A(_11654_),
    .B(_11660_),
    .Y(_11661_));
 NOR2x1_ASAP7_75t_R _28101_ (.A(_01706_),
    .B(_11500_),
    .Y(_11662_));
 AO21x1_ASAP7_75t_R _28102_ (.A1(_11490_),
    .A2(_11661_),
    .B(_11662_),
    .Y(_03921_));
 AND2x2_ASAP7_75t_R _28103_ (.A(_00012_),
    .B(_11479_),
    .Y(_11663_));
 OA222x2_ASAP7_75t_R _28104_ (.A1(_02034_),
    .A2(_05499_),
    .B1(_11478_),
    .B2(_11663_),
    .C1(_05503_),
    .C2(_01936_),
    .Y(_11664_));
 OA21x2_ASAP7_75t_R _28105_ (.A1(_08048_),
    .A2(_11568_),
    .B(_11664_),
    .Y(_11665_));
 OA211x2_ASAP7_75t_R _28106_ (.A1(_04729_),
    .A2(_05477_),
    .B(_05465_),
    .C(_11665_),
    .Y(_11666_));
 AOI21x1_ASAP7_75t_R _28107_ (.A1(_01705_),
    .A2(_05458_),
    .B(_11666_),
    .Y(_11667_));
 AND3x1_ASAP7_75t_R _28108_ (.A(_11653_),
    .B(_11650_),
    .C(_11660_),
    .Y(_11668_));
 XOR2x2_ASAP7_75t_R _28109_ (.A(_11667_),
    .B(_11668_),
    .Y(_11669_));
 NOR2x1_ASAP7_75t_R _28110_ (.A(_01705_),
    .B(_11500_),
    .Y(_11670_));
 AO21x1_ASAP7_75t_R _28111_ (.A1(_11490_),
    .A2(_11669_),
    .B(_11670_),
    .Y(_03922_));
 OA222x2_ASAP7_75t_R _28112_ (.A1(_02033_),
    .A2(_05499_),
    .B1(_05504_),
    .B2(_01935_),
    .C1(_00013_),
    .C2(_11569_),
    .Y(_11671_));
 INVx1_ASAP7_75t_R _28113_ (.A(_11671_),
    .Y(_11672_));
 AO221x1_ASAP7_75t_R _28114_ (.A1(\alu_adder_result_ex[29] ),
    .A2(_10828_),
    .B1(_05476_),
    .B2(net20),
    .C(_11672_),
    .Y(_11673_));
 NAND2x1_ASAP7_75t_R _28115_ (.A(_05465_),
    .B(_11673_),
    .Y(_11674_));
 OA21x2_ASAP7_75t_R _28116_ (.A1(_01704_),
    .A2(_05466_),
    .B(_11674_),
    .Y(_11675_));
 OA211x2_ASAP7_75t_R _28117_ (.A1(_11646_),
    .A2(_11648_),
    .B(_11660_),
    .C(_11667_),
    .Y(_11676_));
 AND3x1_ASAP7_75t_R _28118_ (.A(_11638_),
    .B(_11640_),
    .C(_11676_),
    .Y(_11677_));
 XNOR2x2_ASAP7_75t_R _28119_ (.A(_11675_),
    .B(_11677_),
    .Y(_11678_));
 NOR2x1_ASAP7_75t_R _28120_ (.A(_01704_),
    .B(_11500_),
    .Y(_11679_));
 AO21x1_ASAP7_75t_R _28121_ (.A1(_11490_),
    .A2(_11678_),
    .B(_11679_),
    .Y(_03923_));
 AND3x1_ASAP7_75t_R _28122_ (.A(_01703_),
    .B(_11475_),
    .C(_11472_),
    .Y(_11680_));
 AOI21x1_ASAP7_75t_R _28123_ (.A1(_02330_),
    .A2(_11477_),
    .B(_11680_),
    .Y(_03924_));
 INVx1_ASAP7_75t_R _28124_ (.A(_01702_),
    .Y(_11681_));
 OA222x2_ASAP7_75t_R _28125_ (.A1(_02031_),
    .A2(_05500_),
    .B1(_05504_),
    .B2(_01933_),
    .C1(_00014_),
    .C2(_11569_),
    .Y(_11682_));
 OA211x2_ASAP7_75t_R _28126_ (.A1(_08052_),
    .A2(_11568_),
    .B(_11682_),
    .C(_05466_),
    .Y(_11683_));
 OAI21x1_ASAP7_75t_R _28127_ (.A1(_04983_),
    .A2(_05477_),
    .B(_11683_),
    .Y(_11684_));
 OA21x2_ASAP7_75t_R _28128_ (.A1(_11681_),
    .A2(_05466_),
    .B(_11684_),
    .Y(_11685_));
 INVx1_ASAP7_75t_R _28129_ (.A(_11675_),
    .Y(_11686_));
 AND2x2_ASAP7_75t_R _28130_ (.A(_11686_),
    .B(_11676_),
    .Y(_11687_));
 NAND2x1_ASAP7_75t_R _28131_ (.A(_11650_),
    .B(_11687_),
    .Y(_11688_));
 XNOR2x2_ASAP7_75t_R _28132_ (.A(_11685_),
    .B(_11688_),
    .Y(_11689_));
 AND3x1_ASAP7_75t_R _28133_ (.A(_11681_),
    .B(_05459_),
    .C(_11472_),
    .Y(_11690_));
 AO21x1_ASAP7_75t_R _28134_ (.A1(_11490_),
    .A2(_11689_),
    .B(_11690_),
    .Y(_03925_));
 OA222x2_ASAP7_75t_R _28135_ (.A1(_02030_),
    .A2(_05500_),
    .B1(_05504_),
    .B2(_01932_),
    .C1(_00015_),
    .C2(_11569_),
    .Y(_11691_));
 INVx1_ASAP7_75t_R _28136_ (.A(_11691_),
    .Y(_11692_));
 AO221x1_ASAP7_75t_R _28137_ (.A1(\alu_adder_result_ex[31] ),
    .A2(_10828_),
    .B1(_05476_),
    .B2(net22),
    .C(_11692_),
    .Y(_11693_));
 NAND2x1_ASAP7_75t_R _28138_ (.A(_05466_),
    .B(_11693_),
    .Y(_11694_));
 OA21x2_ASAP7_75t_R _28139_ (.A1(_01701_),
    .A2(_05466_),
    .B(_11694_),
    .Y(_11695_));
 AND4x1_ASAP7_75t_R _28140_ (.A(_11638_),
    .B(_11640_),
    .C(_11685_),
    .D(_11687_),
    .Y(_11696_));
 XNOR2x2_ASAP7_75t_R _28141_ (.A(_11695_),
    .B(_11696_),
    .Y(_11697_));
 NOR2x1_ASAP7_75t_R _28142_ (.A(_01701_),
    .B(_11500_),
    .Y(_11698_));
 AO21x1_ASAP7_75t_R _28143_ (.A1(_11490_),
    .A2(_11697_),
    .B(_11698_),
    .Y(_03926_));
 AND3x1_ASAP7_75t_R _28144_ (.A(_01700_),
    .B(_11475_),
    .C(_11472_),
    .Y(_11699_));
 AOI21x1_ASAP7_75t_R _28145_ (.A1(_02332_),
    .A2(_11477_),
    .B(_11699_),
    .Y(_03927_));
 NOR2x1_ASAP7_75t_R _28146_ (.A(_11440_),
    .B(_11441_),
    .Y(_11700_));
 XNOR2x2_ASAP7_75t_R _28147_ (.A(_11436_),
    .B(_11700_),
    .Y(_11701_));
 NOR2x1_ASAP7_75t_R _28148_ (.A(_01699_),
    .B(_11500_),
    .Y(_11702_));
 AO21x1_ASAP7_75t_R _28149_ (.A1(_11490_),
    .A2(_11701_),
    .B(_11702_),
    .Y(_03928_));
 OR3x1_ASAP7_75t_R _28150_ (.A(_02329_),
    .B(_05521_),
    .C(_11700_),
    .Y(_11703_));
 XNOR2x2_ASAP7_75t_R _28151_ (.A(_11444_),
    .B(_11703_),
    .Y(_11704_));
 NOR2x1_ASAP7_75t_R _28152_ (.A(_01698_),
    .B(_11500_),
    .Y(_11705_));
 AO21x1_ASAP7_75t_R _28153_ (.A1(_11490_),
    .A2(_11704_),
    .B(_11705_),
    .Y(_03929_));
 NAND2x1_ASAP7_75t_R _28154_ (.A(_11436_),
    .B(_11445_),
    .Y(_11706_));
 AND2x4_ASAP7_75t_R _28155_ (.A(_11433_),
    .B(_11449_),
    .Y(_11707_));
 AND2x2_ASAP7_75t_R _28156_ (.A(_11436_),
    .B(_11445_),
    .Y(_11708_));
 NAND2x1_ASAP7_75t_R _28157_ (.A(_18717_),
    .B(_11708_),
    .Y(_11709_));
 AOI21x1_ASAP7_75t_R _28158_ (.A1(_01697_),
    .A2(_18717_),
    .B(_05466_),
    .Y(_11710_));
 OR3x1_ASAP7_75t_R _28159_ (.A(_11706_),
    .B(_11707_),
    .C(_11710_),
    .Y(_11711_));
 INVx1_ASAP7_75t_R _28160_ (.A(_11711_),
    .Y(_11712_));
 AO221x1_ASAP7_75t_R _28161_ (.A1(_11706_),
    .A2(_11707_),
    .B1(_11450_),
    .B2(_11709_),
    .C(_11712_),
    .Y(_03930_));
 XOR2x2_ASAP7_75t_R _28162_ (.A(_11435_),
    .B(_11485_),
    .Y(_11713_));
 NOR2x1_ASAP7_75t_R _28163_ (.A(_01696_),
    .B(_11476_),
    .Y(_11714_));
 AO21x1_ASAP7_75t_R _28164_ (.A1(_11490_),
    .A2(_11713_),
    .B(_11714_),
    .Y(_03931_));
 NAND2x2_ASAP7_75t_R _28165_ (.A(_05467_),
    .B(_11462_),
    .Y(_11715_));
 AOI22x1_ASAP7_75t_R _28166_ (.A1(_11453_),
    .A2(_11715_),
    .B1(_11525_),
    .B2(_01695_),
    .Y(_11716_));
 NAND2x1_ASAP7_75t_R _28167_ (.A(_18717_),
    .B(_11463_),
    .Y(_11717_));
 AO21x1_ASAP7_75t_R _28168_ (.A1(_11715_),
    .A2(_11717_),
    .B(_11453_),
    .Y(_11718_));
 OA21x2_ASAP7_75t_R _28169_ (.A1(_11463_),
    .A2(_11716_),
    .B(_11718_),
    .Y(_03932_));
 AND3x1_ASAP7_75t_R _28170_ (.A(_11435_),
    .B(_11464_),
    .C(_11485_),
    .Y(_11719_));
 XNOR2x2_ASAP7_75t_R _28171_ (.A(_11459_),
    .B(_11719_),
    .Y(_11720_));
 OR3x1_ASAP7_75t_R _28172_ (.A(_01694_),
    .B(_05467_),
    .C(_18717_),
    .Y(_11721_));
 OAI21x1_ASAP7_75t_R _28173_ (.A1(_11525_),
    .A2(_11720_),
    .B(_11721_),
    .Y(_03933_));
 BUFx12f_ASAP7_75t_R _28174_ (.A(_05711_),
    .Y(_11722_));
 BUFx12f_ASAP7_75t_R _28175_ (.A(_11722_),
    .Y(_11723_));
 BUFx6f_ASAP7_75t_R _28176_ (.A(_11723_),
    .Y(_11724_));
 BUFx6f_ASAP7_75t_R _28177_ (.A(_05539_),
    .Y(_11725_));
 OR3x1_ASAP7_75t_R _28178_ (.A(_05543_),
    .B(_05710_),
    .C(_05536_),
    .Y(_11726_));
 AND3x1_ASAP7_75t_R _28179_ (.A(net149),
    .B(_02202_),
    .C(_05709_),
    .Y(_11727_));
 BUFx6f_ASAP7_75t_R _28180_ (.A(_11727_),
    .Y(_11728_));
 OAI21x1_ASAP7_75t_R _28181_ (.A1(_05544_),
    .A2(_05536_),
    .B(_11728_),
    .Y(_11729_));
 NOR2x1_ASAP7_75t_R _28182_ (.A(_05711_),
    .B(_11728_),
    .Y(_11730_));
 NAND2x1_ASAP7_75t_R _28183_ (.A(_05531_),
    .B(_05535_),
    .Y(_11731_));
 AO33x2_ASAP7_75t_R _28184_ (.A1(_11725_),
    .A2(_11726_),
    .A3(_11729_),
    .B1(_11730_),
    .B2(_11731_),
    .B3(_05524_),
    .Y(_11732_));
 OA211x2_ASAP7_75t_R _28185_ (.A1(_10810_),
    .A2(_10812_),
    .B(_05704_),
    .C(_05189_),
    .Y(_11733_));
 OR3x2_ASAP7_75t_R _28186_ (.A(_05406_),
    .B(_10839_),
    .C(_11733_),
    .Y(_11734_));
 OR3x1_ASAP7_75t_R _28187_ (.A(_05545_),
    .B(_11732_),
    .C(_11734_),
    .Y(_11735_));
 INVx1_ASAP7_75t_R _28188_ (.A(_11735_),
    .Y(_11736_));
 AND3x4_ASAP7_75t_R _28189_ (.A(_10848_),
    .B(_10850_),
    .C(_11736_),
    .Y(_11737_));
 AND3x4_ASAP7_75t_R _28190_ (.A(_11724_),
    .B(_10809_),
    .C(_11737_),
    .Y(_11738_));
 INVx1_ASAP7_75t_R _28191_ (.A(_10848_),
    .Y(_11739_));
 AOI21x1_ASAP7_75t_R _28192_ (.A1(_05149_),
    .A2(_05176_),
    .B(_10849_),
    .Y(_11740_));
 OR3x2_ASAP7_75t_R _28193_ (.A(_11739_),
    .B(_11740_),
    .C(_11735_),
    .Y(_11741_));
 BUFx6f_ASAP7_75t_R _28194_ (.A(_11725_),
    .Y(_11742_));
 OA211x2_ASAP7_75t_R _28195_ (.A1(_10824_),
    .A2(_11741_),
    .B(_11728_),
    .C(_11742_),
    .Y(_11743_));
 NOR2x1_ASAP7_75t_R _28196_ (.A(_05545_),
    .B(_11734_),
    .Y(_11744_));
 AND3x1_ASAP7_75t_R _28197_ (.A(_10848_),
    .B(_10850_),
    .C(_11744_),
    .Y(_11745_));
 BUFx6f_ASAP7_75t_R _28198_ (.A(_05537_),
    .Y(_11746_));
 BUFx6f_ASAP7_75t_R _28199_ (.A(_11746_),
    .Y(_11747_));
 AND2x2_ASAP7_75t_R _28200_ (.A(_11747_),
    .B(_11728_),
    .Y(_11748_));
 AND3x1_ASAP7_75t_R _28201_ (.A(_10809_),
    .B(_11745_),
    .C(_11748_),
    .Y(_11749_));
 BUFx6f_ASAP7_75t_R _28202_ (.A(_11749_),
    .Y(_11750_));
 OR3x2_ASAP7_75t_R _28203_ (.A(_11738_),
    .B(_11743_),
    .C(_11750_),
    .Y(_11751_));
 BUFx3_ASAP7_75t_R _28204_ (.A(_11751_),
    .Y(_11752_));
 NAND2x1_ASAP7_75t_R _28205_ (.A(_05533_),
    .B(_05710_),
    .Y(_11753_));
 BUFx12f_ASAP7_75t_R _28206_ (.A(_11724_),
    .Y(_11754_));
 NAND2x1_ASAP7_75t_R _28207_ (.A(_11754_),
    .B(_01692_),
    .Y(_11755_));
 BUFx6f_ASAP7_75t_R _28208_ (.A(_11750_),
    .Y(_11756_));
 NOR2x1_ASAP7_75t_R _28209_ (.A(_01693_),
    .B(_11756_),
    .Y(_11757_));
 NOR2x2_ASAP7_75t_R _28210_ (.A(_11738_),
    .B(_11743_),
    .Y(_11758_));
 BUFx3_ASAP7_75t_R _28211_ (.A(_11758_),
    .Y(_11759_));
 AO32x1_ASAP7_75t_R _28212_ (.A1(_11752_),
    .A2(_11753_),
    .A3(_11755_),
    .B1(_11757_),
    .B2(_11759_),
    .Y(_03934_));
 AND2x4_ASAP7_75t_R _28213_ (.A(_10809_),
    .B(_11737_),
    .Y(_11760_));
 AO21x1_ASAP7_75t_R _28214_ (.A1(_11724_),
    .A2(_11728_),
    .B(_05708_),
    .Y(_11761_));
 OA211x2_ASAP7_75t_R _28215_ (.A1(_10824_),
    .A2(_11741_),
    .B(_11748_),
    .C(_05710_),
    .Y(_11762_));
 AO21x2_ASAP7_75t_R _28216_ (.A1(_11760_),
    .A2(_11761_),
    .B(_11762_),
    .Y(_11763_));
 BUFx3_ASAP7_75t_R _28217_ (.A(_11763_),
    .Y(_11764_));
 BUFx12f_ASAP7_75t_R _28218_ (.A(_05708_),
    .Y(_11765_));
 BUFx6f_ASAP7_75t_R _28219_ (.A(_11765_),
    .Y(_11766_));
 BUFx6f_ASAP7_75t_R _28220_ (.A(_05708_),
    .Y(_11767_));
 NAND2x1_ASAP7_75t_R _28221_ (.A(_01691_),
    .B(_11767_),
    .Y(_11768_));
 OA21x2_ASAP7_75t_R _28222_ (.A1(net115),
    .A2(_11766_),
    .B(_11768_),
    .Y(_11769_));
 AND2x4_ASAP7_75t_R _28223_ (.A(_11723_),
    .B(_11728_),
    .Y(_11770_));
 AOI21x1_ASAP7_75t_R _28224_ (.A1(_11760_),
    .A2(_11770_),
    .B(_11762_),
    .Y(_11771_));
 BUFx6f_ASAP7_75t_R _28225_ (.A(_11771_),
    .Y(_11772_));
 AND3x4_ASAP7_75t_R _28226_ (.A(_05708_),
    .B(_10809_),
    .C(_11737_),
    .Y(_11773_));
 BUFx12f_ASAP7_75t_R _28227_ (.A(_11773_),
    .Y(_11774_));
 NOR2x1_ASAP7_75t_R _28228_ (.A(_01692_),
    .B(_11774_),
    .Y(_11775_));
 AO22x1_ASAP7_75t_R _28229_ (.A1(_11764_),
    .A2(_11769_),
    .B1(_11772_),
    .B2(_11775_),
    .Y(_03935_));
 NAND2x2_ASAP7_75t_R _28230_ (.A(_02205_),
    .B(_11770_),
    .Y(_11776_));
 BUFx12f_ASAP7_75t_R _28231_ (.A(_11776_),
    .Y(_11777_));
 BUFx6f_ASAP7_75t_R _28232_ (.A(_11777_),
    .Y(_11778_));
 BUFx6f_ASAP7_75t_R _28233_ (.A(_11776_),
    .Y(_11779_));
 NAND2x1_ASAP7_75t_R _28234_ (.A(_01691_),
    .B(_11779_),
    .Y(_11780_));
 OA21x2_ASAP7_75t_R _28235_ (.A1(net115),
    .A2(_11778_),
    .B(_11780_),
    .Y(_03936_));
 OA222x2_ASAP7_75t_R _28236_ (.A1(_00749_),
    .A2(_05500_),
    .B1(_07266_),
    .B2(_01945_),
    .C1(_18712_),
    .C2(_05477_),
    .Y(_11781_));
 OR4x1_ASAP7_75t_R _28237_ (.A(_11739_),
    .B(_11740_),
    .C(_11732_),
    .D(_11734_),
    .Y(_11782_));
 BUFx6f_ASAP7_75t_R _28238_ (.A(_11782_),
    .Y(_11783_));
 NOR2x2_ASAP7_75t_R _28239_ (.A(_10824_),
    .B(_11783_),
    .Y(_11784_));
 BUFx6f_ASAP7_75t_R _28240_ (.A(_11784_),
    .Y(_11785_));
 AO21x1_ASAP7_75t_R _28241_ (.A1(_05536_),
    .A2(_11785_),
    .B(_07348_),
    .Y(_11786_));
 AOI21x1_ASAP7_75t_R _28242_ (.A1(_05545_),
    .A2(_11785_),
    .B(_11541_),
    .Y(_11787_));
 AOI22x1_ASAP7_75t_R _28243_ (.A1(_11541_),
    .A2(_11781_),
    .B1(_11786_),
    .B2(_11787_),
    .Y(_03937_));
 BUFx12f_ASAP7_75t_R _28244_ (.A(_05459_),
    .Y(_11788_));
 BUFx6f_ASAP7_75t_R _28245_ (.A(_11783_),
    .Y(_11789_));
 INVx1_ASAP7_75t_R _28246_ (.A(_00267_),
    .Y(_11790_));
 OR2x6_ASAP7_75t_R _28247_ (.A(_00021_),
    .B(_11790_),
    .Y(_11791_));
 OR3x2_ASAP7_75t_R _28248_ (.A(_01668_),
    .B(_01669_),
    .C(_01670_),
    .Y(_11792_));
 OR3x2_ASAP7_75t_R _28249_ (.A(_01666_),
    .B(_01667_),
    .C(_11792_),
    .Y(_11793_));
 OR3x1_ASAP7_75t_R _28250_ (.A(_00022_),
    .B(_01665_),
    .C(_11793_),
    .Y(_11794_));
 OR4x1_ASAP7_75t_R _28251_ (.A(_10825_),
    .B(_11789_),
    .C(_11791_),
    .D(_11794_),
    .Y(_11795_));
 XNOR2x2_ASAP7_75t_R _28252_ (.A(_01690_),
    .B(_11795_),
    .Y(_11796_));
 AOI21x1_ASAP7_75t_R _28253_ (.A1(_11788_),
    .A2(_11796_),
    .B(_11483_),
    .Y(_03938_));
 BUFx6f_ASAP7_75t_R _28254_ (.A(_00750_),
    .Y(_11797_));
 OR3x1_ASAP7_75t_R _28255_ (.A(_11797_),
    .B(_00264_),
    .C(_11731_),
    .Y(_11798_));
 AO21x2_ASAP7_75t_R _28256_ (.A1(_00266_),
    .A2(_11798_),
    .B(_00021_),
    .Y(_11799_));
 OR3x1_ASAP7_75t_R _28257_ (.A(_01690_),
    .B(_11794_),
    .C(_11799_),
    .Y(_11800_));
 OR3x1_ASAP7_75t_R _28258_ (.A(_10825_),
    .B(_11789_),
    .C(_11800_),
    .Y(_11801_));
 XOR2x2_ASAP7_75t_R _28259_ (.A(_07316_),
    .B(_11801_),
    .Y(_11802_));
 OA21x2_ASAP7_75t_R _28260_ (.A1(_11541_),
    .A2(_11802_),
    .B(_11495_),
    .Y(_03939_));
 BUFx12f_ASAP7_75t_R _28261_ (.A(_05459_),
    .Y(_11803_));
 OR2x6_ASAP7_75t_R _28262_ (.A(_10824_),
    .B(_11783_),
    .Y(_11804_));
 BUFx12f_ASAP7_75t_R _28263_ (.A(_11804_),
    .Y(_11805_));
 OR3x2_ASAP7_75t_R _28264_ (.A(_01690_),
    .B(_11791_),
    .C(_11794_),
    .Y(_11806_));
 OR5x1_ASAP7_75t_R _28265_ (.A(_01688_),
    .B(_07316_),
    .C(_11509_),
    .D(_11805_),
    .E(_11806_),
    .Y(_11807_));
 OA21x2_ASAP7_75t_R _28266_ (.A1(_10824_),
    .A2(_11783_),
    .B(_05458_),
    .Y(_11808_));
 NOR2x1_ASAP7_75t_R _28267_ (.A(_07316_),
    .B(_11806_),
    .Y(_11809_));
 NOR2x1_ASAP7_75t_R _28268_ (.A(_11509_),
    .B(_11809_),
    .Y(_11810_));
 OAI21x1_ASAP7_75t_R _28269_ (.A1(_11808_),
    .A2(_11810_),
    .B(_01688_),
    .Y(_11811_));
 OA211x2_ASAP7_75t_R _28270_ (.A1(_11803_),
    .A2(_11509_),
    .B(_11807_),
    .C(_11811_),
    .Y(_03940_));
 OR3x1_ASAP7_75t_R _28271_ (.A(_01688_),
    .B(_07316_),
    .C(_11800_),
    .Y(_11812_));
 BUFx6f_ASAP7_75t_R _28272_ (.A(_11808_),
    .Y(_11813_));
 AO21x1_ASAP7_75t_R _28273_ (.A1(_11520_),
    .A2(_11812_),
    .B(_11813_),
    .Y(_11814_));
 BUFx12f_ASAP7_75t_R _28274_ (.A(_11805_),
    .Y(_11815_));
 OR4x1_ASAP7_75t_R _28275_ (.A(_01687_),
    .B(_01688_),
    .C(_07316_),
    .D(_11800_),
    .Y(_11816_));
 OAI21x1_ASAP7_75t_R _28276_ (.A1(_11815_),
    .A2(_11816_),
    .B(_11803_),
    .Y(_11817_));
 AOI22x1_ASAP7_75t_R _28277_ (.A1(_01687_),
    .A2(_11814_),
    .B1(_11817_),
    .B2(_11520_),
    .Y(_03941_));
 NAND2x1_ASAP7_75t_R _28278_ (.A(_05467_),
    .B(_11530_),
    .Y(_11818_));
 BUFx6f_ASAP7_75t_R _28279_ (.A(_11784_),
    .Y(_11819_));
 OR4x1_ASAP7_75t_R _28280_ (.A(_01687_),
    .B(_01688_),
    .C(_07316_),
    .D(_11806_),
    .Y(_11820_));
 NOR2x1_ASAP7_75t_R _28281_ (.A(_07328_),
    .B(_11820_),
    .Y(_11821_));
 AO21x1_ASAP7_75t_R _28282_ (.A1(_11819_),
    .A2(_11821_),
    .B(_11541_),
    .Y(_11822_));
 AO21x1_ASAP7_75t_R _28283_ (.A1(_11818_),
    .A2(_11820_),
    .B(_11813_),
    .Y(_11823_));
 AOI22x1_ASAP7_75t_R _28284_ (.A1(_11818_),
    .A2(_11822_),
    .B1(_11823_),
    .B2(_07328_),
    .Y(_03942_));
 OR3x2_ASAP7_75t_R _28285_ (.A(_01685_),
    .B(_07328_),
    .C(_11816_),
    .Y(_11824_));
 OAI21x1_ASAP7_75t_R _28286_ (.A1(_11815_),
    .A2(_11824_),
    .B(_11803_),
    .Y(_11825_));
 OA21x2_ASAP7_75t_R _28287_ (.A1(_07328_),
    .A2(_11816_),
    .B(_11551_),
    .Y(_11826_));
 OA21x2_ASAP7_75t_R _28288_ (.A1(_11808_),
    .A2(_11826_),
    .B(_01685_),
    .Y(_11827_));
 AOI21x1_ASAP7_75t_R _28289_ (.A1(_11551_),
    .A2(_11825_),
    .B(_11827_),
    .Y(_03943_));
 OR3x2_ASAP7_75t_R _28290_ (.A(_01685_),
    .B(_07328_),
    .C(_11820_),
    .Y(_11828_));
 AO21x1_ASAP7_75t_R _28291_ (.A1(_11562_),
    .A2(_11828_),
    .B(_11813_),
    .Y(_11829_));
 NOR2x1_ASAP7_75t_R _28292_ (.A(_07335_),
    .B(_11828_),
    .Y(_11830_));
 AO21x1_ASAP7_75t_R _28293_ (.A1(_11785_),
    .A2(_11830_),
    .B(_11541_),
    .Y(_11831_));
 AOI22x1_ASAP7_75t_R _28294_ (.A1(_07335_),
    .A2(_11829_),
    .B1(_11831_),
    .B2(_11562_),
    .Y(_03944_));
 BUFx12f_ASAP7_75t_R _28295_ (.A(_11805_),
    .Y(_11832_));
 NOR3x1_ASAP7_75t_R _28296_ (.A(_07335_),
    .B(_11832_),
    .C(_11824_),
    .Y(_11833_));
 NAND2x1_ASAP7_75t_R _28297_ (.A(_00023_),
    .B(_11475_),
    .Y(_11834_));
 OR5x1_ASAP7_75t_R _28298_ (.A(_00023_),
    .B(_07335_),
    .C(_05467_),
    .D(_11805_),
    .E(_11824_),
    .Y(_11835_));
 OA211x2_ASAP7_75t_R _28299_ (.A1(_11833_),
    .A2(_11834_),
    .B(_11835_),
    .C(_11572_),
    .Y(_03945_));
 OR3x2_ASAP7_75t_R _28300_ (.A(_00023_),
    .B(_07335_),
    .C(_11828_),
    .Y(_11836_));
 OR3x1_ASAP7_75t_R _28301_ (.A(_10825_),
    .B(_11789_),
    .C(_11836_),
    .Y(_11837_));
 XOR2x2_ASAP7_75t_R _28302_ (.A(_01683_),
    .B(_11837_),
    .Y(_11838_));
 AND2x2_ASAP7_75t_R _28303_ (.A(_05467_),
    .B(_11580_),
    .Y(_11839_));
 AO21x1_ASAP7_75t_R _28304_ (.A1(_11788_),
    .A2(_11838_),
    .B(_11839_),
    .Y(_03946_));
 BUFx6f_ASAP7_75t_R _28305_ (.A(_11804_),
    .Y(_11840_));
 OR3x2_ASAP7_75t_R _28306_ (.A(_00023_),
    .B(_07335_),
    .C(_11824_),
    .Y(_11841_));
 OR3x1_ASAP7_75t_R _28307_ (.A(_01682_),
    .B(_01683_),
    .C(_11841_),
    .Y(_11842_));
 OA21x2_ASAP7_75t_R _28308_ (.A1(_11840_),
    .A2(_11842_),
    .B(_11475_),
    .Y(_11843_));
 OA21x2_ASAP7_75t_R _28309_ (.A1(_01683_),
    .A2(_11841_),
    .B(_11594_),
    .Y(_11844_));
 OAI21x1_ASAP7_75t_R _28310_ (.A1(_11813_),
    .A2(_11844_),
    .B(_01682_),
    .Y(_11845_));
 OA21x2_ASAP7_75t_R _28311_ (.A1(_11590_),
    .A2(_11843_),
    .B(_11845_),
    .Y(_03947_));
 BUFx6f_ASAP7_75t_R _28312_ (.A(_10854_),
    .Y(_11846_));
 BUFx6f_ASAP7_75t_R _28313_ (.A(_11783_),
    .Y(_11847_));
 OR3x1_ASAP7_75t_R _28314_ (.A(_00265_),
    .B(_11846_),
    .C(_11847_),
    .Y(_11848_));
 OAI21x1_ASAP7_75t_R _28315_ (.A1(\cs_registers_i.pc_if_i[2] ),
    .A2(_11785_),
    .B(_11848_),
    .Y(_11849_));
 OAI21x1_ASAP7_75t_R _28316_ (.A1(_11541_),
    .A2(_11849_),
    .B(_05507_),
    .Y(_03948_));
 OR5x1_ASAP7_75t_R _28317_ (.A(_01682_),
    .B(_01683_),
    .C(_10854_),
    .D(_11783_),
    .E(_11836_),
    .Y(_11850_));
 XNOR2x2_ASAP7_75t_R _28318_ (.A(_01681_),
    .B(_11850_),
    .Y(_11851_));
 AOI21x1_ASAP7_75t_R _28319_ (.A1(_11788_),
    .A2(_11851_),
    .B(_11602_),
    .Y(_03949_));
 OR3x2_ASAP7_75t_R _28320_ (.A(_01681_),
    .B(_01682_),
    .C(_01683_),
    .Y(_11852_));
 OR2x6_ASAP7_75t_R _28321_ (.A(_11841_),
    .B(_11852_),
    .Y(_11853_));
 OR3x2_ASAP7_75t_R _28322_ (.A(_10854_),
    .B(_11783_),
    .C(_11853_),
    .Y(_11854_));
 XOR2x2_ASAP7_75t_R _28323_ (.A(_01680_),
    .B(_11854_),
    .Y(_11855_));
 AO21x1_ASAP7_75t_R _28324_ (.A1(_11803_),
    .A2(_11855_),
    .B(_11613_),
    .Y(_03950_));
 OR5x1_ASAP7_75t_R _28325_ (.A(_01680_),
    .B(_10854_),
    .C(_11789_),
    .D(_11836_),
    .E(_11852_),
    .Y(_11856_));
 XNOR2x2_ASAP7_75t_R _28326_ (.A(_01679_),
    .B(_11856_),
    .Y(_11857_));
 AOI21x1_ASAP7_75t_R _28327_ (.A1(_11788_),
    .A2(_11857_),
    .B(_11618_),
    .Y(_03951_));
 OR3x1_ASAP7_75t_R _28328_ (.A(_01679_),
    .B(_01680_),
    .C(_11853_),
    .Y(_11858_));
 AO21x1_ASAP7_75t_R _28329_ (.A1(_11628_),
    .A2(_11858_),
    .B(_11813_),
    .Y(_11859_));
 OR3x2_ASAP7_75t_R _28330_ (.A(_01678_),
    .B(_01679_),
    .C(_01680_),
    .Y(_11860_));
 OAI21x1_ASAP7_75t_R _28331_ (.A1(_11854_),
    .A2(_11860_),
    .B(_11803_),
    .Y(_11861_));
 AOI22x1_ASAP7_75t_R _28332_ (.A1(_01678_),
    .A2(_11859_),
    .B1(_11861_),
    .B2(_11628_),
    .Y(_03952_));
 OR5x1_ASAP7_75t_R _28333_ (.A(_10825_),
    .B(_11789_),
    .C(_11836_),
    .D(_11852_),
    .E(_11860_),
    .Y(_11862_));
 XNOR2x2_ASAP7_75t_R _28334_ (.A(_01677_),
    .B(_11862_),
    .Y(_11863_));
 AOI21x1_ASAP7_75t_R _28335_ (.A1(_11788_),
    .A2(_11863_),
    .B(_11637_),
    .Y(_03953_));
 INVx1_ASAP7_75t_R _28336_ (.A(_01676_),
    .Y(_11864_));
 BUFx12f_ASAP7_75t_R _28337_ (.A(_11784_),
    .Y(_11865_));
 OR3x1_ASAP7_75t_R _28338_ (.A(_01677_),
    .B(_11853_),
    .C(_11860_),
    .Y(_11866_));
 INVx1_ASAP7_75t_R _28339_ (.A(_11866_),
    .Y(_11867_));
 OA22x2_ASAP7_75t_R _28340_ (.A1(_05467_),
    .A2(_11865_),
    .B1(_11867_),
    .B2(_11646_),
    .Y(_11868_));
 OR3x2_ASAP7_75t_R _28341_ (.A(_01676_),
    .B(_01677_),
    .C(_11860_),
    .Y(_11869_));
 OA21x2_ASAP7_75t_R _28342_ (.A1(_11854_),
    .A2(_11869_),
    .B(_11475_),
    .Y(_11870_));
 OA22x2_ASAP7_75t_R _28343_ (.A1(_11864_),
    .A2(_11868_),
    .B1(_11870_),
    .B2(_11646_),
    .Y(_03954_));
 OR3x1_ASAP7_75t_R _28344_ (.A(_11836_),
    .B(_11852_),
    .C(_11869_),
    .Y(_11871_));
 OR3x1_ASAP7_75t_R _28345_ (.A(_10854_),
    .B(_11783_),
    .C(_11871_),
    .Y(_11872_));
 XOR2x2_ASAP7_75t_R _28346_ (.A(_01675_),
    .B(_11872_),
    .Y(_11873_));
 INVx1_ASAP7_75t_R _28347_ (.A(_11659_),
    .Y(_11874_));
 AO21x1_ASAP7_75t_R _28348_ (.A1(_11803_),
    .A2(_11873_),
    .B(_11874_),
    .Y(_03955_));
 OR5x1_ASAP7_75t_R _28349_ (.A(_01675_),
    .B(_10854_),
    .C(_11789_),
    .D(_11853_),
    .E(_11869_),
    .Y(_11875_));
 XNOR2x2_ASAP7_75t_R _28350_ (.A(_01674_),
    .B(_11875_),
    .Y(_11876_));
 AOI21x1_ASAP7_75t_R _28351_ (.A1(_11788_),
    .A2(_11876_),
    .B(_11666_),
    .Y(_03956_));
 OR3x1_ASAP7_75t_R _28352_ (.A(_01674_),
    .B(_01675_),
    .C(_11871_),
    .Y(_11877_));
 AO21x1_ASAP7_75t_R _28353_ (.A1(_11674_),
    .A2(_11877_),
    .B(_11813_),
    .Y(_11878_));
 OR3x2_ASAP7_75t_R _28354_ (.A(_01673_),
    .B(_01674_),
    .C(_01675_),
    .Y(_11879_));
 OAI21x1_ASAP7_75t_R _28355_ (.A1(_11872_),
    .A2(_11879_),
    .B(_11803_),
    .Y(_11880_));
 AOI22x1_ASAP7_75t_R _28356_ (.A1(_01673_),
    .A2(_11878_),
    .B1(_11880_),
    .B2(_11674_),
    .Y(_03957_));
 OR5x1_ASAP7_75t_R _28357_ (.A(_10854_),
    .B(_11783_),
    .C(_11853_),
    .D(_11869_),
    .E(_11879_),
    .Y(_11881_));
 XOR2x2_ASAP7_75t_R _28358_ (.A(_01672_),
    .B(_11881_),
    .Y(_11882_));
 OA21x2_ASAP7_75t_R _28359_ (.A1(_11541_),
    .A2(_11882_),
    .B(_11684_),
    .Y(_03958_));
 OR3x1_ASAP7_75t_R _28360_ (.A(_11790_),
    .B(_10825_),
    .C(_11789_),
    .Y(_11883_));
 XNOR2x2_ASAP7_75t_R _28361_ (.A(_00021_),
    .B(_11883_),
    .Y(_11884_));
 OAI21x1_ASAP7_75t_R _28362_ (.A1(_11541_),
    .A2(_11884_),
    .B(_05520_),
    .Y(_03959_));
 OR3x1_ASAP7_75t_R _28363_ (.A(_01672_),
    .B(_11871_),
    .C(_11879_),
    .Y(_11885_));
 NOR2x1_ASAP7_75t_R _28364_ (.A(_01671_),
    .B(_11885_),
    .Y(_11886_));
 AO21x1_ASAP7_75t_R _28365_ (.A1(_11819_),
    .A2(_11886_),
    .B(_05467_),
    .Y(_11887_));
 AO21x1_ASAP7_75t_R _28366_ (.A1(_11694_),
    .A2(_11885_),
    .B(_11813_),
    .Y(_11888_));
 AOI22x1_ASAP7_75t_R _28367_ (.A1(net1964),
    .A2(_11887_),
    .B1(_11888_),
    .B2(_01671_),
    .Y(_03960_));
 INVx1_ASAP7_75t_R _28368_ (.A(_11440_),
    .Y(_11889_));
 AO21x1_ASAP7_75t_R _28369_ (.A1(_11889_),
    .A2(_11799_),
    .B(_11813_),
    .Y(_11890_));
 OR4x1_ASAP7_75t_R _28370_ (.A(_01670_),
    .B(_11846_),
    .C(_11847_),
    .D(_11799_),
    .Y(_11891_));
 AOI21x1_ASAP7_75t_R _28371_ (.A1(_11803_),
    .A2(_11891_),
    .B(_11440_),
    .Y(_11892_));
 AOI21x1_ASAP7_75t_R _28372_ (.A1(_01670_),
    .A2(_11890_),
    .B(_11892_),
    .Y(_03961_));
 OR4x1_ASAP7_75t_R _28373_ (.A(_01670_),
    .B(_10825_),
    .C(_11789_),
    .D(_11791_),
    .Y(_11893_));
 XNOR2x2_ASAP7_75t_R _28374_ (.A(_01669_),
    .B(_11893_),
    .Y(_11894_));
 AOI21x1_ASAP7_75t_R _28375_ (.A1(_11788_),
    .A2(_11894_),
    .B(_11443_),
    .Y(_03962_));
 INVx1_ASAP7_75t_R _28376_ (.A(_11707_),
    .Y(_11895_));
 OR3x1_ASAP7_75t_R _28377_ (.A(_01669_),
    .B(_01670_),
    .C(_11799_),
    .Y(_11896_));
 AO21x1_ASAP7_75t_R _28378_ (.A1(_11895_),
    .A2(_11896_),
    .B(_11813_),
    .Y(_11897_));
 OR4x1_ASAP7_75t_R _28379_ (.A(_11846_),
    .B(_11847_),
    .C(_11792_),
    .D(_11799_),
    .Y(_11898_));
 AOI21x1_ASAP7_75t_R _28380_ (.A1(_11803_),
    .A2(_11898_),
    .B(_11707_),
    .Y(_11899_));
 AOI21x1_ASAP7_75t_R _28381_ (.A1(_01668_),
    .A2(_11897_),
    .B(_11899_),
    .Y(_03963_));
 OR4x1_ASAP7_75t_R _28382_ (.A(_10854_),
    .B(_11789_),
    .C(_11791_),
    .D(_11792_),
    .Y(_11900_));
 XNOR2x2_ASAP7_75t_R _28383_ (.A(_01667_),
    .B(_11900_),
    .Y(_11901_));
 AOI22x1_ASAP7_75t_R _28384_ (.A1(_11433_),
    .A2(_11434_),
    .B1(_11901_),
    .B2(_11788_),
    .Y(_03964_));
 OR3x1_ASAP7_75t_R _28385_ (.A(_01667_),
    .B(_11792_),
    .C(_11799_),
    .Y(_11902_));
 AO21x1_ASAP7_75t_R _28386_ (.A1(_11715_),
    .A2(_11902_),
    .B(_11813_),
    .Y(_11903_));
 OR4x1_ASAP7_75t_R _28387_ (.A(_10825_),
    .B(_11847_),
    .C(_11793_),
    .D(_11799_),
    .Y(_11904_));
 NAND2x1_ASAP7_75t_R _28388_ (.A(_11475_),
    .B(_11904_),
    .Y(_11905_));
 AOI22x1_ASAP7_75t_R _28389_ (.A1(_01666_),
    .A2(_11903_),
    .B1(_11905_),
    .B2(_11715_),
    .Y(_03965_));
 OR4x1_ASAP7_75t_R _28390_ (.A(_10825_),
    .B(_11789_),
    .C(_11791_),
    .D(_11793_),
    .Y(_11906_));
 XNOR2x2_ASAP7_75t_R _28391_ (.A(_01665_),
    .B(_11906_),
    .Y(_11907_));
 AOI21x1_ASAP7_75t_R _28392_ (.A1(_11788_),
    .A2(_11907_),
    .B(_11458_),
    .Y(_03966_));
 OR5x1_ASAP7_75t_R _28393_ (.A(_01665_),
    .B(_10854_),
    .C(_11783_),
    .D(_11793_),
    .E(_11799_),
    .Y(_11908_));
 XOR2x2_ASAP7_75t_R _28394_ (.A(_00022_),
    .B(_11908_),
    .Y(_11909_));
 OA21x2_ASAP7_75t_R _28395_ (.A1(_11541_),
    .A2(_11909_),
    .B(_11469_),
    .Y(_03967_));
 OR2x2_ASAP7_75t_R _28396_ (.A(net117),
    .B(_05711_),
    .Y(_11910_));
 NAND2x1_ASAP7_75t_R _28397_ (.A(_05712_),
    .B(_01639_),
    .Y(_11911_));
 NOR2x1_ASAP7_75t_R _28398_ (.A(_01664_),
    .B(_11756_),
    .Y(_11912_));
 AO32x1_ASAP7_75t_R _28399_ (.A1(_11752_),
    .A2(_11910_),
    .A3(_11911_),
    .B1(_11912_),
    .B2(_11759_),
    .Y(_03968_));
 OR2x2_ASAP7_75t_R _28400_ (.A(net118),
    .B(_05711_),
    .Y(_11913_));
 NAND2x1_ASAP7_75t_R _28401_ (.A(_05712_),
    .B(_01628_),
    .Y(_11914_));
 NOR2x1_ASAP7_75t_R _28402_ (.A(_01663_),
    .B(_11756_),
    .Y(_11915_));
 AO32x1_ASAP7_75t_R _28403_ (.A1(_11752_),
    .A2(_11913_),
    .A3(_11914_),
    .B1(_11915_),
    .B2(_11759_),
    .Y(_03969_));
 OR2x2_ASAP7_75t_R _28404_ (.A(net119),
    .B(_05712_),
    .Y(_11916_));
 NAND2x1_ASAP7_75t_R _28405_ (.A(_05712_),
    .B(_01627_),
    .Y(_11917_));
 NOR2x1_ASAP7_75t_R _28406_ (.A(_01662_),
    .B(_11756_),
    .Y(_11918_));
 AO32x1_ASAP7_75t_R _28407_ (.A1(_11752_),
    .A2(_11916_),
    .A3(_11917_),
    .B1(_11918_),
    .B2(_11759_),
    .Y(_03970_));
 OR2x2_ASAP7_75t_R _28408_ (.A(net120),
    .B(_05712_),
    .Y(_11919_));
 NAND2x1_ASAP7_75t_R _28409_ (.A(_11722_),
    .B(_01626_),
    .Y(_11920_));
 NOR2x1_ASAP7_75t_R _28410_ (.A(_01661_),
    .B(_11756_),
    .Y(_11921_));
 AO32x1_ASAP7_75t_R _28411_ (.A1(_11752_),
    .A2(_11919_),
    .A3(_11920_),
    .B1(_11921_),
    .B2(_11759_),
    .Y(_03971_));
 OR2x2_ASAP7_75t_R _28412_ (.A(net121),
    .B(_05711_),
    .Y(_11922_));
 NAND2x1_ASAP7_75t_R _28413_ (.A(_05712_),
    .B(_01625_),
    .Y(_11923_));
 NOR2x1_ASAP7_75t_R _28414_ (.A(_01660_),
    .B(_11756_),
    .Y(_11924_));
 AO32x1_ASAP7_75t_R _28415_ (.A1(_11752_),
    .A2(_11922_),
    .A3(_11923_),
    .B1(_11924_),
    .B2(_11759_),
    .Y(_03972_));
 NOR2x1_ASAP7_75t_R _28416_ (.A(_01659_),
    .B(_11756_),
    .Y(_11925_));
 NAND2x1_ASAP7_75t_R _28417_ (.A(_11722_),
    .B(_01624_),
    .Y(_11926_));
 OAI21x1_ASAP7_75t_R _28418_ (.A1(net122),
    .A2(_11723_),
    .B(_11926_),
    .Y(_11927_));
 INVx1_ASAP7_75t_R _28419_ (.A(_11927_),
    .Y(_11928_));
 AO22x1_ASAP7_75t_R _28420_ (.A1(_11759_),
    .A2(_11925_),
    .B1(_11928_),
    .B2(_11752_),
    .Y(_03973_));
 BUFx6f_ASAP7_75t_R _28421_ (.A(_11751_),
    .Y(_11929_));
 OR2x2_ASAP7_75t_R _28422_ (.A(net123),
    .B(_11723_),
    .Y(_11930_));
 NAND2x1_ASAP7_75t_R _28423_ (.A(_11723_),
    .B(_01623_),
    .Y(_11931_));
 BUFx12f_ASAP7_75t_R _28424_ (.A(_11750_),
    .Y(_11932_));
 NOR2x1_ASAP7_75t_R _28425_ (.A(_01658_),
    .B(_11932_),
    .Y(_11933_));
 BUFx6f_ASAP7_75t_R _28426_ (.A(_11758_),
    .Y(_11934_));
 AO32x1_ASAP7_75t_R _28427_ (.A1(_11929_),
    .A2(_11930_),
    .A3(_11931_),
    .B1(_11933_),
    .B2(_11934_),
    .Y(_03974_));
 BUFx6f_ASAP7_75t_R _28428_ (.A(_11724_),
    .Y(_11935_));
 OR2x2_ASAP7_75t_R _28429_ (.A(net124),
    .B(_11935_),
    .Y(_11936_));
 NAND2x1_ASAP7_75t_R _28430_ (.A(_11754_),
    .B(_01622_),
    .Y(_11937_));
 NOR2x1_ASAP7_75t_R _28431_ (.A(_01657_),
    .B(_11932_),
    .Y(_11938_));
 AO32x1_ASAP7_75t_R _28432_ (.A1(_11929_),
    .A2(_11936_),
    .A3(_11937_),
    .B1(_11938_),
    .B2(_11934_),
    .Y(_03975_));
 OR2x2_ASAP7_75t_R _28433_ (.A(net125),
    .B(_11935_),
    .Y(_11939_));
 NAND2x1_ASAP7_75t_R _28434_ (.A(_11754_),
    .B(_01621_),
    .Y(_11940_));
 NOR2x1_ASAP7_75t_R _28435_ (.A(_01656_),
    .B(_11932_),
    .Y(_11941_));
 AO32x1_ASAP7_75t_R _28436_ (.A1(_11929_),
    .A2(_11939_),
    .A3(_11940_),
    .B1(_11941_),
    .B2(_11934_),
    .Y(_03976_));
 BUFx6f_ASAP7_75t_R _28437_ (.A(_11724_),
    .Y(_11942_));
 OR2x2_ASAP7_75t_R _28438_ (.A(net126),
    .B(_11942_),
    .Y(_11943_));
 NAND2x1_ASAP7_75t_R _28439_ (.A(_11754_),
    .B(_01619_),
    .Y(_11944_));
 NOR2x1_ASAP7_75t_R _28440_ (.A(_01655_),
    .B(_11932_),
    .Y(_11945_));
 AO32x1_ASAP7_75t_R _28441_ (.A1(_11929_),
    .A2(_11943_),
    .A3(_11944_),
    .B1(_11945_),
    .B2(_11934_),
    .Y(_03977_));
 OR2x2_ASAP7_75t_R _28442_ (.A(net127),
    .B(_11942_),
    .Y(_11946_));
 NAND2x1_ASAP7_75t_R _28443_ (.A(_11754_),
    .B(_01618_),
    .Y(_11947_));
 NOR2x1_ASAP7_75t_R _28444_ (.A(_01654_),
    .B(_11932_),
    .Y(_11948_));
 AO32x1_ASAP7_75t_R _28445_ (.A1(_11929_),
    .A2(_11946_),
    .A3(_11947_),
    .B1(_11948_),
    .B2(_11934_),
    .Y(_03978_));
 OR2x2_ASAP7_75t_R _28446_ (.A(net128),
    .B(_11722_),
    .Y(_11949_));
 NAND2x1_ASAP7_75t_R _28447_ (.A(_11722_),
    .B(_01638_),
    .Y(_11950_));
 NOR2x1_ASAP7_75t_R _28448_ (.A(_01653_),
    .B(_11932_),
    .Y(_11951_));
 AO32x1_ASAP7_75t_R _28449_ (.A1(_11929_),
    .A2(_11949_),
    .A3(_11950_),
    .B1(_11951_),
    .B2(_11934_),
    .Y(_03979_));
 OR2x2_ASAP7_75t_R _28450_ (.A(net129),
    .B(_11942_),
    .Y(_11952_));
 NAND2x1_ASAP7_75t_R _28451_ (.A(_11754_),
    .B(_01617_),
    .Y(_11953_));
 NOR2x1_ASAP7_75t_R _28452_ (.A(_01652_),
    .B(_11932_),
    .Y(_11954_));
 AO32x1_ASAP7_75t_R _28453_ (.A1(_11929_),
    .A2(_11952_),
    .A3(_11953_),
    .B1(_11954_),
    .B2(_11934_),
    .Y(_03980_));
 OR2x2_ASAP7_75t_R _28454_ (.A(net130),
    .B(_11942_),
    .Y(_11955_));
 NAND2x1_ASAP7_75t_R _28455_ (.A(_11754_),
    .B(_01616_),
    .Y(_11956_));
 NOR2x1_ASAP7_75t_R _28456_ (.A(_01651_),
    .B(_11932_),
    .Y(_11957_));
 AO32x1_ASAP7_75t_R _28457_ (.A1(_11929_),
    .A2(_11955_),
    .A3(_11956_),
    .B1(_11957_),
    .B2(_11934_),
    .Y(_03981_));
 OR2x2_ASAP7_75t_R _28458_ (.A(net131),
    .B(_11942_),
    .Y(_11958_));
 NAND2x1_ASAP7_75t_R _28459_ (.A(_11754_),
    .B(_01615_),
    .Y(_11959_));
 NOR2x1_ASAP7_75t_R _28460_ (.A(_01650_),
    .B(_11932_),
    .Y(_11960_));
 AO32x1_ASAP7_75t_R _28461_ (.A1(_11929_),
    .A2(_11958_),
    .A3(_11959_),
    .B1(_11960_),
    .B2(_11934_),
    .Y(_03982_));
 OR2x2_ASAP7_75t_R _28462_ (.A(net132),
    .B(_11942_),
    .Y(_11961_));
 NAND2x1_ASAP7_75t_R _28463_ (.A(_11754_),
    .B(_01614_),
    .Y(_11962_));
 NOR2x1_ASAP7_75t_R _28464_ (.A(_01649_),
    .B(_11932_),
    .Y(_11963_));
 AO32x1_ASAP7_75t_R _28465_ (.A1(_11929_),
    .A2(_11961_),
    .A3(_11962_),
    .B1(_11963_),
    .B2(_11934_),
    .Y(_03983_));
 BUFx6f_ASAP7_75t_R _28466_ (.A(_11751_),
    .Y(_11964_));
 OR2x2_ASAP7_75t_R _28467_ (.A(net133),
    .B(_11942_),
    .Y(_11965_));
 NAND2x1_ASAP7_75t_R _28468_ (.A(_11754_),
    .B(_01613_),
    .Y(_11966_));
 BUFx12f_ASAP7_75t_R _28469_ (.A(_11750_),
    .Y(_11967_));
 NOR2x1_ASAP7_75t_R _28470_ (.A(_01648_),
    .B(_11967_),
    .Y(_11968_));
 BUFx3_ASAP7_75t_R _28471_ (.A(_11758_),
    .Y(_11969_));
 AO32x1_ASAP7_75t_R _28472_ (.A1(_11964_),
    .A2(_11965_),
    .A3(_11966_),
    .B1(_11968_),
    .B2(_11969_),
    .Y(_03984_));
 OR2x2_ASAP7_75t_R _28473_ (.A(net134),
    .B(_11942_),
    .Y(_11970_));
 NAND2x1_ASAP7_75t_R _28474_ (.A(_11935_),
    .B(_01612_),
    .Y(_11971_));
 NOR2x1_ASAP7_75t_R _28475_ (.A(_01647_),
    .B(_11967_),
    .Y(_11972_));
 AO32x1_ASAP7_75t_R _28476_ (.A1(_11964_),
    .A2(_11970_),
    .A3(_11971_),
    .B1(_11972_),
    .B2(_11969_),
    .Y(_03985_));
 OR2x2_ASAP7_75t_R _28477_ (.A(net135),
    .B(_11942_),
    .Y(_11973_));
 NAND2x1_ASAP7_75t_R _28478_ (.A(_11935_),
    .B(_01611_),
    .Y(_11974_));
 NOR2x1_ASAP7_75t_R _28479_ (.A(_01646_),
    .B(_11967_),
    .Y(_11975_));
 AO32x1_ASAP7_75t_R _28480_ (.A1(_11964_),
    .A2(_11973_),
    .A3(_11974_),
    .B1(_11975_),
    .B2(_11969_),
    .Y(_03986_));
 OR2x2_ASAP7_75t_R _28481_ (.A(net136),
    .B(_11942_),
    .Y(_11976_));
 NAND2x1_ASAP7_75t_R _28482_ (.A(_11935_),
    .B(_01610_),
    .Y(_11977_));
 NOR2x1_ASAP7_75t_R _28483_ (.A(_01645_),
    .B(_11967_),
    .Y(_11978_));
 AO32x1_ASAP7_75t_R _28484_ (.A1(_11964_),
    .A2(_11976_),
    .A3(_11977_),
    .B1(_11978_),
    .B2(_11969_),
    .Y(_03987_));
 OR2x2_ASAP7_75t_R _28485_ (.A(net137),
    .B(_11724_),
    .Y(_11979_));
 NAND2x1_ASAP7_75t_R _28486_ (.A(_11935_),
    .B(_01608_),
    .Y(_11980_));
 NOR2x1_ASAP7_75t_R _28487_ (.A(_01644_),
    .B(_11967_),
    .Y(_11981_));
 AO32x1_ASAP7_75t_R _28488_ (.A1(_11964_),
    .A2(_11979_),
    .A3(_11980_),
    .B1(_11981_),
    .B2(_11969_),
    .Y(_03988_));
 OR2x2_ASAP7_75t_R _28489_ (.A(net138),
    .B(_11724_),
    .Y(_11982_));
 NAND2x1_ASAP7_75t_R _28490_ (.A(_11935_),
    .B(_01607_),
    .Y(_11983_));
 NOR2x1_ASAP7_75t_R _28491_ (.A(_01643_),
    .B(_11967_),
    .Y(_11984_));
 AO32x1_ASAP7_75t_R _28492_ (.A1(_11964_),
    .A2(_11982_),
    .A3(_11983_),
    .B1(_11984_),
    .B2(_11969_),
    .Y(_03989_));
 OR2x2_ASAP7_75t_R _28493_ (.A(net139),
    .B(_05712_),
    .Y(_11985_));
 NAND2x1_ASAP7_75t_R _28494_ (.A(_11722_),
    .B(_01637_),
    .Y(_11986_));
 NOR2x1_ASAP7_75t_R _28495_ (.A(_01642_),
    .B(_11967_),
    .Y(_11987_));
 AO32x1_ASAP7_75t_R _28496_ (.A1(_11964_),
    .A2(_11985_),
    .A3(_11986_),
    .B1(_11987_),
    .B2(_11969_),
    .Y(_03990_));
 OR2x2_ASAP7_75t_R _28497_ (.A(net140),
    .B(_11724_),
    .Y(_11988_));
 NAND2x1_ASAP7_75t_R _28498_ (.A(_11935_),
    .B(_01606_),
    .Y(_11989_));
 NOR2x1_ASAP7_75t_R _28499_ (.A(_01641_),
    .B(_11967_),
    .Y(_11990_));
 AO32x1_ASAP7_75t_R _28500_ (.A1(_11964_),
    .A2(_11988_),
    .A3(_11989_),
    .B1(_11990_),
    .B2(_11969_),
    .Y(_03991_));
 OR2x2_ASAP7_75t_R _28501_ (.A(net141),
    .B(_11724_),
    .Y(_11991_));
 NAND2x1_ASAP7_75t_R _28502_ (.A(_11935_),
    .B(_01605_),
    .Y(_11992_));
 NOR2x1_ASAP7_75t_R _28503_ (.A(_01640_),
    .B(_11967_),
    .Y(_11993_));
 AO32x1_ASAP7_75t_R _28504_ (.A1(_11964_),
    .A2(_11991_),
    .A3(_11992_),
    .B1(_11993_),
    .B2(_11969_),
    .Y(_03992_));
 NAND2x1_ASAP7_75t_R _28505_ (.A(_01604_),
    .B(_11767_),
    .Y(_11994_));
 OA21x2_ASAP7_75t_R _28506_ (.A1(net117),
    .A2(_11766_),
    .B(_11994_),
    .Y(_11995_));
 BUFx12f_ASAP7_75t_R _28507_ (.A(_11774_),
    .Y(_11996_));
 NOR2x1_ASAP7_75t_R _28508_ (.A(_01639_),
    .B(_11996_),
    .Y(_11997_));
 AO22x1_ASAP7_75t_R _28509_ (.A1(_11764_),
    .A2(_11995_),
    .B1(_11997_),
    .B2(_11772_),
    .Y(_03993_));
 NAND2x1_ASAP7_75t_R _28510_ (.A(_01603_),
    .B(_11767_),
    .Y(_11998_));
 OA21x2_ASAP7_75t_R _28511_ (.A1(net128),
    .A2(_11766_),
    .B(_11998_),
    .Y(_11999_));
 NOR2x1_ASAP7_75t_R _28512_ (.A(_01638_),
    .B(_11996_),
    .Y(_12000_));
 AO22x1_ASAP7_75t_R _28513_ (.A1(_11764_),
    .A2(_11999_),
    .B1(_12000_),
    .B2(_11772_),
    .Y(_03994_));
 NAND2x1_ASAP7_75t_R _28514_ (.A(_01602_),
    .B(_11767_),
    .Y(_12001_));
 OA21x2_ASAP7_75t_R _28515_ (.A1(net139),
    .A2(_11766_),
    .B(_12001_),
    .Y(_12002_));
 NOR2x1_ASAP7_75t_R _28516_ (.A(_01637_),
    .B(_11996_),
    .Y(_12003_));
 AO22x1_ASAP7_75t_R _28517_ (.A1(_11764_),
    .A2(_12002_),
    .B1(_12003_),
    .B2(_11772_),
    .Y(_03995_));
 NAND2x1_ASAP7_75t_R _28518_ (.A(_01601_),
    .B(_11767_),
    .Y(_12004_));
 OA21x2_ASAP7_75t_R _28519_ (.A1(net142),
    .A2(_11766_),
    .B(_12004_),
    .Y(_12005_));
 NOR2x1_ASAP7_75t_R _28520_ (.A(_01636_),
    .B(_11996_),
    .Y(_12006_));
 AO22x1_ASAP7_75t_R _28521_ (.A1(_11764_),
    .A2(_12005_),
    .B1(_12006_),
    .B2(_11772_),
    .Y(_03996_));
 NAND2x1_ASAP7_75t_R _28522_ (.A(_01600_),
    .B(_11767_),
    .Y(_12007_));
 OA21x2_ASAP7_75t_R _28523_ (.A1(net143),
    .A2(_11766_),
    .B(_12007_),
    .Y(_12008_));
 NOR2x1_ASAP7_75t_R _28524_ (.A(_01635_),
    .B(_11996_),
    .Y(_12009_));
 AO22x1_ASAP7_75t_R _28525_ (.A1(_11764_),
    .A2(_12008_),
    .B1(_12009_),
    .B2(_11772_),
    .Y(_03997_));
 NAND2x1_ASAP7_75t_R _28526_ (.A(_01599_),
    .B(_11767_),
    .Y(_12010_));
 OA21x2_ASAP7_75t_R _28527_ (.A1(net144),
    .A2(_11766_),
    .B(_12010_),
    .Y(_12011_));
 NOR2x1_ASAP7_75t_R _28528_ (.A(_01634_),
    .B(_11996_),
    .Y(_12012_));
 AO22x1_ASAP7_75t_R _28529_ (.A1(_11764_),
    .A2(_12011_),
    .B1(_12012_),
    .B2(_11772_),
    .Y(_03998_));
 BUFx12f_ASAP7_75t_R _28530_ (.A(_11765_),
    .Y(_12013_));
 NAND2x1_ASAP7_75t_R _28531_ (.A(_01597_),
    .B(_12013_),
    .Y(_12014_));
 OA21x2_ASAP7_75t_R _28532_ (.A1(net145),
    .A2(_11766_),
    .B(_12014_),
    .Y(_12015_));
 NOR2x1_ASAP7_75t_R _28533_ (.A(_01633_),
    .B(_11996_),
    .Y(_12016_));
 AO22x1_ASAP7_75t_R _28534_ (.A1(_11764_),
    .A2(_12015_),
    .B1(_12016_),
    .B2(_11772_),
    .Y(_03999_));
 NAND2x1_ASAP7_75t_R _28535_ (.A(_01596_),
    .B(_12013_),
    .Y(_12017_));
 OA21x2_ASAP7_75t_R _28536_ (.A1(net146),
    .A2(_11766_),
    .B(_12017_),
    .Y(_12018_));
 NOR2x1_ASAP7_75t_R _28537_ (.A(_01632_),
    .B(_11996_),
    .Y(_12019_));
 AO22x1_ASAP7_75t_R _28538_ (.A1(_11764_),
    .A2(_12018_),
    .B1(_12019_),
    .B2(_11772_),
    .Y(_04000_));
 OR2x2_ASAP7_75t_R _28539_ (.A(net142),
    .B(_11722_),
    .Y(_12020_));
 NAND2x1_ASAP7_75t_R _28540_ (.A(_11723_),
    .B(_01636_),
    .Y(_12021_));
 NOR2x1_ASAP7_75t_R _28541_ (.A(_01631_),
    .B(_11967_),
    .Y(_12022_));
 AO32x1_ASAP7_75t_R _28542_ (.A1(_11964_),
    .A2(_12020_),
    .A3(_12021_),
    .B1(_12022_),
    .B2(_11969_),
    .Y(_04001_));
 NAND2x1_ASAP7_75t_R _28543_ (.A(_01595_),
    .B(_12013_),
    .Y(_12023_));
 OA21x2_ASAP7_75t_R _28544_ (.A1(net147),
    .A2(_11766_),
    .B(_12023_),
    .Y(_12024_));
 NOR2x1_ASAP7_75t_R _28545_ (.A(_01630_),
    .B(_11996_),
    .Y(_12025_));
 AO22x1_ASAP7_75t_R _28546_ (.A1(_11764_),
    .A2(_12024_),
    .B1(_12025_),
    .B2(_11772_),
    .Y(_04002_));
 BUFx3_ASAP7_75t_R _28547_ (.A(_11763_),
    .Y(_12026_));
 BUFx6f_ASAP7_75t_R _28548_ (.A(_11765_),
    .Y(_12027_));
 NAND2x1_ASAP7_75t_R _28549_ (.A(_01594_),
    .B(_12013_),
    .Y(_12028_));
 OA21x2_ASAP7_75t_R _28550_ (.A1(net148),
    .A2(_12027_),
    .B(_12028_),
    .Y(_12029_));
 NOR2x1_ASAP7_75t_R _28551_ (.A(_01629_),
    .B(_11996_),
    .Y(_12030_));
 BUFx3_ASAP7_75t_R _28552_ (.A(_11771_),
    .Y(_12031_));
 AO22x1_ASAP7_75t_R _28553_ (.A1(_12026_),
    .A2(_12029_),
    .B1(_12030_),
    .B2(_12031_),
    .Y(_04003_));
 NAND2x1_ASAP7_75t_R _28554_ (.A(_01593_),
    .B(_12013_),
    .Y(_12032_));
 OA21x2_ASAP7_75t_R _28555_ (.A1(net118),
    .A2(_12027_),
    .B(_12032_),
    .Y(_12033_));
 BUFx12f_ASAP7_75t_R _28556_ (.A(_11774_),
    .Y(_12034_));
 NOR2x1_ASAP7_75t_R _28557_ (.A(_01628_),
    .B(_12034_),
    .Y(_12035_));
 AO22x1_ASAP7_75t_R _28558_ (.A1(_12026_),
    .A2(_12033_),
    .B1(_12035_),
    .B2(_12031_),
    .Y(_04004_));
 NAND2x1_ASAP7_75t_R _28559_ (.A(_01592_),
    .B(_12013_),
    .Y(_12036_));
 OA21x2_ASAP7_75t_R _28560_ (.A1(net119),
    .A2(_12027_),
    .B(_12036_),
    .Y(_12037_));
 NOR2x1_ASAP7_75t_R _28561_ (.A(_01627_),
    .B(_12034_),
    .Y(_12038_));
 AO22x1_ASAP7_75t_R _28562_ (.A1(_12026_),
    .A2(_12037_),
    .B1(_12038_),
    .B2(_12031_),
    .Y(_04005_));
 NAND2x1_ASAP7_75t_R _28563_ (.A(_01591_),
    .B(_12013_),
    .Y(_12039_));
 OA21x2_ASAP7_75t_R _28564_ (.A1(net120),
    .A2(_12027_),
    .B(_12039_),
    .Y(_12040_));
 NOR2x1_ASAP7_75t_R _28565_ (.A(_01626_),
    .B(_12034_),
    .Y(_12041_));
 AO22x1_ASAP7_75t_R _28566_ (.A1(_12026_),
    .A2(_12040_),
    .B1(_12041_),
    .B2(_12031_),
    .Y(_04006_));
 NAND2x1_ASAP7_75t_R _28567_ (.A(_01590_),
    .B(_12013_),
    .Y(_12042_));
 OA21x2_ASAP7_75t_R _28568_ (.A1(net121),
    .A2(_12027_),
    .B(_12042_),
    .Y(_12043_));
 NOR2x1_ASAP7_75t_R _28569_ (.A(_01625_),
    .B(_12034_),
    .Y(_12044_));
 AO22x1_ASAP7_75t_R _28570_ (.A1(_12026_),
    .A2(_12043_),
    .B1(_12044_),
    .B2(_12031_),
    .Y(_04007_));
 NAND2x1_ASAP7_75t_R _28571_ (.A(_01589_),
    .B(_12013_),
    .Y(_12045_));
 OA21x2_ASAP7_75t_R _28572_ (.A1(net122),
    .A2(_12027_),
    .B(_12045_),
    .Y(_12046_));
 NOR2x1_ASAP7_75t_R _28573_ (.A(_01624_),
    .B(_12034_),
    .Y(_12047_));
 AO22x1_ASAP7_75t_R _28574_ (.A1(_12026_),
    .A2(_12046_),
    .B1(_12047_),
    .B2(_12031_),
    .Y(_04008_));
 NAND2x1_ASAP7_75t_R _28575_ (.A(_01588_),
    .B(_12013_),
    .Y(_12048_));
 OA21x2_ASAP7_75t_R _28576_ (.A1(net123),
    .A2(_12027_),
    .B(_12048_),
    .Y(_12049_));
 NOR2x1_ASAP7_75t_R _28577_ (.A(_01623_),
    .B(_12034_),
    .Y(_12050_));
 AO22x1_ASAP7_75t_R _28578_ (.A1(_12026_),
    .A2(_12049_),
    .B1(_12050_),
    .B2(_12031_),
    .Y(_04009_));
 BUFx12f_ASAP7_75t_R _28579_ (.A(_05708_),
    .Y(_12051_));
 NAND2x1_ASAP7_75t_R _28580_ (.A(_01586_),
    .B(_12051_),
    .Y(_12052_));
 OA21x2_ASAP7_75t_R _28581_ (.A1(net124),
    .A2(_12027_),
    .B(_12052_),
    .Y(_12053_));
 NOR2x1_ASAP7_75t_R _28582_ (.A(_01622_),
    .B(_12034_),
    .Y(_12054_));
 AO22x1_ASAP7_75t_R _28583_ (.A1(_12026_),
    .A2(_12053_),
    .B1(_12054_),
    .B2(_12031_),
    .Y(_04010_));
 NAND2x1_ASAP7_75t_R _28584_ (.A(_01585_),
    .B(_12051_),
    .Y(_12055_));
 OA21x2_ASAP7_75t_R _28585_ (.A1(net125),
    .A2(_12027_),
    .B(_12055_),
    .Y(_12056_));
 NOR2x1_ASAP7_75t_R _28586_ (.A(_01621_),
    .B(_12034_),
    .Y(_12057_));
 AO22x1_ASAP7_75t_R _28587_ (.A1(_12026_),
    .A2(_12056_),
    .B1(_12057_),
    .B2(_12031_),
    .Y(_04011_));
 OR2x2_ASAP7_75t_R _28588_ (.A(net143),
    .B(_05712_),
    .Y(_12058_));
 NAND2x1_ASAP7_75t_R _28589_ (.A(_11722_),
    .B(_01635_),
    .Y(_12059_));
 NOR2x1_ASAP7_75t_R _28590_ (.A(_01620_),
    .B(_11750_),
    .Y(_12060_));
 AO32x1_ASAP7_75t_R _28591_ (.A1(_11751_),
    .A2(_12058_),
    .A3(_12059_),
    .B1(_12060_),
    .B2(_11758_),
    .Y(_04012_));
 NAND2x1_ASAP7_75t_R _28592_ (.A(_01584_),
    .B(_12051_),
    .Y(_12061_));
 OA21x2_ASAP7_75t_R _28593_ (.A1(net126),
    .A2(_12027_),
    .B(_12061_),
    .Y(_12062_));
 NOR2x1_ASAP7_75t_R _28594_ (.A(_01619_),
    .B(_12034_),
    .Y(_12063_));
 AO22x1_ASAP7_75t_R _28595_ (.A1(_12026_),
    .A2(_12062_),
    .B1(_12063_),
    .B2(_12031_),
    .Y(_04013_));
 BUFx3_ASAP7_75t_R _28596_ (.A(_11763_),
    .Y(_12064_));
 BUFx6f_ASAP7_75t_R _28597_ (.A(_11765_),
    .Y(_12065_));
 NAND2x1_ASAP7_75t_R _28598_ (.A(_01583_),
    .B(_12051_),
    .Y(_12066_));
 OA21x2_ASAP7_75t_R _28599_ (.A1(net127),
    .A2(_12065_),
    .B(_12066_),
    .Y(_12067_));
 NOR2x1_ASAP7_75t_R _28600_ (.A(_01618_),
    .B(_12034_),
    .Y(_12068_));
 BUFx3_ASAP7_75t_R _28601_ (.A(_11771_),
    .Y(_12069_));
 AO22x1_ASAP7_75t_R _28602_ (.A1(_12064_),
    .A2(_12067_),
    .B1(_12068_),
    .B2(_12069_),
    .Y(_04014_));
 NAND2x1_ASAP7_75t_R _28603_ (.A(_01582_),
    .B(_12051_),
    .Y(_12070_));
 OA21x2_ASAP7_75t_R _28604_ (.A1(net129),
    .A2(_12065_),
    .B(_12070_),
    .Y(_12071_));
 BUFx12f_ASAP7_75t_R _28605_ (.A(_11774_),
    .Y(_12072_));
 NOR2x1_ASAP7_75t_R _28606_ (.A(_01617_),
    .B(_12072_),
    .Y(_12073_));
 AO22x1_ASAP7_75t_R _28607_ (.A1(_12064_),
    .A2(_12071_),
    .B1(_12073_),
    .B2(_12069_),
    .Y(_04015_));
 NAND2x1_ASAP7_75t_R _28608_ (.A(_01581_),
    .B(_12051_),
    .Y(_12074_));
 OA21x2_ASAP7_75t_R _28609_ (.A1(net130),
    .A2(_12065_),
    .B(_12074_),
    .Y(_12075_));
 NOR2x1_ASAP7_75t_R _28610_ (.A(_01616_),
    .B(_12072_),
    .Y(_12076_));
 AO22x1_ASAP7_75t_R _28611_ (.A1(_12064_),
    .A2(_12075_),
    .B1(_12076_),
    .B2(_12069_),
    .Y(_04016_));
 NAND2x1_ASAP7_75t_R _28612_ (.A(_01580_),
    .B(_12051_),
    .Y(_12077_));
 OA21x2_ASAP7_75t_R _28613_ (.A1(net131),
    .A2(_12065_),
    .B(_12077_),
    .Y(_12078_));
 NOR2x1_ASAP7_75t_R _28614_ (.A(_01615_),
    .B(_12072_),
    .Y(_12079_));
 AO22x1_ASAP7_75t_R _28615_ (.A1(_12064_),
    .A2(_12078_),
    .B1(_12079_),
    .B2(_12069_),
    .Y(_04017_));
 NAND2x1_ASAP7_75t_R _28616_ (.A(_01579_),
    .B(_12051_),
    .Y(_12080_));
 OA21x2_ASAP7_75t_R _28617_ (.A1(net132),
    .A2(_12065_),
    .B(_12080_),
    .Y(_12081_));
 NOR2x1_ASAP7_75t_R _28618_ (.A(_01614_),
    .B(_12072_),
    .Y(_12082_));
 AO22x1_ASAP7_75t_R _28619_ (.A1(_12064_),
    .A2(_12081_),
    .B1(_12082_),
    .B2(_12069_),
    .Y(_04018_));
 NAND2x1_ASAP7_75t_R _28620_ (.A(_01578_),
    .B(_12051_),
    .Y(_12083_));
 OA21x2_ASAP7_75t_R _28621_ (.A1(net133),
    .A2(_12065_),
    .B(_12083_),
    .Y(_12084_));
 NOR2x1_ASAP7_75t_R _28622_ (.A(_01613_),
    .B(_12072_),
    .Y(_12085_));
 AO22x1_ASAP7_75t_R _28623_ (.A1(_12064_),
    .A2(_12084_),
    .B1(_12085_),
    .B2(_12069_),
    .Y(_04019_));
 NAND2x1_ASAP7_75t_R _28624_ (.A(_01577_),
    .B(_12051_),
    .Y(_12086_));
 OA21x2_ASAP7_75t_R _28625_ (.A1(net134),
    .A2(_12065_),
    .B(_12086_),
    .Y(_12087_));
 NOR2x1_ASAP7_75t_R _28626_ (.A(_01612_),
    .B(_12072_),
    .Y(_12088_));
 AO22x1_ASAP7_75t_R _28627_ (.A1(_12064_),
    .A2(_12087_),
    .B1(_12088_),
    .B2(_12069_),
    .Y(_04020_));
 NAND2x1_ASAP7_75t_R _28628_ (.A(_01575_),
    .B(_11765_),
    .Y(_12089_));
 OA21x2_ASAP7_75t_R _28629_ (.A1(net135),
    .A2(_12065_),
    .B(_12089_),
    .Y(_12090_));
 NOR2x1_ASAP7_75t_R _28630_ (.A(_01611_),
    .B(_12072_),
    .Y(_12091_));
 AO22x1_ASAP7_75t_R _28631_ (.A1(_12064_),
    .A2(_12090_),
    .B1(_12091_),
    .B2(_12069_),
    .Y(_04021_));
 NAND2x1_ASAP7_75t_R _28632_ (.A(_01574_),
    .B(_11765_),
    .Y(_12092_));
 OA21x2_ASAP7_75t_R _28633_ (.A1(net136),
    .A2(_12065_),
    .B(_12092_),
    .Y(_12093_));
 NOR2x1_ASAP7_75t_R _28634_ (.A(_01610_),
    .B(_12072_),
    .Y(_12094_));
 AO22x1_ASAP7_75t_R _28635_ (.A1(_12064_),
    .A2(_12093_),
    .B1(_12094_),
    .B2(_12069_),
    .Y(_04022_));
 OR2x2_ASAP7_75t_R _28636_ (.A(net144),
    .B(_11722_),
    .Y(_12095_));
 NAND2x1_ASAP7_75t_R _28637_ (.A(_11723_),
    .B(_01634_),
    .Y(_12096_));
 NOR2x1_ASAP7_75t_R _28638_ (.A(_01609_),
    .B(_11750_),
    .Y(_12097_));
 AO32x1_ASAP7_75t_R _28639_ (.A1(_11751_),
    .A2(_12095_),
    .A3(_12096_),
    .B1(_12097_),
    .B2(_11758_),
    .Y(_04023_));
 NAND2x1_ASAP7_75t_R _28640_ (.A(_01573_),
    .B(_11765_),
    .Y(_12098_));
 OA21x2_ASAP7_75t_R _28641_ (.A1(net137),
    .A2(_12065_),
    .B(_12098_),
    .Y(_12099_));
 NOR2x1_ASAP7_75t_R _28642_ (.A(_01608_),
    .B(_12072_),
    .Y(_12100_));
 AO22x1_ASAP7_75t_R _28643_ (.A1(_12064_),
    .A2(_12099_),
    .B1(_12100_),
    .B2(_12069_),
    .Y(_04024_));
 NAND2x1_ASAP7_75t_R _28644_ (.A(_01572_),
    .B(_11765_),
    .Y(_12101_));
 OA21x2_ASAP7_75t_R _28645_ (.A1(net138),
    .A2(_11767_),
    .B(_12101_),
    .Y(_12102_));
 NOR2x1_ASAP7_75t_R _28646_ (.A(_01607_),
    .B(_12072_),
    .Y(_12103_));
 AO22x1_ASAP7_75t_R _28647_ (.A1(_11763_),
    .A2(_12102_),
    .B1(_12103_),
    .B2(_11771_),
    .Y(_04025_));
 NAND2x1_ASAP7_75t_R _28648_ (.A(_01571_),
    .B(_11765_),
    .Y(_12104_));
 OA21x2_ASAP7_75t_R _28649_ (.A1(net140),
    .A2(_11767_),
    .B(_12104_),
    .Y(_12105_));
 NOR2x1_ASAP7_75t_R _28650_ (.A(_01606_),
    .B(_11774_),
    .Y(_12106_));
 AO22x1_ASAP7_75t_R _28651_ (.A1(_11763_),
    .A2(_12105_),
    .B1(_12106_),
    .B2(_11771_),
    .Y(_04026_));
 NAND2x1_ASAP7_75t_R _28652_ (.A(_01570_),
    .B(_11765_),
    .Y(_12107_));
 OA21x2_ASAP7_75t_R _28653_ (.A1(net141),
    .A2(_11767_),
    .B(_12107_),
    .Y(_12108_));
 NOR2x1_ASAP7_75t_R _28654_ (.A(_01605_),
    .B(_11774_),
    .Y(_12109_));
 AO22x1_ASAP7_75t_R _28655_ (.A1(_11763_),
    .A2(_12108_),
    .B1(_12109_),
    .B2(_11771_),
    .Y(_04027_));
 NAND2x1_ASAP7_75t_R _28656_ (.A(_01604_),
    .B(_11779_),
    .Y(_12110_));
 OA21x2_ASAP7_75t_R _28657_ (.A1(net117),
    .A2(_11778_),
    .B(_12110_),
    .Y(_04028_));
 NAND2x1_ASAP7_75t_R _28658_ (.A(_01603_),
    .B(_11779_),
    .Y(_12111_));
 OA21x2_ASAP7_75t_R _28659_ (.A1(net128),
    .A2(_11778_),
    .B(_12111_),
    .Y(_04029_));
 NAND2x1_ASAP7_75t_R _28660_ (.A(_01602_),
    .B(_11779_),
    .Y(_12112_));
 OA21x2_ASAP7_75t_R _28661_ (.A1(net139),
    .A2(_11778_),
    .B(_12112_),
    .Y(_04030_));
 NAND2x1_ASAP7_75t_R _28662_ (.A(_01601_),
    .B(_11779_),
    .Y(_12113_));
 OA21x2_ASAP7_75t_R _28663_ (.A1(net142),
    .A2(_11778_),
    .B(_12113_),
    .Y(_04031_));
 NAND2x1_ASAP7_75t_R _28664_ (.A(_01600_),
    .B(_11779_),
    .Y(_12114_));
 OA21x2_ASAP7_75t_R _28665_ (.A1(net143),
    .A2(_11778_),
    .B(_12114_),
    .Y(_04032_));
 NAND2x1_ASAP7_75t_R _28666_ (.A(_01599_),
    .B(_11779_),
    .Y(_12115_));
 OA21x2_ASAP7_75t_R _28667_ (.A1(net144),
    .A2(_11778_),
    .B(_12115_),
    .Y(_04033_));
 NOR2x1_ASAP7_75t_R _28668_ (.A(_01598_),
    .B(_11756_),
    .Y(_12116_));
 NAND2x1_ASAP7_75t_R _28669_ (.A(_11723_),
    .B(_01633_),
    .Y(_12117_));
 OAI21x1_ASAP7_75t_R _28670_ (.A1(net145),
    .A2(_11723_),
    .B(_12117_),
    .Y(_12118_));
 INVx1_ASAP7_75t_R _28671_ (.A(_12118_),
    .Y(_12119_));
 AO22x1_ASAP7_75t_R _28672_ (.A1(_11759_),
    .A2(_12116_),
    .B1(_12119_),
    .B2(_11752_),
    .Y(_04034_));
 BUFx12f_ASAP7_75t_R _28673_ (.A(_11777_),
    .Y(_12120_));
 NAND2x1_ASAP7_75t_R _28674_ (.A(_01597_),
    .B(_12120_),
    .Y(_12121_));
 OA21x2_ASAP7_75t_R _28675_ (.A1(net145),
    .A2(_11778_),
    .B(_12121_),
    .Y(_04035_));
 NAND2x1_ASAP7_75t_R _28676_ (.A(_01596_),
    .B(_12120_),
    .Y(_12122_));
 OA21x2_ASAP7_75t_R _28677_ (.A1(net146),
    .A2(_11778_),
    .B(_12122_),
    .Y(_04036_));
 NAND2x1_ASAP7_75t_R _28678_ (.A(_01595_),
    .B(_12120_),
    .Y(_12123_));
 OA21x2_ASAP7_75t_R _28679_ (.A1(net147),
    .A2(_11778_),
    .B(_12123_),
    .Y(_04037_));
 BUFx6f_ASAP7_75t_R _28680_ (.A(_11777_),
    .Y(_12124_));
 NAND2x1_ASAP7_75t_R _28681_ (.A(_01594_),
    .B(_12120_),
    .Y(_12125_));
 OA21x2_ASAP7_75t_R _28682_ (.A1(net148),
    .A2(_12124_),
    .B(_12125_),
    .Y(_04038_));
 NAND2x1_ASAP7_75t_R _28683_ (.A(_01593_),
    .B(_12120_),
    .Y(_12126_));
 OA21x2_ASAP7_75t_R _28684_ (.A1(net118),
    .A2(_12124_),
    .B(_12126_),
    .Y(_04039_));
 NAND2x1_ASAP7_75t_R _28685_ (.A(_01592_),
    .B(_12120_),
    .Y(_12127_));
 OA21x2_ASAP7_75t_R _28686_ (.A1(net119),
    .A2(_12124_),
    .B(_12127_),
    .Y(_04040_));
 NAND2x1_ASAP7_75t_R _28687_ (.A(_01591_),
    .B(_12120_),
    .Y(_12128_));
 OA21x2_ASAP7_75t_R _28688_ (.A1(net120),
    .A2(_12124_),
    .B(_12128_),
    .Y(_04041_));
 NAND2x1_ASAP7_75t_R _28689_ (.A(_01590_),
    .B(_12120_),
    .Y(_12129_));
 OA21x2_ASAP7_75t_R _28690_ (.A1(net121),
    .A2(_12124_),
    .B(_12129_),
    .Y(_04042_));
 NAND2x1_ASAP7_75t_R _28691_ (.A(_01589_),
    .B(_12120_),
    .Y(_12130_));
 OA21x2_ASAP7_75t_R _28692_ (.A1(net122),
    .A2(_12124_),
    .B(_12130_),
    .Y(_04043_));
 NAND2x1_ASAP7_75t_R _28693_ (.A(_01588_),
    .B(_12120_),
    .Y(_12131_));
 OA21x2_ASAP7_75t_R _28694_ (.A1(net123),
    .A2(_12124_),
    .B(_12131_),
    .Y(_04044_));
 NOR2x1_ASAP7_75t_R _28695_ (.A(_01587_),
    .B(_11756_),
    .Y(_12132_));
 NAND2x1_ASAP7_75t_R _28696_ (.A(_11722_),
    .B(_01632_),
    .Y(_12133_));
 OAI21x1_ASAP7_75t_R _28697_ (.A1(net146),
    .A2(_11723_),
    .B(_12133_),
    .Y(_12134_));
 INVx1_ASAP7_75t_R _28698_ (.A(_12134_),
    .Y(_12135_));
 AO22x1_ASAP7_75t_R _28699_ (.A1(_11759_),
    .A2(_12132_),
    .B1(_12135_),
    .B2(_11752_),
    .Y(_04045_));
 BUFx12f_ASAP7_75t_R _28700_ (.A(_11776_),
    .Y(_12136_));
 NAND2x1_ASAP7_75t_R _28701_ (.A(_01586_),
    .B(_12136_),
    .Y(_12137_));
 OA21x2_ASAP7_75t_R _28702_ (.A1(net124),
    .A2(_12124_),
    .B(_12137_),
    .Y(_04046_));
 NAND2x1_ASAP7_75t_R _28703_ (.A(_01585_),
    .B(_12136_),
    .Y(_12138_));
 OA21x2_ASAP7_75t_R _28704_ (.A1(net125),
    .A2(_12124_),
    .B(_12138_),
    .Y(_04047_));
 NAND2x1_ASAP7_75t_R _28705_ (.A(_01584_),
    .B(_12136_),
    .Y(_12139_));
 OA21x2_ASAP7_75t_R _28706_ (.A1(net126),
    .A2(_12124_),
    .B(_12139_),
    .Y(_04048_));
 BUFx6f_ASAP7_75t_R _28707_ (.A(_11777_),
    .Y(_12140_));
 NAND2x1_ASAP7_75t_R _28708_ (.A(_01583_),
    .B(_12136_),
    .Y(_12141_));
 OA21x2_ASAP7_75t_R _28709_ (.A1(net127),
    .A2(_12140_),
    .B(_12141_),
    .Y(_04049_));
 NAND2x1_ASAP7_75t_R _28710_ (.A(_01582_),
    .B(_12136_),
    .Y(_12142_));
 OA21x2_ASAP7_75t_R _28711_ (.A1(net129),
    .A2(_12140_),
    .B(_12142_),
    .Y(_04050_));
 NAND2x1_ASAP7_75t_R _28712_ (.A(_01581_),
    .B(_12136_),
    .Y(_12143_));
 OA21x2_ASAP7_75t_R _28713_ (.A1(net130),
    .A2(_12140_),
    .B(_12143_),
    .Y(_04051_));
 NAND2x1_ASAP7_75t_R _28714_ (.A(_01580_),
    .B(_12136_),
    .Y(_12144_));
 OA21x2_ASAP7_75t_R _28715_ (.A1(net131),
    .A2(_12140_),
    .B(_12144_),
    .Y(_04052_));
 NAND2x1_ASAP7_75t_R _28716_ (.A(_01579_),
    .B(_12136_),
    .Y(_12145_));
 OA21x2_ASAP7_75t_R _28717_ (.A1(net132),
    .A2(_12140_),
    .B(_12145_),
    .Y(_04053_));
 NAND2x1_ASAP7_75t_R _28718_ (.A(_01578_),
    .B(_12136_),
    .Y(_12146_));
 OA21x2_ASAP7_75t_R _28719_ (.A1(net133),
    .A2(_12140_),
    .B(_12146_),
    .Y(_04054_));
 NAND2x1_ASAP7_75t_R _28720_ (.A(_01577_),
    .B(_12136_),
    .Y(_12147_));
 OA21x2_ASAP7_75t_R _28721_ (.A1(net134),
    .A2(_12140_),
    .B(_12147_),
    .Y(_04055_));
 NOR2x1_ASAP7_75t_R _28722_ (.A(_01576_),
    .B(_11756_),
    .Y(_12148_));
 NAND2x1_ASAP7_75t_R _28723_ (.A(_05711_),
    .B(_01630_),
    .Y(_12149_));
 OAI21x1_ASAP7_75t_R _28724_ (.A1(net147),
    .A2(_05711_),
    .B(_12149_),
    .Y(_12150_));
 INVx1_ASAP7_75t_R _28725_ (.A(_12150_),
    .Y(_12151_));
 AO22x1_ASAP7_75t_R _28726_ (.A1(_11759_),
    .A2(_12148_),
    .B1(_12151_),
    .B2(_11752_),
    .Y(_04056_));
 NAND2x1_ASAP7_75t_R _28727_ (.A(_01575_),
    .B(_11777_),
    .Y(_12152_));
 OA21x2_ASAP7_75t_R _28728_ (.A1(net135),
    .A2(_12140_),
    .B(_12152_),
    .Y(_04057_));
 NAND2x1_ASAP7_75t_R _28729_ (.A(_01574_),
    .B(_11777_),
    .Y(_12153_));
 OA21x2_ASAP7_75t_R _28730_ (.A1(net136),
    .A2(_12140_),
    .B(_12153_),
    .Y(_04058_));
 NAND2x1_ASAP7_75t_R _28731_ (.A(_01573_),
    .B(_11777_),
    .Y(_12154_));
 OA21x2_ASAP7_75t_R _28732_ (.A1(net137),
    .A2(_12140_),
    .B(_12154_),
    .Y(_04059_));
 NAND2x1_ASAP7_75t_R _28733_ (.A(_01572_),
    .B(_11777_),
    .Y(_12155_));
 OA21x2_ASAP7_75t_R _28734_ (.A1(net138),
    .A2(_11779_),
    .B(_12155_),
    .Y(_04060_));
 NAND2x1_ASAP7_75t_R _28735_ (.A(_01571_),
    .B(_11777_),
    .Y(_12156_));
 OA21x2_ASAP7_75t_R _28736_ (.A1(net140),
    .A2(_11779_),
    .B(_12156_),
    .Y(_04061_));
 NAND2x1_ASAP7_75t_R _28737_ (.A(_01570_),
    .B(_11777_),
    .Y(_12157_));
 OA21x2_ASAP7_75t_R _28738_ (.A1(net141),
    .A2(_11779_),
    .B(_12157_),
    .Y(_04062_));
 OR2x2_ASAP7_75t_R _28739_ (.A(net148),
    .B(_05711_),
    .Y(_12158_));
 NAND2x1_ASAP7_75t_R _28740_ (.A(_05712_),
    .B(_01629_),
    .Y(_12159_));
 NOR2x1_ASAP7_75t_R _28741_ (.A(_02204_),
    .B(_11750_),
    .Y(_12160_));
 AO32x1_ASAP7_75t_R _28742_ (.A1(_11751_),
    .A2(_12158_),
    .A3(_12159_),
    .B1(_12160_),
    .B2(_11758_),
    .Y(_04063_));
 BUFx6f_ASAP7_75t_R _28743_ (.A(_05460_),
    .Y(_12161_));
 BUFx6f_ASAP7_75t_R _28744_ (.A(_05460_),
    .Y(_12162_));
 NOR2x1_ASAP7_75t_R _28745_ (.A(_12162_),
    .B(_01569_),
    .Y(_12163_));
 AO21x1_ASAP7_75t_R _28746_ (.A1(_12161_),
    .A2(_11486_),
    .B(_12163_),
    .Y(net240));
 OR3x1_ASAP7_75t_R _28747_ (.A(_05703_),
    .B(net116),
    .C(_05715_),
    .Y(_12164_));
 BUFx6f_ASAP7_75t_R _28748_ (.A(_12164_),
    .Y(_12165_));
 BUFx6f_ASAP7_75t_R _28749_ (.A(_12165_),
    .Y(_12166_));
 NAND2x1_ASAP7_75t_R _28750_ (.A(_01569_),
    .B(_12166_),
    .Y(_12167_));
 OA21x2_ASAP7_75t_R _28751_ (.A1(net240),
    .A2(_12166_),
    .B(_12167_),
    .Y(_04064_));
 NOR2x1_ASAP7_75t_R _28752_ (.A(_12162_),
    .B(_01568_),
    .Y(_12168_));
 AO21x1_ASAP7_75t_R _28753_ (.A1(_12161_),
    .A2(_11484_),
    .B(_12168_),
    .Y(net241));
 BUFx6f_ASAP7_75t_R _28754_ (.A(_12165_),
    .Y(_12169_));
 NAND2x1_ASAP7_75t_R _28755_ (.A(_01568_),
    .B(_12166_),
    .Y(_12170_));
 OA21x2_ASAP7_75t_R _28756_ (.A1(_12169_),
    .A2(net241),
    .B(_12170_),
    .Y(_04065_));
 NOR2x1_ASAP7_75t_R _28757_ (.A(_12162_),
    .B(_01567_),
    .Y(_12171_));
 AO21x1_ASAP7_75t_R _28758_ (.A1(_12161_),
    .A2(_11497_),
    .B(_12171_),
    .Y(net242));
 NAND2x1_ASAP7_75t_R _28759_ (.A(_01567_),
    .B(_12166_),
    .Y(_12172_));
 OA21x2_ASAP7_75t_R _28760_ (.A1(_12169_),
    .A2(net242),
    .B(_12172_),
    .Y(_04066_));
 BUFx6f_ASAP7_75t_R _28761_ (.A(_05460_),
    .Y(_12173_));
 INVx1_ASAP7_75t_R _28762_ (.A(_01566_),
    .Y(_12174_));
 BUFx6f_ASAP7_75t_R _28763_ (.A(_05703_),
    .Y(_12175_));
 OR3x1_ASAP7_75t_R _28764_ (.A(_12175_),
    .B(_11502_),
    .C(_11509_),
    .Y(_12176_));
 OA21x2_ASAP7_75t_R _28765_ (.A1(_12173_),
    .A2(_12174_),
    .B(_12176_),
    .Y(net243));
 INVx1_ASAP7_75t_R _28766_ (.A(net116),
    .Y(_12177_));
 AND2x6_ASAP7_75t_R _28767_ (.A(_12177_),
    .B(_05717_),
    .Y(_12178_));
 BUFx6f_ASAP7_75t_R _28768_ (.A(_12178_),
    .Y(_12179_));
 BUFx6f_ASAP7_75t_R _28769_ (.A(_12165_),
    .Y(_12180_));
 AND2x2_ASAP7_75t_R _28770_ (.A(_12174_),
    .B(_12180_),
    .Y(_12181_));
 AO21x1_ASAP7_75t_R _28771_ (.A1(_12179_),
    .A2(net243),
    .B(_12181_),
    .Y(_04067_));
 INVx1_ASAP7_75t_R _28772_ (.A(_01565_),
    .Y(_12182_));
 OR3x1_ASAP7_75t_R _28773_ (.A(_05703_),
    .B(_11514_),
    .C(_11537_),
    .Y(_12183_));
 OA21x2_ASAP7_75t_R _28774_ (.A1(_12173_),
    .A2(_12182_),
    .B(_12183_),
    .Y(net244));
 AND2x2_ASAP7_75t_R _28775_ (.A(_12182_),
    .B(_12180_),
    .Y(_12184_));
 AO21x1_ASAP7_75t_R _28776_ (.A1(_12179_),
    .A2(net244),
    .B(_12184_),
    .Y(_04068_));
 INVx1_ASAP7_75t_R _28777_ (.A(_01564_),
    .Y(_12185_));
 OR3x1_ASAP7_75t_R _28778_ (.A(_05703_),
    .B(_11531_),
    .C(_11532_),
    .Y(_12186_));
 OA21x2_ASAP7_75t_R _28779_ (.A1(_12173_),
    .A2(_12185_),
    .B(_12186_),
    .Y(net245));
 AND2x2_ASAP7_75t_R _28780_ (.A(_12185_),
    .B(_12180_),
    .Y(_12187_));
 AO21x1_ASAP7_75t_R _28781_ (.A1(_12179_),
    .A2(net245),
    .B(_12187_),
    .Y(_04069_));
 NAND2x1_ASAP7_75t_R _28782_ (.A(_12175_),
    .B(_01563_),
    .Y(_12188_));
 OA21x2_ASAP7_75t_R _28783_ (.A1(_12175_),
    .A2(_11555_),
    .B(_12188_),
    .Y(net246));
 BUFx6f_ASAP7_75t_R _28784_ (.A(_12165_),
    .Y(_12189_));
 NAND2x1_ASAP7_75t_R _28785_ (.A(_01563_),
    .B(_12189_),
    .Y(_12190_));
 OA21x2_ASAP7_75t_R _28786_ (.A1(_12169_),
    .A2(net246),
    .B(_12190_),
    .Y(_04070_));
 INVx1_ASAP7_75t_R _28787_ (.A(_01562_),
    .Y(_12191_));
 OR3x1_ASAP7_75t_R _28788_ (.A(_05703_),
    .B(_11554_),
    .C(_11561_),
    .Y(_12192_));
 OA21x2_ASAP7_75t_R _28789_ (.A1(_12173_),
    .A2(_12191_),
    .B(_12192_),
    .Y(net247));
 AND2x2_ASAP7_75t_R _28790_ (.A(_12191_),
    .B(_12180_),
    .Y(_12193_));
 AO21x1_ASAP7_75t_R _28791_ (.A1(_12179_),
    .A2(net247),
    .B(_12193_),
    .Y(_04071_));
 NOR2x1_ASAP7_75t_R _28792_ (.A(_12162_),
    .B(_01561_),
    .Y(_12194_));
 AO21x1_ASAP7_75t_R _28793_ (.A1(_12161_),
    .A2(_11573_),
    .B(_12194_),
    .Y(net248));
 NAND2x1_ASAP7_75t_R _28794_ (.A(_01561_),
    .B(_12189_),
    .Y(_12195_));
 OA21x2_ASAP7_75t_R _28795_ (.A1(_12169_),
    .A2(net248),
    .B(_12195_),
    .Y(_04072_));
 NOR2x1_ASAP7_75t_R _28796_ (.A(_12162_),
    .B(_01560_),
    .Y(_12196_));
 AO21x1_ASAP7_75t_R _28797_ (.A1(_12161_),
    .A2(_11582_),
    .B(_12196_),
    .Y(net249));
 NAND2x1_ASAP7_75t_R _28798_ (.A(_01560_),
    .B(_12189_),
    .Y(_12197_));
 OA21x2_ASAP7_75t_R _28799_ (.A1(_12169_),
    .A2(net249),
    .B(_12197_),
    .Y(_04073_));
 INVx1_ASAP7_75t_R _28800_ (.A(_01559_),
    .Y(_12198_));
 OR3x1_ASAP7_75t_R _28801_ (.A(_05703_),
    .B(_11585_),
    .C(_11590_),
    .Y(_12199_));
 OA21x2_ASAP7_75t_R _28802_ (.A1(_12173_),
    .A2(_12198_),
    .B(_12199_),
    .Y(net250));
 AND2x2_ASAP7_75t_R _28803_ (.A(_12198_),
    .B(_12180_),
    .Y(_12200_));
 AO21x1_ASAP7_75t_R _28804_ (.A1(_12179_),
    .A2(net250),
    .B(_12200_),
    .Y(_04074_));
 NOR2x1_ASAP7_75t_R _28805_ (.A(_12162_),
    .B(_01558_),
    .Y(_12201_));
 AO21x1_ASAP7_75t_R _28806_ (.A1(_12161_),
    .A2(_11606_),
    .B(_12201_),
    .Y(net251));
 NAND2x1_ASAP7_75t_R _28807_ (.A(_01558_),
    .B(_12189_),
    .Y(_12202_));
 OA21x2_ASAP7_75t_R _28808_ (.A1(_12169_),
    .A2(net251),
    .B(_12202_),
    .Y(_04075_));
 INVx1_ASAP7_75t_R _28809_ (.A(_01557_),
    .Y(_12203_));
 OR3x1_ASAP7_75t_R _28810_ (.A(_05703_),
    .B(_11605_),
    .C(_11613_),
    .Y(_12204_));
 OA21x2_ASAP7_75t_R _28811_ (.A1(_12173_),
    .A2(_12203_),
    .B(_12204_),
    .Y(net252));
 AND2x2_ASAP7_75t_R _28812_ (.A(_12203_),
    .B(_12180_),
    .Y(_12205_));
 AO21x1_ASAP7_75t_R _28813_ (.A1(_12179_),
    .A2(net252),
    .B(_12205_),
    .Y(_04076_));
 NOR2x1_ASAP7_75t_R _28814_ (.A(_12162_),
    .B(_01556_),
    .Y(_12206_));
 AO21x1_ASAP7_75t_R _28815_ (.A1(_12161_),
    .A2(_11619_),
    .B(_12206_),
    .Y(net253));
 NAND2x1_ASAP7_75t_R _28816_ (.A(_01556_),
    .B(_12189_),
    .Y(_12207_));
 OA21x2_ASAP7_75t_R _28817_ (.A1(_12169_),
    .A2(net253),
    .B(_12207_),
    .Y(_04077_));
 NAND2x1_ASAP7_75t_R _28818_ (.A(_12175_),
    .B(_01555_),
    .Y(_12208_));
 OA21x2_ASAP7_75t_R _28819_ (.A1(_12175_),
    .A2(_11639_),
    .B(_12208_),
    .Y(net254));
 NAND2x1_ASAP7_75t_R _28820_ (.A(_01555_),
    .B(_12189_),
    .Y(_12209_));
 OA21x2_ASAP7_75t_R _28821_ (.A1(_12169_),
    .A2(net254),
    .B(_12209_),
    .Y(_04078_));
 NOR2x1_ASAP7_75t_R _28822_ (.A(_12162_),
    .B(_01554_),
    .Y(_12210_));
 AO21x1_ASAP7_75t_R _28823_ (.A1(_12161_),
    .A2(_11638_),
    .B(_12210_),
    .Y(net255));
 NAND2x1_ASAP7_75t_R _28824_ (.A(_01554_),
    .B(_12189_),
    .Y(_12211_));
 OA21x2_ASAP7_75t_R _28825_ (.A1(_12169_),
    .A2(net255),
    .B(_12211_),
    .Y(_04079_));
 INVx1_ASAP7_75t_R _28826_ (.A(_01553_),
    .Y(_12212_));
 OR3x1_ASAP7_75t_R _28827_ (.A(_05703_),
    .B(_11646_),
    .C(_11648_),
    .Y(_12213_));
 OA21x2_ASAP7_75t_R _28828_ (.A1(_12173_),
    .A2(_12212_),
    .B(_12213_),
    .Y(net256));
 AND2x2_ASAP7_75t_R _28829_ (.A(_12212_),
    .B(_12165_),
    .Y(_12214_));
 AO21x1_ASAP7_75t_R _28830_ (.A1(_12179_),
    .A2(net256),
    .B(_12214_),
    .Y(_04080_));
 NOR2x1_ASAP7_75t_R _28831_ (.A(_12162_),
    .B(_01552_),
    .Y(_12215_));
 AO21x1_ASAP7_75t_R _28832_ (.A1(_05461_),
    .A2(_11660_),
    .B(_12215_),
    .Y(net257));
 NAND2x1_ASAP7_75t_R _28833_ (.A(_01552_),
    .B(_12189_),
    .Y(_12216_));
 OA21x2_ASAP7_75t_R _28834_ (.A1(_12169_),
    .A2(net257),
    .B(_12216_),
    .Y(_04081_));
 NOR2x1_ASAP7_75t_R _28835_ (.A(_12162_),
    .B(_01551_),
    .Y(_12217_));
 AO21x1_ASAP7_75t_R _28836_ (.A1(_05461_),
    .A2(_11667_),
    .B(_12217_),
    .Y(net258));
 NAND2x1_ASAP7_75t_R _28837_ (.A(_01551_),
    .B(_12189_),
    .Y(_12218_));
 OA21x2_ASAP7_75t_R _28838_ (.A1(_12166_),
    .A2(net258),
    .B(_12218_),
    .Y(_04082_));
 INVx1_ASAP7_75t_R _28839_ (.A(_01550_),
    .Y(_12219_));
 NAND2x1_ASAP7_75t_R _28840_ (.A(_05461_),
    .B(_11675_),
    .Y(_12220_));
 OA21x2_ASAP7_75t_R _28841_ (.A1(_12173_),
    .A2(_12219_),
    .B(_12220_),
    .Y(net259));
 AND2x2_ASAP7_75t_R _28842_ (.A(_12219_),
    .B(_12165_),
    .Y(_12221_));
 AO21x1_ASAP7_75t_R _28843_ (.A1(_12179_),
    .A2(net259),
    .B(_12221_),
    .Y(_04083_));
 AND2x2_ASAP7_75t_R _28844_ (.A(_12175_),
    .B(_01549_),
    .Y(_12222_));
 AOI21x1_ASAP7_75t_R _28845_ (.A1(_12173_),
    .A2(_05508_),
    .B(_12222_),
    .Y(net260));
 NOR2x1_ASAP7_75t_R _28846_ (.A(_01549_),
    .B(_12178_),
    .Y(_12223_));
 AO21x1_ASAP7_75t_R _28847_ (.A1(_12179_),
    .A2(net260),
    .B(_12223_),
    .Y(_04084_));
 NOR2x1_ASAP7_75t_R _28848_ (.A(_05460_),
    .B(_01548_),
    .Y(_12224_));
 AO21x1_ASAP7_75t_R _28849_ (.A1(_05461_),
    .A2(_11685_),
    .B(_12224_),
    .Y(net261));
 NAND2x1_ASAP7_75t_R _28850_ (.A(_01548_),
    .B(_12189_),
    .Y(_12225_));
 OA21x2_ASAP7_75t_R _28851_ (.A1(_12166_),
    .A2(net261),
    .B(_12225_),
    .Y(_04085_));
 INVx1_ASAP7_75t_R _28852_ (.A(_01547_),
    .Y(_12226_));
 NAND2x1_ASAP7_75t_R _28853_ (.A(_05461_),
    .B(_11695_),
    .Y(_12227_));
 OA21x2_ASAP7_75t_R _28854_ (.A1(_12173_),
    .A2(_12226_),
    .B(_12227_),
    .Y(net262));
 AND2x2_ASAP7_75t_R _28855_ (.A(_12226_),
    .B(_12165_),
    .Y(_12228_));
 AO21x1_ASAP7_75t_R _28856_ (.A1(_12179_),
    .A2(net262),
    .B(_12228_),
    .Y(_04086_));
 INVx1_ASAP7_75t_R _28857_ (.A(_01546_),
    .Y(_12229_));
 NAND2x1_ASAP7_75t_R _28858_ (.A(_05461_),
    .B(_05521_),
    .Y(_12230_));
 OA21x2_ASAP7_75t_R _28859_ (.A1(_12161_),
    .A2(_12229_),
    .B(_12230_),
    .Y(net263));
 AND2x2_ASAP7_75t_R _28860_ (.A(_12229_),
    .B(_12165_),
    .Y(_12231_));
 AO21x1_ASAP7_75t_R _28861_ (.A1(_12178_),
    .A2(net263),
    .B(_12231_),
    .Y(_04087_));
 INVx1_ASAP7_75t_R _28862_ (.A(_01545_),
    .Y(_12232_));
 OR3x1_ASAP7_75t_R _28863_ (.A(_05703_),
    .B(_11440_),
    .C(_11441_),
    .Y(_12233_));
 OA21x2_ASAP7_75t_R _28864_ (.A1(_12161_),
    .A2(_12232_),
    .B(_12233_),
    .Y(net264));
 AND2x2_ASAP7_75t_R _28865_ (.A(_12232_),
    .B(_12165_),
    .Y(_12234_));
 AO21x1_ASAP7_75t_R _28866_ (.A1(_12178_),
    .A2(net264),
    .B(_12234_),
    .Y(_04088_));
 NOR2x1_ASAP7_75t_R _28867_ (.A(_05460_),
    .B(_01544_),
    .Y(_12235_));
 AO21x1_ASAP7_75t_R _28868_ (.A1(_05461_),
    .A2(_11444_),
    .B(_12235_),
    .Y(net265));
 NAND2x1_ASAP7_75t_R _28869_ (.A(_01544_),
    .B(_12180_),
    .Y(_12236_));
 OA21x2_ASAP7_75t_R _28870_ (.A1(_12166_),
    .A2(net265),
    .B(_12236_),
    .Y(_04089_));
 NAND2x1_ASAP7_75t_R _28871_ (.A(_12175_),
    .B(_01543_),
    .Y(_12237_));
 OA21x2_ASAP7_75t_R _28872_ (.A1(_12175_),
    .A2(_11451_),
    .B(_12237_),
    .Y(net266));
 INVx1_ASAP7_75t_R _28873_ (.A(_01543_),
    .Y(_12238_));
 AND2x2_ASAP7_75t_R _28874_ (.A(_12238_),
    .B(_12165_),
    .Y(_12239_));
 AO21x1_ASAP7_75t_R _28875_ (.A1(_12178_),
    .A2(net266),
    .B(_12239_),
    .Y(_04090_));
 NOR2x1_ASAP7_75t_R _28876_ (.A(_05460_),
    .B(_01542_),
    .Y(_12240_));
 AO21x1_ASAP7_75t_R _28877_ (.A1(_05461_),
    .A2(_11435_),
    .B(_12240_),
    .Y(net267));
 NAND2x1_ASAP7_75t_R _28878_ (.A(_01542_),
    .B(_12180_),
    .Y(_12241_));
 OA21x2_ASAP7_75t_R _28879_ (.A1(_12166_),
    .A2(net267),
    .B(_12241_),
    .Y(_04091_));
 NAND2x1_ASAP7_75t_R _28880_ (.A(_12175_),
    .B(_01541_),
    .Y(_12242_));
 OA21x2_ASAP7_75t_R _28881_ (.A1(_12175_),
    .A2(_11464_),
    .B(_12242_),
    .Y(net268));
 NAND2x1_ASAP7_75t_R _28882_ (.A(_01541_),
    .B(_12180_),
    .Y(_12243_));
 OA21x2_ASAP7_75t_R _28883_ (.A1(_12166_),
    .A2(net268),
    .B(_12243_),
    .Y(_04092_));
 NOR2x1_ASAP7_75t_R _28884_ (.A(_05460_),
    .B(_02207_),
    .Y(_12244_));
 AO21x1_ASAP7_75t_R _28885_ (.A1(_05461_),
    .A2(_11459_),
    .B(_12244_),
    .Y(net269));
 NAND2x1_ASAP7_75t_R _28886_ (.A(_02207_),
    .B(_12180_),
    .Y(_12245_));
 OA21x2_ASAP7_75t_R _28887_ (.A1(_12166_),
    .A2(net269),
    .B(_12245_),
    .Y(_04093_));
 BUFx6f_ASAP7_75t_R _28888_ (.A(_00375_),
    .Y(_12246_));
 NAND2x1_ASAP7_75t_R _28889_ (.A(net80),
    .B(_05728_),
    .Y(_12247_));
 OR3x1_ASAP7_75t_R _28890_ (.A(_12246_),
    .B(net25),
    .C(_12247_),
    .Y(_12248_));
 NAND2x1_ASAP7_75t_R _28891_ (.A(_05735_),
    .B(_12248_),
    .Y(_12249_));
 AND3x1_ASAP7_75t_R _28892_ (.A(_00375_),
    .B(net26),
    .C(_13256_),
    .Y(_12250_));
 AND4x1_ASAP7_75t_R _28893_ (.A(net80),
    .B(_05182_),
    .C(_05728_),
    .D(_12250_),
    .Y(_12251_));
 AO21x1_ASAP7_75t_R _28894_ (.A1(_01442_),
    .A2(_05736_),
    .B(_12251_),
    .Y(_12252_));
 AO21x2_ASAP7_75t_R _28895_ (.A1(_05180_),
    .A2(_12249_),
    .B(_12252_),
    .Y(_12253_));
 BUFx6f_ASAP7_75t_R _28896_ (.A(_12253_),
    .Y(_12254_));
 BUFx6f_ASAP7_75t_R _28897_ (.A(_12254_),
    .Y(_12255_));
 NOR2x1_ASAP7_75t_R _28898_ (.A(_01477_),
    .B(_12255_),
    .Y(_12256_));
 AO21x1_ASAP7_75t_R _28899_ (.A1(_05255_),
    .A2(_12255_),
    .B(_12256_),
    .Y(_04177_));
 NOR2x1_ASAP7_75t_R _28900_ (.A(_01476_),
    .B(_12255_),
    .Y(_12257_));
 AO21x1_ASAP7_75t_R _28901_ (.A1(\alu_adder_result_ex[10] ),
    .A2(_12255_),
    .B(_12257_),
    .Y(_04178_));
 AOI21x1_ASAP7_75t_R _28902_ (.A1(_05180_),
    .A2(_12249_),
    .B(_12252_),
    .Y(_12258_));
 BUFx12f_ASAP7_75t_R _28903_ (.A(_12258_),
    .Y(_12259_));
 BUFx6f_ASAP7_75t_R _28904_ (.A(_12259_),
    .Y(_12260_));
 BUFx6f_ASAP7_75t_R _28905_ (.A(_12258_),
    .Y(_12261_));
 NAND2x1_ASAP7_75t_R _28906_ (.A(_01475_),
    .B(_12261_),
    .Y(_12262_));
 OA21x2_ASAP7_75t_R _28907_ (.A1(\alu_adder_result_ex[11] ),
    .A2(_12260_),
    .B(_12262_),
    .Y(_04179_));
 AND2x2_ASAP7_75t_R _28908_ (.A(\alu_adder_result_ex[12] ),
    .B(_12254_),
    .Y(_12263_));
 AO21x1_ASAP7_75t_R _28909_ (.A1(_13270_),
    .A2(_12261_),
    .B(_12263_),
    .Y(_04180_));
 NAND2x1_ASAP7_75t_R _28910_ (.A(_01473_),
    .B(_12261_),
    .Y(_12264_));
 OA21x2_ASAP7_75t_R _28911_ (.A1(\alu_adder_result_ex[13] ),
    .A2(_12260_),
    .B(_12264_),
    .Y(_04181_));
 NAND2x1_ASAP7_75t_R _28912_ (.A(_01472_),
    .B(_12261_),
    .Y(_12265_));
 OA21x2_ASAP7_75t_R _28913_ (.A1(\alu_adder_result_ex[14] ),
    .A2(_12260_),
    .B(_12265_),
    .Y(_04182_));
 NAND2x1_ASAP7_75t_R _28914_ (.A(_01471_),
    .B(_12261_),
    .Y(_12266_));
 OA21x2_ASAP7_75t_R _28915_ (.A1(\alu_adder_result_ex[15] ),
    .A2(_12260_),
    .B(_12266_),
    .Y(_04183_));
 NAND2x1_ASAP7_75t_R _28916_ (.A(_01470_),
    .B(_12261_),
    .Y(_12267_));
 OA21x2_ASAP7_75t_R _28917_ (.A1(\alu_adder_result_ex[16] ),
    .A2(_12260_),
    .B(_12267_),
    .Y(_04184_));
 NAND2x1_ASAP7_75t_R _28918_ (.A(_01469_),
    .B(_12261_),
    .Y(_12268_));
 OA21x2_ASAP7_75t_R _28919_ (.A1(\alu_adder_result_ex[17] ),
    .A2(_12260_),
    .B(_12268_),
    .Y(_04185_));
 BUFx6f_ASAP7_75t_R _28920_ (.A(_12259_),
    .Y(_12269_));
 NAND2x1_ASAP7_75t_R _28921_ (.A(_01468_),
    .B(_12269_),
    .Y(_12270_));
 OA21x2_ASAP7_75t_R _28922_ (.A1(\alu_adder_result_ex[18] ),
    .A2(_12260_),
    .B(_12270_),
    .Y(_04186_));
 NAND2x1_ASAP7_75t_R _28923_ (.A(_01467_),
    .B(_12269_),
    .Y(_12271_));
 OA21x2_ASAP7_75t_R _28924_ (.A1(\alu_adder_result_ex[19] ),
    .A2(_12260_),
    .B(_12271_),
    .Y(_04187_));
 NOR2x1_ASAP7_75t_R _28925_ (.A(_01466_),
    .B(_12254_),
    .Y(_12272_));
 AO21x1_ASAP7_75t_R _28926_ (.A1(\alu_adder_result_ex[1] ),
    .A2(_12255_),
    .B(_12272_),
    .Y(_04188_));
 NAND2x1_ASAP7_75t_R _28927_ (.A(_01465_),
    .B(_12269_),
    .Y(_12273_));
 OA21x2_ASAP7_75t_R _28928_ (.A1(\alu_adder_result_ex[20] ),
    .A2(_12260_),
    .B(_12273_),
    .Y(_04189_));
 NAND2x1_ASAP7_75t_R _28929_ (.A(_01464_),
    .B(_12269_),
    .Y(_12274_));
 OA21x2_ASAP7_75t_R _28930_ (.A1(\alu_adder_result_ex[21] ),
    .A2(_12260_),
    .B(_12274_),
    .Y(_04190_));
 BUFx6f_ASAP7_75t_R _28931_ (.A(_12259_),
    .Y(_12275_));
 NAND2x1_ASAP7_75t_R _28932_ (.A(_01463_),
    .B(_12269_),
    .Y(_12276_));
 OA21x2_ASAP7_75t_R _28933_ (.A1(\alu_adder_result_ex[22] ),
    .A2(_12275_),
    .B(_12276_),
    .Y(_04191_));
 NAND2x1_ASAP7_75t_R _28934_ (.A(_01462_),
    .B(_12269_),
    .Y(_12277_));
 OA21x2_ASAP7_75t_R _28935_ (.A1(\alu_adder_result_ex[23] ),
    .A2(_12275_),
    .B(_12277_),
    .Y(_04192_));
 NAND2x1_ASAP7_75t_R _28936_ (.A(_01461_),
    .B(_12269_),
    .Y(_12278_));
 OA21x2_ASAP7_75t_R _28937_ (.A1(\alu_adder_result_ex[24] ),
    .A2(_12275_),
    .B(_12278_),
    .Y(_04193_));
 NAND2x1_ASAP7_75t_R _28938_ (.A(_01460_),
    .B(_12269_),
    .Y(_12279_));
 OA21x2_ASAP7_75t_R _28939_ (.A1(\alu_adder_result_ex[25] ),
    .A2(_12275_),
    .B(_12279_),
    .Y(_04194_));
 NAND2x1_ASAP7_75t_R _28940_ (.A(_01459_),
    .B(_12269_),
    .Y(_12280_));
 OA21x2_ASAP7_75t_R _28941_ (.A1(\alu_adder_result_ex[26] ),
    .A2(_12275_),
    .B(_12280_),
    .Y(_04195_));
 NOR2x1_ASAP7_75t_R _28942_ (.A(_01458_),
    .B(_12254_),
    .Y(_12281_));
 AO21x1_ASAP7_75t_R _28943_ (.A1(\alu_adder_result_ex[27] ),
    .A2(_12255_),
    .B(_12281_),
    .Y(_04196_));
 NAND2x1_ASAP7_75t_R _28944_ (.A(_01457_),
    .B(_12269_),
    .Y(_12282_));
 OA21x2_ASAP7_75t_R _28945_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_12275_),
    .B(_12282_),
    .Y(_04197_));
 NAND2x1_ASAP7_75t_R _28946_ (.A(_01456_),
    .B(_12259_),
    .Y(_12283_));
 OA21x2_ASAP7_75t_R _28947_ (.A1(\alu_adder_result_ex[29] ),
    .A2(_12275_),
    .B(_12283_),
    .Y(_04198_));
 NAND2x1_ASAP7_75t_R _28948_ (.A(_01455_),
    .B(_12259_),
    .Y(_12284_));
 OA21x2_ASAP7_75t_R _28949_ (.A1(\alu_adder_result_ex[2] ),
    .A2(_12275_),
    .B(_12284_),
    .Y(_04199_));
 NAND2x1_ASAP7_75t_R _28950_ (.A(_01454_),
    .B(_12259_),
    .Y(_12285_));
 OA21x2_ASAP7_75t_R _28951_ (.A1(\alu_adder_result_ex[30] ),
    .A2(_12275_),
    .B(_12285_),
    .Y(_04200_));
 NOR2x1_ASAP7_75t_R _28952_ (.A(_01453_),
    .B(_12254_),
    .Y(_12286_));
 AO21x1_ASAP7_75t_R _28953_ (.A1(\alu_adder_result_ex[31] ),
    .A2(_12255_),
    .B(_12286_),
    .Y(_04201_));
 NAND2x1_ASAP7_75t_R _28954_ (.A(_01452_),
    .B(_12259_),
    .Y(_12287_));
 OA21x2_ASAP7_75t_R _28955_ (.A1(\alu_adder_result_ex[3] ),
    .A2(_12275_),
    .B(_12287_),
    .Y(_04202_));
 NOR2x1_ASAP7_75t_R _28956_ (.A(_01451_),
    .B(_12254_),
    .Y(_12288_));
 AO21x1_ASAP7_75t_R _28957_ (.A1(\alu_adder_result_ex[4] ),
    .A2(_12255_),
    .B(_12288_),
    .Y(_04203_));
 NAND2x1_ASAP7_75t_R _28958_ (.A(_01450_),
    .B(_12259_),
    .Y(_12289_));
 OA21x2_ASAP7_75t_R _28959_ (.A1(\alu_adder_result_ex[5] ),
    .A2(_12261_),
    .B(_12289_),
    .Y(_04204_));
 NOR2x1_ASAP7_75t_R _28960_ (.A(_01449_),
    .B(_12254_),
    .Y(_12290_));
 AO21x1_ASAP7_75t_R _28961_ (.A1(\alu_adder_result_ex[6] ),
    .A2(_12255_),
    .B(_12290_),
    .Y(_04205_));
 NAND2x1_ASAP7_75t_R _28962_ (.A(_01448_),
    .B(_12259_),
    .Y(_12291_));
 OA21x2_ASAP7_75t_R _28963_ (.A1(\alu_adder_result_ex[7] ),
    .A2(_12261_),
    .B(_12291_),
    .Y(_04206_));
 NOR2x1_ASAP7_75t_R _28964_ (.A(_01447_),
    .B(_12254_),
    .Y(_12292_));
 AO21x1_ASAP7_75t_R _28965_ (.A1(\alu_adder_result_ex[8] ),
    .A2(_12255_),
    .B(_12292_),
    .Y(_04207_));
 NAND2x1_ASAP7_75t_R _28966_ (.A(_01446_),
    .B(_12259_),
    .Y(_12293_));
 OA21x2_ASAP7_75t_R _28967_ (.A1(\alu_adder_result_ex[9] ),
    .A2(_12261_),
    .B(_12293_),
    .Y(_04208_));
 OR4x1_ASAP7_75t_R _28968_ (.A(_13243_),
    .B(_14265_),
    .C(_13298_),
    .D(_05735_),
    .Y(_12294_));
 OAI21x1_ASAP7_75t_R _28969_ (.A1(_01445_),
    .A2(_05736_),
    .B(_12294_),
    .Y(_04209_));
 AND3x4_ASAP7_75t_R _28970_ (.A(_13243_),
    .B(_05730_),
    .C(_04987_),
    .Y(net239));
 NAND2x1_ASAP7_75t_R _28971_ (.A(_05179_),
    .B(_05735_),
    .Y(_12295_));
 OA21x2_ASAP7_75t_R _28972_ (.A1(_05735_),
    .A2(net239),
    .B(_12295_),
    .Y(_04210_));
 OA21x2_ASAP7_75t_R _28973_ (.A1(_05729_),
    .A2(_05731_),
    .B(net26),
    .Y(_12296_));
 INVx1_ASAP7_75t_R _28974_ (.A(net26),
    .Y(_12297_));
 AOI21x1_ASAP7_75t_R _28975_ (.A1(_12297_),
    .A2(_12247_),
    .B(_05180_),
    .Y(_12298_));
 OA21x2_ASAP7_75t_R _28976_ (.A1(_12296_),
    .A2(_12298_),
    .B(_12246_),
    .Y(_12299_));
 OR2x2_ASAP7_75t_R _28977_ (.A(net26),
    .B(_12247_),
    .Y(_12300_));
 NAND2x1_ASAP7_75t_R _28978_ (.A(_12246_),
    .B(_13253_),
    .Y(_12301_));
 NOR2x1_ASAP7_75t_R _28979_ (.A(_14274_),
    .B(_14135_),
    .Y(_12302_));
 BUFx6f_ASAP7_75t_R _28980_ (.A(_02326_),
    .Y(_12303_));
 OR2x6_ASAP7_75t_R _28981_ (.A(_14274_),
    .B(_14135_),
    .Y(_12304_));
 OR3x1_ASAP7_75t_R _28982_ (.A(_14272_),
    .B(_12303_),
    .C(_12304_),
    .Y(_12305_));
 OA21x2_ASAP7_75t_R _28983_ (.A1(_05209_),
    .A2(_12302_),
    .B(_12305_),
    .Y(_12306_));
 AO32x1_ASAP7_75t_R _28984_ (.A1(_12246_),
    .A2(_13256_),
    .A3(_12300_),
    .B1(_12301_),
    .B2(_12306_),
    .Y(_12307_));
 NAND2x1_ASAP7_75t_R _28985_ (.A(_12299_),
    .B(_12307_),
    .Y(_12308_));
 OA21x2_ASAP7_75t_R _28986_ (.A1(_13255_),
    .A2(_12299_),
    .B(_12308_),
    .Y(_04211_));
 AND2x2_ASAP7_75t_R _28987_ (.A(_05180_),
    .B(_05731_),
    .Y(_12309_));
 AO21x1_ASAP7_75t_R _28988_ (.A1(net80),
    .A2(_13256_),
    .B(_05729_),
    .Y(_12310_));
 OA211x2_ASAP7_75t_R _28989_ (.A1(_12309_),
    .A2(_12310_),
    .B(_12246_),
    .C(_12297_),
    .Y(_04212_));
 INVx1_ASAP7_75t_R _28990_ (.A(_05731_),
    .Y(_12311_));
 OAI21x1_ASAP7_75t_R _28991_ (.A1(_12311_),
    .A2(_12306_),
    .B(_05728_),
    .Y(_12312_));
 AO21x1_ASAP7_75t_R _28992_ (.A1(_05180_),
    .A2(_12312_),
    .B(_12297_),
    .Y(_12313_));
 AND3x1_ASAP7_75t_R _28993_ (.A(_05728_),
    .B(_05731_),
    .C(_12306_),
    .Y(_12314_));
 OR3x1_ASAP7_75t_R _28994_ (.A(net26),
    .B(_13256_),
    .C(_12314_),
    .Y(_12315_));
 AND3x1_ASAP7_75t_R _28995_ (.A(_12246_),
    .B(_12313_),
    .C(_12315_),
    .Y(_04213_));
 INVx1_ASAP7_75t_R _28996_ (.A(net80),
    .Y(_12316_));
 INVx1_ASAP7_75t_R _28997_ (.A(_12246_),
    .Y(_12317_));
 AO21x1_ASAP7_75t_R _28998_ (.A1(_12317_),
    .A2(_05180_),
    .B(_12250_),
    .Y(_12318_));
 AND3x1_ASAP7_75t_R _28999_ (.A(_12316_),
    .B(_05728_),
    .C(_12318_),
    .Y(_04214_));
 XOR2x2_ASAP7_75t_R _29000_ (.A(_12246_),
    .B(_05180_),
    .Y(_12319_));
 AND3x4_ASAP7_75t_R _29001_ (.A(net80),
    .B(_05728_),
    .C(_12319_),
    .Y(_12320_));
 BUFx6f_ASAP7_75t_R _29002_ (.A(_12320_),
    .Y(_12321_));
 AO21x1_ASAP7_75t_R _29003_ (.A1(net80),
    .A2(_12319_),
    .B(_12309_),
    .Y(_12322_));
 AOI21x1_ASAP7_75t_R _29004_ (.A1(_05728_),
    .A2(_12322_),
    .B(_01442_),
    .Y(_12323_));
 AO21x1_ASAP7_75t_R _29005_ (.A1(net25),
    .A2(_12321_),
    .B(_12323_),
    .Y(_04215_));
 OR2x2_ASAP7_75t_R _29006_ (.A(_05255_),
    .B(_05735_),
    .Y(_12324_));
 OA21x2_ASAP7_75t_R _29007_ (.A1(_08290_),
    .A2(_05736_),
    .B(_12324_),
    .Y(_04216_));
 NOR2x1_ASAP7_75t_R _29008_ (.A(_18712_),
    .B(_05735_),
    .Y(_12325_));
 AO21x1_ASAP7_75t_R _29009_ (.A1(_08287_),
    .A2(_05735_),
    .B(_12325_),
    .Y(_04217_));
 NAND2x2_ASAP7_75t_R _29010_ (.A(_05178_),
    .B(_12320_),
    .Y(_12326_));
 BUFx6f_ASAP7_75t_R _29011_ (.A(_12326_),
    .Y(_12327_));
 BUFx6f_ASAP7_75t_R _29012_ (.A(_12326_),
    .Y(_12328_));
 NAND2x1_ASAP7_75t_R _29013_ (.A(_01439_),
    .B(_12328_),
    .Y(_12329_));
 OA21x2_ASAP7_75t_R _29014_ (.A1(net78),
    .A2(_12327_),
    .B(_12329_),
    .Y(_04218_));
 AO21x1_ASAP7_75t_R _29015_ (.A1(_05179_),
    .A2(_12321_),
    .B(_08664_),
    .Y(_12330_));
 OA21x2_ASAP7_75t_R _29016_ (.A1(net57),
    .A2(_12327_),
    .B(_12330_),
    .Y(_04219_));
 AO21x1_ASAP7_75t_R _29017_ (.A1(_05179_),
    .A2(_12321_),
    .B(_08714_),
    .Y(_12331_));
 OA21x2_ASAP7_75t_R _29018_ (.A1(net58),
    .A2(_12327_),
    .B(_12331_),
    .Y(_04220_));
 AO21x1_ASAP7_75t_R _29019_ (.A1(_05179_),
    .A2(_12321_),
    .B(_08984_),
    .Y(_12332_));
 OA21x2_ASAP7_75t_R _29020_ (.A1(net60),
    .A2(_12327_),
    .B(_12332_),
    .Y(_04221_));
 AO21x1_ASAP7_75t_R _29021_ (.A1(_05179_),
    .A2(_12321_),
    .B(_08791_),
    .Y(_12333_));
 OA21x2_ASAP7_75t_R _29022_ (.A1(net61),
    .A2(_12327_),
    .B(_12333_),
    .Y(_04222_));
 AO21x1_ASAP7_75t_R _29023_ (.A1(_05179_),
    .A2(_12321_),
    .B(_08839_),
    .Y(_12334_));
 OA21x2_ASAP7_75t_R _29024_ (.A1(net62),
    .A2(_12327_),
    .B(_12334_),
    .Y(_04223_));
 AO21x1_ASAP7_75t_R _29025_ (.A1(_05179_),
    .A2(_12321_),
    .B(_08856_),
    .Y(_12335_));
 OA21x2_ASAP7_75t_R _29026_ (.A1(net63),
    .A2(_12327_),
    .B(_12335_),
    .Y(_04224_));
 NAND2x1_ASAP7_75t_R _29027_ (.A(_01432_),
    .B(_12328_),
    .Y(_12336_));
 OA21x2_ASAP7_75t_R _29028_ (.A1(net64),
    .A2(_12327_),
    .B(_12336_),
    .Y(_04225_));
 NAND2x1_ASAP7_75t_R _29029_ (.A(_01431_),
    .B(_12328_),
    .Y(_12337_));
 OA21x2_ASAP7_75t_R _29030_ (.A1(net65),
    .A2(_12327_),
    .B(_12337_),
    .Y(_04226_));
 NAND2x1_ASAP7_75t_R _29031_ (.A(_01430_),
    .B(_12328_),
    .Y(_12338_));
 OA21x2_ASAP7_75t_R _29032_ (.A1(net66),
    .A2(_12327_),
    .B(_12338_),
    .Y(_04227_));
 BUFx6f_ASAP7_75t_R _29033_ (.A(_12326_),
    .Y(_12339_));
 NAND2x1_ASAP7_75t_R _29034_ (.A(_01429_),
    .B(_12328_),
    .Y(_12340_));
 OA21x2_ASAP7_75t_R _29035_ (.A1(net67),
    .A2(_12339_),
    .B(_12340_),
    .Y(_04228_));
 AO21x1_ASAP7_75t_R _29036_ (.A1(_05179_),
    .A2(_12321_),
    .B(_09520_),
    .Y(_12341_));
 OA21x2_ASAP7_75t_R _29037_ (.A1(net79),
    .A2(_12339_),
    .B(_12341_),
    .Y(_04229_));
 NAND2x1_ASAP7_75t_R _29038_ (.A(_01427_),
    .B(_12328_),
    .Y(_12342_));
 OA21x2_ASAP7_75t_R _29039_ (.A1(net68),
    .A2(_12339_),
    .B(_12342_),
    .Y(_04230_));
 NAND2x1_ASAP7_75t_R _29040_ (.A(_01426_),
    .B(_12326_),
    .Y(_12343_));
 OA21x2_ASAP7_75t_R _29041_ (.A1(net69),
    .A2(_12339_),
    .B(_12343_),
    .Y(_04231_));
 NAND2x1_ASAP7_75t_R _29042_ (.A(_01425_),
    .B(_12326_),
    .Y(_12344_));
 OA21x2_ASAP7_75t_R _29043_ (.A1(net71),
    .A2(_12339_),
    .B(_12344_),
    .Y(_04232_));
 AO21x1_ASAP7_75t_R _29044_ (.A1(_05178_),
    .A2(_12321_),
    .B(_09127_),
    .Y(_12345_));
 OA21x2_ASAP7_75t_R _29045_ (.A1(net72),
    .A2(_12339_),
    .B(_12345_),
    .Y(_04233_));
 AO21x1_ASAP7_75t_R _29046_ (.A1(_05178_),
    .A2(_12321_),
    .B(_09530_),
    .Y(_12346_));
 OA21x2_ASAP7_75t_R _29047_ (.A1(net28),
    .A2(_12339_),
    .B(_12346_),
    .Y(_04234_));
 AO21x1_ASAP7_75t_R _29048_ (.A1(_05178_),
    .A2(_12320_),
    .B(_09546_),
    .Y(_12347_));
 OA21x2_ASAP7_75t_R _29049_ (.A1(net29),
    .A2(_12339_),
    .B(_12347_),
    .Y(_04235_));
 AO21x1_ASAP7_75t_R _29050_ (.A1(_05178_),
    .A2(_12320_),
    .B(_08985_),
    .Y(_12348_));
 OA21x2_ASAP7_75t_R _29051_ (.A1(net30),
    .A2(_12339_),
    .B(_12348_),
    .Y(_04236_));
 AO21x1_ASAP7_75t_R _29052_ (.A1(_05178_),
    .A2(_12320_),
    .B(_09253_),
    .Y(_12349_));
 OA21x2_ASAP7_75t_R _29053_ (.A1(net31),
    .A2(_12339_),
    .B(_12349_),
    .Y(_04237_));
 AO21x1_ASAP7_75t_R _29054_ (.A1(_05178_),
    .A2(_12320_),
    .B(_09404_),
    .Y(_12350_));
 OA21x2_ASAP7_75t_R _29055_ (.A1(net53),
    .A2(_12328_),
    .B(_12350_),
    .Y(_04238_));
 NAND2x1_ASAP7_75t_R _29056_ (.A(_01418_),
    .B(_12326_),
    .Y(_12351_));
 OA21x2_ASAP7_75t_R _29057_ (.A1(net54),
    .A2(_12328_),
    .B(_12351_),
    .Y(_04239_));
 NAND2x1_ASAP7_75t_R _29058_ (.A(_01417_),
    .B(_12326_),
    .Y(_12352_));
 OA21x2_ASAP7_75t_R _29059_ (.A1(net55),
    .A2(_12328_),
    .B(_12352_),
    .Y(_04240_));
 AO21x1_ASAP7_75t_R _29060_ (.A1(_05178_),
    .A2(_12320_),
    .B(_08600_),
    .Y(_12353_));
 OA21x2_ASAP7_75t_R _29061_ (.A1(net56),
    .A2(_12328_),
    .B(_12353_),
    .Y(_04241_));
 OR5x1_ASAP7_75t_R _29062_ (.A(_05150_),
    .B(_14144_),
    .C(_05935_),
    .D(_05159_),
    .E(_06018_),
    .Y(_12354_));
 NAND2x1_ASAP7_75t_R _29063_ (.A(_07642_),
    .B(_12354_),
    .Y(_12355_));
 OAI21x1_ASAP7_75t_R _29064_ (.A1(_06025_),
    .A2(_06051_),
    .B(_07642_),
    .Y(_12356_));
 NAND2x1_ASAP7_75t_R _29065_ (.A(_12355_),
    .B(_12356_),
    .Y(_12357_));
 NAND2x1_ASAP7_75t_R _29066_ (.A(_00331_),
    .B(_07765_),
    .Y(_12358_));
 OAI22x1_ASAP7_75t_R _29067_ (.A1(_02062_),
    .A2(_07713_),
    .B1(_07504_),
    .B2(_01868_),
    .Y(_12359_));
 AO21x1_ASAP7_75t_R _29068_ (.A1(_12357_),
    .A2(_12358_),
    .B(_12359_),
    .Y(_02708_));
 NAND2x1_ASAP7_75t_R _29069_ (.A(_00332_),
    .B(_07765_),
    .Y(_12360_));
 OAI22x1_ASAP7_75t_R _29070_ (.A1(_18080_),
    .A2(_07713_),
    .B1(_07504_),
    .B2(_01867_),
    .Y(_12361_));
 AO21x1_ASAP7_75t_R _29071_ (.A1(_12357_),
    .A2(_12360_),
    .B(_12361_),
    .Y(_02709_));
 AO21x1_ASAP7_75t_R _29072_ (.A1(_07639_),
    .A2(_01866_),
    .B(_07266_),
    .Y(_12362_));
 AO22x1_ASAP7_75t_R _29073_ (.A1(_00333_),
    .A2(_07765_),
    .B1(_12355_),
    .B2(_07643_),
    .Y(_12363_));
 OA211x2_ASAP7_75t_R _29074_ (.A1(_00759_),
    .A2(_07713_),
    .B(_12362_),
    .C(_12363_),
    .Y(_12364_));
 INVx1_ASAP7_75t_R _29075_ (.A(_12364_),
    .Y(_02710_));
 OA22x2_ASAP7_75t_R _29076_ (.A1(_00333_),
    .A2(_07266_),
    .B1(_07765_),
    .B2(_07956_),
    .Y(_12365_));
 OAI21x1_ASAP7_75t_R _29077_ (.A1(_00759_),
    .A2(_12355_),
    .B(_12365_),
    .Y(_02711_));
 BUFx6f_ASAP7_75t_R _29078_ (.A(_11840_),
    .Y(_12366_));
 AND2x2_ASAP7_75t_R _29079_ (.A(_11797_),
    .B(net123),
    .Y(_12367_));
 AO21x1_ASAP7_75t_R _29080_ (.A1(_05523_),
    .A2(net141),
    .B(_12367_),
    .Y(_12368_));
 INVx1_ASAP7_75t_R _29081_ (.A(_01640_),
    .Y(_12369_));
 NAND2x1_ASAP7_75t_R _29082_ (.A(_11797_),
    .B(_01658_),
    .Y(_12370_));
 OA211x2_ASAP7_75t_R _29083_ (.A1(_05542_),
    .A2(_12369_),
    .B(_12370_),
    .C(_05537_),
    .Y(_12371_));
 AO21x2_ASAP7_75t_R _29084_ (.A1(_05539_),
    .A2(_12368_),
    .B(_12371_),
    .Y(_12372_));
 BUFx6f_ASAP7_75t_R _29085_ (.A(_12372_),
    .Y(_12373_));
 BUFx6f_ASAP7_75t_R _29086_ (.A(_12373_),
    .Y(_12374_));
 BUFx6f_ASAP7_75t_R _29087_ (.A(_12374_),
    .Y(_12375_));
 AND2x2_ASAP7_75t_R _29088_ (.A(_05522_),
    .B(net122),
    .Y(_12376_));
 AO21x1_ASAP7_75t_R _29089_ (.A1(_05523_),
    .A2(net140),
    .B(_12376_),
    .Y(_12377_));
 INVx1_ASAP7_75t_R _29090_ (.A(_01641_),
    .Y(_12378_));
 NAND2x1_ASAP7_75t_R _29091_ (.A(_11797_),
    .B(_01659_),
    .Y(_12379_));
 OA211x2_ASAP7_75t_R _29092_ (.A1(_05542_),
    .A2(_12378_),
    .B(_12379_),
    .C(_05532_),
    .Y(_12380_));
 AO21x2_ASAP7_75t_R _29093_ (.A1(_05539_),
    .A2(_12377_),
    .B(_12380_),
    .Y(_12381_));
 BUFx6f_ASAP7_75t_R _29094_ (.A(_12381_),
    .Y(_12382_));
 BUFx6f_ASAP7_75t_R _29095_ (.A(_12382_),
    .Y(_12383_));
 BUFx6f_ASAP7_75t_R _29096_ (.A(_05522_),
    .Y(_12384_));
 AND2x2_ASAP7_75t_R _29097_ (.A(net120),
    .B(_12384_),
    .Y(_12385_));
 AO21x1_ASAP7_75t_R _29098_ (.A1(net137),
    .A2(_05524_),
    .B(_12385_),
    .Y(_12386_));
 INVx1_ASAP7_75t_R _29099_ (.A(_01644_),
    .Y(_12387_));
 NAND2x1_ASAP7_75t_R _29100_ (.A(_12384_),
    .B(_01661_),
    .Y(_12388_));
 OA211x2_ASAP7_75t_R _29101_ (.A1(_05543_),
    .A2(_12387_),
    .B(_12388_),
    .C(_05537_),
    .Y(_12389_));
 AO21x2_ASAP7_75t_R _29102_ (.A1(_11725_),
    .A2(_12386_),
    .B(_12389_),
    .Y(_12390_));
 BUFx6f_ASAP7_75t_R _29103_ (.A(_12390_),
    .Y(_12391_));
 AND2x2_ASAP7_75t_R _29104_ (.A(_12384_),
    .B(net142),
    .Y(_12392_));
 AO21x1_ASAP7_75t_R _29105_ (.A1(_05524_),
    .A2(net127),
    .B(_12392_),
    .Y(_12393_));
 INVx1_ASAP7_75t_R _29106_ (.A(_01654_),
    .Y(_12394_));
 NAND2x1_ASAP7_75t_R _29107_ (.A(_12384_),
    .B(_01631_),
    .Y(_12395_));
 OA211x2_ASAP7_75t_R _29108_ (.A1(_05543_),
    .A2(_12394_),
    .B(_12395_),
    .C(_05537_),
    .Y(_12396_));
 AO21x2_ASAP7_75t_R _29109_ (.A1(_05539_),
    .A2(_12393_),
    .B(_12396_),
    .Y(_12397_));
 AND2x2_ASAP7_75t_R _29110_ (.A(_05522_),
    .B(net145),
    .Y(_12398_));
 AO21x1_ASAP7_75t_R _29111_ (.A1(_05523_),
    .A2(net131),
    .B(_12398_),
    .Y(_12399_));
 INVx1_ASAP7_75t_R _29112_ (.A(_01650_),
    .Y(_12400_));
 NAND2x1_ASAP7_75t_R _29113_ (.A(_05522_),
    .B(_01598_),
    .Y(_12401_));
 OA211x2_ASAP7_75t_R _29114_ (.A1(_05542_),
    .A2(_12400_),
    .B(_12401_),
    .C(_05532_),
    .Y(_12402_));
 AO21x2_ASAP7_75t_R _29115_ (.A1(_05527_),
    .A2(_12399_),
    .B(_12402_),
    .Y(_12403_));
 AND2x2_ASAP7_75t_R _29116_ (.A(_11797_),
    .B(net144),
    .Y(_12404_));
 AO21x1_ASAP7_75t_R _29117_ (.A1(_05523_),
    .A2(net130),
    .B(_12404_),
    .Y(_12405_));
 INVx1_ASAP7_75t_R _29118_ (.A(_01651_),
    .Y(_12406_));
 NAND2x1_ASAP7_75t_R _29119_ (.A(_11797_),
    .B(_01609_),
    .Y(_12407_));
 OA211x2_ASAP7_75t_R _29120_ (.A1(_05542_),
    .A2(_12406_),
    .B(_12407_),
    .C(_05532_),
    .Y(_12408_));
 AO21x2_ASAP7_75t_R _29121_ (.A1(_05527_),
    .A2(_12405_),
    .B(_12408_),
    .Y(_12409_));
 OR2x6_ASAP7_75t_R _29122_ (.A(_12403_),
    .B(_12409_),
    .Y(_12410_));
 AND2x2_ASAP7_75t_R _29123_ (.A(_12384_),
    .B(net143),
    .Y(_12411_));
 AO21x1_ASAP7_75t_R _29124_ (.A1(_05524_),
    .A2(net129),
    .B(_12411_),
    .Y(_12412_));
 INVx1_ASAP7_75t_R _29125_ (.A(_01652_),
    .Y(_12413_));
 NAND2x1_ASAP7_75t_R _29126_ (.A(_12384_),
    .B(_01620_),
    .Y(_12414_));
 OA211x2_ASAP7_75t_R _29127_ (.A1(_05543_),
    .A2(_12413_),
    .B(_12414_),
    .C(_05537_),
    .Y(_12415_));
 AO21x2_ASAP7_75t_R _29128_ (.A1(_05539_),
    .A2(_12412_),
    .B(_12415_),
    .Y(_12416_));
 AND2x2_ASAP7_75t_R _29129_ (.A(_12384_),
    .B(net139),
    .Y(_12417_));
 AO21x1_ASAP7_75t_R _29130_ (.A1(_05524_),
    .A2(net126),
    .B(_12417_),
    .Y(_12418_));
 INVx1_ASAP7_75t_R _29131_ (.A(_01655_),
    .Y(_12419_));
 NAND2x1_ASAP7_75t_R _29132_ (.A(_12384_),
    .B(_01642_),
    .Y(_12420_));
 OA211x2_ASAP7_75t_R _29133_ (.A1(_05543_),
    .A2(_12419_),
    .B(_12420_),
    .C(_05537_),
    .Y(_12421_));
 AO21x2_ASAP7_75t_R _29134_ (.A1(_05539_),
    .A2(_12418_),
    .B(_12421_),
    .Y(_12422_));
 OR4x1_ASAP7_75t_R _29135_ (.A(_12397_),
    .B(_12410_),
    .C(_12416_),
    .D(_12422_),
    .Y(_12423_));
 BUFx6f_ASAP7_75t_R _29136_ (.A(_12423_),
    .Y(_12424_));
 OR3x1_ASAP7_75t_R _29137_ (.A(_12382_),
    .B(_12391_),
    .C(_12424_),
    .Y(_12425_));
 AND2x2_ASAP7_75t_R _29138_ (.A(net147),
    .B(_05543_),
    .Y(_12426_));
 AO21x1_ASAP7_75t_R _29139_ (.A1(net133),
    .A2(_05524_),
    .B(_12426_),
    .Y(_12427_));
 INVx1_ASAP7_75t_R _29140_ (.A(_01648_),
    .Y(_12428_));
 NAND2x1_ASAP7_75t_R _29141_ (.A(_05543_),
    .B(_01576_),
    .Y(_12429_));
 OA211x2_ASAP7_75t_R _29142_ (.A1(_05543_),
    .A2(_12428_),
    .B(_12429_),
    .C(_05537_),
    .Y(_12430_));
 AO21x2_ASAP7_75t_R _29143_ (.A1(_11725_),
    .A2(_12427_),
    .B(_12430_),
    .Y(_12431_));
 AND2x2_ASAP7_75t_R _29144_ (.A(_11797_),
    .B(net119),
    .Y(_12432_));
 AO21x1_ASAP7_75t_R _29145_ (.A1(_05523_),
    .A2(net136),
    .B(_12432_),
    .Y(_12433_));
 INVx1_ASAP7_75t_R _29146_ (.A(_01645_),
    .Y(_12434_));
 NAND2x1_ASAP7_75t_R _29147_ (.A(_11797_),
    .B(_01662_),
    .Y(_12435_));
 OA211x2_ASAP7_75t_R _29148_ (.A1(_05542_),
    .A2(_12434_),
    .B(_12435_),
    .C(_05532_),
    .Y(_12436_));
 AO21x1_ASAP7_75t_R _29149_ (.A1(_05539_),
    .A2(_12433_),
    .B(_12436_),
    .Y(_12437_));
 AND2x2_ASAP7_75t_R _29150_ (.A(_05522_),
    .B(net118),
    .Y(_12438_));
 AO21x1_ASAP7_75t_R _29151_ (.A1(_05523_),
    .A2(net135),
    .B(_12438_),
    .Y(_12439_));
 INVx1_ASAP7_75t_R _29152_ (.A(_01646_),
    .Y(_12440_));
 NAND2x1_ASAP7_75t_R _29153_ (.A(_05522_),
    .B(_01663_),
    .Y(_12441_));
 OA211x2_ASAP7_75t_R _29154_ (.A1(_05542_),
    .A2(_12440_),
    .B(_12441_),
    .C(_05532_),
    .Y(_12442_));
 AO21x2_ASAP7_75t_R _29155_ (.A1(_05527_),
    .A2(_12439_),
    .B(_12442_),
    .Y(_12443_));
 AND2x2_ASAP7_75t_R _29156_ (.A(_11797_),
    .B(net148),
    .Y(_12444_));
 AO21x1_ASAP7_75t_R _29157_ (.A1(_05523_),
    .A2(net134),
    .B(_12444_),
    .Y(_12445_));
 INVx1_ASAP7_75t_R _29158_ (.A(_01647_),
    .Y(_12446_));
 NAND2x1_ASAP7_75t_R _29159_ (.A(_11797_),
    .B(_02204_),
    .Y(_12447_));
 OA211x2_ASAP7_75t_R _29160_ (.A1(_05542_),
    .A2(_12446_),
    .B(_12447_),
    .C(_05532_),
    .Y(_12448_));
 AO21x1_ASAP7_75t_R _29161_ (.A1(_05527_),
    .A2(_12445_),
    .B(_12448_),
    .Y(_12449_));
 AND2x2_ASAP7_75t_R _29162_ (.A(_05522_),
    .B(net146),
    .Y(_12450_));
 AO21x1_ASAP7_75t_R _29163_ (.A1(_05523_),
    .A2(net132),
    .B(_12450_),
    .Y(_12451_));
 INVx1_ASAP7_75t_R _29164_ (.A(_01649_),
    .Y(_12452_));
 NAND2x1_ASAP7_75t_R _29165_ (.A(_05522_),
    .B(_01587_),
    .Y(_12453_));
 OA211x2_ASAP7_75t_R _29166_ (.A1(_05542_),
    .A2(_12452_),
    .B(_12453_),
    .C(_05532_),
    .Y(_12454_));
 AO21x2_ASAP7_75t_R _29167_ (.A1(_05527_),
    .A2(_12451_),
    .B(_12454_),
    .Y(_12455_));
 OR4x1_ASAP7_75t_R _29168_ (.A(_12437_),
    .B(_12443_),
    .C(_12449_),
    .D(_12455_),
    .Y(_12456_));
 OR2x6_ASAP7_75t_R _29169_ (.A(_12431_),
    .B(_12456_),
    .Y(_12457_));
 AO21x1_ASAP7_75t_R _29170_ (.A1(_12374_),
    .A2(_12425_),
    .B(_12457_),
    .Y(_12458_));
 AND2x2_ASAP7_75t_R _29171_ (.A(_05542_),
    .B(net121),
    .Y(_12459_));
 AO21x1_ASAP7_75t_R _29172_ (.A1(_05524_),
    .A2(net138),
    .B(_12459_),
    .Y(_12460_));
 INVx1_ASAP7_75t_R _29173_ (.A(_01643_),
    .Y(_12461_));
 NAND2x1_ASAP7_75t_R _29174_ (.A(_12384_),
    .B(_01660_),
    .Y(_12462_));
 OA211x2_ASAP7_75t_R _29175_ (.A1(_12384_),
    .A2(_12461_),
    .B(_12462_),
    .C(_05537_),
    .Y(_12463_));
 AOI21x1_ASAP7_75t_R _29176_ (.A1(_11725_),
    .A2(_12460_),
    .B(_12463_),
    .Y(_12464_));
 BUFx12f_ASAP7_75t_R _29177_ (.A(_12464_),
    .Y(_12465_));
 BUFx6f_ASAP7_75t_R _29178_ (.A(_12465_),
    .Y(_12466_));
 BUFx6f_ASAP7_75t_R _29179_ (.A(_12466_),
    .Y(_12467_));
 OA211x2_ASAP7_75t_R _29180_ (.A1(_12375_),
    .A2(_12383_),
    .B(_12458_),
    .C(_12467_),
    .Y(_12468_));
 INVx1_ASAP7_75t_R _29181_ (.A(_12468_),
    .Y(_12469_));
 BUFx6f_ASAP7_75t_R _29182_ (.A(_12391_),
    .Y(_12470_));
 BUFx6f_ASAP7_75t_R _29183_ (.A(_12470_),
    .Y(_12471_));
 AO21x2_ASAP7_75t_R _29184_ (.A1(_05539_),
    .A2(_12460_),
    .B(_12463_),
    .Y(_12472_));
 OR3x2_ASAP7_75t_R _29185_ (.A(_12373_),
    .B(_12382_),
    .C(_12472_),
    .Y(_12473_));
 BUFx6f_ASAP7_75t_R _29186_ (.A(_12473_),
    .Y(_12474_));
 BUFx6f_ASAP7_75t_R _29187_ (.A(_11725_),
    .Y(_12475_));
 AND2x2_ASAP7_75t_R _29188_ (.A(_05544_),
    .B(net117),
    .Y(_12476_));
 AO21x1_ASAP7_75t_R _29189_ (.A1(_05524_),
    .A2(net124),
    .B(_12476_),
    .Y(_12477_));
 NAND2x1_ASAP7_75t_R _29190_ (.A(_05543_),
    .B(_01664_),
    .Y(_12478_));
 OA211x2_ASAP7_75t_R _29191_ (.A1(_05544_),
    .A2(_05530_),
    .B(_12478_),
    .C(_11746_),
    .Y(_12479_));
 AOI21x1_ASAP7_75t_R _29192_ (.A1(_12475_),
    .A2(_12477_),
    .B(_12479_),
    .Y(_12480_));
 AND2x2_ASAP7_75t_R _29193_ (.A(_05544_),
    .B(net128),
    .Y(_12481_));
 AO21x1_ASAP7_75t_R _29194_ (.A1(_05524_),
    .A2(net125),
    .B(_12481_),
    .Y(_12482_));
 INVx1_ASAP7_75t_R _29195_ (.A(_01656_),
    .Y(_12483_));
 NAND2x1_ASAP7_75t_R _29196_ (.A(_05544_),
    .B(_01653_),
    .Y(_12484_));
 OA211x2_ASAP7_75t_R _29197_ (.A1(_05544_),
    .A2(_12483_),
    .B(_12484_),
    .C(_11746_),
    .Y(_12485_));
 AO21x1_ASAP7_75t_R _29198_ (.A1(_12475_),
    .A2(_12482_),
    .B(_12485_),
    .Y(_12486_));
 BUFx6f_ASAP7_75t_R _29199_ (.A(_12486_),
    .Y(_12487_));
 AND2x6_ASAP7_75t_R _29200_ (.A(_12480_),
    .B(_12487_),
    .Y(_12488_));
 OA21x2_ASAP7_75t_R _29201_ (.A1(_12471_),
    .A2(_12474_),
    .B(_12488_),
    .Y(_12489_));
 NAND2x1_ASAP7_75t_R _29202_ (.A(_12382_),
    .B(_12465_),
    .Y(_12490_));
 AOI21x1_ASAP7_75t_R _29203_ (.A1(_11742_),
    .A2(_12482_),
    .B(_12485_),
    .Y(_12491_));
 AND2x4_ASAP7_75t_R _29204_ (.A(_12480_),
    .B(_12491_),
    .Y(_12492_));
 AND2x6_ASAP7_75t_R _29205_ (.A(_12490_),
    .B(_12492_),
    .Y(_12493_));
 AOI21x1_ASAP7_75t_R _29206_ (.A1(_05539_),
    .A2(_12368_),
    .B(_12371_),
    .Y(_12494_));
 AND2x4_ASAP7_75t_R _29207_ (.A(_12494_),
    .B(_12465_),
    .Y(_12495_));
 BUFx6f_ASAP7_75t_R _29208_ (.A(_12495_),
    .Y(_12496_));
 OR3x1_ASAP7_75t_R _29209_ (.A(_12457_),
    .B(_12471_),
    .C(_12410_),
    .Y(_12497_));
 NAND2x1_ASAP7_75t_R _29210_ (.A(_12496_),
    .B(_12497_),
    .Y(_12498_));
 AOI21x1_ASAP7_75t_R _29211_ (.A1(_11725_),
    .A2(_12377_),
    .B(_12380_),
    .Y(_12499_));
 BUFx6f_ASAP7_75t_R _29212_ (.A(_12499_),
    .Y(_12500_));
 AND2x4_ASAP7_75t_R _29213_ (.A(_12500_),
    .B(_12465_),
    .Y(_12501_));
 BUFx6f_ASAP7_75t_R _29214_ (.A(_12437_),
    .Y(_12502_));
 INVx2_ASAP7_75t_R _29215_ (.A(_12502_),
    .Y(_12503_));
 BUFx6f_ASAP7_75t_R _29216_ (.A(_12443_),
    .Y(_12504_));
 OA211x2_ASAP7_75t_R _29217_ (.A1(_12503_),
    .A2(_12504_),
    .B(_12375_),
    .C(_12470_),
    .Y(_12505_));
 AOI21x1_ASAP7_75t_R _29218_ (.A1(_12475_),
    .A2(_12386_),
    .B(_12389_),
    .Y(_12506_));
 INVx1_ASAP7_75t_R _29219_ (.A(_12424_),
    .Y(_12507_));
 BUFx6f_ASAP7_75t_R _29220_ (.A(_12472_),
    .Y(_12508_));
 BUFx6f_ASAP7_75t_R _29221_ (.A(_12508_),
    .Y(_12509_));
 AND2x6_ASAP7_75t_R _29222_ (.A(_12494_),
    .B(_12381_),
    .Y(_12510_));
 AND4x1_ASAP7_75t_R _29223_ (.A(_12506_),
    .B(_12507_),
    .C(_12509_),
    .D(_12510_),
    .Y(_12511_));
 AO21x1_ASAP7_75t_R _29224_ (.A1(_12501_),
    .A2(_12505_),
    .B(_12511_),
    .Y(_12512_));
 AO21x2_ASAP7_75t_R _29225_ (.A1(_11742_),
    .A2(_12477_),
    .B(_12479_),
    .Y(_12513_));
 AND2x4_ASAP7_75t_R _29226_ (.A(_12513_),
    .B(_12491_),
    .Y(_12514_));
 BUFx6f_ASAP7_75t_R _29227_ (.A(_12514_),
    .Y(_12515_));
 AO222x2_ASAP7_75t_R _29228_ (.A1(_12469_),
    .A2(_12489_),
    .B1(_12493_),
    .B2(_12498_),
    .C1(_12512_),
    .C2(_12515_),
    .Y(_12516_));
 NAND2x1_ASAP7_75t_R _29229_ (.A(_01540_),
    .B(_11815_),
    .Y(_12517_));
 OA21x2_ASAP7_75t_R _29230_ (.A1(_12366_),
    .A2(_12516_),
    .B(_12517_),
    .Y(_04094_));
 BUFx6f_ASAP7_75t_R _29231_ (.A(_11805_),
    .Y(_12518_));
 OA21x2_ASAP7_75t_R _29232_ (.A1(_05533_),
    .A2(_05531_),
    .B(_05710_),
    .Y(_12519_));
 OAI21x1_ASAP7_75t_R _29233_ (.A1(_07348_),
    .A2(_12519_),
    .B(_05535_),
    .Y(_12520_));
 INVx1_ASAP7_75t_R _29234_ (.A(_01693_),
    .Y(_12521_));
 NOR2x1_ASAP7_75t_R _29235_ (.A(_01692_),
    .B(_05536_),
    .Y(_12522_));
 OR4x1_ASAP7_75t_R _29236_ (.A(_07348_),
    .B(_05710_),
    .C(_12521_),
    .D(_12522_),
    .Y(_12523_));
 AND3x4_ASAP7_75t_R _29237_ (.A(_11865_),
    .B(_12520_),
    .C(_12523_),
    .Y(_12524_));
 AO21x1_ASAP7_75t_R _29238_ (.A1(_05152_),
    .A2(_12518_),
    .B(_12524_),
    .Y(_04095_));
 BUFx6f_ASAP7_75t_R _29239_ (.A(_11865_),
    .Y(_12525_));
 OR3x1_ASAP7_75t_R _29240_ (.A(_11742_),
    .B(_05533_),
    .C(_11724_),
    .Y(_12526_));
 OA21x2_ASAP7_75t_R _29241_ (.A1(_05710_),
    .A2(_01692_),
    .B(_12526_),
    .Y(_12527_));
 OR4x1_ASAP7_75t_R _29242_ (.A(_07348_),
    .B(_12521_),
    .C(_11840_),
    .D(_12527_),
    .Y(_12528_));
 OAI21x1_ASAP7_75t_R _29243_ (.A1(_07790_),
    .A2(_12525_),
    .B(_12528_),
    .Y(_04096_));
 BUFx6f_ASAP7_75t_R _29244_ (.A(_12513_),
    .Y(_12529_));
 BUFx6f_ASAP7_75t_R _29245_ (.A(_12487_),
    .Y(_12530_));
 AND2x4_ASAP7_75t_R _29246_ (.A(_12529_),
    .B(_12530_),
    .Y(_12531_));
 NAND2x1_ASAP7_75t_R _29247_ (.A(_11785_),
    .B(_12531_),
    .Y(_12532_));
 OA21x2_ASAP7_75t_R _29248_ (.A1(_07774_),
    .A2(_12525_),
    .B(_12532_),
    .Y(_04097_));
 NAND2x1_ASAP7_75t_R _29249_ (.A(_01537_),
    .B(_11815_),
    .Y(_12533_));
 OA21x2_ASAP7_75t_R _29250_ (.A1(_12366_),
    .A2(_12529_),
    .B(_12533_),
    .Y(_04098_));
 NAND2x1_ASAP7_75t_R _29251_ (.A(_01536_),
    .B(_11815_),
    .Y(_12534_));
 OA21x2_ASAP7_75t_R _29252_ (.A1(_12366_),
    .A2(_12504_),
    .B(_12534_),
    .Y(_04099_));
 NAND2x1_ASAP7_75t_R _29253_ (.A(_01535_),
    .B(_11815_),
    .Y(_12535_));
 OA21x2_ASAP7_75t_R _29254_ (.A1(_12366_),
    .A2(_12502_),
    .B(_12535_),
    .Y(_04100_));
 NAND2x1_ASAP7_75t_R _29255_ (.A(_01534_),
    .B(_11815_),
    .Y(_12536_));
 OA21x2_ASAP7_75t_R _29256_ (.A1(_12366_),
    .A2(_12471_),
    .B(_12536_),
    .Y(_04101_));
 NAND2x1_ASAP7_75t_R _29257_ (.A(_01533_),
    .B(_11815_),
    .Y(_12537_));
 OA21x2_ASAP7_75t_R _29258_ (.A1(_12366_),
    .A2(_12509_),
    .B(_12537_),
    .Y(_04102_));
 NAND2x1_ASAP7_75t_R _29259_ (.A(_01532_),
    .B(_11815_),
    .Y(_12538_));
 OA21x2_ASAP7_75t_R _29260_ (.A1(_12366_),
    .A2(_12383_),
    .B(_12538_),
    .Y(_04103_));
 NAND2x1_ASAP7_75t_R _29261_ (.A(_01531_),
    .B(_11815_),
    .Y(_12539_));
 OA21x2_ASAP7_75t_R _29262_ (.A1(_12366_),
    .A2(_12375_),
    .B(_12539_),
    .Y(_04104_));
 BUFx12f_ASAP7_75t_R _29263_ (.A(_11805_),
    .Y(_12540_));
 NAND2x1_ASAP7_75t_R _29264_ (.A(_01530_),
    .B(_12540_),
    .Y(_12541_));
 OA21x2_ASAP7_75t_R _29265_ (.A1(_12366_),
    .A2(_12530_),
    .B(_12541_),
    .Y(_04105_));
 BUFx6f_ASAP7_75t_R _29266_ (.A(_12422_),
    .Y(_12542_));
 NAND2x1_ASAP7_75t_R _29267_ (.A(_01529_),
    .B(_12540_),
    .Y(_12543_));
 OA21x2_ASAP7_75t_R _29268_ (.A1(_12366_),
    .A2(_12542_),
    .B(_12543_),
    .Y(_04106_));
 BUFx6f_ASAP7_75t_R _29269_ (.A(_12397_),
    .Y(_12544_));
 NAND2x1_ASAP7_75t_R _29270_ (.A(_01528_),
    .B(_12540_),
    .Y(_12545_));
 OA21x2_ASAP7_75t_R _29271_ (.A1(_12518_),
    .A2(_12544_),
    .B(_12545_),
    .Y(_04107_));
 BUFx6f_ASAP7_75t_R _29272_ (.A(_12416_),
    .Y(_12546_));
 NAND2x1_ASAP7_75t_R _29273_ (.A(_01527_),
    .B(_12540_),
    .Y(_12547_));
 OA21x2_ASAP7_75t_R _29274_ (.A1(_12518_),
    .A2(_12546_),
    .B(_12547_),
    .Y(_04108_));
 BUFx6f_ASAP7_75t_R _29275_ (.A(_12409_),
    .Y(_12548_));
 NAND2x1_ASAP7_75t_R _29276_ (.A(_01526_),
    .B(_12540_),
    .Y(_12549_));
 OA21x2_ASAP7_75t_R _29277_ (.A1(_12518_),
    .A2(_12548_),
    .B(_12549_),
    .Y(_04109_));
 BUFx6f_ASAP7_75t_R _29278_ (.A(_12403_),
    .Y(_12550_));
 NAND2x1_ASAP7_75t_R _29279_ (.A(_01525_),
    .B(_12540_),
    .Y(_12551_));
 OA21x2_ASAP7_75t_R _29280_ (.A1(_12518_),
    .A2(_12550_),
    .B(_12551_),
    .Y(_04110_));
 BUFx6f_ASAP7_75t_R _29281_ (.A(_12455_),
    .Y(_12552_));
 NAND2x1_ASAP7_75t_R _29282_ (.A(_01524_),
    .B(_12540_),
    .Y(_12553_));
 OA21x2_ASAP7_75t_R _29283_ (.A1(_12518_),
    .A2(_12552_),
    .B(_12553_),
    .Y(_04111_));
 NAND2x1_ASAP7_75t_R _29284_ (.A(_01523_),
    .B(_12540_),
    .Y(_12554_));
 OA21x2_ASAP7_75t_R _29285_ (.A1(_12518_),
    .A2(_12431_),
    .B(_12554_),
    .Y(_04112_));
 BUFx6f_ASAP7_75t_R _29286_ (.A(_12449_),
    .Y(_12555_));
 NAND2x1_ASAP7_75t_R _29287_ (.A(_01522_),
    .B(_12540_),
    .Y(_12556_));
 OA21x2_ASAP7_75t_R _29288_ (.A1(_12518_),
    .A2(_12555_),
    .B(_12556_),
    .Y(_04113_));
 BUFx12f_ASAP7_75t_R _29289_ (.A(_11832_),
    .Y(_12557_));
 BUFx6f_ASAP7_75t_R _29290_ (.A(_11784_),
    .Y(_12558_));
 BUFx6f_ASAP7_75t_R _29291_ (.A(_12480_),
    .Y(_12559_));
 BUFx6f_ASAP7_75t_R _29292_ (.A(_12559_),
    .Y(_12560_));
 AND2x4_ASAP7_75t_R _29293_ (.A(_12500_),
    .B(_12491_),
    .Y(_12561_));
 AO21x1_ASAP7_75t_R _29294_ (.A1(_12375_),
    .A2(_12561_),
    .B(_12509_),
    .Y(_12562_));
 AND3x1_ASAP7_75t_R _29295_ (.A(_12558_),
    .B(_12560_),
    .C(_12562_),
    .Y(_12563_));
 AOI21x1_ASAP7_75t_R _29296_ (.A1(_13238_),
    .A2(_12557_),
    .B(_12563_),
    .Y(_04114_));
 OR3x2_ASAP7_75t_R _29297_ (.A(_12494_),
    .B(_12382_),
    .C(_12472_),
    .Y(_12564_));
 NOR2x1_ASAP7_75t_R _29298_ (.A(_12424_),
    .B(_12564_),
    .Y(_12565_));
 BUFx6f_ASAP7_75t_R _29299_ (.A(_12500_),
    .Y(_12566_));
 BUFx6f_ASAP7_75t_R _29300_ (.A(_12491_),
    .Y(_12567_));
 BUFx6f_ASAP7_75t_R _29301_ (.A(_12567_),
    .Y(_12568_));
 AOI21x1_ASAP7_75t_R _29302_ (.A1(_11742_),
    .A2(_12439_),
    .B(_12442_),
    .Y(_12569_));
 AO21x1_ASAP7_75t_R _29303_ (.A1(_12566_),
    .A2(_12568_),
    .B(_12569_),
    .Y(_12570_));
 AO21x1_ASAP7_75t_R _29304_ (.A1(_12568_),
    .A2(_12496_),
    .B(_12504_),
    .Y(_12571_));
 AND2x4_ASAP7_75t_R _29305_ (.A(_12373_),
    .B(_12500_),
    .Y(_12572_));
 AO21x1_ASAP7_75t_R _29306_ (.A1(_12572_),
    .A2(_12515_),
    .B(_12504_),
    .Y(_12573_));
 AOI22x1_ASAP7_75t_R _29307_ (.A1(_12560_),
    .A2(_12571_),
    .B1(_12573_),
    .B2(_12467_),
    .Y(_12574_));
 AO221x1_ASAP7_75t_R _29308_ (.A1(_12488_),
    .A2(_12565_),
    .B1(_12570_),
    .B2(_12574_),
    .C(_11832_),
    .Y(_12575_));
 OAI21x1_ASAP7_75t_R _29309_ (.A1(_13685_),
    .A2(_12525_),
    .B(_12575_),
    .Y(_04115_));
 AND2x6_ASAP7_75t_R _29310_ (.A(_12502_),
    .B(_12443_),
    .Y(_12576_));
 NAND2x2_ASAP7_75t_R _29311_ (.A(_12391_),
    .B(_12576_),
    .Y(_12577_));
 AO21x1_ASAP7_75t_R _29312_ (.A1(_12374_),
    .A2(_12577_),
    .B(_12508_),
    .Y(_12578_));
 AND3x1_ASAP7_75t_R _29313_ (.A(_12566_),
    .B(_12529_),
    .C(_12578_),
    .Y(_12579_));
 AO21x1_ASAP7_75t_R _29314_ (.A1(_12560_),
    .A2(_12496_),
    .B(_12579_),
    .Y(_12580_));
 OR3x1_ASAP7_75t_R _29315_ (.A(_12424_),
    .B(_12529_),
    .C(_12564_),
    .Y(_12581_));
 NOR2x1_ASAP7_75t_R _29316_ (.A(_12568_),
    .B(_12581_),
    .Y(_12582_));
 AO21x1_ASAP7_75t_R _29317_ (.A1(_12568_),
    .A2(_12580_),
    .B(_12582_),
    .Y(_12583_));
 OR3x1_ASAP7_75t_R _29318_ (.A(_11832_),
    .B(_12503_),
    .C(_12583_),
    .Y(_12584_));
 OAI21x1_ASAP7_75t_R _29319_ (.A1(_07799_),
    .A2(_12525_),
    .B(_12584_),
    .Y(_04116_));
 AND2x4_ASAP7_75t_R _29320_ (.A(_12473_),
    .B(_12514_),
    .Y(_12585_));
 BUFx6f_ASAP7_75t_R _29321_ (.A(_12585_),
    .Y(_12586_));
 AND2x6_ASAP7_75t_R _29322_ (.A(_12372_),
    .B(_12381_),
    .Y(_12587_));
 AO21x1_ASAP7_75t_R _29323_ (.A1(_12500_),
    .A2(_12391_),
    .B(_12587_),
    .Y(_12588_));
 NAND2x1_ASAP7_75t_R _29324_ (.A(_12502_),
    .B(_12504_),
    .Y(_12589_));
 AO21x1_ASAP7_75t_R _29325_ (.A1(_12550_),
    .A2(_12409_),
    .B(_12589_),
    .Y(_12590_));
 AO21x1_ASAP7_75t_R _29326_ (.A1(_12466_),
    .A2(_12590_),
    .B(_12470_),
    .Y(_12591_));
 AOI21x1_ASAP7_75t_R _29327_ (.A1(_11725_),
    .A2(_12427_),
    .B(_12430_),
    .Y(_12592_));
 OA211x2_ASAP7_75t_R _29328_ (.A1(_12592_),
    .A2(_12456_),
    .B(_12472_),
    .C(_12510_),
    .Y(_12593_));
 BUFx6f_ASAP7_75t_R _29329_ (.A(_12593_),
    .Y(_12594_));
 AO222x2_ASAP7_75t_R _29330_ (.A1(_12508_),
    .A2(_12588_),
    .B1(_12591_),
    .B2(_12572_),
    .C1(_12594_),
    .C2(_12542_),
    .Y(_12595_));
 AND3x1_ASAP7_75t_R _29331_ (.A(_12373_),
    .B(_12391_),
    .C(_12491_),
    .Y(_12596_));
 AO21x1_ASAP7_75t_R _29332_ (.A1(_12487_),
    .A2(_12496_),
    .B(_12596_),
    .Y(_12597_));
 AO22x1_ASAP7_75t_R _29333_ (.A1(_12471_),
    .A2(_12509_),
    .B1(_12597_),
    .B2(_12566_),
    .Y(_12598_));
 AO222x2_ASAP7_75t_R _29334_ (.A1(_12471_),
    .A2(_12531_),
    .B1(_12586_),
    .B2(_12595_),
    .C1(_12598_),
    .C2(_12560_),
    .Y(_12599_));
 OR3x1_ASAP7_75t_R _29335_ (.A(_11846_),
    .B(_11847_),
    .C(_12599_),
    .Y(_12600_));
 OA21x2_ASAP7_75t_R _29336_ (.A1(_14117_),
    .A2(_12525_),
    .B(_12600_),
    .Y(_04117_));
 AND2x6_ASAP7_75t_R _29337_ (.A(_12499_),
    .B(_12472_),
    .Y(_12601_));
 AND3x4_ASAP7_75t_R _29338_ (.A(_12373_),
    .B(_12499_),
    .C(_12464_),
    .Y(_12602_));
 AND2x6_ASAP7_75t_R _29339_ (.A(_12502_),
    .B(_12602_),
    .Y(_12603_));
 AO21x1_ASAP7_75t_R _29340_ (.A1(_12506_),
    .A2(_12550_),
    .B(_12569_),
    .Y(_12604_));
 AO222x2_ASAP7_75t_R _29341_ (.A1(_12471_),
    .A2(_12601_),
    .B1(_12603_),
    .B2(_12604_),
    .C1(_12594_),
    .C2(_12544_),
    .Y(_12605_));
 AO21x1_ASAP7_75t_R _29342_ (.A1(_12383_),
    .A2(_12560_),
    .B(_12509_),
    .Y(_12606_));
 NAND2x1_ASAP7_75t_R _29343_ (.A(_12529_),
    .B(_12567_),
    .Y(_12607_));
 AO221x1_ASAP7_75t_R _29344_ (.A1(_12586_),
    .A2(_12605_),
    .B1(_12606_),
    .B2(_12607_),
    .C(_11840_),
    .Y(_12608_));
 OA21x2_ASAP7_75t_R _29345_ (.A1(_14274_),
    .A2(_12525_),
    .B(_12608_),
    .Y(_04118_));
 NAND2x2_ASAP7_75t_R _29346_ (.A(_12465_),
    .B(_12480_),
    .Y(_12609_));
 BUFx6f_ASAP7_75t_R _29347_ (.A(_12602_),
    .Y(_12610_));
 AO21x1_ASAP7_75t_R _29348_ (.A1(_12506_),
    .A2(_12410_),
    .B(_12589_),
    .Y(_12611_));
 AO222x2_ASAP7_75t_R _29349_ (.A1(_12470_),
    .A2(_12601_),
    .B1(_12610_),
    .B2(_12611_),
    .C1(_12594_),
    .C2(_12546_),
    .Y(_12612_));
 AO32x1_ASAP7_75t_R _29350_ (.A1(_12383_),
    .A2(_12607_),
    .A3(_12609_),
    .B1(_12612_),
    .B2(_12586_),
    .Y(_12613_));
 OR3x1_ASAP7_75t_R _29351_ (.A(_11846_),
    .B(_11847_),
    .C(_12613_),
    .Y(_12614_));
 OA21x2_ASAP7_75t_R _29352_ (.A1(_14541_),
    .A2(_12525_),
    .B(_12614_),
    .Y(_04119_));
 OR3x1_ASAP7_75t_R _29353_ (.A(_12383_),
    .B(_12470_),
    .C(_12466_),
    .Y(_12615_));
 AO21x1_ASAP7_75t_R _29354_ (.A1(_12455_),
    .A2(_12374_),
    .B(_12500_),
    .Y(_12616_));
 BUFx6f_ASAP7_75t_R _29355_ (.A(_12494_),
    .Y(_12617_));
 OA21x2_ASAP7_75t_R _29356_ (.A1(_12508_),
    .A2(_12576_),
    .B(_12391_),
    .Y(_12618_));
 OR3x1_ASAP7_75t_R _29357_ (.A(_12455_),
    .B(_12617_),
    .C(_12618_),
    .Y(_12619_));
 AO32x1_ASAP7_75t_R _29358_ (.A1(_12615_),
    .A2(_12616_),
    .A3(_12619_),
    .B1(_12594_),
    .B2(_12548_),
    .Y(_12620_));
 OA211x2_ASAP7_75t_R _29359_ (.A1(_12552_),
    .A2(_12474_),
    .B(_12515_),
    .C(_12620_),
    .Y(_12621_));
 NAND2x1_ASAP7_75t_R _29360_ (.A(_12506_),
    .B(_12424_),
    .Y(_12622_));
 OR2x6_ASAP7_75t_R _29361_ (.A(_12617_),
    .B(_12622_),
    .Y(_12623_));
 AND3x1_ASAP7_75t_R _29362_ (.A(_12566_),
    .B(_12530_),
    .C(_12623_),
    .Y(_12624_));
 AO21x1_ASAP7_75t_R _29363_ (.A1(_12383_),
    .A2(_12568_),
    .B(_12624_),
    .Y(_12625_));
 AND3x1_ASAP7_75t_R _29364_ (.A(_12552_),
    .B(_12467_),
    .C(_12559_),
    .Y(_12626_));
 AND2x6_ASAP7_75t_R _29365_ (.A(_12487_),
    .B(_12609_),
    .Y(_12627_));
 OA21x2_ASAP7_75t_R _29366_ (.A1(_12493_),
    .A2(_12627_),
    .B(_12375_),
    .Y(_12628_));
 AO21x1_ASAP7_75t_R _29367_ (.A1(_12625_),
    .A2(_12626_),
    .B(_12628_),
    .Y(_12629_));
 OR3x2_ASAP7_75t_R _29368_ (.A(_11832_),
    .B(_12621_),
    .C(_12629_),
    .Y(_12630_));
 OA21x2_ASAP7_75t_R _29369_ (.A1(_14363_),
    .A2(_12525_),
    .B(_12630_),
    .Y(_04120_));
 BUFx12f_ASAP7_75t_R _29370_ (.A(_11805_),
    .Y(_12631_));
 BUFx6f_ASAP7_75t_R _29371_ (.A(_12492_),
    .Y(_12632_));
 AND3x1_ASAP7_75t_R _29372_ (.A(_05525_),
    .B(_11910_),
    .C(_11911_),
    .Y(_12633_));
 NOR2x1_ASAP7_75t_R _29373_ (.A(_12475_),
    .B(_01657_),
    .Y(_12634_));
 OA21x2_ASAP7_75t_R _29374_ (.A1(_05528_),
    .A2(_12634_),
    .B(_05544_),
    .Y(_12635_));
 NOR2x1_ASAP7_75t_R _29375_ (.A(_12633_),
    .B(_12635_),
    .Y(_12636_));
 AO21x2_ASAP7_75t_R _29376_ (.A1(_12373_),
    .A2(_12500_),
    .B(_12472_),
    .Y(_12637_));
 AO32x1_ASAP7_75t_R _29377_ (.A1(_12592_),
    .A2(_12383_),
    .A3(_12467_),
    .B1(_12636_),
    .B2(_12637_),
    .Y(_12638_));
 NAND2x1_ASAP7_75t_R _29378_ (.A(_12431_),
    .B(_12623_),
    .Y(_12639_));
 AO32x1_ASAP7_75t_R _29379_ (.A1(_12559_),
    .A2(_12501_),
    .A3(_12639_),
    .B1(_12636_),
    .B2(_12509_),
    .Y(_12640_));
 NOR2x1_ASAP7_75t_R _29380_ (.A(_12592_),
    .B(_12456_),
    .Y(_12641_));
 AND3x4_ASAP7_75t_R _29381_ (.A(_12472_),
    .B(_12510_),
    .C(_12641_),
    .Y(_12642_));
 AO22x1_ASAP7_75t_R _29382_ (.A1(_12499_),
    .A2(_12390_),
    .B1(_12403_),
    .B2(_12510_),
    .Y(_12643_));
 AND3x1_ASAP7_75t_R _29383_ (.A(_12494_),
    .B(_12499_),
    .C(_12464_),
    .Y(_12644_));
 AO221x1_ASAP7_75t_R _29384_ (.A1(_12431_),
    .A2(_12587_),
    .B1(_12643_),
    .B2(_12472_),
    .C(_12644_),
    .Y(_12645_));
 NOR2x1_ASAP7_75t_R _29385_ (.A(_12642_),
    .B(_12645_),
    .Y(_12646_));
 BUFx6f_ASAP7_75t_R _29386_ (.A(_12644_),
    .Y(_12647_));
 AO21x1_ASAP7_75t_R _29387_ (.A1(_12577_),
    .A2(_12646_),
    .B(_12647_),
    .Y(_12648_));
 AND3x4_ASAP7_75t_R _29388_ (.A(_12502_),
    .B(_12443_),
    .C(_12390_),
    .Y(_12649_));
 AO21x1_ASAP7_75t_R _29389_ (.A1(_12649_),
    .A2(_12636_),
    .B(_12564_),
    .Y(_12650_));
 AO221x1_ASAP7_75t_R _29390_ (.A1(_12592_),
    .A2(_12648_),
    .B1(_12650_),
    .B2(_12646_),
    .C(_12487_),
    .Y(_12651_));
 OA211x2_ASAP7_75t_R _29391_ (.A1(_12567_),
    .A2(_12636_),
    .B(_12651_),
    .C(_12529_),
    .Y(_12652_));
 AO221x1_ASAP7_75t_R _29392_ (.A1(_12632_),
    .A2(_12638_),
    .B1(_12640_),
    .B2(_12530_),
    .C(_12652_),
    .Y(_12653_));
 NOR2x2_ASAP7_75t_R _29393_ (.A(_11832_),
    .B(_12653_),
    .Y(_12654_));
 AO21x1_ASAP7_75t_R _29394_ (.A1(_14286_),
    .A2(_12631_),
    .B(_12654_),
    .Y(_04121_));
 OR2x2_ASAP7_75t_R _29395_ (.A(_12555_),
    .B(_12474_),
    .Y(_12655_));
 AO21x1_ASAP7_75t_R _29396_ (.A1(_11742_),
    .A2(net125),
    .B(_05529_),
    .Y(_12656_));
 AND3x1_ASAP7_75t_R _29397_ (.A(_05526_),
    .B(_11949_),
    .C(_11950_),
    .Y(_12657_));
 AO21x2_ASAP7_75t_R _29398_ (.A1(_07348_),
    .A2(_12656_),
    .B(_12657_),
    .Y(_12658_));
 AND2x4_ASAP7_75t_R _29399_ (.A(_12602_),
    .B(_12649_),
    .Y(_12659_));
 AO21x1_ASAP7_75t_R _29400_ (.A1(_12610_),
    .A2(_12577_),
    .B(_12587_),
    .Y(_12660_));
 OR2x2_ASAP7_75t_R _29401_ (.A(_12601_),
    .B(_12594_),
    .Y(_12661_));
 AO21x2_ASAP7_75t_R _29402_ (.A1(_12391_),
    .A2(_12661_),
    .B(_12647_),
    .Y(_12662_));
 AO221x1_ASAP7_75t_R _29403_ (.A1(_12658_),
    .A2(_12659_),
    .B1(_12660_),
    .B2(_12555_),
    .C(_12662_),
    .Y(_12663_));
 AND2x4_ASAP7_75t_R _29404_ (.A(_12382_),
    .B(_12465_),
    .Y(_12664_));
 AO21x1_ASAP7_75t_R _29405_ (.A1(_12555_),
    .A2(_12622_),
    .B(_12617_),
    .Y(_12665_));
 AO22x1_ASAP7_75t_R _29406_ (.A1(_12508_),
    .A2(_12658_),
    .B1(_12665_),
    .B2(_12501_),
    .Y(_12666_));
 AO32x1_ASAP7_75t_R _29407_ (.A1(_12555_),
    .A2(_12664_),
    .A3(_12632_),
    .B1(_12666_),
    .B2(_12488_),
    .Y(_12667_));
 AO21x1_ASAP7_75t_R _29408_ (.A1(_12515_),
    .A2(_12663_),
    .B(_12667_),
    .Y(_12668_));
 BUFx6f_ASAP7_75t_R _29409_ (.A(_12637_),
    .Y(_12669_));
 AO21x1_ASAP7_75t_R _29410_ (.A1(_12632_),
    .A2(_12669_),
    .B(_12531_),
    .Y(_12670_));
 AO221x1_ASAP7_75t_R _29411_ (.A1(_12655_),
    .A2(_12668_),
    .B1(_12670_),
    .B2(_12658_),
    .C(_11840_),
    .Y(_12671_));
 OA21x2_ASAP7_75t_R _29412_ (.A1(_14307_),
    .A2(_12525_),
    .B(_12671_),
    .Y(_04122_));
 AND2x2_ASAP7_75t_R _29413_ (.A(_12475_),
    .B(net126),
    .Y(_12672_));
 AO21x1_ASAP7_75t_R _29414_ (.A1(_11747_),
    .A2(_12419_),
    .B(_12672_),
    .Y(_12673_));
 AND3x1_ASAP7_75t_R _29415_ (.A(_05525_),
    .B(_11985_),
    .C(_11986_),
    .Y(_12674_));
 AOI21x1_ASAP7_75t_R _29416_ (.A1(_07347_),
    .A2(_12673_),
    .B(_12674_),
    .Y(_12675_));
 INVx1_ASAP7_75t_R _29417_ (.A(_12675_),
    .Y(_12676_));
 OA21x2_ASAP7_75t_R _29418_ (.A1(_12577_),
    .A2(_12676_),
    .B(_12602_),
    .Y(_12677_));
 OR3x1_ASAP7_75t_R _29419_ (.A(_12587_),
    .B(_12662_),
    .C(_12677_),
    .Y(_12678_));
 OA211x2_ASAP7_75t_R _29420_ (.A1(_12504_),
    .A2(_12474_),
    .B(_12515_),
    .C(_12678_),
    .Y(_12679_));
 AND3x1_ASAP7_75t_R _29421_ (.A(_12504_),
    .B(_12501_),
    .C(_12623_),
    .Y(_12680_));
 OA21x2_ASAP7_75t_R _29422_ (.A1(_12567_),
    .A2(_12680_),
    .B(_12559_),
    .Y(_12681_));
 AO21x1_ASAP7_75t_R _29423_ (.A1(_12627_),
    .A2(_12676_),
    .B(_12681_),
    .Y(_12682_));
 OAI21x1_ASAP7_75t_R _29424_ (.A1(_12496_),
    .A2(_12675_),
    .B(_12493_),
    .Y(_12683_));
 OA211x2_ASAP7_75t_R _29425_ (.A1(_12679_),
    .A2(_12682_),
    .B(_12683_),
    .C(_11784_),
    .Y(_12684_));
 AO21x1_ASAP7_75t_R _29426_ (.A1(_14283_),
    .A2(_12631_),
    .B(_12684_),
    .Y(_04123_));
 NAND2x1_ASAP7_75t_R _29427_ (.A(_12503_),
    .B(_12647_),
    .Y(_12685_));
 AND2x2_ASAP7_75t_R _29428_ (.A(_11742_),
    .B(net127),
    .Y(_12686_));
 AO21x1_ASAP7_75t_R _29429_ (.A1(_11747_),
    .A2(_12394_),
    .B(_12686_),
    .Y(_12687_));
 AND3x1_ASAP7_75t_R _29430_ (.A(_05526_),
    .B(_12020_),
    .C(_12021_),
    .Y(_12688_));
 AO21x1_ASAP7_75t_R _29431_ (.A1(_07348_),
    .A2(_12687_),
    .B(_12688_),
    .Y(_12689_));
 AO221x1_ASAP7_75t_R _29432_ (.A1(_12603_),
    .A2(_12622_),
    .B1(_12689_),
    .B2(_12509_),
    .C(_12647_),
    .Y(_12690_));
 AO22x1_ASAP7_75t_R _29433_ (.A1(_12515_),
    .A2(_12662_),
    .B1(_12690_),
    .B2(_12488_),
    .Y(_12691_));
 OA21x2_ASAP7_75t_R _29434_ (.A1(_12487_),
    .A2(_12659_),
    .B(_12529_),
    .Y(_12692_));
 AO21x1_ASAP7_75t_R _29435_ (.A1(_12492_),
    .A2(_12637_),
    .B(_12692_),
    .Y(_12693_));
 AO221x1_ASAP7_75t_R _29436_ (.A1(_12685_),
    .A2(_12691_),
    .B1(_12693_),
    .B2(_12689_),
    .C(_11840_),
    .Y(_12694_));
 OA21x2_ASAP7_75t_R _29437_ (.A1(_14281_),
    .A2(_12525_),
    .B(_12694_),
    .Y(_04124_));
 AND3x1_ASAP7_75t_R _29438_ (.A(_12529_),
    .B(_12610_),
    .C(_12649_),
    .Y(_12695_));
 AO21x1_ASAP7_75t_R _29439_ (.A1(_12560_),
    .A2(_12669_),
    .B(_12695_),
    .Y(_12696_));
 AND3x1_ASAP7_75t_R _29440_ (.A(_12558_),
    .B(_12568_),
    .C(_12696_),
    .Y(_12697_));
 AOI21x1_ASAP7_75t_R _29441_ (.A1(_13237_),
    .A2(_12557_),
    .B(_12697_),
    .Y(_04125_));
 BUFx6f_ASAP7_75t_R _29442_ (.A(_11865_),
    .Y(_12698_));
 AND2x2_ASAP7_75t_R _29443_ (.A(_12475_),
    .B(net129),
    .Y(_12699_));
 AO21x1_ASAP7_75t_R _29444_ (.A1(_11747_),
    .A2(_12413_),
    .B(_12699_),
    .Y(_12700_));
 AND3x1_ASAP7_75t_R _29445_ (.A(_05525_),
    .B(_12058_),
    .C(_12059_),
    .Y(_12701_));
 AOI21x1_ASAP7_75t_R _29446_ (.A1(_07347_),
    .A2(_12700_),
    .B(_12701_),
    .Y(_12702_));
 INVx1_ASAP7_75t_R _29447_ (.A(_12702_),
    .Y(_12703_));
 AO22x1_ASAP7_75t_R _29448_ (.A1(_12542_),
    .A2(_12664_),
    .B1(_12703_),
    .B2(_12500_),
    .Y(_12704_));
 NOR2x1_ASAP7_75t_R _29449_ (.A(_12466_),
    .B(_12702_),
    .Y(_12705_));
 AO21x1_ASAP7_75t_R _29450_ (.A1(_12375_),
    .A2(_12704_),
    .B(_12705_),
    .Y(_12706_));
 AO22x1_ASAP7_75t_R _29451_ (.A1(_12531_),
    .A2(_12703_),
    .B1(_12706_),
    .B2(_12632_),
    .Y(_12707_));
 AND3x4_ASAP7_75t_R _29452_ (.A(_12617_),
    .B(_12382_),
    .C(_12465_),
    .Y(_12708_));
 AO21x1_ASAP7_75t_R _29453_ (.A1(_12602_),
    .A2(_12577_),
    .B(_12708_),
    .Y(_12709_));
 AO221x1_ASAP7_75t_R _29454_ (.A1(_12659_),
    .A2(_12703_),
    .B1(_12709_),
    .B2(_12542_),
    .C(_12662_),
    .Y(_12710_));
 OR3x2_ASAP7_75t_R _29455_ (.A(_12431_),
    .B(_12456_),
    .C(_12506_),
    .Y(_12711_));
 NOR2x1_ASAP7_75t_R _29456_ (.A(_12424_),
    .B(_12711_),
    .Y(_12712_));
 AO21x1_ASAP7_75t_R _29457_ (.A1(_12373_),
    .A2(_12422_),
    .B(_12499_),
    .Y(_12713_));
 OA211x2_ASAP7_75t_R _29458_ (.A1(_12422_),
    .A2(_12712_),
    .B(_12713_),
    .C(_12465_),
    .Y(_12714_));
 OA21x2_ASAP7_75t_R _29459_ (.A1(_12705_),
    .A2(_12714_),
    .B(_12488_),
    .Y(_12715_));
 AO21x1_ASAP7_75t_R _29460_ (.A1(_12515_),
    .A2(_12710_),
    .B(_12715_),
    .Y(_12716_));
 OA21x2_ASAP7_75t_R _29461_ (.A1(_12542_),
    .A2(_12474_),
    .B(_12716_),
    .Y(_12717_));
 OR3x2_ASAP7_75t_R _29462_ (.A(_11832_),
    .B(_12707_),
    .C(_12717_),
    .Y(_12718_));
 OA21x2_ASAP7_75t_R _29463_ (.A1(_16337_),
    .A2(_12698_),
    .B(_12718_),
    .Y(_04126_));
 AND2x2_ASAP7_75t_R _29464_ (.A(_12471_),
    .B(_12594_),
    .Y(_12719_));
 AND2x2_ASAP7_75t_R _29465_ (.A(_11742_),
    .B(net130),
    .Y(_12720_));
 AO21x1_ASAP7_75t_R _29466_ (.A1(_11747_),
    .A2(_12406_),
    .B(_12720_),
    .Y(_12721_));
 AND3x1_ASAP7_75t_R _29467_ (.A(_05526_),
    .B(_12095_),
    .C(_12096_),
    .Y(_12722_));
 AO21x1_ASAP7_75t_R _29468_ (.A1(_07348_),
    .A2(_12721_),
    .B(_12722_),
    .Y(_12723_));
 AO32x1_ASAP7_75t_R _29469_ (.A1(_12610_),
    .A2(_12649_),
    .A3(_12723_),
    .B1(_12709_),
    .B2(_12544_),
    .Y(_12724_));
 OA21x2_ASAP7_75t_R _29470_ (.A1(_12719_),
    .A2(_12724_),
    .B(_12586_),
    .Y(_12725_));
 AO32x1_ASAP7_75t_R _29471_ (.A1(_12375_),
    .A2(_12544_),
    .A3(_12664_),
    .B1(_12637_),
    .B2(_12723_),
    .Y(_12726_));
 NOR2x1_ASAP7_75t_R _29472_ (.A(_12510_),
    .B(_12609_),
    .Y(_12727_));
 AO22x1_ASAP7_75t_R _29473_ (.A1(_12609_),
    .A2(_12723_),
    .B1(_12727_),
    .B2(_12544_),
    .Y(_12728_));
 NAND2x1_ASAP7_75t_R _29474_ (.A(_12374_),
    .B(_12466_),
    .Y(_12729_));
 AND4x1_ASAP7_75t_R _29475_ (.A(_12544_),
    .B(_12529_),
    .C(_12729_),
    .D(_12561_),
    .Y(_12730_));
 AO221x1_ASAP7_75t_R _29476_ (.A1(_12632_),
    .A2(_12726_),
    .B1(_12728_),
    .B2(_12530_),
    .C(_12730_),
    .Y(_12731_));
 OR3x2_ASAP7_75t_R _29477_ (.A(_11840_),
    .B(_12725_),
    .C(_12731_),
    .Y(_12732_));
 OA21x2_ASAP7_75t_R _29478_ (.A1(_15436_),
    .A2(_12698_),
    .B(_12732_),
    .Y(_04127_));
 NAND2x1_ASAP7_75t_R _29479_ (.A(_12374_),
    .B(_12383_),
    .Y(_12733_));
 AND3x1_ASAP7_75t_R _29480_ (.A(_12466_),
    .B(_12559_),
    .C(_12487_),
    .Y(_12734_));
 AO32x1_ASAP7_75t_R _29481_ (.A1(_12566_),
    .A2(_12729_),
    .A3(_12515_),
    .B1(_12733_),
    .B2(_12734_),
    .Y(_12735_));
 NAND2x1_ASAP7_75t_R _29482_ (.A(_11747_),
    .B(_01650_),
    .Y(_12736_));
 OA211x2_ASAP7_75t_R _29483_ (.A1(_11747_),
    .A2(net131),
    .B(_12736_),
    .C(_07347_),
    .Y(_12737_));
 AO21x2_ASAP7_75t_R _29484_ (.A1(_05526_),
    .A2(_12119_),
    .B(_12737_),
    .Y(_12738_));
 AO32x1_ASAP7_75t_R _29485_ (.A1(_12550_),
    .A2(_12496_),
    .A3(_12632_),
    .B1(_12627_),
    .B2(_12738_),
    .Y(_12739_));
 AO21x1_ASAP7_75t_R _29486_ (.A1(_12546_),
    .A2(_12735_),
    .B(_12739_),
    .Y(_12740_));
 AND5x1_ASAP7_75t_R _29487_ (.A(_12374_),
    .B(_12383_),
    .C(_12546_),
    .D(_12466_),
    .E(_12488_),
    .Y(_12741_));
 AO32x1_ASAP7_75t_R _29488_ (.A1(_12546_),
    .A2(_12467_),
    .A3(_12587_),
    .B1(_12637_),
    .B2(_12738_),
    .Y(_12742_));
 OA21x2_ASAP7_75t_R _29489_ (.A1(_12632_),
    .A2(_12741_),
    .B(_12742_),
    .Y(_12743_));
 AO21x1_ASAP7_75t_R _29490_ (.A1(_12610_),
    .A2(_12577_),
    .B(_12495_),
    .Y(_12744_));
 AO32x1_ASAP7_75t_R _29491_ (.A1(_12610_),
    .A2(_12649_),
    .A3(_12738_),
    .B1(_12744_),
    .B2(_12546_),
    .Y(_12745_));
 OA21x2_ASAP7_75t_R _29492_ (.A1(_12719_),
    .A2(_12745_),
    .B(_12586_),
    .Y(_12746_));
 OR4x1_ASAP7_75t_R _29493_ (.A(_11805_),
    .B(_12740_),
    .C(_12743_),
    .D(_12746_),
    .Y(_12747_));
 OA21x2_ASAP7_75t_R _29494_ (.A1(_16218_),
    .A2(_12698_),
    .B(_12747_),
    .Y(_04128_));
 NAND2x1_ASAP7_75t_R _29495_ (.A(_11742_),
    .B(net132),
    .Y(_12748_));
 OR2x2_ASAP7_75t_R _29496_ (.A(_12475_),
    .B(_01649_),
    .Y(_12749_));
 AO21x1_ASAP7_75t_R _29497_ (.A1(_12748_),
    .A2(_12749_),
    .B(_05526_),
    .Y(_12750_));
 OA21x2_ASAP7_75t_R _29498_ (.A1(_07348_),
    .A2(_12134_),
    .B(_12750_),
    .Y(_12751_));
 NAND2x1_ASAP7_75t_R _29499_ (.A(_12470_),
    .B(_12751_),
    .Y(_12752_));
 AO21x1_ASAP7_75t_R _29500_ (.A1(_12610_),
    .A2(_12589_),
    .B(_12708_),
    .Y(_12753_));
 AO32x1_ASAP7_75t_R _29501_ (.A1(_12610_),
    .A2(_12576_),
    .A3(_12752_),
    .B1(_12753_),
    .B2(_12548_),
    .Y(_12754_));
 OA21x2_ASAP7_75t_R _29502_ (.A1(_12719_),
    .A2(_12754_),
    .B(_12586_),
    .Y(_12755_));
 INVx1_ASAP7_75t_R _29503_ (.A(_12751_),
    .Y(_12756_));
 NAND2x2_ASAP7_75t_R _29504_ (.A(_12480_),
    .B(_12567_),
    .Y(_12757_));
 AOI221x1_ASAP7_75t_R _29505_ (.A1(_12569_),
    .A2(_12708_),
    .B1(_12751_),
    .B2(_12637_),
    .C(_12757_),
    .Y(_12758_));
 AO32x1_ASAP7_75t_R _29506_ (.A1(_12530_),
    .A2(_12609_),
    .A3(_12756_),
    .B1(_12758_),
    .B2(_12474_),
    .Y(_12759_));
 AO32x1_ASAP7_75t_R _29507_ (.A1(_12566_),
    .A2(_12729_),
    .A3(_12514_),
    .B1(_12466_),
    .B2(_12488_),
    .Y(_12760_));
 OA21x2_ASAP7_75t_R _29508_ (.A1(_12758_),
    .A2(_12760_),
    .B(_12548_),
    .Y(_12761_));
 OR4x1_ASAP7_75t_R _29509_ (.A(_11805_),
    .B(_12755_),
    .C(_12759_),
    .D(_12761_),
    .Y(_12762_));
 OA21x2_ASAP7_75t_R _29510_ (.A1(_15588_),
    .A2(_12698_),
    .B(_12762_),
    .Y(_04129_));
 NAND2x1_ASAP7_75t_R _29511_ (.A(_05537_),
    .B(_01648_),
    .Y(_12763_));
 OA211x2_ASAP7_75t_R _29512_ (.A1(_11746_),
    .A2(net133),
    .B(_05544_),
    .C(_12763_),
    .Y(_12764_));
 AO21x2_ASAP7_75t_R _29513_ (.A1(_05525_),
    .A2(_12151_),
    .B(_12764_),
    .Y(_12765_));
 AND3x1_ASAP7_75t_R _29514_ (.A(_12390_),
    .B(_12576_),
    .C(_12765_),
    .Y(_12766_));
 AO21x1_ASAP7_75t_R _29515_ (.A1(_12403_),
    .A2(_12589_),
    .B(_12766_),
    .Y(_12767_));
 AO21x1_ASAP7_75t_R _29516_ (.A1(_12390_),
    .A2(_12594_),
    .B(_12647_),
    .Y(_12768_));
 AO221x1_ASAP7_75t_R _29517_ (.A1(_12502_),
    .A2(_12601_),
    .B1(_12602_),
    .B2(_12767_),
    .C(_12768_),
    .Y(_12769_));
 OR3x1_ASAP7_75t_R _29518_ (.A(_12642_),
    .B(_12708_),
    .C(_12769_),
    .Y(_12770_));
 AO21x1_ASAP7_75t_R _29519_ (.A1(_12474_),
    .A2(_12769_),
    .B(_12550_),
    .Y(_12771_));
 AO21x1_ASAP7_75t_R _29520_ (.A1(_12770_),
    .A2(_12771_),
    .B(_12530_),
    .Y(_12772_));
 OA21x2_ASAP7_75t_R _29521_ (.A1(_12568_),
    .A2(_12765_),
    .B(_12772_),
    .Y(_12773_));
 OA22x2_ASAP7_75t_R _29522_ (.A1(_12550_),
    .A2(_12609_),
    .B1(_12765_),
    .B2(_12467_),
    .Y(_12774_));
 AO221x1_ASAP7_75t_R _29523_ (.A1(_12502_),
    .A2(_12496_),
    .B1(_12637_),
    .B2(_12765_),
    .C(_12757_),
    .Y(_12775_));
 OA21x2_ASAP7_75t_R _29524_ (.A1(_12568_),
    .A2(_12774_),
    .B(_12775_),
    .Y(_12776_));
 OA211x2_ASAP7_75t_R _29525_ (.A1(_12560_),
    .A2(_12773_),
    .B(_12776_),
    .C(_11784_),
    .Y(_12777_));
 AO21x1_ASAP7_75t_R _29526_ (.A1(_15434_),
    .A2(_12631_),
    .B(_12777_),
    .Y(_04130_));
 AND2x2_ASAP7_75t_R _29527_ (.A(_11725_),
    .B(net134),
    .Y(_12778_));
 AO21x1_ASAP7_75t_R _29528_ (.A1(_11746_),
    .A2(_12446_),
    .B(_12778_),
    .Y(_12779_));
 AND3x1_ASAP7_75t_R _29529_ (.A(_05525_),
    .B(_12158_),
    .C(_12159_),
    .Y(_12780_));
 AOI21x1_ASAP7_75t_R _29530_ (.A1(_07347_),
    .A2(_12779_),
    .B(_12780_),
    .Y(_12781_));
 NAND2x1_ASAP7_75t_R _29531_ (.A(_12669_),
    .B(_12781_),
    .Y(_12782_));
 OA21x2_ASAP7_75t_R _29532_ (.A1(_12471_),
    .A2(_12669_),
    .B(_12782_),
    .Y(_12783_));
 OA21x2_ASAP7_75t_R _29533_ (.A1(_12470_),
    .A2(_12474_),
    .B(_12515_),
    .Y(_12784_));
 OR2x6_ASAP7_75t_R _29534_ (.A(_12587_),
    .B(_12601_),
    .Y(_12785_));
 OA21x2_ASAP7_75t_R _29535_ (.A1(_12785_),
    .A2(_12642_),
    .B(_12542_),
    .Y(_12786_));
 INVx1_ASAP7_75t_R _29536_ (.A(_12781_),
    .Y(_12787_));
 OA21x2_ASAP7_75t_R _29537_ (.A1(_12569_),
    .A2(_12787_),
    .B(_12603_),
    .Y(_12788_));
 OA21x2_ASAP7_75t_R _29538_ (.A1(_12496_),
    .A2(_12788_),
    .B(_12470_),
    .Y(_12789_));
 OR3x1_ASAP7_75t_R _29539_ (.A(_12768_),
    .B(_12786_),
    .C(_12789_),
    .Y(_12790_));
 AND2x4_ASAP7_75t_R _29540_ (.A(_12382_),
    .B(_12390_),
    .Y(_12791_));
 AO21x1_ASAP7_75t_R _29541_ (.A1(_12466_),
    .A2(_12791_),
    .B(_12567_),
    .Y(_12792_));
 AO32x1_ASAP7_75t_R _29542_ (.A1(_12607_),
    .A2(_12609_),
    .A3(_12787_),
    .B1(_12792_),
    .B2(_12559_),
    .Y(_12793_));
 AO21x1_ASAP7_75t_R _29543_ (.A1(_12784_),
    .A2(_12790_),
    .B(_12793_),
    .Y(_12794_));
 OA211x2_ASAP7_75t_R _29544_ (.A1(_12757_),
    .A2(_12783_),
    .B(_12794_),
    .C(_11784_),
    .Y(_12795_));
 AO21x1_ASAP7_75t_R _29545_ (.A1(_13832_),
    .A2(_12631_),
    .B(_12795_),
    .Y(_04131_));
 AO21x1_ASAP7_75t_R _29546_ (.A1(_12548_),
    .A2(_12587_),
    .B(_12647_),
    .Y(_12796_));
 AND2x2_ASAP7_75t_R _29547_ (.A(_12475_),
    .B(net135),
    .Y(_12797_));
 AO21x1_ASAP7_75t_R _29548_ (.A1(_11746_),
    .A2(_12440_),
    .B(_12797_),
    .Y(_12798_));
 AND3x1_ASAP7_75t_R _29549_ (.A(_05525_),
    .B(_11913_),
    .C(_11914_),
    .Y(_12799_));
 AO21x1_ASAP7_75t_R _29550_ (.A1(_07347_),
    .A2(_12798_),
    .B(_12799_),
    .Y(_12800_));
 OA21x2_ASAP7_75t_R _29551_ (.A1(_12569_),
    .A2(_12800_),
    .B(_12603_),
    .Y(_12801_));
 OR3x1_ASAP7_75t_R _29552_ (.A(_12594_),
    .B(_12708_),
    .C(_12801_),
    .Y(_12802_));
 AND3x1_ASAP7_75t_R _29553_ (.A(_12382_),
    .B(_12548_),
    .C(_12641_),
    .Y(_12803_));
 AO21x1_ASAP7_75t_R _29554_ (.A1(_12552_),
    .A2(_12500_),
    .B(_12803_),
    .Y(_12804_));
 AO22x1_ASAP7_75t_R _29555_ (.A1(_12471_),
    .A2(_12802_),
    .B1(_12804_),
    .B2(_12509_),
    .Y(_12805_));
 OA21x2_ASAP7_75t_R _29556_ (.A1(_12796_),
    .A2(_12805_),
    .B(_12784_),
    .Y(_12806_));
 AND2x2_ASAP7_75t_R _29557_ (.A(_12455_),
    .B(_12374_),
    .Y(_12807_));
 AO21x1_ASAP7_75t_R _29558_ (.A1(_12617_),
    .A2(_12542_),
    .B(_12807_),
    .Y(_12808_));
 AND3x1_ASAP7_75t_R _29559_ (.A(_12488_),
    .B(_12664_),
    .C(_12808_),
    .Y(_12809_));
 OA21x2_ASAP7_75t_R _29560_ (.A1(_12548_),
    .A2(_12490_),
    .B(_12492_),
    .Y(_12810_));
 OA21x2_ASAP7_75t_R _29561_ (.A1(_12552_),
    .A2(_12473_),
    .B(_12810_),
    .Y(_12811_));
 NOR2x1_ASAP7_75t_R _29562_ (.A(_12508_),
    .B(_12572_),
    .Y(_12812_));
 AO21x1_ASAP7_75t_R _29563_ (.A1(_12812_),
    .A2(_12811_),
    .B(_12800_),
    .Y(_12813_));
 OA21x2_ASAP7_75t_R _29564_ (.A1(_12627_),
    .A2(_12811_),
    .B(_12813_),
    .Y(_12814_));
 OR4x1_ASAP7_75t_R _29565_ (.A(_11805_),
    .B(_12806_),
    .C(_12809_),
    .D(_12814_),
    .Y(_12815_));
 OA21x2_ASAP7_75t_R _29566_ (.A1(_13838_),
    .A2(_12698_),
    .B(_12815_),
    .Y(_04132_));
 AND2x2_ASAP7_75t_R _29567_ (.A(_12475_),
    .B(net136),
    .Y(_12816_));
 AO21x1_ASAP7_75t_R _29568_ (.A1(_11746_),
    .A2(_12434_),
    .B(_12816_),
    .Y(_12817_));
 AND3x1_ASAP7_75t_R _29569_ (.A(_05525_),
    .B(_11916_),
    .C(_11917_),
    .Y(_12818_));
 AOI21x1_ASAP7_75t_R _29570_ (.A1(_07347_),
    .A2(_12817_),
    .B(_12818_),
    .Y(_12819_));
 INVx2_ASAP7_75t_R _29571_ (.A(_12819_),
    .Y(_12820_));
 AO221x1_ASAP7_75t_R _29572_ (.A1(_12431_),
    .A2(_12647_),
    .B1(_12669_),
    .B2(_12820_),
    .C(_12757_),
    .Y(_12821_));
 OA21x2_ASAP7_75t_R _29573_ (.A1(_12569_),
    .A2(_12820_),
    .B(_12603_),
    .Y(_12822_));
 OR3x1_ASAP7_75t_R _29574_ (.A(_12594_),
    .B(_12708_),
    .C(_12822_),
    .Y(_12823_));
 AO221x1_ASAP7_75t_R _29575_ (.A1(_12550_),
    .A2(_12785_),
    .B1(_12642_),
    .B2(_12544_),
    .C(_12647_),
    .Y(_12824_));
 AO21x1_ASAP7_75t_R _29576_ (.A1(_12471_),
    .A2(_12823_),
    .B(_12824_),
    .Y(_12825_));
 AND2x2_ASAP7_75t_R _29577_ (.A(_12431_),
    .B(_12373_),
    .Y(_12826_));
 AO21x1_ASAP7_75t_R _29578_ (.A1(_12617_),
    .A2(_12397_),
    .B(_12826_),
    .Y(_12827_));
 AO21x1_ASAP7_75t_R _29579_ (.A1(_12664_),
    .A2(_12827_),
    .B(_12567_),
    .Y(_12828_));
 AO32x1_ASAP7_75t_R _29580_ (.A1(_12607_),
    .A2(_12609_),
    .A3(_12820_),
    .B1(_12828_),
    .B2(_12559_),
    .Y(_12829_));
 AO21x1_ASAP7_75t_R _29581_ (.A1(_12784_),
    .A2(_12825_),
    .B(_12829_),
    .Y(_12830_));
 AND3x4_ASAP7_75t_R _29582_ (.A(_11865_),
    .B(_12821_),
    .C(_12830_),
    .Y(_12831_));
 AO21x1_ASAP7_75t_R _29583_ (.A1(_13910_),
    .A2(_12631_),
    .B(_12831_),
    .Y(_04133_));
 AND2x2_ASAP7_75t_R _29584_ (.A(_12475_),
    .B(net137),
    .Y(_12832_));
 AO21x1_ASAP7_75t_R _29585_ (.A1(_11746_),
    .A2(_12387_),
    .B(_12832_),
    .Y(_12833_));
 AND3x1_ASAP7_75t_R _29586_ (.A(_05525_),
    .B(_11919_),
    .C(_11920_),
    .Y(_12834_));
 AO21x2_ASAP7_75t_R _29587_ (.A1(_07347_),
    .A2(_12833_),
    .B(_12834_),
    .Y(_12835_));
 AO221x1_ASAP7_75t_R _29588_ (.A1(_12555_),
    .A2(_12647_),
    .B1(_12669_),
    .B2(_12835_),
    .C(_12757_),
    .Y(_12836_));
 OA21x2_ASAP7_75t_R _29589_ (.A1(_12373_),
    .A2(_12465_),
    .B(_12791_),
    .Y(_12837_));
 AO21x1_ASAP7_75t_R _29590_ (.A1(_12555_),
    .A2(_12601_),
    .B(_12837_),
    .Y(_12838_));
 OA211x2_ASAP7_75t_R _29591_ (.A1(_12569_),
    .A2(_12835_),
    .B(_12603_),
    .C(_12391_),
    .Y(_12839_));
 AND2x2_ASAP7_75t_R _29592_ (.A(_12416_),
    .B(_12642_),
    .Y(_12840_));
 OR4x1_ASAP7_75t_R _29593_ (.A(_12768_),
    .B(_12838_),
    .C(_12839_),
    .D(_12840_),
    .Y(_12841_));
 AO221x1_ASAP7_75t_R _29594_ (.A1(_12627_),
    .A2(_12835_),
    .B1(_12841_),
    .B2(_12784_),
    .C(_12632_),
    .Y(_12842_));
 AND3x4_ASAP7_75t_R _29595_ (.A(_11865_),
    .B(_12836_),
    .C(_12842_),
    .Y(_12843_));
 AO21x1_ASAP7_75t_R _29596_ (.A1(_13970_),
    .A2(_12631_),
    .B(_12843_),
    .Y(_04134_));
 AND2x2_ASAP7_75t_R _29597_ (.A(_11725_),
    .B(net138),
    .Y(_12844_));
 AO21x1_ASAP7_75t_R _29598_ (.A1(_11746_),
    .A2(_12461_),
    .B(_12844_),
    .Y(_12845_));
 AND3x1_ASAP7_75t_R _29599_ (.A(_05525_),
    .B(_11922_),
    .C(_11923_),
    .Y(_12846_));
 AO21x2_ASAP7_75t_R _29600_ (.A1(_07347_),
    .A2(_12845_),
    .B(_12846_),
    .Y(_12847_));
 AO221x1_ASAP7_75t_R _29601_ (.A1(_12504_),
    .A2(_12647_),
    .B1(_12669_),
    .B2(_12847_),
    .C(_12757_),
    .Y(_12848_));
 OA21x2_ASAP7_75t_R _29602_ (.A1(_12569_),
    .A2(_12847_),
    .B(_12603_),
    .Y(_12849_));
 OR3x1_ASAP7_75t_R _29603_ (.A(_12382_),
    .B(_12495_),
    .C(_12849_),
    .Y(_12850_));
 AO32x1_ASAP7_75t_R _29604_ (.A1(_12504_),
    .A2(_12566_),
    .A3(_12509_),
    .B1(_12850_),
    .B2(_12470_),
    .Y(_12851_));
 AO221x1_ASAP7_75t_R _29605_ (.A1(_12627_),
    .A2(_12847_),
    .B1(_12851_),
    .B2(_12515_),
    .C(_12632_),
    .Y(_12852_));
 AND3x1_ASAP7_75t_R _29606_ (.A(_11865_),
    .B(_12848_),
    .C(_12852_),
    .Y(_12853_));
 AO21x1_ASAP7_75t_R _29607_ (.A1(_14027_),
    .A2(_12631_),
    .B(_12853_),
    .Y(_04135_));
 AO32x1_ASAP7_75t_R _29608_ (.A1(_12507_),
    .A2(_12610_),
    .A3(_12711_),
    .B1(_12508_),
    .B2(_12542_),
    .Y(_12854_));
 AO32x1_ASAP7_75t_R _29609_ (.A1(_12488_),
    .A2(_12474_),
    .A3(_12854_),
    .B1(_12693_),
    .B2(_12542_),
    .Y(_12855_));
 AO21x1_ASAP7_75t_R _29610_ (.A1(_12586_),
    .A2(_12661_),
    .B(_12855_),
    .Y(_12856_));
 OR3x2_ASAP7_75t_R _29611_ (.A(_11846_),
    .B(_11847_),
    .C(_12856_),
    .Y(_12857_));
 OA21x2_ASAP7_75t_R _29612_ (.A1(_14124_),
    .A2(_12698_),
    .B(_12857_),
    .Y(_04136_));
 OA21x2_ASAP7_75t_R _29613_ (.A1(_12391_),
    .A2(_12410_),
    .B(_12502_),
    .Y(_12858_));
 NOR2x1_ASAP7_75t_R _29614_ (.A(_12569_),
    .B(_12858_),
    .Y(_12859_));
 NAND2x1_ASAP7_75t_R _29615_ (.A(_11746_),
    .B(_01641_),
    .Y(_12860_));
 OA211x2_ASAP7_75t_R _29616_ (.A1(_11747_),
    .A2(net140),
    .B(_12860_),
    .C(_07347_),
    .Y(_12861_));
 AO21x2_ASAP7_75t_R _29617_ (.A1(_05526_),
    .A2(_11928_),
    .B(_12861_),
    .Y(_12862_));
 OA211x2_ASAP7_75t_R _29618_ (.A1(_12569_),
    .A2(_12862_),
    .B(_12470_),
    .C(_12502_),
    .Y(_12863_));
 OR3x1_ASAP7_75t_R _29619_ (.A(_12729_),
    .B(_12859_),
    .C(_12863_),
    .Y(_12864_));
 OA21x2_ASAP7_75t_R _29620_ (.A1(_12431_),
    .A2(_12467_),
    .B(_12566_),
    .Y(_12865_));
 AO21x1_ASAP7_75t_R _29621_ (.A1(_12864_),
    .A2(_12865_),
    .B(_12791_),
    .Y(_12866_));
 AOI21x1_ASAP7_75t_R _29622_ (.A1(_12632_),
    .A2(_12637_),
    .B(_12627_),
    .Y(_12867_));
 INVx1_ASAP7_75t_R _29623_ (.A(_12867_),
    .Y(_12868_));
 AO221x1_ASAP7_75t_R _29624_ (.A1(_12784_),
    .A2(_12866_),
    .B1(_12868_),
    .B2(_12862_),
    .C(_11840_),
    .Y(_12869_));
 OA21x2_ASAP7_75t_R _29625_ (.A1(_14202_),
    .A2(_12698_),
    .B(_12869_),
    .Y(_04137_));
 AND2x2_ASAP7_75t_R _29626_ (.A(_11742_),
    .B(net141),
    .Y(_12870_));
 AO21x1_ASAP7_75t_R _29627_ (.A1(_11747_),
    .A2(_12369_),
    .B(_12870_),
    .Y(_12871_));
 AND3x1_ASAP7_75t_R _29628_ (.A(_05526_),
    .B(_11930_),
    .C(_11931_),
    .Y(_12872_));
 AOI21x1_ASAP7_75t_R _29629_ (.A1(_07348_),
    .A2(_12871_),
    .B(_12872_),
    .Y(_12873_));
 AO21x1_ASAP7_75t_R _29630_ (.A1(_12504_),
    .A2(_12873_),
    .B(_12503_),
    .Y(_12874_));
 OR3x1_ASAP7_75t_R _29631_ (.A(_12506_),
    .B(_12559_),
    .C(_12530_),
    .Y(_12875_));
 AO21x1_ASAP7_75t_R _29632_ (.A1(_12610_),
    .A2(_12874_),
    .B(_12875_),
    .Y(_12876_));
 OA211x2_ASAP7_75t_R _29633_ (.A1(_12867_),
    .A2(_12873_),
    .B(_12876_),
    .C(_11865_),
    .Y(_12877_));
 AOI21x1_ASAP7_75t_R _29634_ (.A1(_14099_),
    .A2(_12557_),
    .B(_12877_),
    .Y(_04138_));
 AO21x1_ASAP7_75t_R _29635_ (.A1(_12586_),
    .A2(_12659_),
    .B(_12868_),
    .Y(_12878_));
 AO221x1_ASAP7_75t_R _29636_ (.A1(_12601_),
    .A2(_12586_),
    .B1(_12878_),
    .B2(_12544_),
    .C(_11840_),
    .Y(_12879_));
 OA21x2_ASAP7_75t_R _29637_ (.A1(_13230_),
    .A2(_12698_),
    .B(_12879_),
    .Y(_04139_));
 INVx1_ASAP7_75t_R _29638_ (.A(_12546_),
    .Y(_12880_));
 AND3x1_ASAP7_75t_R _29639_ (.A(_12375_),
    .B(_12880_),
    .C(_12649_),
    .Y(_12881_));
 OR3x1_ASAP7_75t_R _29640_ (.A(_12607_),
    .B(_12785_),
    .C(_12881_),
    .Y(_12882_));
 NAND2x1_ASAP7_75t_R _29641_ (.A(_12617_),
    .B(_12467_),
    .Y(_12883_));
 AOI21x1_ASAP7_75t_R _29642_ (.A1(_12546_),
    .A2(_12627_),
    .B(_12493_),
    .Y(_12884_));
 AO21x1_ASAP7_75t_R _29643_ (.A1(_12880_),
    .A2(_12883_),
    .B(_12884_),
    .Y(_12885_));
 NAND2x1_ASAP7_75t_R _29644_ (.A(_12559_),
    .B(_12530_),
    .Y(_12886_));
 AND3x1_ASAP7_75t_R _29645_ (.A(_12375_),
    .B(_12507_),
    .C(_12711_),
    .Y(_12887_));
 OR4x1_ASAP7_75t_R _29646_ (.A(_12383_),
    .B(_12509_),
    .C(_12886_),
    .D(_12887_),
    .Y(_12888_));
 AND4x1_ASAP7_75t_R _29647_ (.A(_11865_),
    .B(_12882_),
    .C(_12885_),
    .D(_12888_),
    .Y(_12889_));
 AOI21x1_ASAP7_75t_R _29648_ (.A1(_13280_),
    .A2(_12557_),
    .B(_12889_),
    .Y(_04140_));
 OA211x2_ASAP7_75t_R _29649_ (.A1(_12506_),
    .A2(_12548_),
    .B(_12576_),
    .C(_12374_),
    .Y(_12890_));
 OR3x1_ASAP7_75t_R _29650_ (.A(_12785_),
    .B(_12594_),
    .C(_12890_),
    .Y(_12891_));
 AO21x1_ASAP7_75t_R _29651_ (.A1(_12548_),
    .A2(_12530_),
    .B(_12559_),
    .Y(_12892_));
 OA21x2_ASAP7_75t_R _29652_ (.A1(_12529_),
    .A2(_12883_),
    .B(_12892_),
    .Y(_12893_));
 INVx1_ASAP7_75t_R _29653_ (.A(_12561_),
    .Y(_12894_));
 AO21x1_ASAP7_75t_R _29654_ (.A1(_12467_),
    .A2(_12894_),
    .B(_12548_),
    .Y(_12895_));
 AO221x1_ASAP7_75t_R _29655_ (.A1(_12586_),
    .A2(_12891_),
    .B1(_12893_),
    .B2(_12895_),
    .C(_11840_),
    .Y(_12896_));
 OA21x2_ASAP7_75t_R _29656_ (.A1(_13243_),
    .A2(_12698_),
    .B(_12896_),
    .Y(_04141_));
 AO21x1_ASAP7_75t_R _29657_ (.A1(_12550_),
    .A2(_12508_),
    .B(_12565_),
    .Y(_12897_));
 AO32x1_ASAP7_75t_R _29658_ (.A1(_12488_),
    .A2(_12474_),
    .A3(_12897_),
    .B1(_12585_),
    .B2(_12785_),
    .Y(_12898_));
 AO21x1_ASAP7_75t_R _29659_ (.A1(_12550_),
    .A2(_12693_),
    .B(_12898_),
    .Y(_12899_));
 OR3x1_ASAP7_75t_R _29660_ (.A(_11846_),
    .B(_11847_),
    .C(_12899_),
    .Y(_12900_));
 OA21x2_ASAP7_75t_R _29661_ (.A1(_13244_),
    .A2(_12698_),
    .B(_12900_),
    .Y(_04142_));
 AO221x1_ASAP7_75t_R _29662_ (.A1(_12542_),
    .A2(_12496_),
    .B1(_12669_),
    .B2(_12552_),
    .C(_12757_),
    .Y(_12901_));
 AND3x1_ASAP7_75t_R _29663_ (.A(_12617_),
    .B(_12508_),
    .C(_12567_),
    .Y(_12902_));
 AO21x1_ASAP7_75t_R _29664_ (.A1(_12552_),
    .A2(_12466_),
    .B(_12902_),
    .Y(_12903_));
 OR3x1_ASAP7_75t_R _29665_ (.A(_12617_),
    .B(_12487_),
    .C(_12791_),
    .Y(_12904_));
 AO21x1_ASAP7_75t_R _29666_ (.A1(_12375_),
    .A2(_12567_),
    .B(_12552_),
    .Y(_12905_));
 AO221x1_ASAP7_75t_R _29667_ (.A1(_12566_),
    .A2(_12903_),
    .B1(_12904_),
    .B2(_12905_),
    .C(_12560_),
    .Y(_12906_));
 AND5x1_ASAP7_75t_R _29668_ (.A(_12457_),
    .B(_12373_),
    .C(_12391_),
    .D(_12507_),
    .E(_12465_),
    .Y(_12907_));
 AO21x1_ASAP7_75t_R _29669_ (.A1(_12552_),
    .A2(_12424_),
    .B(_12907_),
    .Y(_12908_));
 AO221x1_ASAP7_75t_R _29670_ (.A1(_12552_),
    .A2(_12729_),
    .B1(_12908_),
    .B2(_12566_),
    .C(_12886_),
    .Y(_12909_));
 AND4x1_ASAP7_75t_R _29671_ (.A(_11784_),
    .B(_12901_),
    .C(_12906_),
    .D(_12909_),
    .Y(_12910_));
 AO21x1_ASAP7_75t_R _29672_ (.A1(_09617_),
    .A2(_12631_),
    .B(_12910_),
    .Y(_04143_));
 AO21x1_ASAP7_75t_R _29673_ (.A1(_12544_),
    .A2(_12587_),
    .B(_12560_),
    .Y(_12911_));
 OAI22x1_ASAP7_75t_R _29674_ (.A1(_12424_),
    .A2(_12609_),
    .B1(_12627_),
    .B2(_12500_),
    .Y(_12912_));
 AO221x1_ASAP7_75t_R _29675_ (.A1(_12508_),
    .A2(_12561_),
    .B1(_12912_),
    .B2(_12374_),
    .C(_12592_),
    .Y(_12913_));
 INVx1_ASAP7_75t_R _29676_ (.A(_12913_),
    .Y(_12914_));
 AO21x1_ASAP7_75t_R _29677_ (.A1(_12568_),
    .A2(_12911_),
    .B(_12914_),
    .Y(_12915_));
 AO221x1_ASAP7_75t_R _29678_ (.A1(_12544_),
    .A2(_12496_),
    .B1(_12669_),
    .B2(_12431_),
    .C(_12757_),
    .Y(_12916_));
 AND3x4_ASAP7_75t_R _29679_ (.A(_11865_),
    .B(_12915_),
    .C(_12916_),
    .Y(_12917_));
 AO21x1_ASAP7_75t_R _29680_ (.A1(_13456_),
    .A2(_12631_),
    .B(_12917_),
    .Y(_04144_));
 NAND2x1_ASAP7_75t_R _29681_ (.A(_12567_),
    .B(_12785_),
    .Y(_12918_));
 AO221x1_ASAP7_75t_R _29682_ (.A1(_12546_),
    .A2(_12587_),
    .B1(_12918_),
    .B2(_12555_),
    .C(_12560_),
    .Y(_12919_));
 AO22x1_ASAP7_75t_R _29683_ (.A1(_12617_),
    .A2(_12546_),
    .B1(_12587_),
    .B2(_12550_),
    .Y(_12920_));
 AO221x1_ASAP7_75t_R _29684_ (.A1(_12555_),
    .A2(_12669_),
    .B1(_12920_),
    .B2(_12467_),
    .C(_12757_),
    .Y(_12921_));
 AO21x1_ASAP7_75t_R _29685_ (.A1(_12555_),
    .A2(_12581_),
    .B(_12568_),
    .Y(_12922_));
 AND4x1_ASAP7_75t_R _29686_ (.A(_11784_),
    .B(_12919_),
    .C(_12921_),
    .D(_12922_),
    .Y(_12923_));
 AO21x1_ASAP7_75t_R _29687_ (.A1(_13603_),
    .A2(_12631_),
    .B(_12923_),
    .Y(_04145_));
 AND2x2_ASAP7_75t_R _29688_ (.A(_00022_),
    .B(_11819_),
    .Y(_12924_));
 AOI21x1_ASAP7_75t_R _29689_ (.A1(_00019_),
    .A2(_12557_),
    .B(_12924_),
    .Y(_04146_));
 AND2x2_ASAP7_75t_R _29690_ (.A(_01690_),
    .B(_11819_),
    .Y(_12925_));
 AOI21x1_ASAP7_75t_R _29691_ (.A1(_14379_),
    .A2(_12557_),
    .B(_12925_),
    .Y(_04147_));
 NAND2x1_ASAP7_75t_R _29692_ (.A(_07316_),
    .B(_11785_),
    .Y(_12926_));
 OA21x2_ASAP7_75t_R _29693_ (.A1(_13274_),
    .A2(_11785_),
    .B(_12926_),
    .Y(_04148_));
 INVx1_ASAP7_75t_R _29694_ (.A(_01688_),
    .Y(_12927_));
 NAND2x1_ASAP7_75t_R _29695_ (.A(_01502_),
    .B(_12540_),
    .Y(_12928_));
 OA21x2_ASAP7_75t_R _29696_ (.A1(_12927_),
    .A2(_12518_),
    .B(_12928_),
    .Y(_04149_));
 AND2x2_ASAP7_75t_R _29697_ (.A(_01687_),
    .B(_11819_),
    .Y(_12929_));
 AOI21x1_ASAP7_75t_R _29698_ (.A1(_01501_),
    .A2(_12557_),
    .B(_12929_),
    .Y(_04150_));
 AND2x2_ASAP7_75t_R _29699_ (.A(_07328_),
    .B(_11819_),
    .Y(_12930_));
 AOI21x1_ASAP7_75t_R _29700_ (.A1(_15708_),
    .A2(_12557_),
    .B(_12930_),
    .Y(_04151_));
 AND2x2_ASAP7_75t_R _29701_ (.A(_01685_),
    .B(_11819_),
    .Y(_12931_));
 AOI21x1_ASAP7_75t_R _29702_ (.A1(_15832_),
    .A2(_12557_),
    .B(_12931_),
    .Y(_04152_));
 AND2x2_ASAP7_75t_R _29703_ (.A(_07335_),
    .B(_11819_),
    .Y(_12932_));
 AOI21x1_ASAP7_75t_R _29704_ (.A1(_01498_),
    .A2(_12557_),
    .B(_12932_),
    .Y(_04153_));
 BUFx12f_ASAP7_75t_R _29705_ (.A(_11832_),
    .Y(_12933_));
 AND2x2_ASAP7_75t_R _29706_ (.A(_00023_),
    .B(_11819_),
    .Y(_12934_));
 AOI21x1_ASAP7_75t_R _29707_ (.A1(_16079_),
    .A2(_12933_),
    .B(_12934_),
    .Y(_04154_));
 AND2x2_ASAP7_75t_R _29708_ (.A(_01683_),
    .B(_11819_),
    .Y(_12935_));
 AOI21x1_ASAP7_75t_R _29709_ (.A1(_16192_),
    .A2(_12933_),
    .B(_12935_),
    .Y(_04155_));
 OR3x1_ASAP7_75t_R _29710_ (.A(_05526_),
    .B(_11846_),
    .C(_11847_),
    .Y(_12936_));
 OA21x2_ASAP7_75t_R _29711_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(_11785_),
    .B(_12936_),
    .Y(_04156_));
 BUFx6f_ASAP7_75t_R _29712_ (.A(_11784_),
    .Y(_12937_));
 AND2x2_ASAP7_75t_R _29713_ (.A(_01682_),
    .B(_12937_),
    .Y(_12938_));
 AOI21x1_ASAP7_75t_R _29714_ (.A1(_01495_),
    .A2(_12933_),
    .B(_12938_),
    .Y(_04157_));
 AND2x2_ASAP7_75t_R _29715_ (.A(_01681_),
    .B(_12937_),
    .Y(_12939_));
 AOI21x1_ASAP7_75t_R _29716_ (.A1(_01494_),
    .A2(_12933_),
    .B(_12939_),
    .Y(_04158_));
 AND2x2_ASAP7_75t_R _29717_ (.A(_01680_),
    .B(_12937_),
    .Y(_12940_));
 AOI21x1_ASAP7_75t_R _29718_ (.A1(_01493_),
    .A2(_12933_),
    .B(_12940_),
    .Y(_04159_));
 AND2x2_ASAP7_75t_R _29719_ (.A(_01679_),
    .B(_12937_),
    .Y(_12941_));
 AOI21x1_ASAP7_75t_R _29720_ (.A1(_16698_),
    .A2(_12933_),
    .B(_12941_),
    .Y(_04160_));
 AND2x2_ASAP7_75t_R _29721_ (.A(_01678_),
    .B(_12937_),
    .Y(_12942_));
 AOI21x1_ASAP7_75t_R _29722_ (.A1(_01491_),
    .A2(_12933_),
    .B(_12942_),
    .Y(_04161_));
 AND2x2_ASAP7_75t_R _29723_ (.A(_01677_),
    .B(_12937_),
    .Y(_12943_));
 AOI21x1_ASAP7_75t_R _29724_ (.A1(_01490_),
    .A2(_12933_),
    .B(_12943_),
    .Y(_04162_));
 NAND2x1_ASAP7_75t_R _29725_ (.A(_04306_),
    .B(_11832_),
    .Y(_12944_));
 OA21x2_ASAP7_75t_R _29726_ (.A1(_11864_),
    .A2(_12518_),
    .B(_12944_),
    .Y(_04163_));
 AND2x2_ASAP7_75t_R _29727_ (.A(_01675_),
    .B(_12937_),
    .Y(_12945_));
 AOI21x1_ASAP7_75t_R _29728_ (.A1(_04419_),
    .A2(_12933_),
    .B(_12945_),
    .Y(_04164_));
 AND2x2_ASAP7_75t_R _29729_ (.A(_01674_),
    .B(_12937_),
    .Y(_12946_));
 AOI21x1_ASAP7_75t_R _29730_ (.A1(_01487_),
    .A2(_12933_),
    .B(_12946_),
    .Y(_04165_));
 BUFx12f_ASAP7_75t_R _29731_ (.A(_11832_),
    .Y(_12947_));
 AND2x2_ASAP7_75t_R _29732_ (.A(_01673_),
    .B(_12937_),
    .Y(_12948_));
 AOI21x1_ASAP7_75t_R _29733_ (.A1(_04667_),
    .A2(_12947_),
    .B(_12948_),
    .Y(_04166_));
 OR3x1_ASAP7_75t_R _29734_ (.A(\cs_registers_i.pc_if_i[2] ),
    .B(_11846_),
    .C(_11847_),
    .Y(_12949_));
 OA21x2_ASAP7_75t_R _29735_ (.A1(\cs_registers_i.pc_id_i[2] ),
    .A2(_11785_),
    .B(_12949_),
    .Y(_04167_));
 AND2x2_ASAP7_75t_R _29736_ (.A(_01672_),
    .B(_12937_),
    .Y(_12950_));
 AOI21x1_ASAP7_75t_R _29737_ (.A1(_01485_),
    .A2(_12947_),
    .B(_12950_),
    .Y(_04168_));
 AND2x2_ASAP7_75t_R _29738_ (.A(_01671_),
    .B(_12558_),
    .Y(_12951_));
 AOI21x1_ASAP7_75t_R _29739_ (.A1(_01484_),
    .A2(_12947_),
    .B(_12951_),
    .Y(_04169_));
 AND2x2_ASAP7_75t_R _29740_ (.A(_00021_),
    .B(_12558_),
    .Y(_12952_));
 AOI21x1_ASAP7_75t_R _29741_ (.A1(_14773_),
    .A2(_12947_),
    .B(_12952_),
    .Y(_04170_));
 AND2x2_ASAP7_75t_R _29742_ (.A(_01670_),
    .B(_12558_),
    .Y(_12953_));
 AOI21x1_ASAP7_75t_R _29743_ (.A1(_14837_),
    .A2(_12947_),
    .B(_12953_),
    .Y(_04171_));
 AND2x2_ASAP7_75t_R _29744_ (.A(_01669_),
    .B(_12558_),
    .Y(_12954_));
 AOI21x1_ASAP7_75t_R _29745_ (.A1(_14900_),
    .A2(_12947_),
    .B(_12954_),
    .Y(_04172_));
 AND2x2_ASAP7_75t_R _29746_ (.A(_01668_),
    .B(_12558_),
    .Y(_12955_));
 AOI21x1_ASAP7_75t_R _29747_ (.A1(_14966_),
    .A2(_12947_),
    .B(_12955_),
    .Y(_04173_));
 AND2x2_ASAP7_75t_R _29748_ (.A(_01667_),
    .B(_12558_),
    .Y(_12956_));
 AOI21x1_ASAP7_75t_R _29749_ (.A1(_01480_),
    .A2(_12947_),
    .B(_12956_),
    .Y(_04174_));
 AND2x2_ASAP7_75t_R _29750_ (.A(_01666_),
    .B(_12558_),
    .Y(_12957_));
 AOI21x1_ASAP7_75t_R _29751_ (.A1(_15099_),
    .A2(_12947_),
    .B(_12957_),
    .Y(_04175_));
 AND2x2_ASAP7_75t_R _29752_ (.A(_01665_),
    .B(_12558_),
    .Y(_12958_));
 AOI21x1_ASAP7_75t_R _29753_ (.A1(_15158_),
    .A2(_12947_),
    .B(_12958_),
    .Y(_04176_));
 INVx1_ASAP7_75t_R _29754_ (.A(_18314_),
    .Y(_17485_));
 INVx1_ASAP7_75t_R _29755_ (.A(_02269_),
    .Y(_18226_));
 INVx1_ASAP7_75t_R _29756_ (.A(_18153_),
    .Y(_17118_));
 INVx1_ASAP7_75t_R _29757_ (.A(_18141_),
    .Y(_17096_));
 INVx1_ASAP7_75t_R _29758_ (.A(_18152_),
    .Y(_17095_));
 INVx1_ASAP7_75t_R _29759_ (.A(_18133_),
    .Y(_17068_));
 INVx1_ASAP7_75t_R _29760_ (.A(_18475_),
    .Y(_17829_));
 INVx1_ASAP7_75t_R _29761_ (.A(_18491_),
    .Y(_17828_));
 INVx1_ASAP7_75t_R _29762_ (.A(_18443_),
    .Y(_17709_));
 INVx1_ASAP7_75t_R _29763_ (.A(_18425_),
    .Y(_17710_));
 INVx1_ASAP7_75t_R _29764_ (.A(_18423_),
    .Y(_17662_));
 INVx1_ASAP7_75t_R _29765_ (.A(_18404_),
    .Y(_17663_));
 INVx1_ASAP7_75t_R _29766_ (.A(_18440_),
    .Y(_17703_));
 INVx1_ASAP7_75t_R _29767_ (.A(_18140_),
    .Y(_17067_));
 INVx1_ASAP7_75t_R _29768_ (.A(_18424_),
    .Y(_17704_));
 INVx1_ASAP7_75t_R _29769_ (.A(_18170_),
    .Y(_17158_));
 INVx1_ASAP7_75t_R _29770_ (.A(_18355_),
    .Y(_17519_));
 INVx1_ASAP7_75t_R _29771_ (.A(_18333_),
    .Y(_17520_));
 INVx1_ASAP7_75t_R _29772_ (.A(_18358_),
    .Y(_17572_));
 INVx1_ASAP7_75t_R _29773_ (.A(_18385_),
    .Y(_17571_));
 INVx1_ASAP7_75t_R _29774_ (.A(_18357_),
    .Y(_17524_));
 INVx1_ASAP7_75t_R _29775_ (.A(_18334_),
    .Y(_17525_));
 INVx1_ASAP7_75t_R _29776_ (.A(_18378_),
    .Y(_17568_));
 INVx1_ASAP7_75t_R _29777_ (.A(_18356_),
    .Y(_17569_));
 INVx1_ASAP7_75t_R _29778_ (.A(_17738_),
    .Y(_17689_));
 INVx1_ASAP7_75t_R _29779_ (.A(_18439_),
    .Y(_17698_));
 INVx1_ASAP7_75t_R _29780_ (.A(_18422_),
    .Y(_17699_));
 INVx1_ASAP7_75t_R _29781_ (.A(_18419_),
    .Y(_17649_));
 INVx1_ASAP7_75t_R _29782_ (.A(_18399_),
    .Y(_17650_));
 INVx1_ASAP7_75t_R _29783_ (.A(_18442_),
    .Y(_17695_));
 INVx1_ASAP7_75t_R _29784_ (.A(_18420_),
    .Y(_17696_));
 INVx1_ASAP7_75t_R _29785_ (.A(_18362_),
    .Y(_17580_));
 INVx1_ASAP7_75t_R _29786_ (.A(_18401_),
    .Y(_17616_));
 INVx1_ASAP7_75t_R _29787_ (.A(_18381_),
    .Y(_17617_));
 INVx1_ASAP7_75t_R _29788_ (.A(_18386_),
    .Y(_17585_));
 INVx1_ASAP7_75t_R _29789_ (.A(_02276_),
    .Y(_17551_));
 INVx1_ASAP7_75t_R _29790_ (.A(_18382_),
    .Y(_17579_));
 INVx1_ASAP7_75t_R _29791_ (.A(_18406_),
    .Y(_17613_));
 INVx1_ASAP7_75t_R _29792_ (.A(_18379_),
    .Y(_17614_));
 INVx1_ASAP7_75t_R _29793_ (.A(_18387_),
    .Y(_17629_));
 INVx1_ASAP7_75t_R _29794_ (.A(_18384_),
    .Y(_17628_));
 INVx1_ASAP7_75t_R _29795_ (.A(_18403_),
    .Y(_17621_));
 INVx1_ASAP7_75t_R _29796_ (.A(_18383_),
    .Y(_17622_));
 INVx1_ASAP7_75t_R _29797_ (.A(_18398_),
    .Y(_17606_));
 INVx1_ASAP7_75t_R _29798_ (.A(_18377_),
    .Y(_17607_));
 INVx1_ASAP7_75t_R _29799_ (.A(_18380_),
    .Y(_17574_));
 INVx1_ASAP7_75t_R _29800_ (.A(_18360_),
    .Y(_17575_));
 INVx1_ASAP7_75t_R _29801_ (.A(_18389_),
    .Y(_17631_));
 INVx1_ASAP7_75t_R _29802_ (.A(_02279_),
    .Y(_17679_));
 INVx1_ASAP7_75t_R _29803_ (.A(_18169_),
    .Y(_17128_));
 INVx1_ASAP7_75t_R _29804_ (.A(_00215_),
    .Y(_17639_));
 INVx1_ASAP7_75t_R _29805_ (.A(_18415_),
    .Y(_17642_));
 INVx1_ASAP7_75t_R _29806_ (.A(_18394_),
    .Y(_17643_));
 INVx1_ASAP7_75t_R _29807_ (.A(_18388_),
    .Y(_17588_));
 INVx1_ASAP7_75t_R _29808_ (.A(_18368_),
    .Y(_17589_));
 INVx1_ASAP7_75t_R _29809_ (.A(_18369_),
    .Y(_17594_));
 INVx1_ASAP7_75t_R _29810_ (.A(_18332_),
    .Y(_17474_));
 INVx1_ASAP7_75t_R _29811_ (.A(_18309_),
    .Y(_17475_));
 INVx1_ASAP7_75t_R _29812_ (.A(_18366_),
    .Y(_17587_));
 INVx1_ASAP7_75t_R _29813_ (.A(_18364_),
    .Y(_17527_));
 INVx1_ASAP7_75t_R _29814_ (.A(_18336_),
    .Y(_17528_));
 INVx1_ASAP7_75t_R _29815_ (.A(_18335_),
    .Y(_17479_));
 INVx1_ASAP7_75t_R _29816_ (.A(_18310_),
    .Y(_17480_));
 INVx1_ASAP7_75t_R _29817_ (.A(_18435_),
    .Y(_17683_));
 INVx1_ASAP7_75t_R _29818_ (.A(_18416_),
    .Y(_17684_));
 INVx1_ASAP7_75t_R _29819_ (.A(_18429_),
    .Y(_17671_));
 INVx1_ASAP7_75t_R _29820_ (.A(_18410_),
    .Y(_17672_));
 INVx1_ASAP7_75t_R _29821_ (.A(_18408_),
    .Y(_17670_));
 INVx1_ASAP7_75t_R _29822_ (.A(_18427_),
    .Y(_17668_));
 INVx1_ASAP7_75t_R _29823_ (.A(_18405_),
    .Y(_17669_));
 INVx1_ASAP7_75t_R _29824_ (.A(_18421_),
    .Y(_17657_));
 INVx1_ASAP7_75t_R _29825_ (.A(_18402_),
    .Y(_17658_));
 INVx1_ASAP7_75t_R _29826_ (.A(_18426_),
    .Y(_17655_));
 INVx1_ASAP7_75t_R _29827_ (.A(_18400_),
    .Y(_17656_));
 INVx1_ASAP7_75t_R _29828_ (.A(_02260_),
    .Y(_17165_));
 INVx1_ASAP7_75t_R _29829_ (.A(_18142_),
    .Y(_17074_));
 INVx1_ASAP7_75t_R _29830_ (.A(_18135_),
    .Y(_17075_));
 INVx1_ASAP7_75t_R _29831_ (.A(_17739_),
    .Y(_17731_));
 INVx1_ASAP7_75t_R _29832_ (.A(_17773_),
    .Y(_17730_));
 INVx1_ASAP7_75t_R _29833_ (.A(_18432_),
    .Y(_17676_));
 INVx1_ASAP7_75t_R _29834_ (.A(_18411_),
    .Y(_17677_));
 INVx1_ASAP7_75t_R _29835_ (.A(_18412_),
    .Y(_17635_));
 INVx1_ASAP7_75t_R _29836_ (.A(_18390_),
    .Y(_17636_));
 INVx1_ASAP7_75t_R _29837_ (.A(_18168_),
    .Y(_17156_));
 INVx1_ASAP7_75t_R _29838_ (.A(_18182_),
    .Y(_17155_));
 INVx1_ASAP7_75t_R _29839_ (.A(_18391_),
    .Y(_17593_));
 INVx1_ASAP7_75t_R _29840_ (.A(_02211_),
    .Y(_17131_));
 INVx1_ASAP7_75t_R _29841_ (.A(_18179_),
    .Y(_17150_));
 INVx1_ASAP7_75t_R _29842_ (.A(_18167_),
    .Y(_17151_));
 INVx1_ASAP7_75t_R _29843_ (.A(_18190_),
    .Y(_17179_));
 INVx1_ASAP7_75t_R _29844_ (.A(_18180_),
    .Y(_17180_));
 INVx1_ASAP7_75t_R _29845_ (.A(_02212_),
    .Y(_17273_));
 INVx1_ASAP7_75t_R _29846_ (.A(_18178_),
    .Y(_17174_));
 INVx1_ASAP7_75t_R _29847_ (.A(_02274_),
    .Y(_17416_));
 INVx1_ASAP7_75t_R _29848_ (.A(_18363_),
    .Y(_17586_));
 INVx1_ASAP7_75t_R _29849_ (.A(_18407_),
    .Y(_17627_));
 INVx1_ASAP7_75t_R _29850_ (.A(_18409_),
    .Y(_17630_));
 INVx1_ASAP7_75t_R _29851_ (.A(_18155_),
    .Y(_17124_));
 INVx1_ASAP7_75t_R _29852_ (.A(_02213_),
    .Y(_17314_));
 INVx1_ASAP7_75t_R _29853_ (.A(_18338_),
    .Y(_17530_));
 INVx1_ASAP7_75t_R _29854_ (.A(_18359_),
    .Y(_17529_));
 INVx1_ASAP7_75t_R _29855_ (.A(_02275_),
    .Y(_17506_));
 INVx1_ASAP7_75t_R _29856_ (.A(_18154_),
    .Y(_17102_));
 INVx1_ASAP7_75t_R _29857_ (.A(_02251_),
    .Y(_17079_));
 INVx1_ASAP7_75t_R _29858_ (.A(_18122_),
    .Y(_17043_));
 INVx1_ASAP7_75t_R _29859_ (.A(_18112_),
    .Y(_17044_));
 INVx1_ASAP7_75t_R _29860_ (.A(_00123_),
    .Y(_18126_));
 INVx1_ASAP7_75t_R _29861_ (.A(_18108_),
    .Y(_17021_));
 INVx1_ASAP7_75t_R _29862_ (.A(_18104_),
    .Y(_17022_));
 INVx1_ASAP7_75t_R _29863_ (.A(_18365_),
    .Y(_17540_));
 INVx1_ASAP7_75t_R _29864_ (.A(_18341_),
    .Y(_17541_));
 INVx1_ASAP7_75t_R _29865_ (.A(_18110_),
    .Y(_17042_));
 INVx1_ASAP7_75t_R _29866_ (.A(_00137_),
    .Y(_17072_));
 INVx1_ASAP7_75t_R _29867_ (.A(_00236_),
    .Y(_17894_));
 INVx1_ASAP7_75t_R _29868_ (.A(_02286_),
    .Y(_17921_));
 INVx1_ASAP7_75t_R _29869_ (.A(_18181_),
    .Y(_17185_));
 INVx1_ASAP7_75t_R _29870_ (.A(_18193_),
    .Y(_17184_));
 INVx1_ASAP7_75t_R _29871_ (.A(_18183_),
    .Y(_17188_));
 INVx1_ASAP7_75t_R _29872_ (.A(_18203_),
    .Y(_17187_));
 INVx1_ASAP7_75t_R _29873_ (.A(_00138_),
    .Y(_17081_));
 INVx1_ASAP7_75t_R _29874_ (.A(_18143_),
    .Y(_17103_));
 INVx1_ASAP7_75t_R _29875_ (.A(_18165_),
    .Y(_17145_));
 INVx1_ASAP7_75t_R _29876_ (.A(_00140_),
    .Y(_18149_));
 INVx1_ASAP7_75t_R _29877_ (.A(_17563_),
    .Y(_17559_));
 INVx1_ASAP7_75t_R _29878_ (.A(_18166_),
    .Y(_17123_));
 INVx1_ASAP7_75t_R _29879_ (.A(_18132_),
    .Y(_17049_));
 INVx1_ASAP7_75t_R _29880_ (.A(_18144_),
    .Y(_17083_));
 INVx1_ASAP7_75t_R _29881_ (.A(_17935_),
    .Y(_17932_));
 INVx5_ASAP7_75t_R _29882_ (.A(_18456_),
    .Y(_17735_));
 INVx1_ASAP7_75t_R _29883_ (.A(_02266_),
    .Y(_18201_));
 INVx1_ASAP7_75t_R _29884_ (.A(_18519_),
    .Y(_17914_));
 INVx1_ASAP7_75t_R _29885_ (.A(_18540_),
    .Y(_17950_));
 INVx1_ASAP7_75t_R _29886_ (.A(_18518_),
    .Y(_17885_));
 INVx1_ASAP7_75t_R _29887_ (.A(_18172_),
    .Y(_17160_));
 INVx1_ASAP7_75t_R _29888_ (.A(_18184_),
    .Y(_17159_));
 INVx1_ASAP7_75t_R _29889_ (.A(_02268_),
    .Y(_17320_));
 INVx1_ASAP7_75t_R _29890_ (.A(_18246_),
    .Y(_17328_));
 INVx1_ASAP7_75t_R _29891_ (.A(_02271_),
    .Y(_17360_));
 INVx1_ASAP7_75t_R _29892_ (.A(_18134_),
    .Y(_17056_));
 INVx1_ASAP7_75t_R _29893_ (.A(_18339_),
    .Y(_17489_));
 INVx1_ASAP7_75t_R _29894_ (.A(_18316_),
    .Y(_17490_));
 INVx1_ASAP7_75t_R _29895_ (.A(_18123_),
    .Y(_17057_));
 INVx1_ASAP7_75t_R _29896_ (.A(_18177_),
    .Y(_17144_));
 INVx1_ASAP7_75t_R _29897_ (.A(_18521_),
    .Y(_17890_));
 INVx1_ASAP7_75t_R _29898_ (.A(_00149_),
    .Y(_18163_));
 INVx1_ASAP7_75t_R _29899_ (.A(_02261_),
    .Y(_18162_));
 INVx1_ASAP7_75t_R _29900_ (.A(_18471_),
    .Y(_17783_));
 INVx1_ASAP7_75t_R _29901_ (.A(_18541_),
    .Y(_17977_));
 INVx1_ASAP7_75t_R _29902_ (.A(_02257_),
    .Y(_18148_));
 INVx1_ASAP7_75t_R _29903_ (.A(_18340_),
    .Y(_17535_));
 INVx1_ASAP7_75t_R _29904_ (.A(_18361_),
    .Y(_17534_));
 INVx1_ASAP7_75t_R _29905_ (.A(_18109_),
    .Y(_17038_));
 INVx1_ASAP7_75t_R _29906_ (.A(_18120_),
    .Y(_17037_));
 INVx1_ASAP7_75t_R _29907_ (.A(_18509_),
    .Y(_17867_));
 INVx1_ASAP7_75t_R _29908_ (.A(_18490_),
    .Y(_17861_));
 INVx1_ASAP7_75t_R _29909_ (.A(_18506_),
    .Y(_17860_));
 INVx1_ASAP7_75t_R _29910_ (.A(_18121_),
    .Y(_17050_));
 INVx1_ASAP7_75t_R _29911_ (.A(_00155_),
    .Y(_17169_));
 INVx1_ASAP7_75t_R _29912_ (.A(_00164_),
    .Y(_17168_));
 INVx1_ASAP7_75t_R _29913_ (.A(_00209_),
    .Y(_17552_));
 INVx1_ASAP7_75t_R _29914_ (.A(_02277_),
    .Y(_17596_));
 INVx1_ASAP7_75t_R _29915_ (.A(_02247_),
    .Y(_17059_));
 INVx1_ASAP7_75t_R _29916_ (.A(_00250_),
    .Y(_17968_));
 INVx1_ASAP7_75t_R _29917_ (.A(_17961_),
    .Y(_17957_));
 INVx1_ASAP7_75t_R _29918_ (.A(_17984_),
    .Y(_17956_));
 INVx1_ASAP7_75t_R _29919_ (.A(_18374_),
    .Y(_17601_));
 INVx1_ASAP7_75t_R _29920_ (.A(_18395_),
    .Y(_17600_));
 INVx1_ASAP7_75t_R _29921_ (.A(_17960_),
    .Y(_17931_));
 INVx1_ASAP7_75t_R _29922_ (.A(_18277_),
    .Y(_17389_));
 INVx1_ASAP7_75t_R _29923_ (.A(_18291_),
    .Y(_17388_));
 INVx1_ASAP7_75t_R _29924_ (.A(_17965_),
    .Y(_17959_));
 INVx1_ASAP7_75t_R _29925_ (.A(_17987_),
    .Y(_17958_));
 INVx1_ASAP7_75t_R _29926_ (.A(_02217_),
    .Y(_17991_));
 INVx1_ASAP7_75t_R _29927_ (.A(_18285_),
    .Y(_17430_));
 INVx2_ASAP7_75t_R _29928_ (.A(_18515_),
    .Y(_17911_));
 INVx1_ASAP7_75t_R _29929_ (.A(_18308_),
    .Y(_17429_));
 INVx1_ASAP7_75t_R _29930_ (.A(_18528_),
    .Y(_17910_));
 INVx1_ASAP7_75t_R _29931_ (.A(_18293_),
    .Y(_17451_));
 INVx1_ASAP7_75t_R _29932_ (.A(_18319_),
    .Y(_17450_));
 INVx2_ASAP7_75t_R _29933_ (.A(_17937_),
    .Y(_17936_));
 INVx1_ASAP7_75t_R _29934_ (.A(_17964_),
    .Y(_17934_));
 INVx1_ASAP7_75t_R _29935_ (.A(_18537_),
    .Y(_17963_));
 INVx1_ASAP7_75t_R _29936_ (.A(_18544_),
    .Y(_17962_));
 INVx1_ASAP7_75t_R _29937_ (.A(_18271_),
    .Y(_17379_));
 INVx1_ASAP7_75t_R _29938_ (.A(_18287_),
    .Y(_17378_));
 INVx1_ASAP7_75t_R _29939_ (.A(_18288_),
    .Y(_17438_));
 INVx1_ASAP7_75t_R _29940_ (.A(_18318_),
    .Y(_17437_));
 INVx1_ASAP7_75t_R _29941_ (.A(_18500_),
    .Y(_17883_));
 INVx1_ASAP7_75t_R _29942_ (.A(_18516_),
    .Y(_17882_));
 INVx1_ASAP7_75t_R _29943_ (.A(_18517_),
    .Y(_17912_));
 INVx1_ASAP7_75t_R _29944_ (.A(_18514_),
    .Y(_17906_));
 INVx1_ASAP7_75t_R _29945_ (.A(_18513_),
    .Y(_17877_));
 INVx1_ASAP7_75t_R _29946_ (.A(_18499_),
    .Y(_17878_));
 INVx1_ASAP7_75t_R _29947_ (.A(_18320_),
    .Y(_17497_));
 INVx1_ASAP7_75t_R _29948_ (.A(_18529_),
    .Y(_17913_));
 INVx1_ASAP7_75t_R _29949_ (.A(_18534_),
    .Y(_17951_));
 INVx1_ASAP7_75t_R _29950_ (.A(_18485_),
    .Y(_17853_));
 INVx1_ASAP7_75t_R _29951_ (.A(_18501_),
    .Y(_17852_));
 INVx1_ASAP7_75t_R _29952_ (.A(_18502_),
    .Y(_17884_));
 INVx1_ASAP7_75t_R _29953_ (.A(_18484_),
    .Y(_17846_));
 INVx1_ASAP7_75t_R _29954_ (.A(_18498_),
    .Y(_17845_));
 INVx1_ASAP7_75t_R _29955_ (.A(_18504_),
    .Y(_17886_));
 INVx1_ASAP7_75t_R _29956_ (.A(_18525_),
    .Y(_17926_));
 INVx1_ASAP7_75t_R _29957_ (.A(_18533_),
    .Y(_17925_));
 INVx1_ASAP7_75t_R _29958_ (.A(_18367_),
    .Y(_17543_));
 INVx1_ASAP7_75t_R _29959_ (.A(_18346_),
    .Y(_17544_));
 INVx1_ASAP7_75t_R _29960_ (.A(_18530_),
    .Y(_17918_));
 INVx1_ASAP7_75t_R _29961_ (.A(_18520_),
    .Y(_17919_));
 INVx1_ASAP7_75t_R _29962_ (.A(_18095_),
    .Y(_17006_));
 INVx1_ASAP7_75t_R _29963_ (.A(_18268_),
    .Y(_17327_));
 INVx1_ASAP7_75t_R _29964_ (.A(_02267_),
    .Y(_18208_));
 INVx1_ASAP7_75t_R _29965_ (.A(_00171_),
    .Y(_18209_));
 INVx1_ASAP7_75t_R _29966_ (.A(_18270_),
    .Y(_17374_));
 INVx1_ASAP7_75t_R _29967_ (.A(_00132_),
    .Y(_17062_));
 INVx1_ASAP7_75t_R _29968_ (.A(_18284_),
    .Y(_17373_));
 INVx1_ASAP7_75t_R _29969_ (.A(_18197_),
    .Y(_17194_));
 INVx1_ASAP7_75t_R _29970_ (.A(_18290_),
    .Y(_17440_));
 INVx1_ASAP7_75t_R _29971_ (.A(_18313_),
    .Y(_17439_));
 INVx1_ASAP7_75t_R _29972_ (.A(_18322_),
    .Y(_17499_));
 INVx1_ASAP7_75t_R _29973_ (.A(_00112_),
    .Y(_18106_));
 INVx1_ASAP7_75t_R _29974_ (.A(_18345_),
    .Y(_17498_));
 INVx1_ASAP7_75t_R _29975_ (.A(_00118_),
    .Y(_18116_));
 INVx1_ASAP7_75t_R _29976_ (.A(_02248_),
    .Y(_18115_));
 INVx1_ASAP7_75t_R _29977_ (.A(_00119_),
    .Y(_18118_));
 INVx1_ASAP7_75t_R _29978_ (.A(_02249_),
    .Y(_18117_));
 INVx1_ASAP7_75t_R _29979_ (.A(_00125_),
    .Y(_18129_));
 INVx1_ASAP7_75t_R _29980_ (.A(_02253_),
    .Y(_18128_));
 INVx1_ASAP7_75t_R _29981_ (.A(_17091_),
    .Y(_18139_));
 INVx1_ASAP7_75t_R _29982_ (.A(_02255_),
    .Y(_18138_));
 INVx1_ASAP7_75t_R _29983_ (.A(_00133_),
    .Y(_18137_));
 INVx1_ASAP7_75t_R _29984_ (.A(_02254_),
    .Y(_18136_));
 INVx1_ASAP7_75t_R _29985_ (.A(_00141_),
    .Y(_18151_));
 INVx1_ASAP7_75t_R _29986_ (.A(_02258_),
    .Y(_18150_));
 INVx1_ASAP7_75t_R _29987_ (.A(_00102_),
    .Y(_17011_));
 INVx1_ASAP7_75t_R _29988_ (.A(_00106_),
    .Y(_17010_));
 INVx1_ASAP7_75t_R _29989_ (.A(_18470_),
    .Y(_17820_));
 INVx1_ASAP7_75t_R _29990_ (.A(_18486_),
    .Y(_17819_));
 INVx1_ASAP7_75t_R _29991_ (.A(_18487_),
    .Y(_17854_));
 INVx1_ASAP7_75t_R _29992_ (.A(_18469_),
    .Y(_17811_));
 INVx1_ASAP7_75t_R _29993_ (.A(_18483_),
    .Y(_17810_));
 INVx1_ASAP7_75t_R _29994_ (.A(_18489_),
    .Y(_17856_));
 INVx1_ASAP7_75t_R _29995_ (.A(_18503_),
    .Y(_17855_));
 INVx1_ASAP7_75t_R _29996_ (.A(_18510_),
    .Y(_17898_));
 INVx1_ASAP7_75t_R _29997_ (.A(_18524_),
    .Y(_17897_));
 INVx1_ASAP7_75t_R _29998_ (.A(_18505_),
    .Y(_17891_));
 INVx1_ASAP7_75t_R _29999_ (.A(_18352_),
    .Y(_17556_));
 INVx1_ASAP7_75t_R _30000_ (.A(_18373_),
    .Y(_17555_));
 INVx1_ASAP7_75t_R _30001_ (.A(_17944_),
    .Y(_17908_));
 INVx1_ASAP7_75t_R _30002_ (.A(_17903_),
    .Y(_17901_));
 INVx1_ASAP7_75t_R _30003_ (.A(_18455_),
    .Y(_17784_));
 INVx1_ASAP7_75t_R _30004_ (.A(_18472_),
    .Y(_17821_));
 INVx1_ASAP7_75t_R _30005_ (.A(_18474_),
    .Y(_17824_));
 INVx1_ASAP7_75t_R _30006_ (.A(_18488_),
    .Y(_17823_));
 INVx1_ASAP7_75t_R _30007_ (.A(_18495_),
    .Y(_17868_));
 INVx1_ASAP7_75t_R _30008_ (.A(_18312_),
    .Y(_17483_));
 INVx1_ASAP7_75t_R _30009_ (.A(_18347_),
    .Y(_17549_));
 INVx1_ASAP7_75t_R _30010_ (.A(_18441_),
    .Y(_17749_));
 INVx2_ASAP7_75t_R _30011_ (.A(_18457_),
    .Y(_17748_));
 INVx1_ASAP7_75t_R _30012_ (.A(_18458_),
    .Y(_17785_));
 INVx1_ASAP7_75t_R _30013_ (.A(_18370_),
    .Y(_17548_));
 INVx1_ASAP7_75t_R _30014_ (.A(_18460_),
    .Y(_17789_));
 INVx1_ASAP7_75t_R _30015_ (.A(_18473_),
    .Y(_17788_));
 INVx1_ASAP7_75t_R _30016_ (.A(_18480_),
    .Y(_17836_));
 INVx1_ASAP7_75t_R _30017_ (.A(_18494_),
    .Y(_17835_));
 INVx1_ASAP7_75t_R _30018_ (.A(_00212_),
    .Y(_17597_));
 INVx1_ASAP7_75t_R _30019_ (.A(_02278_),
    .Y(_17638_));
 INVx1_ASAP7_75t_R _30020_ (.A(_02284_),
    .Y(_17863_));
 INVx1_ASAP7_75t_R _30021_ (.A(_18444_),
    .Y(_17750_));
 INVx1_ASAP7_75t_R _30022_ (.A(_18446_),
    .Y(_17753_));
 INVx1_ASAP7_75t_R _30023_ (.A(_18459_),
    .Y(_17752_));
 INVx2_ASAP7_75t_R _30024_ (.A(_18476_),
    .Y(_17793_));
 INVx1_ASAP7_75t_R _30025_ (.A(_18461_),
    .Y(_17794_));
 INVx2_ASAP7_75t_R _30026_ (.A(_02283_),
    .Y(_17831_));
 INVx1_ASAP7_75t_R _30027_ (.A(_18479_),
    .Y(_17800_));
 INVx1_ASAP7_75t_R _30028_ (.A(_18466_),
    .Y(_17801_));
 INVx1_ASAP7_75t_R _30029_ (.A(_18428_),
    .Y(_17711_));
 INVx1_ASAP7_75t_R _30030_ (.A(_18430_),
    .Y(_17713_));
 INVx1_ASAP7_75t_R _30031_ (.A(_18445_),
    .Y(_17712_));
 INVx1_ASAP7_75t_R _30032_ (.A(_18452_),
    .Y(_17765_));
 INVx1_ASAP7_75t_R _30033_ (.A(_18465_),
    .Y(_17764_));
 INVx1_ASAP7_75t_R _30034_ (.A(_02282_),
    .Y(_17796_));
 INVx1_ASAP7_75t_R _30035_ (.A(_18447_),
    .Y(_17758_));
 INVx1_ASAP7_75t_R _30036_ (.A(_18462_),
    .Y(_17757_));
 INVx1_ASAP7_75t_R _30037_ (.A(_18436_),
    .Y(_17725_));
 INVx1_ASAP7_75t_R _30038_ (.A(_18451_),
    .Y(_17724_));
 INVx1_ASAP7_75t_R _30039_ (.A(_00239_),
    .Y(_17922_));
 INVx1_ASAP7_75t_R _30040_ (.A(_02287_),
    .Y(_17945_));
 INVx1_ASAP7_75t_R _30041_ (.A(_18448_),
    .Y(_17717_));
 INVx1_ASAP7_75t_R _30042_ (.A(_18431_),
    .Y(_17718_));
 INVx1_ASAP7_75t_R _30043_ (.A(_02281_),
    .Y(_17760_));
 INVx1_ASAP7_75t_R _30044_ (.A(_02263_),
    .Y(_17203_));
 INVx1_ASAP7_75t_R _30045_ (.A(_00242_),
    .Y(_17946_));
 INVx1_ASAP7_75t_R _30046_ (.A(_02288_),
    .Y(_17971_));
 INVx1_ASAP7_75t_R _30047_ (.A(_18145_),
    .Y(_17112_));
 INVx1_ASAP7_75t_R _30048_ (.A(_18156_),
    .Y(_17111_));
 INVx1_ASAP7_75t_R _30049_ (.A(_02210_),
    .Y(_17109_));
 INVx1_ASAP7_75t_R _30050_ (.A(_00233_),
    .Y(_17864_));
 INVx1_ASAP7_75t_R _30051_ (.A(_02285_),
    .Y(_17893_));
 INVx1_ASAP7_75t_R _30052_ (.A(_17733_),
    .Y(_17729_));
 INVx1_ASAP7_75t_R _30053_ (.A(_17771_),
    .Y(_17728_));
 INVx1_ASAP7_75t_R _30054_ (.A(_00218_),
    .Y(_17680_));
 INVx1_ASAP7_75t_R _30055_ (.A(_02280_),
    .Y(_17720_));
 INVx1_ASAP7_75t_R _30056_ (.A(_17985_),
    .Y(_17982_));
 INVx1_ASAP7_75t_R _30057_ (.A(_17988_),
    .Y(_17983_));
 INVx1_ASAP7_75t_R _30058_ (.A(_18545_),
    .Y(_17986_));
 INVx1_ASAP7_75t_R _30059_ (.A(_18548_),
    .Y(_17995_));
 INVx1_ASAP7_75t_R _30060_ (.A(_00146_),
    .Y(_17100_));
 INVx1_ASAP7_75t_R _30061_ (.A(_18547_),
    .Y(_17976_));
 INVx1_ASAP7_75t_R _30062_ (.A(_02252_),
    .Y(_17084_));
 INVx1_ASAP7_75t_R _30063_ (.A(_00131_),
    .Y(_17088_));
 INVx1_ASAP7_75t_R _30064_ (.A(_00130_),
    .Y(_17054_));
 INVx1_ASAP7_75t_R _30065_ (.A(_18096_),
    .Y(_17016_));
 INVx1_ASAP7_75t_R _30066_ (.A(_18103_),
    .Y(_17015_));
 INVx1_ASAP7_75t_R _30067_ (.A(_18111_),
    .Y(_17028_));
 INVx1_ASAP7_75t_R _30068_ (.A(_02242_),
    .Y(_17029_));
 INVx1_ASAP7_75t_R _30069_ (.A(_00165_),
    .Y(_18187_));
 INVx1_ASAP7_75t_R _30070_ (.A(_02265_),
    .Y(_18186_));
 INVx1_ASAP7_75t_R _30071_ (.A(_00111_),
    .Y(_17033_));
 INVx1_ASAP7_75t_R _30072_ (.A(_00117_),
    .Y(_17032_));
 INVx1_ASAP7_75t_R _30073_ (.A(_00116_),
    .Y(_17026_));
 INVx1_ASAP7_75t_R _30074_ (.A(_02256_),
    .Y(_17136_));
 INVx1_ASAP7_75t_R _30075_ (.A(_17691_),
    .Y(_17688_));
 INVx1_ASAP7_75t_R _30076_ (.A(_18337_),
    .Y(_17484_));
 INVx1_ASAP7_75t_R _30077_ (.A(_18323_),
    .Y(_17504_));
 INVx1_ASAP7_75t_R _30078_ (.A(_18348_),
    .Y(_17503_));
 INVx1_ASAP7_75t_R _30079_ (.A(_17732_),
    .Y(_17687_));
 INVx1_ASAP7_75t_R _30080_ (.A(_00107_),
    .Y(_18101_));
 INVx1_ASAP7_75t_R _30081_ (.A(_02243_),
    .Y(_18100_));
 INVx1_ASAP7_75t_R _30082_ (.A(_02245_),
    .Y(_18105_));
 INVx1_ASAP7_75t_R _30083_ (.A(_00126_),
    .Y(_18131_));
 INVx1_ASAP7_75t_R _30084_ (.A(_17090_),
    .Y(_18130_));
 INVx1_ASAP7_75t_R _30085_ (.A(_00189_),
    .Y(_18265_));
 INVx1_ASAP7_75t_R _30086_ (.A(_02272_),
    .Y(_17404_));
 INVx1_ASAP7_75t_R _30087_ (.A(_18256_),
    .Y(_17348_));
 INVx1_ASAP7_75t_R _30088_ (.A(_18276_),
    .Y(_17347_));
 INVx1_ASAP7_75t_R _30089_ (.A(_18278_),
    .Y(_17395_));
 INVx1_ASAP7_75t_R _30090_ (.A(_18295_),
    .Y(_17394_));
 INVx1_ASAP7_75t_R _30091_ (.A(_18249_),
    .Y(_17339_));
 INVx1_ASAP7_75t_R _30092_ (.A(_18272_),
    .Y(_17338_));
 INVx1_ASAP7_75t_R _30093_ (.A(_02239_),
    .Y(_18091_));
 INVx1_ASAP7_75t_R _30094_ (.A(_02240_),
    .Y(_18093_));
 INVx1_ASAP7_75t_R _30095_ (.A(_18273_),
    .Y(_17382_));
 INVx1_ASAP7_75t_R _30096_ (.A(_18294_),
    .Y(_17381_));
 INVx1_ASAP7_75t_R _30097_ (.A(_02241_),
    .Y(_18094_));
 INVx1_ASAP7_75t_R _30098_ (.A(_18296_),
    .Y(_17452_));
 INVx1_ASAP7_75t_R _30099_ (.A(_18229_),
    .Y(_17282_));
 INVx1_ASAP7_75t_R _30100_ (.A(_18245_),
    .Y(_17281_));
 INVx1_ASAP7_75t_R _30101_ (.A(_18248_),
    .Y(_17334_));
 INVx1_ASAP7_75t_R _30102_ (.A(_18269_),
    .Y(_17333_));
 INVx1_ASAP7_75t_R _30103_ (.A(_02244_),
    .Y(_18102_));
 INVx1_ASAP7_75t_R _30104_ (.A(_18275_),
    .Y(_17384_));
 INVx1_ASAP7_75t_R _30105_ (.A(_02246_),
    .Y(_18107_));
 INVx1_ASAP7_75t_R _30106_ (.A(_02250_),
    .Y(_18119_));
 INVx1_ASAP7_75t_R _30107_ (.A(_18292_),
    .Y(_17445_));
 INVx1_ASAP7_75t_R _30108_ (.A(_18315_),
    .Y(_17444_));
 INVx1_ASAP7_75t_R _30109_ (.A(_18317_),
    .Y(_17496_));
 INVx1_ASAP7_75t_R _30110_ (.A(_18343_),
    .Y(_17495_));
 INVx1_ASAP7_75t_R _30111_ (.A(_18286_),
    .Y(_17435_));
 INVx1_ASAP7_75t_R _30112_ (.A(_18311_),
    .Y(_17434_));
 INVx1_ASAP7_75t_R _30113_ (.A(_18289_),
    .Y(_17383_));
 INVx1_ASAP7_75t_R _30114_ (.A(_18342_),
    .Y(_17482_));
 INVx1_ASAP7_75t_R _30115_ (.A(_18298_),
    .Y(_17454_));
 INVx1_ASAP7_75t_R _30116_ (.A(_18321_),
    .Y(_17453_));
 INVx1_ASAP7_75t_R _30117_ (.A(_18328_),
    .Y(_17511_));
 INVx1_ASAP7_75t_R _30118_ (.A(_18351_),
    .Y(_17510_));
 INVx1_ASAP7_75t_R _30119_ (.A(_18344_),
    .Y(_17542_));
 INVx1_ASAP7_75t_R _30120_ (.A(_00148_),
    .Y(_17140_));
 INVx1_ASAP7_75t_R _30121_ (.A(_00156_),
    .Y(_17139_));
 INVx1_ASAP7_75t_R _30122_ (.A(_18157_),
    .Y(_17134_));
 INVx1_ASAP7_75t_R _30123_ (.A(_18171_),
    .Y(_17133_));
 INVx1_ASAP7_75t_R _30124_ (.A(_02264_),
    .Y(_18175_));
 INVx1_ASAP7_75t_R _30125_ (.A(_00183_),
    .Y(_18244_));
 INVx1_ASAP7_75t_R _30126_ (.A(_02270_),
    .Y(_18243_));
 INVx1_ASAP7_75t_R _30127_ (.A(_00191_),
    .Y(_18267_));
 INVx1_ASAP7_75t_R _30128_ (.A(_02273_),
    .Y(_17411_));
 INVx1_ASAP7_75t_R _30129_ (.A(_00124_),
    .Y(_17063_));
 INVx1_ASAP7_75t_R _30130_ (.A(_18164_),
    .Y(_17117_));
 INVx1_ASAP7_75t_R _30131_ (.A(_18188_),
    .Y(_17173_));
 INVx1_ASAP7_75t_R _30132_ (.A(_00245_),
    .Y(_17972_));
 INVx1_ASAP7_75t_R _30133_ (.A(_02289_),
    .Y(_17992_));
 INVx1_ASAP7_75t_R _30134_ (.A(_17562_),
    .Y(_17513_));
 INVx1_ASAP7_75t_R _30135_ (.A(_18303_),
    .Y(_17410_));
 INVx1_ASAP7_75t_R _30136_ (.A(_18239_),
    .Y(_17304_));
 INVx1_ASAP7_75t_R _30137_ (.A(_18255_),
    .Y(_17303_));
 INVx1_ASAP7_75t_R _30138_ (.A(_18257_),
    .Y(_17355_));
 INVx1_ASAP7_75t_R _30139_ (.A(_18280_),
    .Y(_17354_));
 INVx1_ASAP7_75t_R _30140_ (.A(_18233_),
    .Y(_17294_));
 INVx1_ASAP7_75t_R _30141_ (.A(_18251_),
    .Y(_17293_));
 INVx1_ASAP7_75t_R _30142_ (.A(_18230_),
    .Y(_17287_));
 INVx1_ASAP7_75t_R _30143_ (.A(_18250_),
    .Y(_17286_));
 INVx1_ASAP7_75t_R _30144_ (.A(_18252_),
    .Y(_17341_));
 INVx1_ASAP7_75t_R _30145_ (.A(_18279_),
    .Y(_17340_));
 INVx1_ASAP7_75t_R _30146_ (.A(_18281_),
    .Y(_17397_));
 INVx1_ASAP7_75t_R _30147_ (.A(_18302_),
    .Y(_17396_));
 INVx1_ASAP7_75t_R _30148_ (.A(_18304_),
    .Y(_17463_));
 INVx1_ASAP7_75t_R _30149_ (.A(_18329_),
    .Y(_17462_));
 INVx1_ASAP7_75t_R _30150_ (.A(_18211_),
    .Y(_17244_));
 INVx1_ASAP7_75t_R _30151_ (.A(_18228_),
    .Y(_17243_));
 INVx1_ASAP7_75t_R _30152_ (.A(_18232_),
    .Y(_17289_));
 INVx1_ASAP7_75t_R _30153_ (.A(_18247_),
    .Y(_17288_));
 INVx1_ASAP7_75t_R _30154_ (.A(_18254_),
    .Y(_17343_));
 INVx1_ASAP7_75t_R _30155_ (.A(_18274_),
    .Y(_17342_));
 INVx1_ASAP7_75t_R _30156_ (.A(_18283_),
    .Y(_17399_));
 INVx1_ASAP7_75t_R _30157_ (.A(_18297_),
    .Y(_17398_));
 INVx1_ASAP7_75t_R _30158_ (.A(_18306_),
    .Y(_17465_));
 INVx1_ASAP7_75t_R _30159_ (.A(_18327_),
    .Y(_17464_));
 INVx1_ASAP7_75t_R _30160_ (.A(_18299_),
    .Y(_17459_));
 INVx1_ASAP7_75t_R _30161_ (.A(_18324_),
    .Y(_17458_));
 INVx1_ASAP7_75t_R _30162_ (.A(_18220_),
    .Y(_17264_));
 INVx1_ASAP7_75t_R _30163_ (.A(_18238_),
    .Y(_17263_));
 INVx1_ASAP7_75t_R _30164_ (.A(_18259_),
    .Y(_17310_));
 INVx1_ASAP7_75t_R _30165_ (.A(_18214_),
    .Y(_17255_));
 INVx1_ASAP7_75t_R _30166_ (.A(_18234_),
    .Y(_17254_));
 INVx1_ASAP7_75t_R _30167_ (.A(_18235_),
    .Y(_17297_));
 INVx1_ASAP7_75t_R _30168_ (.A(_18258_),
    .Y(_17296_));
 INVx1_ASAP7_75t_R _30169_ (.A(_18260_),
    .Y(_17356_));
 INVx1_ASAP7_75t_R _30170_ (.A(_18189_),
    .Y(_17212_));
 INVx1_ASAP7_75t_R _30171_ (.A(_18210_),
    .Y(_17211_));
 INVx1_ASAP7_75t_R _30172_ (.A(_18213_),
    .Y(_17250_));
 INVx1_ASAP7_75t_R _30173_ (.A(_18231_),
    .Y(_17249_));
 INVx1_ASAP7_75t_R _30174_ (.A(_18237_),
    .Y(_17299_));
 INVx1_ASAP7_75t_R _30175_ (.A(_18253_),
    .Y(_17298_));
 INVx1_ASAP7_75t_R _30176_ (.A(_18262_),
    .Y(_17358_));
 INVx1_ASAP7_75t_R _30177_ (.A(_18282_),
    .Y(_17357_));
 INVx1_ASAP7_75t_R _30178_ (.A(_18305_),
    .Y(_17415_));
 INVx1_ASAP7_75t_R _30179_ (.A(_18300_),
    .Y(_17403_));
 INVx1_ASAP7_75t_R _30180_ (.A(_18192_),
    .Y(_17223_));
 INVx1_ASAP7_75t_R _30181_ (.A(_18215_),
    .Y(_17222_));
 INVx1_ASAP7_75t_R _30182_ (.A(_18216_),
    .Y(_17257_));
 INVx1_ASAP7_75t_R _30183_ (.A(_18191_),
    .Y(_17218_));
 INVx1_ASAP7_75t_R _30184_ (.A(_18212_),
    .Y(_17217_));
 INVx1_ASAP7_75t_R _30185_ (.A(_18218_),
    .Y(_17259_));
 INVx1_ASAP7_75t_R _30186_ (.A(_18236_),
    .Y(_17258_));
 INVx1_ASAP7_75t_R _30187_ (.A(_18241_),
    .Y(_17317_));
 INVx1_ASAP7_75t_R _30188_ (.A(_18261_),
    .Y(_17316_));
 INVx1_ASAP7_75t_R _30189_ (.A(_02259_),
    .Y(_18160_));
 INVx1_ASAP7_75t_R _30190_ (.A(_00147_),
    .Y(_18161_));
 INVx1_ASAP7_75t_R _30191_ (.A(_00154_),
    .Y(_18174_));
 INVx1_ASAP7_75t_R _30192_ (.A(_02262_),
    .Y(_17199_));
 INVx1_ASAP7_75t_R _30193_ (.A(_18194_),
    .Y(_17225_));
 INVx1_ASAP7_75t_R _30194_ (.A(_18196_),
    .Y(_17227_));
 INVx1_ASAP7_75t_R _30195_ (.A(_18217_),
    .Y(_17226_));
 INVx1_ASAP7_75t_R _30196_ (.A(_18221_),
    .Y(_17276_));
 INVx1_ASAP7_75t_R _30197_ (.A(_18240_),
    .Y(_17275_));
 INVx1_ASAP7_75t_R _30198_ (.A(_00188_),
    .Y(_17308_));
 INVx1_ASAP7_75t_R _30199_ (.A(_18198_),
    .Y(_17232_));
 INVx1_ASAP7_75t_R _30200_ (.A(_18219_),
    .Y(_17231_));
 INVx1_ASAP7_75t_R _30201_ (.A(_18202_),
    .Y(_17234_));
 INVx1_ASAP7_75t_R _30202_ (.A(_18204_),
    .Y(_17236_));
 INVx1_ASAP7_75t_R _30203_ (.A(_18185_),
    .Y(_17190_));
 INVx1_ASAP7_75t_R _30204_ (.A(_18195_),
    .Y(_17189_));
 INVx1_ASAP7_75t_R _30205_ (.A(_18206_),
    .Y(_17238_));
 INVx1_ASAP7_75t_R _30206_ (.A(_18222_),
    .Y(_17237_));
 INVx1_ASAP7_75t_R _30207_ (.A(_00182_),
    .Y(_17268_));
 INVx1_ASAP7_75t_R _30208_ (.A(_18205_),
    .Y(_17202_));
 INVx1_ASAP7_75t_R _30209_ (.A(_00163_),
    .Y(_17207_));
 AND2x6_ASAP7_75t_R _30210_ (.A(_05460_),
    .B(_05715_),
    .Y(_12959_));
 AND5x2_ASAP7_75t_R _30211_ (.A(_12246_),
    .B(_00261_),
    .C(_05180_),
    .D(_05728_),
    .E(_02206_),
    .Y(_12960_));
 OA211x2_ASAP7_75t_R _30212_ (.A1(_05154_),
    .A2(_10838_),
    .B(_10839_),
    .C(_12960_),
    .Y(_12961_));
 NAND2x1_ASAP7_75t_R _30213_ (.A(_12959_),
    .B(_12961_),
    .Y(core_busy_d));
 AND2x2_ASAP7_75t_R _30214_ (.A(clknet_1_0__leaf_clk_i),
    .B(\core_clock_gate_i.en_latch ),
    .Y(clk));
 BUFx6f_ASAP7_75t_R _30215_ (.A(_05209_),
    .Y(_12962_));
 AND2x2_ASAP7_75t_R _30216_ (.A(_14117_),
    .B(_02324_),
    .Y(_12963_));
 AO21x1_ASAP7_75t_R _30217_ (.A1(_14273_),
    .A2(_12962_),
    .B(_12963_),
    .Y(_12964_));
 NAND2x1_ASAP7_75t_R _30218_ (.A(_02325_),
    .B(_12304_),
    .Y(_12965_));
 OA21x2_ASAP7_75t_R _30219_ (.A1(_12304_),
    .A2(_12964_),
    .B(_12965_),
    .Y(net202));
 AND3x1_ASAP7_75t_R _30220_ (.A(_14112_),
    .B(_14273_),
    .C(_05730_),
    .Y(_12966_));
 BUFx6f_ASAP7_75t_R _30221_ (.A(_02327_),
    .Y(_12967_));
 BUFx6f_ASAP7_75t_R _30222_ (.A(_12303_),
    .Y(_12968_));
 AO21x1_ASAP7_75t_R _30223_ (.A1(_12967_),
    .A2(_12968_),
    .B(_12302_),
    .Y(_12969_));
 BUFx6f_ASAP7_75t_R _30224_ (.A(_02328_),
    .Y(_12970_));
 AO21x1_ASAP7_75t_R _30225_ (.A1(_05208_),
    .A2(_12970_),
    .B(_13255_),
    .Y(_12971_));
 OA211x2_ASAP7_75t_R _30226_ (.A1(_18707_),
    .A2(_12969_),
    .B(_12971_),
    .C(_05739_),
    .Y(_12972_));
 AOI21x1_ASAP7_75t_R _30227_ (.A1(_00335_),
    .A2(_12966_),
    .B(_12972_),
    .Y(net203));
 OR3x1_ASAP7_75t_R _30228_ (.A(_00338_),
    .B(_14273_),
    .C(_12304_),
    .Y(_12973_));
 INVx1_ASAP7_75t_R _30229_ (.A(_12973_),
    .Y(_12974_));
 AO21x1_ASAP7_75t_R _30230_ (.A1(_00336_),
    .A2(_12304_),
    .B(_12974_),
    .Y(_12975_));
 INVx1_ASAP7_75t_R _30231_ (.A(_12303_),
    .Y(_12976_));
 BUFx6f_ASAP7_75t_R _30232_ (.A(_12976_),
    .Y(_12977_));
 INVx1_ASAP7_75t_R _30233_ (.A(_00337_),
    .Y(_12978_));
 AO32x1_ASAP7_75t_R _30234_ (.A1(_13255_),
    .A2(_12977_),
    .A3(_12304_),
    .B1(_12966_),
    .B2(_12978_),
    .Y(_12979_));
 AO21x2_ASAP7_75t_R _30235_ (.A1(_18707_),
    .A2(_12975_),
    .B(_12979_),
    .Y(net204));
 BUFx6f_ASAP7_75t_R _30236_ (.A(_02327_),
    .Y(_12980_));
 BUFx6f_ASAP7_75t_R _30237_ (.A(_12303_),
    .Y(_12981_));
 OA211x2_ASAP7_75t_R _30238_ (.A1(_14273_),
    .A2(_12980_),
    .B(_12981_),
    .C(_12302_),
    .Y(_12982_));
 AOI21x1_ASAP7_75t_R _30239_ (.A1(_13255_),
    .A2(_05739_),
    .B(_12982_),
    .Y(net205));
 AO21x2_ASAP7_75t_R _30240_ (.A1(_12246_),
    .A2(_13253_),
    .B(_05731_),
    .Y(net206));
 BUFx6f_ASAP7_75t_R _30241_ (.A(_05208_),
    .Y(_12983_));
 BUFx6f_ASAP7_75t_R _30242_ (.A(_05208_),
    .Y(_12984_));
 BUFx6f_ASAP7_75t_R _30243_ (.A(_12970_),
    .Y(_12985_));
 OA222x2_ASAP7_75t_R _30244_ (.A1(_12980_),
    .A2(_15884_),
    .B1(_16871_),
    .B2(_12985_),
    .C1(_12981_),
    .C2(_04996_),
    .Y(_12986_));
 NAND2x1_ASAP7_75t_R _30245_ (.A(_12984_),
    .B(_12986_),
    .Y(_12987_));
 OA21x2_ASAP7_75t_R _30246_ (.A1(_12983_),
    .A2(_13420_),
    .B(_12987_),
    .Y(net207));
 BUFx12f_ASAP7_75t_R _30247_ (.A(_12962_),
    .Y(_12988_));
 INVx3_ASAP7_75t_R _30248_ (.A(_12970_),
    .Y(_12989_));
 INVx1_ASAP7_75t_R _30249_ (.A(_02327_),
    .Y(_12990_));
 BUFx6f_ASAP7_75t_R _30250_ (.A(_12990_),
    .Y(_12991_));
 AOI22x1_ASAP7_75t_R _30251_ (.A1(_12989_),
    .A2(_13601_),
    .B1(_04357_),
    .B2(_12991_),
    .Y(_12992_));
 BUFx6f_ASAP7_75t_R _30252_ (.A(_05208_),
    .Y(_12993_));
 OA211x2_ASAP7_75t_R _30253_ (.A1(_12981_),
    .A2(net1965),
    .B(_12992_),
    .C(_12993_),
    .Y(_12994_));
 AOI21x1_ASAP7_75t_R _30254_ (.A1(_12988_),
    .A2(_05002_),
    .B(_12994_),
    .Y(net208));
 OA222x2_ASAP7_75t_R _30255_ (.A1(_12970_),
    .A2(_05572_),
    .B1(_16242_),
    .B2(_12968_),
    .C1(_04468_),
    .C2(_02327_),
    .Y(_12995_));
 NOR2x1_ASAP7_75t_R _30256_ (.A(_12962_),
    .B(_12995_),
    .Y(_12996_));
 AO21x2_ASAP7_75t_R _30257_ (.A1(_12962_),
    .A2(_14260_),
    .B(_12996_),
    .Y(net209));
 AO222x2_ASAP7_75t_R _30258_ (.A1(_12989_),
    .A2(_13762_),
    .B1(_16384_),
    .B2(_12977_),
    .C1(_04605_),
    .C2(_12991_),
    .Y(_12997_));
 AND3x1_ASAP7_75t_R _30259_ (.A(_05209_),
    .B(_15315_),
    .C(_15362_),
    .Y(_12998_));
 AO21x2_ASAP7_75t_R _30260_ (.A1(_12984_),
    .A2(_12997_),
    .B(_12998_),
    .Y(net210));
 AO222x2_ASAP7_75t_R _30261_ (.A1(_12989_),
    .A2(_13830_),
    .B1(_16498_),
    .B2(_12977_),
    .C1(_04717_),
    .C2(_12991_),
    .Y(_12999_));
 AND3x1_ASAP7_75t_R _30262_ (.A(_05209_),
    .B(_15465_),
    .C(_15501_),
    .Y(_13000_));
 AO21x2_ASAP7_75t_R _30263_ (.A1(_12984_),
    .A2(_12999_),
    .B(_13000_),
    .Y(net211));
 AO33x2_ASAP7_75t_R _30264_ (.A1(_12976_),
    .A2(_16613_),
    .A3(_16636_),
    .B1(_04813_),
    .B2(_04836_),
    .B3(_12990_),
    .Y(_13001_));
 AO21x1_ASAP7_75t_R _30265_ (.A1(_12989_),
    .A2(_13908_),
    .B(_13001_),
    .Y(_13002_));
 BUFx6f_ASAP7_75t_R _30266_ (.A(_05208_),
    .Y(_13003_));
 NOR2x1_ASAP7_75t_R _30267_ (.A(_13003_),
    .B(net1946),
    .Y(_13004_));
 AO21x2_ASAP7_75t_R _30268_ (.A1(_12984_),
    .A2(_13002_),
    .B(_13004_),
    .Y(net212));
 AOI22x1_ASAP7_75t_R _30269_ (.A1(_12989_),
    .A2(_13968_),
    .B1(_04963_),
    .B2(_12991_),
    .Y(_13005_));
 OA211x2_ASAP7_75t_R _30270_ (.A1(_12981_),
    .A2(_16747_),
    .B(_13005_),
    .C(_12993_),
    .Y(_13006_));
 AOI21x1_ASAP7_75t_R _30271_ (.A1(_12988_),
    .A2(_15759_),
    .B(_13006_),
    .Y(net213));
 OA222x2_ASAP7_75t_R _30272_ (.A1(_12980_),
    .A2(_10872_),
    .B1(_04996_),
    .B2(_12985_),
    .C1(_16871_),
    .C2(_12968_),
    .Y(_13007_));
 NAND2x1_ASAP7_75t_R _30273_ (.A(_12984_),
    .B(_13007_),
    .Y(_13008_));
 OA21x2_ASAP7_75t_R _30274_ (.A1(_12983_),
    .A2(_05261_),
    .B(_13008_),
    .Y(net214));
 AO222x2_ASAP7_75t_R _30275_ (.A1(_12991_),
    .A2(_05354_),
    .B1(_14089_),
    .B2(_12989_),
    .C1(_16983_),
    .C2(_12977_),
    .Y(_13009_));
 NOR2x1_ASAP7_75t_R _30276_ (.A(_12993_),
    .B(_15995_),
    .Y(_13010_));
 AO21x2_ASAP7_75t_R _30277_ (.A1(_12984_),
    .A2(_13009_),
    .B(_13010_),
    .Y(net215));
 BUFx6f_ASAP7_75t_R _30278_ (.A(_12970_),
    .Y(_13011_));
 AOI22x1_ASAP7_75t_R _30279_ (.A1(_12991_),
    .A2(_13601_),
    .B1(_04357_),
    .B2(_12977_),
    .Y(_13012_));
 OA211x2_ASAP7_75t_R _30280_ (.A1(_13011_),
    .A2(_05002_),
    .B(_13012_),
    .C(_12993_),
    .Y(_13013_));
 AOI21x1_ASAP7_75t_R _30281_ (.A1(_12988_),
    .A2(net1965),
    .B(_13013_),
    .Y(net216));
 INVx1_ASAP7_75t_R _30282_ (.A(_14260_),
    .Y(_13014_));
 OA222x2_ASAP7_75t_R _30283_ (.A1(_12980_),
    .A2(_05572_),
    .B1(_13014_),
    .B2(_13011_),
    .C1(_04468_),
    .C2(_12981_),
    .Y(_13015_));
 OR2x2_ASAP7_75t_R _30284_ (.A(_12993_),
    .B(_16242_),
    .Y(_13016_));
 OAI21x1_ASAP7_75t_R _30285_ (.A1(_12988_),
    .A2(_13015_),
    .B(_13016_),
    .Y(net217));
 NOR2x1_ASAP7_75t_R _30286_ (.A(_12967_),
    .B(_15995_),
    .Y(_13017_));
 AO221x1_ASAP7_75t_R _30287_ (.A1(_12977_),
    .A2(_14089_),
    .B1(_16983_),
    .B2(_12989_),
    .C(_13017_),
    .Y(_13018_));
 AND2x2_ASAP7_75t_R _30288_ (.A(_05209_),
    .B(_05354_),
    .Y(_13019_));
 AO21x2_ASAP7_75t_R _30289_ (.A1(_12984_),
    .A2(_13018_),
    .B(_13019_),
    .Y(net218));
 OA222x2_ASAP7_75t_R _30290_ (.A1(_12980_),
    .A2(_05578_),
    .B1(_15363_),
    .B2(_12985_),
    .C1(_04606_),
    .C2(_12968_),
    .Y(_13020_));
 NAND2x1_ASAP7_75t_R _30291_ (.A(_13003_),
    .B(_13020_),
    .Y(_13021_));
 OA21x2_ASAP7_75t_R _30292_ (.A1(_12983_),
    .A2(_16384_),
    .B(_13021_),
    .Y(net219));
 INVx1_ASAP7_75t_R _30293_ (.A(_13830_),
    .Y(_13022_));
 OA222x2_ASAP7_75t_R _30294_ (.A1(_12980_),
    .A2(_13022_),
    .B1(_15502_),
    .B2(_12985_),
    .C1(_04718_),
    .C2(_12968_),
    .Y(_13023_));
 NAND2x1_ASAP7_75t_R _30295_ (.A(_13003_),
    .B(_13023_),
    .Y(_13024_));
 OA21x2_ASAP7_75t_R _30296_ (.A1(_12983_),
    .A2(_16498_),
    .B(_13024_),
    .Y(net220));
 OAI22x1_ASAP7_75t_R _30297_ (.A1(_13011_),
    .A2(net1946),
    .B1(_04837_),
    .B2(_12981_),
    .Y(_13025_));
 AO21x1_ASAP7_75t_R _30298_ (.A1(_12991_),
    .A2(_13908_),
    .B(_13025_),
    .Y(_13026_));
 AND3x1_ASAP7_75t_R _30299_ (.A(_05209_),
    .B(_16613_),
    .C(_16636_),
    .Y(_13027_));
 AO21x2_ASAP7_75t_R _30300_ (.A1(_12984_),
    .A2(_13026_),
    .B(_13027_),
    .Y(net221));
 AOI22x1_ASAP7_75t_R _30301_ (.A1(_12991_),
    .A2(_13968_),
    .B1(_04963_),
    .B2(_12977_),
    .Y(_13028_));
 OA211x2_ASAP7_75t_R _30302_ (.A1(_13011_),
    .A2(_15759_),
    .B(_13028_),
    .C(_12993_),
    .Y(_13029_));
 AOI21x1_ASAP7_75t_R _30303_ (.A1(_12988_),
    .A2(_16747_),
    .B(_13029_),
    .Y(net222));
 OA222x2_ASAP7_75t_R _30304_ (.A1(_12967_),
    .A2(_04996_),
    .B1(_15884_),
    .B2(_12970_),
    .C1(_12303_),
    .C2(_10872_),
    .Y(_13030_));
 NOR2x1_ASAP7_75t_R _30305_ (.A(_12962_),
    .B(_13030_),
    .Y(_13031_));
 AO21x2_ASAP7_75t_R _30306_ (.A1(_12962_),
    .A2(_16870_),
    .B(_13031_),
    .Y(net223));
 AOI22x1_ASAP7_75t_R _30307_ (.A1(_12977_),
    .A2(_05354_),
    .B1(_14089_),
    .B2(_12991_),
    .Y(_13032_));
 OA211x2_ASAP7_75t_R _30308_ (.A1(_13011_),
    .A2(_15995_),
    .B(_13032_),
    .C(_12993_),
    .Y(_13033_));
 AOI21x1_ASAP7_75t_R _30309_ (.A1(_12988_),
    .A2(_16984_),
    .B(_13033_),
    .Y(net224));
 AOI22x1_ASAP7_75t_R _30310_ (.A1(_12977_),
    .A2(_13601_),
    .B1(_14201_),
    .B2(_12991_),
    .Y(_13034_));
 OA211x2_ASAP7_75t_R _30311_ (.A1(_13011_),
    .A2(net1965),
    .B(_13034_),
    .C(_12993_),
    .Y(_13035_));
 AOI21x1_ASAP7_75t_R _30312_ (.A1(_12988_),
    .A2(_04358_),
    .B(_13035_),
    .Y(net225));
 OA222x2_ASAP7_75t_R _30313_ (.A1(_12980_),
    .A2(_13014_),
    .B1(_16242_),
    .B2(_13011_),
    .C1(_12981_),
    .C2(_05572_),
    .Y(_13036_));
 OR2x2_ASAP7_75t_R _30314_ (.A(_12993_),
    .B(_04468_),
    .Y(_13037_));
 OAI21x1_ASAP7_75t_R _30315_ (.A1(_12988_),
    .A2(_13036_),
    .B(_13037_),
    .Y(net226));
 OA222x2_ASAP7_75t_R _30316_ (.A1(_12980_),
    .A2(_15363_),
    .B1(_16385_),
    .B2(_12985_),
    .C1(_12981_),
    .C2(_05578_),
    .Y(_13038_));
 NAND2x1_ASAP7_75t_R _30317_ (.A(_13003_),
    .B(_13038_),
    .Y(_13039_));
 OA21x2_ASAP7_75t_R _30318_ (.A1(_12983_),
    .A2(_04605_),
    .B(_13039_),
    .Y(net227));
 OA222x2_ASAP7_75t_R _30319_ (.A1(_12967_),
    .A2(_15502_),
    .B1(_16499_),
    .B2(_12985_),
    .C1(_12968_),
    .C2(_13022_),
    .Y(_13040_));
 NAND2x1_ASAP7_75t_R _30320_ (.A(_13003_),
    .B(_13040_),
    .Y(_13041_));
 OA21x2_ASAP7_75t_R _30321_ (.A1(_12983_),
    .A2(_04717_),
    .B(_13041_),
    .Y(net228));
 OA222x2_ASAP7_75t_R _30322_ (.A1(_12967_),
    .A2(net1965),
    .B1(_04358_),
    .B2(_12985_),
    .C1(_12968_),
    .C2(_05002_),
    .Y(_13042_));
 NAND2x1_ASAP7_75t_R _30323_ (.A(_13003_),
    .B(_13042_),
    .Y(_13043_));
 OA21x2_ASAP7_75t_R _30324_ (.A1(_12983_),
    .A2(_13601_),
    .B(_13043_),
    .Y(net229));
 OAI22x1_ASAP7_75t_R _30325_ (.A1(_12980_),
    .A2(net1946),
    .B1(_16637_),
    .B2(_13011_),
    .Y(_13044_));
 AO21x1_ASAP7_75t_R _30326_ (.A1(_12977_),
    .A2(_13908_),
    .B(_13044_),
    .Y(_13045_));
 AND3x1_ASAP7_75t_R _30327_ (.A(_05209_),
    .B(_04813_),
    .C(_04836_),
    .Y(_13046_));
 AO21x2_ASAP7_75t_R _30328_ (.A1(_12984_),
    .A2(_13045_),
    .B(_13046_),
    .Y(net230));
 INVx1_ASAP7_75t_R _30329_ (.A(_04963_),
    .Y(_13047_));
 OA22x2_ASAP7_75t_R _30330_ (.A1(_12303_),
    .A2(_05038_),
    .B1(_15759_),
    .B2(_02327_),
    .Y(_13048_));
 OA211x2_ASAP7_75t_R _30331_ (.A1(_13011_),
    .A2(_16747_),
    .B(_13048_),
    .C(_05208_),
    .Y(_13049_));
 AOI21x1_ASAP7_75t_R _30332_ (.A1(_12988_),
    .A2(_13047_),
    .B(_13049_),
    .Y(net231));
 OA222x2_ASAP7_75t_R _30333_ (.A1(_12967_),
    .A2(_16242_),
    .B1(_04468_),
    .B2(_12985_),
    .C1(_12968_),
    .C2(_13014_),
    .Y(_13050_));
 NAND2x1_ASAP7_75t_R _30334_ (.A(_13003_),
    .B(_13050_),
    .Y(_13051_));
 OA21x2_ASAP7_75t_R _30335_ (.A1(_12983_),
    .A2(_13684_),
    .B(_13051_),
    .Y(net232));
 OA222x2_ASAP7_75t_R _30336_ (.A1(_12967_),
    .A2(_16385_),
    .B1(_04606_),
    .B2(_12985_),
    .C1(_12968_),
    .C2(_15363_),
    .Y(_13052_));
 NAND2x1_ASAP7_75t_R _30337_ (.A(_13003_),
    .B(_13052_),
    .Y(_13053_));
 OA21x2_ASAP7_75t_R _30338_ (.A1(_12983_),
    .A2(_13762_),
    .B(_13053_),
    .Y(net233));
 OA222x2_ASAP7_75t_R _30339_ (.A1(_12967_),
    .A2(_16499_),
    .B1(_04718_),
    .B2(_12970_),
    .C1(_12968_),
    .C2(_15502_),
    .Y(_13054_));
 NAND2x1_ASAP7_75t_R _30340_ (.A(_13003_),
    .B(_13054_),
    .Y(_13055_));
 OA21x2_ASAP7_75t_R _30341_ (.A1(_12983_),
    .A2(_13830_),
    .B(_13055_),
    .Y(net234));
 OA222x2_ASAP7_75t_R _30342_ (.A1(_12967_),
    .A2(_16637_),
    .B1(_04837_),
    .B2(_12970_),
    .C1(_12303_),
    .C2(_15646_),
    .Y(_13056_));
 NOR2x1_ASAP7_75t_R _30343_ (.A(_12962_),
    .B(_13056_),
    .Y(_13057_));
 AO21x2_ASAP7_75t_R _30344_ (.A1(_12962_),
    .A2(_13908_),
    .B(_13057_),
    .Y(net235));
 OA222x2_ASAP7_75t_R _30345_ (.A1(_02327_),
    .A2(_16747_),
    .B1(_13047_),
    .B2(_12970_),
    .C1(_12303_),
    .C2(_15759_),
    .Y(_13058_));
 NOR2x1_ASAP7_75t_R _30346_ (.A(_12962_),
    .B(_13058_),
    .Y(_13059_));
 AO21x2_ASAP7_75t_R _30347_ (.A1(_12962_),
    .A2(_13968_),
    .B(_13059_),
    .Y(net236));
 OA222x2_ASAP7_75t_R _30348_ (.A1(_13011_),
    .A2(_10872_),
    .B1(_15884_),
    .B2(_12981_),
    .C1(_16871_),
    .C2(_12980_),
    .Y(_13060_));
 OR3x2_ASAP7_75t_R _30349_ (.A(_12993_),
    .B(_05059_),
    .C(_05064_),
    .Y(_13061_));
 OAI21x1_ASAP7_75t_R _30350_ (.A1(_12988_),
    .A2(_13060_),
    .B(_13061_),
    .Y(net237));
 OA222x2_ASAP7_75t_R _30351_ (.A1(_12985_),
    .A2(_05556_),
    .B1(_15995_),
    .B2(_12981_),
    .C1(_16984_),
    .C2(_12967_),
    .Y(_13062_));
 NAND2x1_ASAP7_75t_R _30352_ (.A(_13003_),
    .B(_13062_),
    .Y(_13063_));
 OA21x2_ASAP7_75t_R _30353_ (.A1(_12984_),
    .A2(_14089_),
    .B(_13063_),
    .Y(net238));
 NOR2x1_ASAP7_75t_R _30354_ (.A(_06883_),
    .B(_07156_),
    .Y(\id_stage_i.branch_set_d ));
 INVx1_ASAP7_75t_R _30355_ (.A(net149),
    .Y(_13064_));
 AO21x1_ASAP7_75t_R _30356_ (.A1(_13064_),
    .A2(_05459_),
    .B(_02206_),
    .Y(_13065_));
 OA21x2_ASAP7_75t_R _30357_ (.A1(_00261_),
    .A2(_05459_),
    .B(_02203_),
    .Y(_13066_));
 AND2x4_ASAP7_75t_R _30358_ (.A(net149),
    .B(_05709_),
    .Y(_13067_));
 AOI22x1_ASAP7_75t_R _30359_ (.A1(_02202_),
    .A2(_13065_),
    .B1(_13066_),
    .B2(_13067_),
    .Y(_13068_));
 AO21x1_ASAP7_75t_R _30360_ (.A1(net116),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .B(_13068_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ));
 NAND3x1_ASAP7_75t_R _30361_ (.A(net116),
    .B(_05709_),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .Y(_13069_));
 AOI21x1_ASAP7_75t_R _30362_ (.A1(_13066_),
    .A2(_13069_),
    .B(_13067_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ));
 NAND2x1_ASAP7_75t_R _30363_ (.A(_10809_),
    .B(_11737_),
    .Y(_13070_));
 AO21x1_ASAP7_75t_R _30364_ (.A1(_11728_),
    .A2(_13070_),
    .B(_11738_),
    .Y(_13071_));
 NAND2x1_ASAP7_75t_R _30365_ (.A(_11730_),
    .B(_11760_),
    .Y(_13072_));
 OA211x2_ASAP7_75t_R _30366_ (.A1(_11747_),
    .A2(_13071_),
    .B(_13072_),
    .C(_11475_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ));
 OR3x1_ASAP7_75t_R _30367_ (.A(_10825_),
    .B(_11728_),
    .C(_11741_),
    .Y(_13073_));
 AO221x1_ASAP7_75t_R _30368_ (.A1(_13070_),
    .A2(_11748_),
    .B1(_13073_),
    .B2(_11935_),
    .C(_11774_),
    .Y(_13074_));
 AND2x2_ASAP7_75t_R _30369_ (.A(_11788_),
    .B(_13074_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ));
 AND3x1_ASAP7_75t_R _30370_ (.A(_11475_),
    .B(_13070_),
    .C(_11761_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ));
 INVx2_ASAP7_75t_R _30371_ (.A(_12959_),
    .Y(net270));
 OA21x2_ASAP7_75t_R _30372_ (.A1(_05714_),
    .A2(_13064_),
    .B(_05709_),
    .Y(_13075_));
 AO21x1_ASAP7_75t_R _30373_ (.A1(net116),
    .A2(net270),
    .B(_13075_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ));
 OR3x1_ASAP7_75t_R _30374_ (.A(_12177_),
    .B(_02206_),
    .C(_12959_),
    .Y(_13076_));
 AOI21x1_ASAP7_75t_R _30375_ (.A1(_00261_),
    .A2(_13076_),
    .B(_13067_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ));
 AND2x2_ASAP7_75t_R _30376_ (.A(_12177_),
    .B(net270),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ));
 INVx1_ASAP7_75t_R _30377_ (.A(_10864_),
    .Y(_13077_));
 OR3x1_ASAP7_75t_R _30378_ (.A(_13233_),
    .B(_10839_),
    .C(_13077_),
    .Y(_13078_));
 AOI21x1_ASAP7_75t_R _30379_ (.A1(_05406_),
    .A2(_05417_),
    .B(_13078_),
    .Y(_13079_));
 OA21x2_ASAP7_75t_R _30380_ (.A1(_11846_),
    .A2(_10851_),
    .B(_13079_),
    .Y(_13080_));
 AO21x1_ASAP7_75t_R _30381_ (.A1(_11803_),
    .A2(_11785_),
    .B(_13080_),
    .Y(\if_stage_i.instr_valid_id_d ));
 INVx6_ASAP7_75t_R _30382_ (.A(_00340_),
    .Y(_13081_));
 BUFx6f_ASAP7_75t_R _30383_ (.A(_13081_),
    .Y(_13082_));
 INVx2_ASAP7_75t_R _30384_ (.A(_00341_),
    .Y(_13083_));
 BUFx12f_ASAP7_75t_R _30385_ (.A(_13083_),
    .Y(_13084_));
 BUFx12f_ASAP7_75t_R _30386_ (.A(_13084_),
    .Y(_13085_));
 BUFx6f_ASAP7_75t_R _30387_ (.A(_13085_),
    .Y(_13086_));
 BUFx12f_ASAP7_75t_R _30388_ (.A(_00344_),
    .Y(_13087_));
 BUFx12f_ASAP7_75t_R _30389_ (.A(_13087_),
    .Y(_13088_));
 BUFx12f_ASAP7_75t_R _30390_ (.A(_13088_),
    .Y(_13089_));
 BUFx12f_ASAP7_75t_R _30391_ (.A(_13089_),
    .Y(_13090_));
 INVx4_ASAP7_75t_R _30392_ (.A(_00343_),
    .Y(_13091_));
 BUFx6f_ASAP7_75t_R _30393_ (.A(_13091_),
    .Y(_13092_));
 BUFx12f_ASAP7_75t_R _30394_ (.A(_00343_),
    .Y(_13093_));
 BUFx12f_ASAP7_75t_R _30395_ (.A(_13093_),
    .Y(_13094_));
 BUFx12f_ASAP7_75t_R _30396_ (.A(_13094_),
    .Y(_13095_));
 BUFx12f_ASAP7_75t_R _30397_ (.A(_13095_),
    .Y(_13096_));
 BUFx12f_ASAP7_75t_R _30398_ (.A(_13096_),
    .Y(_13097_));
 AND2x2_ASAP7_75t_R _30399_ (.A(_13097_),
    .B(_01784_),
    .Y(_13098_));
 AO21x1_ASAP7_75t_R _30400_ (.A1(_00346_),
    .A2(_13092_),
    .B(_13098_),
    .Y(_13099_));
 BUFx12f_ASAP7_75t_R _30401_ (.A(_13087_),
    .Y(_13100_));
 NAND2x2_ASAP7_75t_R _30402_ (.A(_13100_),
    .B(_13091_),
    .Y(_13101_));
 BUFx12f_ASAP7_75t_R _30403_ (.A(_13101_),
    .Y(_13102_));
 OAI22x1_ASAP7_75t_R _30404_ (.A1(_13090_),
    .A2(_13099_),
    .B1(_13102_),
    .B2(_00345_),
    .Y(_13103_));
 BUFx12f_ASAP7_75t_R _30405_ (.A(_00341_),
    .Y(_13104_));
 BUFx12f_ASAP7_75t_R _30406_ (.A(_13104_),
    .Y(_13105_));
 BUFx12f_ASAP7_75t_R _30407_ (.A(_13095_),
    .Y(_13106_));
 BUFx12f_ASAP7_75t_R _30408_ (.A(_13106_),
    .Y(_13107_));
 INVx2_ASAP7_75t_R _30409_ (.A(_00354_),
    .Y(_13108_));
 BUFx12f_ASAP7_75t_R _30410_ (.A(_13094_),
    .Y(_13109_));
 BUFx12f_ASAP7_75t_R _30411_ (.A(_13109_),
    .Y(_13110_));
 NAND2x1_ASAP7_75t_R _30412_ (.A(_13110_),
    .B(_00352_),
    .Y(_13111_));
 INVx2_ASAP7_75t_R _30413_ (.A(_00344_),
    .Y(_13112_));
 BUFx12f_ASAP7_75t_R _30414_ (.A(_13112_),
    .Y(_13113_));
 BUFx12f_ASAP7_75t_R _30415_ (.A(_13113_),
    .Y(_13114_));
 BUFx12f_ASAP7_75t_R _30416_ (.A(_13114_),
    .Y(_13115_));
 OA211x2_ASAP7_75t_R _30417_ (.A1(_13107_),
    .A2(_13108_),
    .B(_13111_),
    .C(_13115_),
    .Y(_13116_));
 INVx1_ASAP7_75t_R _30418_ (.A(_00353_),
    .Y(_13117_));
 BUFx12f_ASAP7_75t_R _30419_ (.A(_13109_),
    .Y(_13118_));
 NAND2x1_ASAP7_75t_R _30420_ (.A(_13118_),
    .B(_00351_),
    .Y(_13119_));
 BUFx12f_ASAP7_75t_R _30421_ (.A(_13100_),
    .Y(_13120_));
 OA211x2_ASAP7_75t_R _30422_ (.A1(_13107_),
    .A2(_13117_),
    .B(_13119_),
    .C(_13120_),
    .Y(_13121_));
 OR3x1_ASAP7_75t_R _30423_ (.A(_13105_),
    .B(_13116_),
    .C(_13121_),
    .Y(_13122_));
 BUFx6f_ASAP7_75t_R _30424_ (.A(_00342_),
    .Y(_13123_));
 BUFx12f_ASAP7_75t_R _30425_ (.A(_13123_),
    .Y(_13124_));
 BUFx12f_ASAP7_75t_R _30426_ (.A(_13124_),
    .Y(_13125_));
 OA211x2_ASAP7_75t_R _30427_ (.A1(_13086_),
    .A2(_13103_),
    .B(_13122_),
    .C(_13125_),
    .Y(_13126_));
 INVx2_ASAP7_75t_R _30428_ (.A(_13123_),
    .Y(_13127_));
 BUFx12f_ASAP7_75t_R _30429_ (.A(_13127_),
    .Y(_13128_));
 BUFx12f_ASAP7_75t_R _30430_ (.A(_13128_),
    .Y(_13129_));
 BUFx12f_ASAP7_75t_R _30431_ (.A(_13084_),
    .Y(_13130_));
 BUFx12f_ASAP7_75t_R _30432_ (.A(_13130_),
    .Y(_13131_));
 BUFx12f_ASAP7_75t_R _30433_ (.A(_13095_),
    .Y(_13132_));
 BUFx6f_ASAP7_75t_R _30434_ (.A(_13132_),
    .Y(_13133_));
 INVx2_ASAP7_75t_R _30435_ (.A(_00350_),
    .Y(_13134_));
 BUFx12f_ASAP7_75t_R _30436_ (.A(_13094_),
    .Y(_13135_));
 BUFx12f_ASAP7_75t_R _30437_ (.A(_13135_),
    .Y(_13136_));
 BUFx12f_ASAP7_75t_R _30438_ (.A(_13136_),
    .Y(_13137_));
 NAND2x1_ASAP7_75t_R _30439_ (.A(_13137_),
    .B(_00348_),
    .Y(_13138_));
 BUFx12f_ASAP7_75t_R _30440_ (.A(_13113_),
    .Y(_13139_));
 BUFx6f_ASAP7_75t_R _30441_ (.A(_13139_),
    .Y(_13140_));
 OA211x2_ASAP7_75t_R _30442_ (.A1(_13133_),
    .A2(_13134_),
    .B(_13138_),
    .C(_13140_),
    .Y(_13141_));
 BUFx12f_ASAP7_75t_R _30443_ (.A(_13109_),
    .Y(_13142_));
 BUFx6f_ASAP7_75t_R _30444_ (.A(_13142_),
    .Y(_13143_));
 INVx2_ASAP7_75t_R _30445_ (.A(_00349_),
    .Y(_13144_));
 BUFx12f_ASAP7_75t_R _30446_ (.A(_13094_),
    .Y(_13145_));
 BUFx12f_ASAP7_75t_R _30447_ (.A(_13145_),
    .Y(_13146_));
 NAND2x1_ASAP7_75t_R _30448_ (.A(_13146_),
    .B(_00347_),
    .Y(_13147_));
 BUFx12f_ASAP7_75t_R _30449_ (.A(_13087_),
    .Y(_13148_));
 BUFx12f_ASAP7_75t_R _30450_ (.A(_13148_),
    .Y(_13149_));
 OA211x2_ASAP7_75t_R _30451_ (.A1(_13143_),
    .A2(_13144_),
    .B(_13147_),
    .C(_13149_),
    .Y(_13150_));
 OR3x1_ASAP7_75t_R _30452_ (.A(_13131_),
    .B(_13141_),
    .C(_13150_),
    .Y(_13151_));
 BUFx12f_ASAP7_75t_R _30453_ (.A(_13104_),
    .Y(_13152_));
 BUFx12f_ASAP7_75t_R _30454_ (.A(_13152_),
    .Y(_13153_));
 INVx2_ASAP7_75t_R _30455_ (.A(_00358_),
    .Y(_13154_));
 NAND2x1_ASAP7_75t_R _30456_ (.A(_13146_),
    .B(_00356_),
    .Y(_13155_));
 OA211x2_ASAP7_75t_R _30457_ (.A1(_13143_),
    .A2(_13154_),
    .B(_13155_),
    .C(_13140_),
    .Y(_13156_));
 INVx2_ASAP7_75t_R _30458_ (.A(_00357_),
    .Y(_13157_));
 NAND2x1_ASAP7_75t_R _30459_ (.A(_13146_),
    .B(_00355_),
    .Y(_13158_));
 OA211x2_ASAP7_75t_R _30460_ (.A1(_13143_),
    .A2(_13157_),
    .B(_13158_),
    .C(_13149_),
    .Y(_13159_));
 OR3x1_ASAP7_75t_R _30461_ (.A(_13153_),
    .B(_13156_),
    .C(_13159_),
    .Y(_13160_));
 AND3x4_ASAP7_75t_R _30462_ (.A(_13129_),
    .B(_13151_),
    .C(_13160_),
    .Y(_13161_));
 OR3x2_ASAP7_75t_R _30463_ (.A(_13082_),
    .B(_13126_),
    .C(_13161_),
    .Y(_13162_));
 BUFx12f_ASAP7_75t_R _30464_ (.A(_00340_),
    .Y(_13163_));
 BUFx6f_ASAP7_75t_R _30465_ (.A(_13163_),
    .Y(_13164_));
 BUFx12f_ASAP7_75t_R _30466_ (.A(_13095_),
    .Y(_13165_));
 BUFx12f_ASAP7_75t_R _30467_ (.A(_13165_),
    .Y(_13166_));
 INVx2_ASAP7_75t_R _30468_ (.A(_00366_),
    .Y(_13167_));
 BUFx12f_ASAP7_75t_R _30469_ (.A(_13136_),
    .Y(_13168_));
 NAND2x1_ASAP7_75t_R _30470_ (.A(_13168_),
    .B(_00364_),
    .Y(_13169_));
 OA211x2_ASAP7_75t_R _30471_ (.A1(_13166_),
    .A2(_13167_),
    .B(_13169_),
    .C(_13140_),
    .Y(_13170_));
 INVx2_ASAP7_75t_R _30472_ (.A(_00365_),
    .Y(_13171_));
 NAND2x1_ASAP7_75t_R _30473_ (.A(_13137_),
    .B(_00363_),
    .Y(_13172_));
 BUFx12f_ASAP7_75t_R _30474_ (.A(_13087_),
    .Y(_13173_));
 BUFx6f_ASAP7_75t_R _30475_ (.A(_13173_),
    .Y(_13174_));
 OA211x2_ASAP7_75t_R _30476_ (.A1(_13143_),
    .A2(_13171_),
    .B(_13172_),
    .C(_13174_),
    .Y(_13175_));
 OR3x1_ASAP7_75t_R _30477_ (.A(_13131_),
    .B(_13170_),
    .C(_13175_),
    .Y(_13176_));
 INVx1_ASAP7_75t_R _30478_ (.A(_00374_),
    .Y(_13177_));
 NAND2x1_ASAP7_75t_R _30479_ (.A(_13168_),
    .B(_00372_),
    .Y(_13178_));
 OA211x2_ASAP7_75t_R _30480_ (.A1(_13133_),
    .A2(_13177_),
    .B(_13178_),
    .C(_13140_),
    .Y(_13179_));
 INVx2_ASAP7_75t_R _30481_ (.A(_00373_),
    .Y(_13180_));
 NAND2x1_ASAP7_75t_R _30482_ (.A(_13146_),
    .B(_00371_),
    .Y(_13181_));
 OA211x2_ASAP7_75t_R _30483_ (.A1(_13143_),
    .A2(_13180_),
    .B(_13181_),
    .C(_13149_),
    .Y(_13182_));
 OR3x1_ASAP7_75t_R _30484_ (.A(_13153_),
    .B(_13179_),
    .C(_13182_),
    .Y(_13183_));
 AND3x1_ASAP7_75t_R _30485_ (.A(_13129_),
    .B(_13176_),
    .C(_13183_),
    .Y(_13184_));
 BUFx12f_ASAP7_75t_R _30486_ (.A(_13104_),
    .Y(_13185_));
 BUFx6f_ASAP7_75t_R _30487_ (.A(_13185_),
    .Y(_13186_));
 BUFx12f_ASAP7_75t_R _30488_ (.A(_13149_),
    .Y(_13187_));
 BUFx12f_ASAP7_75t_R _30489_ (.A(_13094_),
    .Y(_13188_));
 BUFx12f_ASAP7_75t_R _30490_ (.A(_13188_),
    .Y(_13189_));
 BUFx6f_ASAP7_75t_R _30491_ (.A(_13189_),
    .Y(_13190_));
 INVx2_ASAP7_75t_R _30492_ (.A(_00367_),
    .Y(_13191_));
 BUFx12f_ASAP7_75t_R _30493_ (.A(_13095_),
    .Y(_13192_));
 BUFx12f_ASAP7_75t_R _30494_ (.A(_13192_),
    .Y(_13193_));
 NOR2x1_ASAP7_75t_R _30495_ (.A(_13193_),
    .B(_00369_),
    .Y(_13194_));
 AO21x1_ASAP7_75t_R _30496_ (.A1(_13190_),
    .A2(_13191_),
    .B(_13194_),
    .Y(_13195_));
 BUFx12f_ASAP7_75t_R _30497_ (.A(_13109_),
    .Y(_13196_));
 BUFx12f_ASAP7_75t_R _30498_ (.A(_13196_),
    .Y(_13197_));
 INVx2_ASAP7_75t_R _30499_ (.A(_00370_),
    .Y(_13198_));
 BUFx12f_ASAP7_75t_R _30500_ (.A(_13135_),
    .Y(_13199_));
 BUFx12f_ASAP7_75t_R _30501_ (.A(_13199_),
    .Y(_13200_));
 NAND2x1_ASAP7_75t_R _30502_ (.A(_13200_),
    .B(_00368_),
    .Y(_13201_));
 BUFx6f_ASAP7_75t_R _30503_ (.A(_13139_),
    .Y(_13202_));
 OA211x2_ASAP7_75t_R _30504_ (.A1(_13197_),
    .A2(_13198_),
    .B(_13201_),
    .C(_13202_),
    .Y(_13203_));
 AO21x1_ASAP7_75t_R _30505_ (.A1(_13187_),
    .A2(_13195_),
    .B(_13203_),
    .Y(_13204_));
 BUFx12f_ASAP7_75t_R _30506_ (.A(_13135_),
    .Y(_13205_));
 BUFx12f_ASAP7_75t_R _30507_ (.A(_13205_),
    .Y(_13206_));
 INVx2_ASAP7_75t_R _30508_ (.A(_00362_),
    .Y(_13207_));
 NAND2x1_ASAP7_75t_R _30509_ (.A(_13118_),
    .B(_00360_),
    .Y(_13208_));
 OA211x2_ASAP7_75t_R _30510_ (.A1(_13206_),
    .A2(_13207_),
    .B(_13208_),
    .C(_13115_),
    .Y(_13209_));
 INVx2_ASAP7_75t_R _30511_ (.A(_00361_),
    .Y(_13210_));
 BUFx6f_ASAP7_75t_R _30512_ (.A(_13109_),
    .Y(_13211_));
 NAND2x1_ASAP7_75t_R _30513_ (.A(_13211_),
    .B(_00359_),
    .Y(_13212_));
 OA211x2_ASAP7_75t_R _30514_ (.A1(_13206_),
    .A2(_13210_),
    .B(_13212_),
    .C(_13120_),
    .Y(_13213_));
 OR3x1_ASAP7_75t_R _30515_ (.A(_13085_),
    .B(_13209_),
    .C(_13213_),
    .Y(_13214_));
 OA211x2_ASAP7_75t_R _30516_ (.A1(_13186_),
    .A2(_13204_),
    .B(_13214_),
    .C(_13125_),
    .Y(_13215_));
 OR3x2_ASAP7_75t_R _30517_ (.A(_13164_),
    .B(_13184_),
    .C(_13215_),
    .Y(_13216_));
 BUFx6f_ASAP7_75t_R _30518_ (.A(_01511_),
    .Y(_13217_));
 BUFx6f_ASAP7_75t_R _30519_ (.A(_01508_),
    .Y(_13218_));
 INVx2_ASAP7_75t_R _30520_ (.A(_13218_),
    .Y(_13219_));
 BUFx6f_ASAP7_75t_R _30521_ (.A(_13219_),
    .Y(_13220_));
 BUFx6f_ASAP7_75t_R _30522_ (.A(_01509_),
    .Y(_13221_));
 BUFx6f_ASAP7_75t_R _30523_ (.A(_00376_),
    .Y(_13222_));
 OR2x6_ASAP7_75t_R _30524_ (.A(_13222_),
    .B(_01507_),
    .Y(_13223_));
 OR3x1_ASAP7_75t_R _30525_ (.A(_13220_),
    .B(_13221_),
    .C(_13223_),
    .Y(_13224_));
 NAND2x1_ASAP7_75t_R _30526_ (.A(_13222_),
    .B(_01507_),
    .Y(_13225_));
 BUFx12f_ASAP7_75t_R _30527_ (.A(_00377_),
    .Y(_13226_));
 BUFx12f_ASAP7_75t_R _30528_ (.A(_00413_),
    .Y(_13227_));
 AND3x4_ASAP7_75t_R _30529_ (.A(_13226_),
    .B(_13227_),
    .C(_01519_),
    .Y(_13228_));
 OR4x1_ASAP7_75t_R _30530_ (.A(_13219_),
    .B(_13221_),
    .C(_13225_),
    .D(_13228_),
    .Y(_13229_));
 INVx2_ASAP7_75t_R _30531_ (.A(_13221_),
    .Y(_13230_));
 OR3x1_ASAP7_75t_R _30532_ (.A(_13218_),
    .B(_13230_),
    .C(_13225_),
    .Y(_13231_));
 AND3x1_ASAP7_75t_R _30533_ (.A(_13224_),
    .B(_13229_),
    .C(_13231_),
    .Y(_13232_));
 BUFx12f_ASAP7_75t_R _30534_ (.A(_00760_),
    .Y(_13233_));
 INVx5_ASAP7_75t_R _30535_ (.A(_13233_),
    .Y(_13234_));
 BUFx12f_ASAP7_75t_R _30536_ (.A(_01757_),
    .Y(_13235_));
 AO211x2_ASAP7_75t_R _30537_ (.A1(_13234_),
    .A2(_13235_),
    .B(_13219_),
    .C(_13223_),
    .Y(_13236_));
 BUFx6f_ASAP7_75t_R _30538_ (.A(_01518_),
    .Y(_13237_));
 BUFx6f_ASAP7_75t_R _30539_ (.A(_01521_),
    .Y(_13238_));
 NOR2x1_ASAP7_75t_R _30540_ (.A(_13237_),
    .B(_13238_),
    .Y(_13239_));
 BUFx6f_ASAP7_75t_R _30541_ (.A(_13239_),
    .Y(_13240_));
 OA21x2_ASAP7_75t_R _30542_ (.A1(_13230_),
    .A2(_13236_),
    .B(_13240_),
    .Y(_13241_));
 BUFx6f_ASAP7_75t_R _30543_ (.A(_01507_),
    .Y(_13242_));
 INVx3_ASAP7_75t_R _30544_ (.A(_13242_),
    .Y(_13243_));
 INVx2_ASAP7_75t_R _30545_ (.A(_13222_),
    .Y(_13244_));
 AO21x1_ASAP7_75t_R _30546_ (.A1(_13244_),
    .A2(_13218_),
    .B(_13217_),
    .Y(_13245_));
 NOR2x1_ASAP7_75t_R _30547_ (.A(_13221_),
    .B(_01511_),
    .Y(_13246_));
 AND2x2_ASAP7_75t_R _30548_ (.A(_01507_),
    .B(_13218_),
    .Y(_13247_));
 AND2x6_ASAP7_75t_R _30549_ (.A(_13221_),
    .B(_01511_),
    .Y(_13248_));
 AO21x1_ASAP7_75t_R _30550_ (.A1(_13246_),
    .A2(_13247_),
    .B(_13248_),
    .Y(_13249_));
 AO32x1_ASAP7_75t_R _30551_ (.A1(_13243_),
    .A2(_13221_),
    .A3(_13245_),
    .B1(_13249_),
    .B2(_13222_),
    .Y(_13250_));
 OA211x2_ASAP7_75t_R _30552_ (.A1(_13217_),
    .A2(_13232_),
    .B(_13241_),
    .C(_13250_),
    .Y(_13251_));
 BUFx6f_ASAP7_75t_R _30553_ (.A(_13251_),
    .Y(_13252_));
 NAND2x1_ASAP7_75t_R _30554_ (.A(_01443_),
    .B(_01444_),
    .Y(_13253_));
 NOR2x2_ASAP7_75t_R _30555_ (.A(_00375_),
    .B(_13253_),
    .Y(_13254_));
 INVx2_ASAP7_75t_R _30556_ (.A(_18707_),
    .Y(_13255_));
 INVx2_ASAP7_75t_R _30557_ (.A(_01443_),
    .Y(_13256_));
 OA211x2_ASAP7_75t_R _30558_ (.A1(_13255_),
    .A2(_01444_),
    .B(_13256_),
    .C(_00375_),
    .Y(_13257_));
 NOR2x2_ASAP7_75t_R _30559_ (.A(_13254_),
    .B(_13257_),
    .Y(_13258_));
 BUFx12f_ASAP7_75t_R _30560_ (.A(_13258_),
    .Y(_13259_));
 BUFx12f_ASAP7_75t_R _30561_ (.A(_13259_),
    .Y(_13260_));
 INVx2_ASAP7_75t_R _30562_ (.A(_13226_),
    .Y(_13261_));
 BUFx12f_ASAP7_75t_R _30563_ (.A(_13261_),
    .Y(_13262_));
 BUFx6f_ASAP7_75t_R _30564_ (.A(_13221_),
    .Y(_13263_));
 NOR2x2_ASAP7_75t_R _30565_ (.A(_13222_),
    .B(_01507_),
    .Y(_13264_));
 AND5x2_ASAP7_75t_R _30566_ (.A(_13220_),
    .B(_13263_),
    .C(_13217_),
    .D(_13239_),
    .E(_13264_),
    .Y(_13265_));
 NAND2x2_ASAP7_75t_R _30567_ (.A(_13262_),
    .B(_13265_),
    .Y(_13266_));
 NAND3x2_ASAP7_75t_R _30568_ (.B(_13260_),
    .C(_13266_),
    .Y(_13267_),
    .A(_13252_));
 BUFx6f_ASAP7_75t_R _30569_ (.A(_13267_),
    .Y(_13268_));
 AO21x2_ASAP7_75t_R _30570_ (.A1(_13162_),
    .A2(_13216_),
    .B(_13268_),
    .Y(_13269_));
 INVx1_ASAP7_75t_R _30571_ (.A(_01474_),
    .Y(_13270_));
 OR2x6_ASAP7_75t_R _30572_ (.A(_13254_),
    .B(_13257_),
    .Y(_13271_));
 BUFx6f_ASAP7_75t_R _30573_ (.A(_13271_),
    .Y(_13272_));
 AO21x1_ASAP7_75t_R _30574_ (.A1(_13252_),
    .A2(_13266_),
    .B(_13272_),
    .Y(_13273_));
 INVx2_ASAP7_75t_R _30575_ (.A(_01503_),
    .Y(_13274_));
 AO211x2_ASAP7_75t_R _30576_ (.A1(_13252_),
    .A2(_13266_),
    .B(_13272_),
    .C(_13274_),
    .Y(_13275_));
 NAND2x2_ASAP7_75t_R _30577_ (.A(_13221_),
    .B(_01511_),
    .Y(_13276_));
 BUFx6f_ASAP7_75t_R _30578_ (.A(_13222_),
    .Y(_13277_));
 OR3x1_ASAP7_75t_R _30579_ (.A(_13277_),
    .B(_13220_),
    .C(_13217_),
    .Y(_13278_));
 AO21x2_ASAP7_75t_R _30580_ (.A1(_13276_),
    .A2(_13278_),
    .B(_13242_),
    .Y(_13279_));
 BUFx6f_ASAP7_75t_R _30581_ (.A(_13218_),
    .Y(_13280_));
 AND2x2_ASAP7_75t_R _30582_ (.A(_13280_),
    .B(_13246_),
    .Y(_13281_));
 AO21x1_ASAP7_75t_R _30583_ (.A1(_13220_),
    .A2(_13263_),
    .B(_13248_),
    .Y(_13282_));
 OA21x2_ASAP7_75t_R _30584_ (.A1(_13242_),
    .A2(_13248_),
    .B(_13277_),
    .Y(_13283_));
 OAI21x1_ASAP7_75t_R _30585_ (.A1(_13281_),
    .A2(_13282_),
    .B(_13283_),
    .Y(_13284_));
 OR2x6_ASAP7_75t_R _30586_ (.A(_13237_),
    .B(_13238_),
    .Y(_13285_));
 OR3x2_ASAP7_75t_R _30587_ (.A(_13285_),
    .B(_13254_),
    .C(_13257_),
    .Y(_13286_));
 BUFx6f_ASAP7_75t_R _30588_ (.A(_13226_),
    .Y(_13287_));
 OR4x1_ASAP7_75t_R _30589_ (.A(_13287_),
    .B(_13280_),
    .C(_13276_),
    .D(_13223_),
    .Y(_13288_));
 AO21x1_ASAP7_75t_R _30590_ (.A1(_13226_),
    .A2(_13227_),
    .B(_13217_),
    .Y(_13289_));
 OR4x1_ASAP7_75t_R _30591_ (.A(_13220_),
    .B(_13263_),
    .C(_13225_),
    .D(_13289_),
    .Y(_13290_));
 NAND2x1_ASAP7_75t_R _30592_ (.A(_13288_),
    .B(_13290_),
    .Y(_13291_));
 AOI211x1_ASAP7_75t_R _30593_ (.A1(_13279_),
    .A2(_13284_),
    .B(_13286_),
    .C(_13291_),
    .Y(_13292_));
 AO22x2_ASAP7_75t_R _30594_ (.A1(_13270_),
    .A2(_13273_),
    .B1(_13275_),
    .B2(_13292_),
    .Y(_13293_));
 AND2x4_ASAP7_75t_R _30595_ (.A(_13269_),
    .B(_13293_),
    .Y(_18615_));
 INVx3_ASAP7_75t_R _30596_ (.A(_18615_),
    .Y(_18613_));
 INVx2_ASAP7_75t_R _30597_ (.A(_01757_),
    .Y(_13294_));
 OA211x2_ASAP7_75t_R _30598_ (.A1(_13233_),
    .A2(_13294_),
    .B(_13218_),
    .C(_13264_),
    .Y(_13295_));
 BUFx6f_ASAP7_75t_R _30599_ (.A(_13295_),
    .Y(_13296_));
 OR3x2_ASAP7_75t_R _30600_ (.A(_13242_),
    .B(_13276_),
    .C(_13285_),
    .Y(_13297_));
 NAND3x1_ASAP7_75t_R _30601_ (.A(_13222_),
    .B(_13226_),
    .C(_13218_),
    .Y(_13298_));
 OAI21x1_ASAP7_75t_R _30602_ (.A1(_13277_),
    .A2(_13280_),
    .B(_13298_),
    .Y(_13299_));
 NOR3x1_ASAP7_75t_R _30603_ (.A(_13296_),
    .B(_13297_),
    .C(_13299_),
    .Y(_13300_));
 AND2x6_ASAP7_75t_R _30604_ (.A(_13259_),
    .B(_13300_),
    .Y(_13301_));
 BUFx12f_ASAP7_75t_R _30605_ (.A(_13301_),
    .Y(_13302_));
 BUFx12f_ASAP7_75t_R _30606_ (.A(_00378_),
    .Y(_13303_));
 BUFx12f_ASAP7_75t_R _30607_ (.A(_13303_),
    .Y(_13304_));
 BUFx12f_ASAP7_75t_R _30608_ (.A(_13304_),
    .Y(_13305_));
 BUFx12f_ASAP7_75t_R _30609_ (.A(_13305_),
    .Y(_13306_));
 BUFx12f_ASAP7_75t_R _30610_ (.A(_01516_),
    .Y(_13307_));
 BUFx12f_ASAP7_75t_R _30611_ (.A(_13307_),
    .Y(_13308_));
 BUFx12f_ASAP7_75t_R _30612_ (.A(_00379_),
    .Y(_13309_));
 AND2x6_ASAP7_75t_R _30613_ (.A(_13308_),
    .B(_13309_),
    .Y(_13310_));
 BUFx12f_ASAP7_75t_R _30614_ (.A(_01517_),
    .Y(_13311_));
 INVx3_ASAP7_75t_R _30615_ (.A(_13311_),
    .Y(_13312_));
 BUFx12f_ASAP7_75t_R _30616_ (.A(_13312_),
    .Y(_13313_));
 BUFx12f_ASAP7_75t_R _30617_ (.A(_13313_),
    .Y(_13314_));
 BUFx12f_ASAP7_75t_R _30618_ (.A(_13311_),
    .Y(_13315_));
 BUFx12f_ASAP7_75t_R _30619_ (.A(_13315_),
    .Y(_13316_));
 BUFx6f_ASAP7_75t_R _30620_ (.A(_13316_),
    .Y(_13317_));
 AND2x2_ASAP7_75t_R _30621_ (.A(_13317_),
    .B(_01796_),
    .Y(_13318_));
 AO21x1_ASAP7_75t_R _30622_ (.A1(_00382_),
    .A2(_13314_),
    .B(_13318_),
    .Y(_13319_));
 BUFx12f_ASAP7_75t_R _30623_ (.A(_00380_),
    .Y(_13320_));
 BUFx12f_ASAP7_75t_R _30624_ (.A(_13320_),
    .Y(_13321_));
 BUFx12f_ASAP7_75t_R _30625_ (.A(_13321_),
    .Y(_13322_));
 BUFx12f_ASAP7_75t_R _30626_ (.A(_13322_),
    .Y(_13323_));
 AO21x1_ASAP7_75t_R _30627_ (.A1(_13310_),
    .A2(_13319_),
    .B(_13323_),
    .Y(_13324_));
 NAND2x1_ASAP7_75t_R _30628_ (.A(_13306_),
    .B(_13324_),
    .Y(_13325_));
 BUFx12f_ASAP7_75t_R _30629_ (.A(_13312_),
    .Y(_13326_));
 BUFx12f_ASAP7_75t_R _30630_ (.A(_13326_),
    .Y(_13327_));
 BUFx12f_ASAP7_75t_R _30631_ (.A(_13327_),
    .Y(_13328_));
 INVx5_ASAP7_75t_R _30632_ (.A(_00379_),
    .Y(_13329_));
 INVx4_ASAP7_75t_R _30633_ (.A(_13307_),
    .Y(_13330_));
 BUFx12f_ASAP7_75t_R _30634_ (.A(_13330_),
    .Y(_13331_));
 BUFx12f_ASAP7_75t_R _30635_ (.A(_13331_),
    .Y(_13332_));
 BUFx12f_ASAP7_75t_R _30636_ (.A(_13307_),
    .Y(_13333_));
 BUFx12f_ASAP7_75t_R _30637_ (.A(_13333_),
    .Y(_13334_));
 AND2x2_ASAP7_75t_R _30638_ (.A(_13334_),
    .B(_00389_),
    .Y(_13335_));
 AO21x1_ASAP7_75t_R _30639_ (.A1(_13332_),
    .A2(_00393_),
    .B(_13335_),
    .Y(_13336_));
 AND3x1_ASAP7_75t_R _30640_ (.A(_13328_),
    .B(_13329_),
    .C(_13336_),
    .Y(_13337_));
 BUFx12f_ASAP7_75t_R _30641_ (.A(_13315_),
    .Y(_13338_));
 BUFx12f_ASAP7_75t_R _30642_ (.A(_13338_),
    .Y(_13339_));
 BUFx6f_ASAP7_75t_R _30643_ (.A(_13339_),
    .Y(_13340_));
 AND2x2_ASAP7_75t_R _30644_ (.A(_13334_),
    .B(_00387_),
    .Y(_13341_));
 AO21x1_ASAP7_75t_R _30645_ (.A1(_13332_),
    .A2(_00391_),
    .B(_13341_),
    .Y(_13342_));
 INVx2_ASAP7_75t_R _30646_ (.A(_00380_),
    .Y(_13343_));
 BUFx6f_ASAP7_75t_R _30647_ (.A(_13343_),
    .Y(_13344_));
 BUFx6f_ASAP7_75t_R _30648_ (.A(_13344_),
    .Y(_13345_));
 BUFx6f_ASAP7_75t_R _30649_ (.A(_13345_),
    .Y(_13346_));
 BUFx12f_ASAP7_75t_R _30650_ (.A(_13315_),
    .Y(_13347_));
 BUFx12f_ASAP7_75t_R _30651_ (.A(_13347_),
    .Y(_13348_));
 OR3x1_ASAP7_75t_R _30652_ (.A(_00381_),
    .B(_13346_),
    .C(_13348_),
    .Y(_13349_));
 AO32x1_ASAP7_75t_R _30653_ (.A1(_13340_),
    .A2(_13329_),
    .A3(_13342_),
    .B1(_13349_),
    .B2(_13310_),
    .Y(_13350_));
 NOR2x1_ASAP7_75t_R _30654_ (.A(_13337_),
    .B(_13350_),
    .Y(_13351_));
 BUFx6f_ASAP7_75t_R _30655_ (.A(_13321_),
    .Y(_13352_));
 BUFx6f_ASAP7_75t_R _30656_ (.A(_13352_),
    .Y(_13353_));
 BUFx6f_ASAP7_75t_R _30657_ (.A(_13308_),
    .Y(_13354_));
 INVx1_ASAP7_75t_R _30658_ (.A(_00410_),
    .Y(_13355_));
 BUFx12f_ASAP7_75t_R _30659_ (.A(_13307_),
    .Y(_13356_));
 NAND2x1_ASAP7_75t_R _30660_ (.A(_13356_),
    .B(_00406_),
    .Y(_13357_));
 OA211x2_ASAP7_75t_R _30661_ (.A1(_13354_),
    .A2(_13355_),
    .B(_13357_),
    .C(_13326_),
    .Y(_13358_));
 INVx1_ASAP7_75t_R _30662_ (.A(_00408_),
    .Y(_13359_));
 NAND2x1_ASAP7_75t_R _30663_ (.A(_13356_),
    .B(_00404_),
    .Y(_13360_));
 BUFx3_ASAP7_75t_R rebuffer40 (.A(_00751_),
    .Y(net1975));
 BUFx12f_ASAP7_75t_R _30665_ (.A(_01517_),
    .Y(_13362_));
 BUFx12f_ASAP7_75t_R _30666_ (.A(_13362_),
    .Y(_13363_));
 OA211x2_ASAP7_75t_R _30667_ (.A1(_13354_),
    .A2(_13359_),
    .B(_13360_),
    .C(_13363_),
    .Y(_13364_));
 OR2x6_ASAP7_75t_R _30668_ (.A(_00379_),
    .B(_13303_),
    .Y(_13365_));
 OR4x1_ASAP7_75t_R _30669_ (.A(_13353_),
    .B(_13358_),
    .C(_13364_),
    .D(_13365_),
    .Y(_13366_));
 INVx1_ASAP7_75t_R _30670_ (.A(_00386_),
    .Y(_13367_));
 NAND2x1_ASAP7_75t_R _30671_ (.A(_13347_),
    .B(_00384_),
    .Y(_13368_));
 BUFx6f_ASAP7_75t_R _30672_ (.A(_13344_),
    .Y(_13369_));
 OA211x2_ASAP7_75t_R _30673_ (.A1(_13317_),
    .A2(_13367_),
    .B(_13368_),
    .C(_13369_),
    .Y(_13370_));
 INVx1_ASAP7_75t_R _30674_ (.A(_00385_),
    .Y(_13371_));
 NAND2x1_ASAP7_75t_R _30675_ (.A(_13347_),
    .B(_00383_),
    .Y(_13372_));
 OA211x2_ASAP7_75t_R _30676_ (.A1(_13317_),
    .A2(_13371_),
    .B(_13372_),
    .C(_13352_),
    .Y(_13373_));
 AND2x6_ASAP7_75t_R _30677_ (.A(_00379_),
    .B(_00378_),
    .Y(_13374_));
 NAND2x2_ASAP7_75t_R _30678_ (.A(_13330_),
    .B(_13374_),
    .Y(_13375_));
 OR3x1_ASAP7_75t_R _30679_ (.A(_13370_),
    .B(_13373_),
    .C(_13375_),
    .Y(_13376_));
 AND2x2_ASAP7_75t_R _30680_ (.A(_13366_),
    .B(_13376_),
    .Y(_13377_));
 BUFx12f_ASAP7_75t_R _30681_ (.A(_13362_),
    .Y(_13378_));
 INVx2_ASAP7_75t_R _30682_ (.A(_00402_),
    .Y(_13379_));
 NAND2x1_ASAP7_75t_R _30683_ (.A(_13338_),
    .B(_00400_),
    .Y(_13380_));
 OA211x2_ASAP7_75t_R _30684_ (.A1(_13378_),
    .A2(_13379_),
    .B(_13380_),
    .C(_13369_),
    .Y(_13381_));
 INVx1_ASAP7_75t_R _30685_ (.A(_00401_),
    .Y(_13382_));
 NAND2x1_ASAP7_75t_R _30686_ (.A(_13338_),
    .B(_00399_),
    .Y(_13383_));
 OA211x2_ASAP7_75t_R _30687_ (.A1(_13378_),
    .A2(_13382_),
    .B(_13383_),
    .C(_13352_),
    .Y(_13384_));
 OR3x1_ASAP7_75t_R _30688_ (.A(_13307_),
    .B(_13329_),
    .C(_00378_),
    .Y(_13385_));
 BUFx6f_ASAP7_75t_R _30689_ (.A(_13385_),
    .Y(_13386_));
 OR3x1_ASAP7_75t_R _30690_ (.A(_13381_),
    .B(_13384_),
    .C(_13386_),
    .Y(_13387_));
 BUFx6f_ASAP7_75t_R _30691_ (.A(_13303_),
    .Y(_13388_));
 NAND2x2_ASAP7_75t_R _30692_ (.A(_13307_),
    .B(_13309_),
    .Y(_13389_));
 INVx2_ASAP7_75t_R _30693_ (.A(_00397_),
    .Y(_13390_));
 BUFx12f_ASAP7_75t_R _30694_ (.A(net1976),
    .Y(_13391_));
 NAND2x1_ASAP7_75t_R _30695_ (.A(_13391_),
    .B(_00395_),
    .Y(_13392_));
 BUFx6f_ASAP7_75t_R _30696_ (.A(_13320_),
    .Y(_13393_));
 OA211x2_ASAP7_75t_R _30697_ (.A1(_13347_),
    .A2(_13390_),
    .B(_13392_),
    .C(_13393_),
    .Y(_13394_));
 INVx2_ASAP7_75t_R _30698_ (.A(_00398_),
    .Y(_13395_));
 NAND2x1_ASAP7_75t_R _30699_ (.A(_13391_),
    .B(_00396_),
    .Y(_13396_));
 OA211x2_ASAP7_75t_R _30700_ (.A1(_13347_),
    .A2(_13395_),
    .B(_13396_),
    .C(_13345_),
    .Y(_13397_));
 OR4x1_ASAP7_75t_R _30701_ (.A(_13388_),
    .B(_13389_),
    .C(_13394_),
    .D(_13397_),
    .Y(_13398_));
 INVx1_ASAP7_75t_R _30702_ (.A(_00407_),
    .Y(_13399_));
 BUFx12f_ASAP7_75t_R _30703_ (.A(_13307_),
    .Y(_13400_));
 NAND2x1_ASAP7_75t_R _30704_ (.A(_13400_),
    .B(_00403_),
    .Y(_13401_));
 BUFx6f_ASAP7_75t_R _30705_ (.A(net1977),
    .Y(_13402_));
 OA211x2_ASAP7_75t_R _30706_ (.A1(_13354_),
    .A2(_13399_),
    .B(_13401_),
    .C(_13402_),
    .Y(_13403_));
 INVx2_ASAP7_75t_R _30707_ (.A(_00409_),
    .Y(_13404_));
 NAND2x1_ASAP7_75t_R _30708_ (.A(_13400_),
    .B(_00405_),
    .Y(_13405_));
 OA211x2_ASAP7_75t_R _30709_ (.A1(_13354_),
    .A2(_13404_),
    .B(_13405_),
    .C(_13313_),
    .Y(_13406_));
 NOR2x2_ASAP7_75t_R _30710_ (.A(_13309_),
    .B(_13303_),
    .Y(_13407_));
 NAND2x1_ASAP7_75t_R _30711_ (.A(_13352_),
    .B(_13407_),
    .Y(_13408_));
 OR3x1_ASAP7_75t_R _30712_ (.A(_13403_),
    .B(_13406_),
    .C(_13408_),
    .Y(_13409_));
 INVx2_ASAP7_75t_R _30713_ (.A(_00394_),
    .Y(_13410_));
 NAND2x1_ASAP7_75t_R _30714_ (.A(_13400_),
    .B(_00390_),
    .Y(_13411_));
 OA211x2_ASAP7_75t_R _30715_ (.A1(_13354_),
    .A2(_13410_),
    .B(_13411_),
    .C(_13313_),
    .Y(_13412_));
 INVx1_ASAP7_75t_R _30716_ (.A(_00392_),
    .Y(_13413_));
 NAND2x1_ASAP7_75t_R _30717_ (.A(_13356_),
    .B(_00388_),
    .Y(_13414_));
 OA211x2_ASAP7_75t_R _30718_ (.A1(_13354_),
    .A2(_13413_),
    .B(_13414_),
    .C(_13363_),
    .Y(_13415_));
 NOR2x2_ASAP7_75t_R _30719_ (.A(_13320_),
    .B(_13309_),
    .Y(_13416_));
 NAND2x2_ASAP7_75t_R _30720_ (.A(_13303_),
    .B(_13416_),
    .Y(_13417_));
 OR3x1_ASAP7_75t_R _30721_ (.A(_13412_),
    .B(_13415_),
    .C(_13417_),
    .Y(_13418_));
 AND4x1_ASAP7_75t_R _30722_ (.A(_13387_),
    .B(_13398_),
    .C(_13409_),
    .D(_13418_),
    .Y(_13419_));
 OA211x2_ASAP7_75t_R _30723_ (.A1(_13325_),
    .A2(_13351_),
    .B(_13377_),
    .C(_13419_),
    .Y(_13420_));
 BUFx6f_ASAP7_75t_R _30724_ (.A(_01519_),
    .Y(_13421_));
 NAND2x2_ASAP7_75t_R _30725_ (.A(_13226_),
    .B(_13227_),
    .Y(_13422_));
 OR5x2_ASAP7_75t_R _30726_ (.A(_13219_),
    .B(_13221_),
    .C(_13421_),
    .D(_13225_),
    .E(_13422_),
    .Y(_13423_));
 OR3x2_ASAP7_75t_R _30727_ (.A(_01511_),
    .B(_13237_),
    .C(_13238_),
    .Y(_13424_));
 AO21x1_ASAP7_75t_R _30728_ (.A1(_13236_),
    .A2(_13423_),
    .B(_13424_),
    .Y(_13425_));
 BUFx6f_ASAP7_75t_R _30729_ (.A(_13425_),
    .Y(_13426_));
 OR4x1_ASAP7_75t_R _30730_ (.A(_13244_),
    .B(_13218_),
    .C(_13230_),
    .D(_13424_),
    .Y(_13427_));
 OA21x2_ASAP7_75t_R _30731_ (.A1(_13298_),
    .A2(_13297_),
    .B(_13427_),
    .Y(_13428_));
 BUFx6f_ASAP7_75t_R _30732_ (.A(_13428_),
    .Y(_13429_));
 BUFx12f_ASAP7_75t_R _30733_ (.A(_01506_),
    .Y(_13430_));
 AOI211x1_ASAP7_75t_R _30734_ (.A1(_13426_),
    .A2(_13429_),
    .B(_13430_),
    .C(_13272_),
    .Y(_13431_));
 AND2x2_ASAP7_75t_R _30735_ (.A(_13236_),
    .B(_13423_),
    .Y(_13432_));
 OR3x1_ASAP7_75t_R _30736_ (.A(_13254_),
    .B(_13257_),
    .C(_13424_),
    .Y(_13433_));
 BUFx12f_ASAP7_75t_R _30737_ (.A(_13369_),
    .Y(_13434_));
 OA21x2_ASAP7_75t_R _30738_ (.A1(_13297_),
    .A2(_13299_),
    .B(_13434_),
    .Y(_13435_));
 OA221x2_ASAP7_75t_R _30739_ (.A1(_13432_),
    .A2(_13433_),
    .B1(_13429_),
    .B2(_13272_),
    .C(_13435_),
    .Y(_13436_));
 AND2x6_ASAP7_75t_R _30740_ (.A(_13248_),
    .B(_13240_),
    .Y(_13437_));
 NAND2x1_ASAP7_75t_R _30741_ (.A(_13296_),
    .B(_13437_),
    .Y(_13438_));
 AND3x4_ASAP7_75t_R _30742_ (.A(_13258_),
    .B(_13427_),
    .C(_13438_),
    .Y(_13439_));
 NOR3x1_ASAP7_75t_R _30743_ (.A(_13217_),
    .B(_13237_),
    .C(_13238_),
    .Y(_13440_));
 NAND2x1_ASAP7_75t_R _30744_ (.A(_13280_),
    .B(_13264_),
    .Y(_13441_));
 AND3x1_ASAP7_75t_R _30745_ (.A(_13234_),
    .B(_13235_),
    .C(_13263_),
    .Y(_13442_));
 OAI21x1_ASAP7_75t_R _30746_ (.A1(_13441_),
    .A2(_13442_),
    .B(_13423_),
    .Y(_13443_));
 NAND2x1_ASAP7_75t_R _30747_ (.A(_13440_),
    .B(_13443_),
    .Y(_13444_));
 OA211x2_ASAP7_75t_R _30748_ (.A1(_13431_),
    .A2(_13436_),
    .B(_13439_),
    .C(_13444_),
    .Y(_13445_));
 AOI21x1_ASAP7_75t_R _30749_ (.A1(_13302_),
    .A2(_13420_),
    .B(_13445_),
    .Y(_13446_));
 INVx5_ASAP7_75t_R _30750_ (.A(_13446_),
    .Y(_13447_));
 BUFx12f_ASAP7_75t_R _30751_ (.A(_13447_),
    .Y(_13448_));
 BUFx12f_ASAP7_75t_R _30752_ (.A(_13448_),
    .Y(_13449_));
 BUFx6f_ASAP7_75t_R _30753_ (.A(_13449_),
    .Y(_13450_));
 BUFx6f_ASAP7_75t_R _30754_ (.A(_13450_),
    .Y(_18555_));
 BUFx12f_ASAP7_75t_R _30755_ (.A(_13446_),
    .Y(_13451_));
 BUFx12f_ASAP7_75t_R _30756_ (.A(_13451_),
    .Y(_13452_));
 BUFx12f_ASAP7_75t_R _30757_ (.A(_13452_),
    .Y(_13453_));
 BUFx6f_ASAP7_75t_R _30758_ (.A(_13453_),
    .Y(_13454_));
 BUFx6f_ASAP7_75t_R _30759_ (.A(_13454_),
    .Y(_18553_));
 BUFx12f_ASAP7_75t_R _30760_ (.A(_01505_),
    .Y(_13455_));
 INVx3_ASAP7_75t_R _30761_ (.A(_13455_),
    .Y(_13456_));
 NAND2x1_ASAP7_75t_R _30762_ (.A(_13426_),
    .B(_13429_),
    .Y(_13457_));
 AO32x2_ASAP7_75t_R _30763_ (.A1(_13439_),
    .A2(_13444_),
    .A3(_13457_),
    .B1(_13437_),
    .B2(_13296_),
    .Y(_13458_));
 BUFx12f_ASAP7_75t_R _30764_ (.A(_13309_),
    .Y(_13459_));
 INVx5_ASAP7_75t_R _30765_ (.A(_13303_),
    .Y(_13460_));
 BUFx12f_ASAP7_75t_R _30766_ (.A(_13460_),
    .Y(_13461_));
 INVx2_ASAP7_75t_R _30767_ (.A(_00427_),
    .Y(_13462_));
 NOR2x1_ASAP7_75t_R _30768_ (.A(_13321_),
    .B(_13338_),
    .Y(_13463_));
 NAND2x1_ASAP7_75t_R _30769_ (.A(_13400_),
    .B(_00423_),
    .Y(_13464_));
 OA211x2_ASAP7_75t_R _30770_ (.A1(_13354_),
    .A2(_13462_),
    .B(_13463_),
    .C(_13464_),
    .Y(_13465_));
 OR3x1_ASAP7_75t_R _30771_ (.A(_13459_),
    .B(_13461_),
    .C(_13465_),
    .Y(_13466_));
 AND2x6_ASAP7_75t_R _30772_ (.A(_13345_),
    .B(_13363_),
    .Y(_13467_));
 OR2x2_ASAP7_75t_R _30773_ (.A(_13333_),
    .B(_00425_),
    .Y(_13468_));
 OAI21x1_ASAP7_75t_R _30774_ (.A1(_13331_),
    .A2(_00421_),
    .B(_13468_),
    .Y(_13469_));
 AND2x6_ASAP7_75t_R _30775_ (.A(_13393_),
    .B(_13363_),
    .Y(_13470_));
 OR2x2_ASAP7_75t_R _30776_ (.A(_13333_),
    .B(_00424_),
    .Y(_13471_));
 OAI21x1_ASAP7_75t_R _30777_ (.A1(_13331_),
    .A2(_00420_),
    .B(_13471_),
    .Y(_13472_));
 INVx1_ASAP7_75t_R _30778_ (.A(_00422_),
    .Y(_13473_));
 NOR2x1_ASAP7_75t_R _30779_ (.A(_13400_),
    .B(_00426_),
    .Y(_13474_));
 AO21x1_ASAP7_75t_R _30780_ (.A1(_13334_),
    .A2(_13473_),
    .B(_13474_),
    .Y(_13475_));
 AND2x6_ASAP7_75t_R _30781_ (.A(_13320_),
    .B(_13312_),
    .Y(_13476_));
 AO222x2_ASAP7_75t_R _30782_ (.A1(_13467_),
    .A2(_13469_),
    .B1(_13470_),
    .B2(_13472_),
    .C1(_13475_),
    .C2(_13476_),
    .Y(_13477_));
 INVx1_ASAP7_75t_R _30783_ (.A(_00414_),
    .Y(_13478_));
 BUFx12f_ASAP7_75t_R _30784_ (.A(_13362_),
    .Y(_13479_));
 INVx1_ASAP7_75t_R _30785_ (.A(_00415_),
    .Y(_13480_));
 BUFx12f_ASAP7_75t_R _30786_ (.A(_13315_),
    .Y(_13481_));
 NAND2x1_ASAP7_75t_R _30787_ (.A(_13481_),
    .B(_01795_),
    .Y(_13482_));
 OA21x2_ASAP7_75t_R _30788_ (.A1(_13479_),
    .A2(_13480_),
    .B(_13482_),
    .Y(_13483_));
 AND3x4_ASAP7_75t_R _30789_ (.A(_13308_),
    .B(_13309_),
    .C(_13303_),
    .Y(_13484_));
 INVx2_ASAP7_75t_R _30790_ (.A(_13484_),
    .Y(_13485_));
 AO221x1_ASAP7_75t_R _30791_ (.A1(_13478_),
    .A2(_13476_),
    .B1(_13483_),
    .B2(_13346_),
    .C(_13485_),
    .Y(_13486_));
 BUFx12f_ASAP7_75t_R _30792_ (.A(_13400_),
    .Y(_13487_));
 INVx1_ASAP7_75t_R _30793_ (.A(_00442_),
    .Y(_13488_));
 NAND2x1_ASAP7_75t_R _30794_ (.A(_13391_),
    .B(_00440_),
    .Y(_13489_));
 OA211x2_ASAP7_75t_R _30795_ (.A1(_13481_),
    .A2(_13488_),
    .B(_13489_),
    .C(_13321_),
    .Y(_13490_));
 INVx1_ASAP7_75t_R _30796_ (.A(_00443_),
    .Y(_13491_));
 NAND2x1_ASAP7_75t_R _30797_ (.A(_13391_),
    .B(_00441_),
    .Y(_13492_));
 OA211x2_ASAP7_75t_R _30798_ (.A1(_13481_),
    .A2(_13491_),
    .B(_13492_),
    .C(_13344_),
    .Y(_13493_));
 OR4x1_ASAP7_75t_R _30799_ (.A(_13487_),
    .B(_13365_),
    .C(_13490_),
    .D(_13493_),
    .Y(_13494_));
 OA211x2_ASAP7_75t_R _30800_ (.A1(_13466_),
    .A2(_13477_),
    .B(_13486_),
    .C(_13494_),
    .Y(_13495_));
 BUFx6f_ASAP7_75t_R _30801_ (.A(_13354_),
    .Y(_13496_));
 INVx1_ASAP7_75t_R _30802_ (.A(_00419_),
    .Y(_13497_));
 BUFx6f_ASAP7_75t_R _30803_ (.A(_13315_),
    .Y(_13498_));
 NAND2x1_ASAP7_75t_R _30804_ (.A(_13498_),
    .B(_00417_),
    .Y(_13499_));
 OA211x2_ASAP7_75t_R _30805_ (.A1(_13479_),
    .A2(_13497_),
    .B(_13499_),
    .C(_13345_),
    .Y(_13500_));
 INVx1_ASAP7_75t_R _30806_ (.A(_00418_),
    .Y(_13501_));
 NAND2x1_ASAP7_75t_R _30807_ (.A(_13498_),
    .B(_00416_),
    .Y(_13502_));
 OA211x2_ASAP7_75t_R _30808_ (.A1(_13402_),
    .A2(_13501_),
    .B(_13502_),
    .C(_13393_),
    .Y(_13503_));
 OR4x1_ASAP7_75t_R _30809_ (.A(_13496_),
    .B(_13461_),
    .C(_13500_),
    .D(_13503_),
    .Y(_13504_));
 INVx2_ASAP7_75t_R _30810_ (.A(_00431_),
    .Y(_13505_));
 NAND2x1_ASAP7_75t_R _30811_ (.A(_13498_),
    .B(_00429_),
    .Y(_13506_));
 OA211x2_ASAP7_75t_R _30812_ (.A1(_13402_),
    .A2(_13505_),
    .B(_13506_),
    .C(_13345_),
    .Y(_13507_));
 INVx1_ASAP7_75t_R _30813_ (.A(_00430_),
    .Y(_13508_));
 NAND2x1_ASAP7_75t_R _30814_ (.A(_13316_),
    .B(_00428_),
    .Y(_13509_));
 OA211x2_ASAP7_75t_R _30815_ (.A1(_13402_),
    .A2(_13508_),
    .B(_13509_),
    .C(_13393_),
    .Y(_13510_));
 OR4x1_ASAP7_75t_R _30816_ (.A(_13332_),
    .B(_13305_),
    .C(_13507_),
    .D(_13510_),
    .Y(_13511_));
 AO21x2_ASAP7_75t_R _30817_ (.A1(_13504_),
    .A2(_13511_),
    .B(_13329_),
    .Y(_13512_));
 NAND2x1_ASAP7_75t_R _30818_ (.A(_13331_),
    .B(_13459_),
    .Y(_13513_));
 INVx1_ASAP7_75t_R _30819_ (.A(_00435_),
    .Y(_13514_));
 NAND2x1_ASAP7_75t_R _30820_ (.A(_13347_),
    .B(_00433_),
    .Y(_13515_));
 OA211x2_ASAP7_75t_R _30821_ (.A1(_13317_),
    .A2(_13514_),
    .B(_13515_),
    .C(_13369_),
    .Y(_13516_));
 BUFx12f_ASAP7_75t_R _30822_ (.A(_13315_),
    .Y(_13517_));
 BUFx12f_ASAP7_75t_R _30823_ (.A(_13517_),
    .Y(_13518_));
 INVx1_ASAP7_75t_R _30824_ (.A(_00434_),
    .Y(_13519_));
 NAND2x1_ASAP7_75t_R _30825_ (.A(_13347_),
    .B(_00432_),
    .Y(_13520_));
 OA211x2_ASAP7_75t_R _30826_ (.A1(_13518_),
    .A2(_13519_),
    .B(_13520_),
    .C(_13352_),
    .Y(_13521_));
 OR3x1_ASAP7_75t_R _30827_ (.A(_13513_),
    .B(_13516_),
    .C(_13521_),
    .Y(_13522_));
 INVx2_ASAP7_75t_R _30828_ (.A(_00439_),
    .Y(_13523_));
 NAND2x1_ASAP7_75t_R _30829_ (.A(_13498_),
    .B(_00437_),
    .Y(_13524_));
 OA211x2_ASAP7_75t_R _30830_ (.A1(_13402_),
    .A2(_13523_),
    .B(_13524_),
    .C(_13345_),
    .Y(_13525_));
 INVx1_ASAP7_75t_R _30831_ (.A(_00438_),
    .Y(_13526_));
 NAND2x1_ASAP7_75t_R _30832_ (.A(_13316_),
    .B(_00436_),
    .Y(_13527_));
 OA211x2_ASAP7_75t_R _30833_ (.A1(_13402_),
    .A2(_13526_),
    .B(_13527_),
    .C(_13393_),
    .Y(_13528_));
 OR4x1_ASAP7_75t_R _30834_ (.A(_13332_),
    .B(_13459_),
    .C(_13525_),
    .D(_13528_),
    .Y(_13529_));
 AO21x2_ASAP7_75t_R _30835_ (.A1(_13522_),
    .A2(_13529_),
    .B(_13306_),
    .Y(_13530_));
 NAND2x2_ASAP7_75t_R _30836_ (.A(_13259_),
    .B(_13300_),
    .Y(_13531_));
 AO31x2_ASAP7_75t_R _30837_ (.A1(_13495_),
    .A2(_13512_),
    .A3(_13530_),
    .B(_13531_),
    .Y(_13532_));
 BUFx6f_ASAP7_75t_R _30838_ (.A(_00444_),
    .Y(_13533_));
 INVx4_ASAP7_75t_R _30839_ (.A(_13533_),
    .Y(_13534_));
 AOI21x1_ASAP7_75t_R _30840_ (.A1(_13236_),
    .A2(_13423_),
    .B(_13424_),
    .Y(_13535_));
 AND2x2_ASAP7_75t_R _30841_ (.A(_13259_),
    .B(_13535_),
    .Y(_13536_));
 AND4x1_ASAP7_75t_R _30842_ (.A(_13258_),
    .B(_13427_),
    .C(_13438_),
    .D(_13429_),
    .Y(_13537_));
 OA21x2_ASAP7_75t_R _30843_ (.A1(_13271_),
    .A2(_13426_),
    .B(_13328_),
    .Y(_13538_));
 AO221x1_ASAP7_75t_R _30844_ (.A1(_13534_),
    .A2(_13536_),
    .B1(_13537_),
    .B2(_13538_),
    .C(_13301_),
    .Y(_13539_));
 AO32x2_ASAP7_75t_R _30845_ (.A1(_13456_),
    .A2(_13260_),
    .A3(_13458_),
    .B1(_13532_),
    .B2(_13539_),
    .Y(_13540_));
 BUFx12f_ASAP7_75t_R _30846_ (.A(_13540_),
    .Y(_13541_));
 BUFx12f_ASAP7_75t_R _30847_ (.A(_13541_),
    .Y(_13542_));
 BUFx12f_ASAP7_75t_R _30848_ (.A(_13542_),
    .Y(_13543_));
 BUFx12f_ASAP7_75t_R _30849_ (.A(_13543_),
    .Y(_18559_));
 INVx3_ASAP7_75t_R _30850_ (.A(_13542_),
    .Y(_18552_));
 OR3x2_ASAP7_75t_R _30851_ (.A(_13344_),
    .B(_13309_),
    .C(_13460_),
    .Y(_13544_));
 INVx1_ASAP7_75t_R _30852_ (.A(_00455_),
    .Y(_13545_));
 NAND2x1_ASAP7_75t_R _30853_ (.A(_13308_),
    .B(_00451_),
    .Y(_13546_));
 OA211x2_ASAP7_75t_R _30854_ (.A1(_13356_),
    .A2(_13545_),
    .B(_13546_),
    .C(_13316_),
    .Y(_13547_));
 INVx1_ASAP7_75t_R _30855_ (.A(_00457_),
    .Y(_13548_));
 NAND2x1_ASAP7_75t_R _30856_ (.A(_13308_),
    .B(_00453_),
    .Y(_13549_));
 OA211x2_ASAP7_75t_R _30857_ (.A1(_13356_),
    .A2(_13548_),
    .B(_13549_),
    .C(_13326_),
    .Y(_13550_));
 OR3x1_ASAP7_75t_R _30858_ (.A(_13544_),
    .B(_13547_),
    .C(_13550_),
    .Y(_13551_));
 NAND2x1_ASAP7_75t_R _30859_ (.A(_13326_),
    .B(_00446_),
    .Y(_13552_));
 NAND2x1_ASAP7_75t_R _30860_ (.A(_13391_),
    .B(_01794_),
    .Y(_13553_));
 INVx1_ASAP7_75t_R _30861_ (.A(_00445_),
    .Y(_13554_));
 AO32x1_ASAP7_75t_R _30862_ (.A1(_13344_),
    .A2(_13552_),
    .A3(_13553_),
    .B1(_13554_),
    .B2(_13476_),
    .Y(_13555_));
 INVx1_ASAP7_75t_R _30863_ (.A(_00449_),
    .Y(_13556_));
 NAND2x1_ASAP7_75t_R _30864_ (.A(net1959),
    .B(_00447_),
    .Y(_13557_));
 OA211x2_ASAP7_75t_R _30865_ (.A1(_13315_),
    .A2(_13556_),
    .B(_13557_),
    .C(_13320_),
    .Y(_13558_));
 INVx1_ASAP7_75t_R _30866_ (.A(_00450_),
    .Y(_13559_));
 NAND2x1_ASAP7_75t_R _30867_ (.A(net1959),
    .B(_00448_),
    .Y(_13560_));
 OA211x2_ASAP7_75t_R _30868_ (.A1(_13315_),
    .A2(_13559_),
    .B(_13560_),
    .C(_13343_),
    .Y(_13561_));
 OR3x2_ASAP7_75t_R _30869_ (.A(_13375_),
    .B(_13558_),
    .C(_13561_),
    .Y(_13562_));
 OA21x2_ASAP7_75t_R _30870_ (.A1(_13485_),
    .A2(_13555_),
    .B(_13562_),
    .Y(_13563_));
 INVx1_ASAP7_75t_R _30871_ (.A(_00456_),
    .Y(_13564_));
 NAND2x1_ASAP7_75t_R _30872_ (.A(_13308_),
    .B(_00452_),
    .Y(_13565_));
 OA211x2_ASAP7_75t_R _30873_ (.A1(_13356_),
    .A2(_13564_),
    .B(_13565_),
    .C(_13316_),
    .Y(_13566_));
 INVx1_ASAP7_75t_R _30874_ (.A(_00458_),
    .Y(_13567_));
 NAND2x1_ASAP7_75t_R _30875_ (.A(_13308_),
    .B(_00454_),
    .Y(_13568_));
 OA211x2_ASAP7_75t_R _30876_ (.A1(_13333_),
    .A2(_13567_),
    .B(_13568_),
    .C(_13326_),
    .Y(_13569_));
 OR3x1_ASAP7_75t_R _30877_ (.A(_13417_),
    .B(_13566_),
    .C(_13569_),
    .Y(_13570_));
 INVx2_ASAP7_75t_R _30878_ (.A(_00466_),
    .Y(_13571_));
 NAND2x1_ASAP7_75t_R _30879_ (.A(_13311_),
    .B(_00464_),
    .Y(_13572_));
 OA211x2_ASAP7_75t_R _30880_ (.A1(_13315_),
    .A2(_13571_),
    .B(_13572_),
    .C(_13343_),
    .Y(_13573_));
 INVx1_ASAP7_75t_R _30881_ (.A(_00465_),
    .Y(_13574_));
 NAND2x1_ASAP7_75t_R _30882_ (.A(_13311_),
    .B(_00463_),
    .Y(_13575_));
 OA211x2_ASAP7_75t_R _30883_ (.A1(_13315_),
    .A2(_13574_),
    .B(_13575_),
    .C(_13320_),
    .Y(_13576_));
 OR3x1_ASAP7_75t_R _30884_ (.A(_13386_),
    .B(_13573_),
    .C(_13576_),
    .Y(_13577_));
 INVx1_ASAP7_75t_R _30885_ (.A(_00462_),
    .Y(_13578_));
 NAND2x1_ASAP7_75t_R _30886_ (.A(_13311_),
    .B(_00460_),
    .Y(_13579_));
 OA211x2_ASAP7_75t_R _30887_ (.A1(net1959),
    .A2(_13578_),
    .B(_13579_),
    .C(_13343_),
    .Y(_13580_));
 INVx1_ASAP7_75t_R _30888_ (.A(_00461_),
    .Y(_13581_));
 NAND2x1_ASAP7_75t_R _30889_ (.A(_13311_),
    .B(_00459_),
    .Y(_13582_));
 OA211x2_ASAP7_75t_R _30890_ (.A1(net1959),
    .A2(_13581_),
    .B(_13582_),
    .C(_13320_),
    .Y(_13583_));
 OR4x1_ASAP7_75t_R _30891_ (.A(_13303_),
    .B(_13389_),
    .C(_13580_),
    .D(_13583_),
    .Y(_13584_));
 INVx2_ASAP7_75t_R _30892_ (.A(_00473_),
    .Y(_13585_));
 NAND2x1_ASAP7_75t_R _30893_ (.A(_13311_),
    .B(_00471_),
    .Y(_13586_));
 OA211x2_ASAP7_75t_R _30894_ (.A1(net1959),
    .A2(_13585_),
    .B(_13586_),
    .C(_13320_),
    .Y(_13587_));
 INVx1_ASAP7_75t_R _30895_ (.A(_00474_),
    .Y(_13588_));
 NAND2x1_ASAP7_75t_R _30896_ (.A(_13311_),
    .B(_00472_),
    .Y(_13589_));
 OA211x2_ASAP7_75t_R _30897_ (.A1(net1959),
    .A2(_13588_),
    .B(_13589_),
    .C(_13343_),
    .Y(_13590_));
 OR4x1_ASAP7_75t_R _30898_ (.A(_13333_),
    .B(_13365_),
    .C(_13587_),
    .D(_13590_),
    .Y(_13591_));
 INVx1_ASAP7_75t_R _30899_ (.A(_00469_),
    .Y(_13592_));
 NAND2x1_ASAP7_75t_R _30900_ (.A(_13311_),
    .B(_00467_),
    .Y(_13593_));
 OA211x2_ASAP7_75t_R _30901_ (.A1(net1959),
    .A2(_13592_),
    .B(_13593_),
    .C(_13320_),
    .Y(_13594_));
 INVx2_ASAP7_75t_R _30902_ (.A(_00470_),
    .Y(_13595_));
 NAND2x1_ASAP7_75t_R _30903_ (.A(_13311_),
    .B(_00468_),
    .Y(_13596_));
 OA211x2_ASAP7_75t_R _30904_ (.A1(net1959),
    .A2(_13595_),
    .B(_13596_),
    .C(_13343_),
    .Y(_13597_));
 OR4x1_ASAP7_75t_R _30905_ (.A(_13330_),
    .B(_13365_),
    .C(_13594_),
    .D(_13597_),
    .Y(_13598_));
 AND4x1_ASAP7_75t_R _30906_ (.A(_13577_),
    .B(_13584_),
    .C(_13591_),
    .D(_13598_),
    .Y(_13599_));
 AND4x1_ASAP7_75t_R _30907_ (.A(_13551_),
    .B(_13563_),
    .C(_13570_),
    .D(_13599_),
    .Y(_13600_));
 BUFx12f_ASAP7_75t_R _30908_ (.A(_13600_),
    .Y(_13601_));
 BUFx12f_ASAP7_75t_R _30909_ (.A(_02208_),
    .Y(_13602_));
 INVx4_ASAP7_75t_R _30910_ (.A(_13602_),
    .Y(_13603_));
 AND4x1_ASAP7_75t_R _30911_ (.A(_13603_),
    .B(_13439_),
    .C(_13444_),
    .D(_13457_),
    .Y(_13604_));
 AO21x1_ASAP7_75t_R _30912_ (.A1(_13426_),
    .A2(_13429_),
    .B(_13271_),
    .Y(_13605_));
 AND4x1_ASAP7_75t_R _30913_ (.A(_13332_),
    .B(_13258_),
    .C(_13427_),
    .D(_13438_),
    .Y(_13606_));
 OR3x1_ASAP7_75t_R _30914_ (.A(_13242_),
    .B(_13296_),
    .C(_13299_),
    .Y(_13607_));
 OAI21x1_ASAP7_75t_R _30915_ (.A1(_13602_),
    .A2(_13236_),
    .B(_13607_),
    .Y(_13608_));
 AO21x1_ASAP7_75t_R _30916_ (.A1(_13533_),
    .A2(_13535_),
    .B(_13271_),
    .Y(_13609_));
 AO221x1_ASAP7_75t_R _30917_ (.A1(_13605_),
    .A2(_13606_),
    .B1(_13608_),
    .B2(_13437_),
    .C(_13609_),
    .Y(_13610_));
 OA22x2_ASAP7_75t_R _30918_ (.A1(_13531_),
    .A2(_13601_),
    .B1(_13604_),
    .B2(_13610_),
    .Y(_13611_));
 BUFx6f_ASAP7_75t_R _30919_ (.A(_13611_),
    .Y(_13612_));
 INVx1_ASAP7_75t_R _30920_ (.A(_13612_),
    .Y(_13613_));
 BUFx6f_ASAP7_75t_R _30921_ (.A(_13613_),
    .Y(_13614_));
 BUFx12f_ASAP7_75t_R _30922_ (.A(_13614_),
    .Y(_18565_));
 BUFx12f_ASAP7_75t_R _30923_ (.A(_13612_),
    .Y(_18563_));
 NOR2x1_ASAP7_75t_R _30924_ (.A(_13496_),
    .B(_13305_),
    .Y(_13615_));
 BUFx6f_ASAP7_75t_R _30925_ (.A(net1977),
    .Y(_13616_));
 INVx2_ASAP7_75t_R _30926_ (.A(_00503_),
    .Y(_13617_));
 NAND2x1_ASAP7_75t_R _30927_ (.A(_13517_),
    .B(_00501_),
    .Y(_13618_));
 OA211x2_ASAP7_75t_R _30928_ (.A1(_13616_),
    .A2(_13617_),
    .B(_13618_),
    .C(_13329_),
    .Y(_13619_));
 INVx2_ASAP7_75t_R _30929_ (.A(_00495_),
    .Y(_13620_));
 NAND2x1_ASAP7_75t_R _30930_ (.A(_13517_),
    .B(_00493_),
    .Y(_13621_));
 OA211x2_ASAP7_75t_R _30931_ (.A1(_13616_),
    .A2(_13620_),
    .B(_13621_),
    .C(_13309_),
    .Y(_13622_));
 OR3x1_ASAP7_75t_R _30932_ (.A(_13346_),
    .B(_13619_),
    .C(_13622_),
    .Y(_13623_));
 INVx2_ASAP7_75t_R _30933_ (.A(_00504_),
    .Y(_13624_));
 NAND2x1_ASAP7_75t_R _30934_ (.A(_13517_),
    .B(_00502_),
    .Y(_13625_));
 OA211x2_ASAP7_75t_R _30935_ (.A1(_13616_),
    .A2(_13624_),
    .B(_13625_),
    .C(_13329_),
    .Y(_13626_));
 INVx2_ASAP7_75t_R _30936_ (.A(_00496_),
    .Y(_13627_));
 NAND2x1_ASAP7_75t_R _30937_ (.A(_13517_),
    .B(_00494_),
    .Y(_13628_));
 OA211x2_ASAP7_75t_R _30938_ (.A1(_13616_),
    .A2(_13627_),
    .B(_13628_),
    .C(_13309_),
    .Y(_13629_));
 OR3x1_ASAP7_75t_R _30939_ (.A(_13322_),
    .B(_13626_),
    .C(_13629_),
    .Y(_13630_));
 AND3x1_ASAP7_75t_R _30940_ (.A(_13615_),
    .B(_13623_),
    .C(_13630_),
    .Y(_13631_));
 AND2x6_ASAP7_75t_R _30941_ (.A(_13321_),
    .B(_13330_),
    .Y(_13632_));
 INVx2_ASAP7_75t_R _30942_ (.A(_00485_),
    .Y(_13633_));
 NOR2x1_ASAP7_75t_R _30943_ (.A(_13481_),
    .B(_00487_),
    .Y(_13634_));
 AO21x1_ASAP7_75t_R _30944_ (.A1(_13479_),
    .A2(_13633_),
    .B(_13634_),
    .Y(_13635_));
 INVx2_ASAP7_75t_R _30945_ (.A(_00488_),
    .Y(_13636_));
 NOR2x2_ASAP7_75t_R _30946_ (.A(_13321_),
    .B(_13308_),
    .Y(_13637_));
 NAND2x1_ASAP7_75t_R _30947_ (.A(_13517_),
    .B(_00486_),
    .Y(_13638_));
 OA211x2_ASAP7_75t_R _30948_ (.A1(_13616_),
    .A2(_13636_),
    .B(_13637_),
    .C(_13638_),
    .Y(_13639_));
 AO21x1_ASAP7_75t_R _30949_ (.A1(_13632_),
    .A2(_13635_),
    .B(_13639_),
    .Y(_13640_));
 AND2x6_ASAP7_75t_R _30950_ (.A(_13344_),
    .B(_13308_),
    .Y(_13641_));
 INVx1_ASAP7_75t_R _30951_ (.A(_00482_),
    .Y(_13642_));
 NOR2x1_ASAP7_75t_R _30952_ (.A(_13338_),
    .B(_00484_),
    .Y(_13643_));
 AO21x1_ASAP7_75t_R _30953_ (.A1(_13479_),
    .A2(_13642_),
    .B(_13643_),
    .Y(_13644_));
 INVx2_ASAP7_75t_R _30954_ (.A(_00483_),
    .Y(_13645_));
 AND2x6_ASAP7_75t_R _30955_ (.A(_13320_),
    .B(_13307_),
    .Y(_13646_));
 NAND2x1_ASAP7_75t_R _30956_ (.A(_13391_),
    .B(_00481_),
    .Y(_13647_));
 OA211x2_ASAP7_75t_R _30957_ (.A1(_13616_),
    .A2(_13645_),
    .B(_13646_),
    .C(_13647_),
    .Y(_13648_));
 AO21x1_ASAP7_75t_R _30958_ (.A1(_13641_),
    .A2(_13644_),
    .B(_13648_),
    .Y(_13649_));
 OA211x2_ASAP7_75t_R _30959_ (.A1(_13640_),
    .A2(_13649_),
    .B(_13329_),
    .C(_13305_),
    .Y(_13650_));
 BUFx6f_ASAP7_75t_R _30960_ (.A(_13400_),
    .Y(_13651_));
 AND2x2_ASAP7_75t_R _30961_ (.A(_13651_),
    .B(_13407_),
    .Y(_13652_));
 INVx2_ASAP7_75t_R _30962_ (.A(_00497_),
    .Y(_13653_));
 NOR2x1_ASAP7_75t_R _30963_ (.A(_13363_),
    .B(_00499_),
    .Y(_13654_));
 AO21x1_ASAP7_75t_R _30964_ (.A1(_13317_),
    .A2(_13653_),
    .B(_13654_),
    .Y(_13655_));
 INVx2_ASAP7_75t_R _30965_ (.A(_00500_),
    .Y(_13656_));
 NAND2x1_ASAP7_75t_R _30966_ (.A(_13498_),
    .B(_00498_),
    .Y(_13657_));
 OA211x2_ASAP7_75t_R _30967_ (.A1(_13479_),
    .A2(_13656_),
    .B(_13657_),
    .C(_13369_),
    .Y(_13658_));
 AO21x1_ASAP7_75t_R _30968_ (.A1(_13353_),
    .A2(_13655_),
    .B(_13658_),
    .Y(_13659_));
 INVx2_ASAP7_75t_R _30969_ (.A(_00492_),
    .Y(_13660_));
 NAND2x1_ASAP7_75t_R _30970_ (.A(_13316_),
    .B(_00490_),
    .Y(_13661_));
 OA211x2_ASAP7_75t_R _30971_ (.A1(_13402_),
    .A2(_13660_),
    .B(_13661_),
    .C(_13345_),
    .Y(_13662_));
 INVx2_ASAP7_75t_R _30972_ (.A(_00491_),
    .Y(_13663_));
 NAND2x1_ASAP7_75t_R _30973_ (.A(_13316_),
    .B(_00489_),
    .Y(_13664_));
 OA211x2_ASAP7_75t_R _30974_ (.A1(_13402_),
    .A2(_13663_),
    .B(_13664_),
    .C(_13393_),
    .Y(_13665_));
 AND2x6_ASAP7_75t_R _30975_ (.A(_13460_),
    .B(_13310_),
    .Y(_13666_));
 OA21x2_ASAP7_75t_R _30976_ (.A1(_13662_),
    .A2(_13665_),
    .B(_13666_),
    .Y(_13667_));
 AO21x1_ASAP7_75t_R _30977_ (.A1(_13652_),
    .A2(_13659_),
    .B(_13667_),
    .Y(_13668_));
 BUFx12f_ASAP7_75t_R _30978_ (.A(_13331_),
    .Y(_13669_));
 NAND2x2_ASAP7_75t_R _30979_ (.A(_13321_),
    .B(_13326_),
    .Y(_13670_));
 AND2x2_ASAP7_75t_R _30980_ (.A(_13316_),
    .B(_01793_),
    .Y(_13671_));
 AO21x1_ASAP7_75t_R _30981_ (.A1(_13313_),
    .A2(_00476_),
    .B(_13671_),
    .Y(_13672_));
 BUFx6f_ASAP7_75t_R _30982_ (.A(_13352_),
    .Y(_13673_));
 OAI22x1_ASAP7_75t_R _30983_ (.A1(_00475_),
    .A2(_13670_),
    .B1(_13672_),
    .B2(_13673_),
    .Y(_13674_));
 BUFx12f_ASAP7_75t_R _30984_ (.A(_13400_),
    .Y(_13675_));
 INVx2_ASAP7_75t_R _30985_ (.A(_00480_),
    .Y(_13676_));
 NAND2x1_ASAP7_75t_R _30986_ (.A(_13362_),
    .B(_00478_),
    .Y(_13677_));
 OA211x2_ASAP7_75t_R _30987_ (.A1(_13498_),
    .A2(_13676_),
    .B(_13677_),
    .C(_13344_),
    .Y(_13678_));
 INVx2_ASAP7_75t_R _30988_ (.A(_00479_),
    .Y(_13679_));
 NAND2x1_ASAP7_75t_R _30989_ (.A(_13362_),
    .B(_00477_),
    .Y(_13680_));
 OA211x2_ASAP7_75t_R _30990_ (.A1(_13498_),
    .A2(_13679_),
    .B(_13680_),
    .C(_13321_),
    .Y(_13681_));
 OR3x1_ASAP7_75t_R _30991_ (.A(_13675_),
    .B(_13678_),
    .C(_13681_),
    .Y(_13682_));
 OA211x2_ASAP7_75t_R _30992_ (.A1(_13669_),
    .A2(_13674_),
    .B(_13682_),
    .C(_13374_),
    .Y(_13683_));
 OR4x1_ASAP7_75t_R _30993_ (.A(_13631_),
    .B(_13650_),
    .C(_13668_),
    .D(_13683_),
    .Y(_13684_));
 BUFx12f_ASAP7_75t_R _30994_ (.A(_01520_),
    .Y(_13685_));
 INVx3_ASAP7_75t_R _30995_ (.A(_13685_),
    .Y(_13686_));
 AND2x2_ASAP7_75t_R _30996_ (.A(_13686_),
    .B(_13259_),
    .Y(_13687_));
 BUFx12f_ASAP7_75t_R _30997_ (.A(_13329_),
    .Y(_13688_));
 AND4x1_ASAP7_75t_R _30998_ (.A(_13688_),
    .B(_13439_),
    .C(_13605_),
    .D(_13531_),
    .Y(_13689_));
 AOI221x1_ASAP7_75t_R _30999_ (.A1(_13301_),
    .A2(_13684_),
    .B1(_13687_),
    .B2(_13458_),
    .C(_13689_),
    .Y(_13690_));
 INVx3_ASAP7_75t_R _31000_ (.A(_13690_),
    .Y(_13691_));
 BUFx12f_ASAP7_75t_R _31001_ (.A(_13691_),
    .Y(_18568_));
 BUFx12f_ASAP7_75t_R _31002_ (.A(_13690_),
    .Y(_18570_));
 INVx2_ASAP7_75t_R _31003_ (.A(_00339_),
    .Y(_13692_));
 AND2x2_ASAP7_75t_R _31004_ (.A(_13692_),
    .B(_13260_),
    .Y(_13693_));
 AND2x6_ASAP7_75t_R _31005_ (.A(_13331_),
    .B(_13309_),
    .Y(_13694_));
 BUFx12f_ASAP7_75t_R _31006_ (.A(_13338_),
    .Y(_13695_));
 AND2x2_ASAP7_75t_R _31007_ (.A(_13695_),
    .B(_00507_),
    .Y(_13696_));
 AO21x1_ASAP7_75t_R _31008_ (.A1(_13314_),
    .A2(_00509_),
    .B(_13696_),
    .Y(_13697_));
 NAND2x1_ASAP7_75t_R _31009_ (.A(_13694_),
    .B(_13697_),
    .Y(_13698_));
 INVx1_ASAP7_75t_R _31010_ (.A(_00515_),
    .Y(_13699_));
 NAND2x1_ASAP7_75t_R _31011_ (.A(_13334_),
    .B(_00511_),
    .Y(_13700_));
 BUFx12f_ASAP7_75t_R _31012_ (.A(_13481_),
    .Y(_13701_));
 OA211x2_ASAP7_75t_R _31013_ (.A1(_13487_),
    .A2(_13699_),
    .B(_13700_),
    .C(_13701_),
    .Y(_13702_));
 INVx1_ASAP7_75t_R _31014_ (.A(_00517_),
    .Y(_13703_));
 NAND2x1_ASAP7_75t_R _31015_ (.A(_13334_),
    .B(_00513_),
    .Y(_13704_));
 OA211x2_ASAP7_75t_R _31016_ (.A1(_13487_),
    .A2(_13703_),
    .B(_13704_),
    .C(_13327_),
    .Y(_13705_));
 OR3x1_ASAP7_75t_R _31017_ (.A(_13459_),
    .B(_13702_),
    .C(_13705_),
    .Y(_13706_));
 AO21x1_ASAP7_75t_R _31018_ (.A1(_13698_),
    .A2(_13706_),
    .B(_13434_),
    .Y(_13707_));
 AND2x2_ASAP7_75t_R _31019_ (.A(_13317_),
    .B(_01792_),
    .Y(_13708_));
 AO21x1_ASAP7_75t_R _31020_ (.A1(_13314_),
    .A2(_00506_),
    .B(_13708_),
    .Y(_13709_));
 OA22x2_ASAP7_75t_R _31021_ (.A1(_00505_),
    .A2(_13670_),
    .B1(_13709_),
    .B2(_13323_),
    .Y(_13710_));
 BUFx12f_ASAP7_75t_R _31022_ (.A(_13333_),
    .Y(_13711_));
 BUFx6f_ASAP7_75t_R _31023_ (.A(_13711_),
    .Y(_13712_));
 INVx1_ASAP7_75t_R _31024_ (.A(_00516_),
    .Y(_13713_));
 NAND2x1_ASAP7_75t_R _31025_ (.A(_13712_),
    .B(_00512_),
    .Y(_13714_));
 OA21x2_ASAP7_75t_R _31026_ (.A1(_13712_),
    .A2(_13713_),
    .B(_13714_),
    .Y(_13715_));
 NAND2x1_ASAP7_75t_R _31027_ (.A(_13340_),
    .B(_13416_),
    .Y(_13716_));
 OAI21x1_ASAP7_75t_R _31028_ (.A1(_13715_),
    .A2(_13716_),
    .B(_13306_),
    .Y(_13717_));
 AND2x2_ASAP7_75t_R _31029_ (.A(_13334_),
    .B(_00514_),
    .Y(_13718_));
 AO21x1_ASAP7_75t_R _31030_ (.A1(_13332_),
    .A2(_00518_),
    .B(_13718_),
    .Y(_13719_));
 AND2x2_ASAP7_75t_R _31031_ (.A(_13378_),
    .B(_00508_),
    .Y(_13720_));
 AO21x1_ASAP7_75t_R _31032_ (.A1(_13327_),
    .A2(_00510_),
    .B(_13720_),
    .Y(_13721_));
 AO33x2_ASAP7_75t_R _31033_ (.A1(_13328_),
    .A2(_13416_),
    .A3(_13719_),
    .B1(_13721_),
    .B2(_13637_),
    .B3(_13459_),
    .Y(_13722_));
 AOI211x1_ASAP7_75t_R _31034_ (.A1(_13310_),
    .A2(_13710_),
    .B(_13717_),
    .C(_13722_),
    .Y(_13723_));
 BUFx12f_ASAP7_75t_R _31035_ (.A(_13459_),
    .Y(_13724_));
 BUFx12f_ASAP7_75t_R _31036_ (.A(_13363_),
    .Y(_13725_));
 INVx1_ASAP7_75t_R _31037_ (.A(_00524_),
    .Y(_13726_));
 NOR2x1_ASAP7_75t_R _31038_ (.A(_13317_),
    .B(_00526_),
    .Y(_13727_));
 AO21x1_ASAP7_75t_R _31039_ (.A1(_13725_),
    .A2(_13726_),
    .B(_13727_),
    .Y(_13728_));
 INVx1_ASAP7_75t_R _31040_ (.A(_00525_),
    .Y(_13729_));
 NAND2x1_ASAP7_75t_R _31041_ (.A(_13479_),
    .B(_00523_),
    .Y(_13730_));
 OA211x2_ASAP7_75t_R _31042_ (.A1(_13695_),
    .A2(_13729_),
    .B(_13730_),
    .C(_13322_),
    .Y(_13731_));
 AO21x1_ASAP7_75t_R _31043_ (.A1(_13434_),
    .A2(_13728_),
    .B(_13731_),
    .Y(_13732_));
 INVx1_ASAP7_75t_R _31044_ (.A(_00531_),
    .Y(_13733_));
 BUFx6f_ASAP7_75t_R _31045_ (.A(_13378_),
    .Y(_13734_));
 NOR2x1_ASAP7_75t_R _31046_ (.A(_13734_),
    .B(_00533_),
    .Y(_13735_));
 AO21x1_ASAP7_75t_R _31047_ (.A1(_13340_),
    .A2(_13733_),
    .B(_13735_),
    .Y(_13736_));
 AND2x2_ASAP7_75t_R _31048_ (.A(_13353_),
    .B(_13329_),
    .Y(_13737_));
 BUFx12f_ASAP7_75t_R _31049_ (.A(_13518_),
    .Y(_13738_));
 INVx1_ASAP7_75t_R _31050_ (.A(_00534_),
    .Y(_13739_));
 NAND2x1_ASAP7_75t_R _31051_ (.A(_13725_),
    .B(_00532_),
    .Y(_13740_));
 OA211x2_ASAP7_75t_R _31052_ (.A1(_13738_),
    .A2(_13739_),
    .B(_13416_),
    .C(_13740_),
    .Y(_13741_));
 AO221x1_ASAP7_75t_R _31053_ (.A1(_13724_),
    .A2(_13732_),
    .B1(_13736_),
    .B2(_13737_),
    .C(_13741_),
    .Y(_13742_));
 INVx2_ASAP7_75t_R _31054_ (.A(_00527_),
    .Y(_13743_));
 NOR2x1_ASAP7_75t_R _31055_ (.A(_13725_),
    .B(_00529_),
    .Y(_13744_));
 AO21x1_ASAP7_75t_R _31056_ (.A1(_13738_),
    .A2(_13743_),
    .B(_13744_),
    .Y(_13745_));
 BUFx6f_ASAP7_75t_R _31057_ (.A(_13479_),
    .Y(_13746_));
 INVx2_ASAP7_75t_R _31058_ (.A(_00530_),
    .Y(_13747_));
 BUFx12f_ASAP7_75t_R _31059_ (.A(_13338_),
    .Y(_13748_));
 NAND2x1_ASAP7_75t_R _31060_ (.A(_13748_),
    .B(_00528_),
    .Y(_13749_));
 BUFx6f_ASAP7_75t_R _31061_ (.A(_13369_),
    .Y(_13750_));
 OA211x2_ASAP7_75t_R _31062_ (.A1(_13746_),
    .A2(_13747_),
    .B(_13749_),
    .C(_13750_),
    .Y(_13751_));
 AO21x1_ASAP7_75t_R _31063_ (.A1(_13323_),
    .A2(_13745_),
    .B(_13751_),
    .Y(_13752_));
 BUFx6f_ASAP7_75t_R _31064_ (.A(_13363_),
    .Y(_13753_));
 INVx2_ASAP7_75t_R _31065_ (.A(_00522_),
    .Y(_13754_));
 NAND2x1_ASAP7_75t_R _31066_ (.A(_13339_),
    .B(_00520_),
    .Y(_13755_));
 OA211x2_ASAP7_75t_R _31067_ (.A1(_13753_),
    .A2(_13754_),
    .B(_13755_),
    .C(_13346_),
    .Y(_13756_));
 INVx2_ASAP7_75t_R _31068_ (.A(_00521_),
    .Y(_13757_));
 NAND2x1_ASAP7_75t_R _31069_ (.A(_13339_),
    .B(_00519_),
    .Y(_13758_));
 OA211x2_ASAP7_75t_R _31070_ (.A1(_13753_),
    .A2(_13757_),
    .B(_13758_),
    .C(_13322_),
    .Y(_13759_));
 OA21x2_ASAP7_75t_R _31071_ (.A1(_13756_),
    .A2(_13759_),
    .B(_13666_),
    .Y(_13760_));
 AO21x1_ASAP7_75t_R _31072_ (.A1(_13652_),
    .A2(_13752_),
    .B(_13760_),
    .Y(_13761_));
 AO221x1_ASAP7_75t_R _31073_ (.A1(_13707_),
    .A2(_13723_),
    .B1(_13742_),
    .B2(_13615_),
    .C(_13761_),
    .Y(_13762_));
 BUFx12f_ASAP7_75t_R _31074_ (.A(_13531_),
    .Y(_13763_));
 BUFx12f_ASAP7_75t_R _31075_ (.A(_13461_),
    .Y(_13764_));
 AND4x1_ASAP7_75t_R _31076_ (.A(_13764_),
    .B(_13259_),
    .C(_13426_),
    .D(_13429_),
    .Y(_13765_));
 AND3x1_ASAP7_75t_R _31077_ (.A(_13439_),
    .B(_13763_),
    .C(_13765_),
    .Y(_13766_));
 AOI221x1_ASAP7_75t_R _31078_ (.A1(_13458_),
    .A2(_13693_),
    .B1(_13762_),
    .B2(_13302_),
    .C(_13766_),
    .Y(_13767_));
 INVx4_ASAP7_75t_R _31079_ (.A(_13767_),
    .Y(_13768_));
 BUFx12f_ASAP7_75t_R _31080_ (.A(_13768_),
    .Y(_18573_));
 BUFx6f_ASAP7_75t_R _31081_ (.A(_13767_),
    .Y(_13769_));
 BUFx12f_ASAP7_75t_R _31082_ (.A(_13769_),
    .Y(_18575_));
 INVx2_ASAP7_75t_R _31083_ (.A(_00540_),
    .Y(_13770_));
 NAND2x1_ASAP7_75t_R _31084_ (.A(_13348_),
    .B(_00538_),
    .Y(_13771_));
 OA21x2_ASAP7_75t_R _31085_ (.A1(_13734_),
    .A2(_13770_),
    .B(_13771_),
    .Y(_13772_));
 BUFx6f_ASAP7_75t_R _31086_ (.A(_13378_),
    .Y(_13773_));
 INVx2_ASAP7_75t_R _31087_ (.A(_00539_),
    .Y(_13774_));
 NAND2x1_ASAP7_75t_R _31088_ (.A(_13339_),
    .B(_00537_),
    .Y(_13775_));
 OA211x2_ASAP7_75t_R _31089_ (.A1(_13773_),
    .A2(_13774_),
    .B(_13775_),
    .C(_13673_),
    .Y(_13776_));
 AO21x1_ASAP7_75t_R _31090_ (.A1(_13434_),
    .A2(_13772_),
    .B(_13776_),
    .Y(_13777_));
 INVx1_ASAP7_75t_R _31091_ (.A(_00553_),
    .Y(_13778_));
 NOR2x1_ASAP7_75t_R _31092_ (.A(_13725_),
    .B(_00555_),
    .Y(_13779_));
 AO21x1_ASAP7_75t_R _31093_ (.A1(_13738_),
    .A2(_13778_),
    .B(_13779_),
    .Y(_13780_));
 INVx2_ASAP7_75t_R _31094_ (.A(_00556_),
    .Y(_13781_));
 NAND2x1_ASAP7_75t_R _31095_ (.A(_13748_),
    .B(_00554_),
    .Y(_13782_));
 OA211x2_ASAP7_75t_R _31096_ (.A1(_13746_),
    .A2(_13781_),
    .B(_13782_),
    .C(_13750_),
    .Y(_13783_));
 AO21x2_ASAP7_75t_R _31097_ (.A1(_13323_),
    .A2(_13780_),
    .B(_13783_),
    .Y(_13784_));
 OA22x2_ASAP7_75t_R _31098_ (.A1(_13375_),
    .A2(_13777_),
    .B1(_13784_),
    .B2(_13386_),
    .Y(_13785_));
 AND2x2_ASAP7_75t_R _31099_ (.A(_13348_),
    .B(_01791_),
    .Y(_13786_));
 AO21x1_ASAP7_75t_R _31100_ (.A1(_13314_),
    .A2(_00536_),
    .B(_13786_),
    .Y(_13787_));
 OA22x2_ASAP7_75t_R _31101_ (.A1(_00535_),
    .A2(_13670_),
    .B1(_13787_),
    .B2(_13323_),
    .Y(_13788_));
 INVx2_ASAP7_75t_R _31102_ (.A(_00552_),
    .Y(_13789_));
 NAND2x1_ASAP7_75t_R _31103_ (.A(_13753_),
    .B(_00550_),
    .Y(_13790_));
 OA211x2_ASAP7_75t_R _31104_ (.A1(_13340_),
    .A2(_13789_),
    .B(_13790_),
    .C(_13750_),
    .Y(_13791_));
 INVx2_ASAP7_75t_R _31105_ (.A(_00551_),
    .Y(_13792_));
 NAND2x1_ASAP7_75t_R _31106_ (.A(_13773_),
    .B(_00549_),
    .Y(_13793_));
 OA211x2_ASAP7_75t_R _31107_ (.A1(_13340_),
    .A2(_13792_),
    .B(_13793_),
    .C(_13353_),
    .Y(_13794_));
 NOR2x1_ASAP7_75t_R _31108_ (.A(_13791_),
    .B(_13794_),
    .Y(_13795_));
 AOI22x1_ASAP7_75t_R _31109_ (.A1(_13484_),
    .A2(_13788_),
    .B1(_13795_),
    .B2(_13666_),
    .Y(_13796_));
 AND2x2_ASAP7_75t_R _31110_ (.A(_13339_),
    .B(_13461_),
    .Y(_13797_));
 OR2x2_ASAP7_75t_R _31111_ (.A(_13487_),
    .B(_00562_),
    .Y(_13798_));
 OAI21x1_ASAP7_75t_R _31112_ (.A1(_13669_),
    .A2(_00558_),
    .B(_13798_),
    .Y(_13799_));
 INVx1_ASAP7_75t_R _31113_ (.A(_00546_),
    .Y(_13800_));
 AND2x2_ASAP7_75t_R _31114_ (.A(_13616_),
    .B(_13304_),
    .Y(_13801_));
 NAND2x1_ASAP7_75t_R _31115_ (.A(_13487_),
    .B(_00542_),
    .Y(_13802_));
 OA211x2_ASAP7_75t_R _31116_ (.A1(_13712_),
    .A2(_13800_),
    .B(_13801_),
    .C(_13802_),
    .Y(_13803_));
 INVx2_ASAP7_75t_R _31117_ (.A(_00564_),
    .Y(_13804_));
 NOR2x1_ASAP7_75t_R _31118_ (.A(_13701_),
    .B(_13388_),
    .Y(_13805_));
 NAND2x1_ASAP7_75t_R _31119_ (.A(_13651_),
    .B(_00560_),
    .Y(_13806_));
 OA211x2_ASAP7_75t_R _31120_ (.A1(_13712_),
    .A2(_13804_),
    .B(_13805_),
    .C(_13806_),
    .Y(_13807_));
 AOI211x1_ASAP7_75t_R _31121_ (.A1(_13797_),
    .A2(_13799_),
    .B(_13803_),
    .C(_13807_),
    .Y(_13808_));
 NAND2x1_ASAP7_75t_R _31122_ (.A(_13314_),
    .B(_13305_),
    .Y(_13809_));
 AND2x2_ASAP7_75t_R _31123_ (.A(_13675_),
    .B(_00544_),
    .Y(_13810_));
 AO21x1_ASAP7_75t_R _31124_ (.A1(_13669_),
    .A2(_00548_),
    .B(_13810_),
    .Y(_13811_));
 OA21x2_ASAP7_75t_R _31125_ (.A1(_13809_),
    .A2(_13811_),
    .B(_13416_),
    .Y(_13812_));
 BUFx12f_ASAP7_75t_R _31126_ (.A(_13725_),
    .Y(_13813_));
 BUFx12f_ASAP7_75t_R _31127_ (.A(_13487_),
    .Y(_13814_));
 INVx2_ASAP7_75t_R _31128_ (.A(_00557_),
    .Y(_13815_));
 NOR2x1_ASAP7_75t_R _31129_ (.A(_13496_),
    .B(_00561_),
    .Y(_13816_));
 AO21x1_ASAP7_75t_R _31130_ (.A1(_13814_),
    .A2(_13815_),
    .B(_13816_),
    .Y(_13817_));
 INVx2_ASAP7_75t_R _31131_ (.A(_00563_),
    .Y(_13818_));
 NAND2x1_ASAP7_75t_R _31132_ (.A(_13651_),
    .B(_00559_),
    .Y(_13819_));
 OA211x2_ASAP7_75t_R _31133_ (.A1(_13712_),
    .A2(_13818_),
    .B(_13819_),
    .C(_13314_),
    .Y(_13820_));
 AOI211x1_ASAP7_75t_R _31134_ (.A1(_13813_),
    .A2(_13817_),
    .B(_13820_),
    .C(_13408_),
    .Y(_13821_));
 INVx2_ASAP7_75t_R _31135_ (.A(_00547_),
    .Y(_13822_));
 NAND2x1_ASAP7_75t_R _31136_ (.A(_13651_),
    .B(_00543_),
    .Y(_13823_));
 OA21x2_ASAP7_75t_R _31137_ (.A1(_13712_),
    .A2(_13822_),
    .B(_13823_),
    .Y(_13824_));
 INVx1_ASAP7_75t_R _31138_ (.A(_00545_),
    .Y(_13825_));
 NAND2x1_ASAP7_75t_R _31139_ (.A(_13651_),
    .B(_00541_),
    .Y(_13826_));
 OA211x2_ASAP7_75t_R _31140_ (.A1(_13712_),
    .A2(_13825_),
    .B(_13826_),
    .C(_13738_),
    .Y(_13827_));
 AOI211x1_ASAP7_75t_R _31141_ (.A1(_13328_),
    .A2(_13824_),
    .B(_13827_),
    .C(_13544_),
    .Y(_13828_));
 AOI211x1_ASAP7_75t_R _31142_ (.A1(_13808_),
    .A2(_13812_),
    .B(_13821_),
    .C(_13828_),
    .Y(_13829_));
 AND3x4_ASAP7_75t_R _31143_ (.A(_13785_),
    .B(_13796_),
    .C(_13829_),
    .Y(_13830_));
 BUFx12f_ASAP7_75t_R _31144_ (.A(_01515_),
    .Y(_13831_));
 INVx3_ASAP7_75t_R _31145_ (.A(_13831_),
    .Y(_13832_));
 OR3x1_ASAP7_75t_R _31146_ (.A(_13296_),
    .B(_13297_),
    .C(_13299_),
    .Y(_13833_));
 AND4x1_ASAP7_75t_R _31147_ (.A(_13259_),
    .B(_13427_),
    .C(_13426_),
    .D(_13833_),
    .Y(_13834_));
 AND2x2_ASAP7_75t_R _31148_ (.A(_13832_),
    .B(_13834_),
    .Y(_13835_));
 AOI21x1_ASAP7_75t_R _31149_ (.A1(_13302_),
    .A2(_13830_),
    .B(_13835_),
    .Y(_13836_));
 INVx4_ASAP7_75t_R _31150_ (.A(_13836_),
    .Y(_18578_));
 BUFx6f_ASAP7_75t_R _31151_ (.A(_13836_),
    .Y(_18580_));
 BUFx12f_ASAP7_75t_R _31152_ (.A(_00411_),
    .Y(_13837_));
 INVx2_ASAP7_75t_R _31153_ (.A(_13837_),
    .Y(_13838_));
 BUFx12f_ASAP7_75t_R _31154_ (.A(_13834_),
    .Y(_13839_));
 AND3x4_ASAP7_75t_R _31155_ (.A(_13673_),
    .B(_13329_),
    .C(_13388_),
    .Y(_13840_));
 INVx2_ASAP7_75t_R _31156_ (.A(_00577_),
    .Y(_13841_));
 BUFx12f_ASAP7_75t_R _31157_ (.A(_13308_),
    .Y(_13842_));
 NAND2x1_ASAP7_75t_R _31158_ (.A(_13842_),
    .B(_00573_),
    .Y(_13843_));
 OA211x2_ASAP7_75t_R _31159_ (.A1(_13711_),
    .A2(_13841_),
    .B(_13843_),
    .C(_13313_),
    .Y(_13844_));
 INVx1_ASAP7_75t_R _31160_ (.A(_00575_),
    .Y(_13845_));
 NAND2x1_ASAP7_75t_R _31161_ (.A(_13842_),
    .B(_00571_),
    .Y(_13846_));
 OA211x2_ASAP7_75t_R _31162_ (.A1(_13711_),
    .A2(_13845_),
    .B(_13846_),
    .C(_13317_),
    .Y(_13847_));
 NOR2x1_ASAP7_75t_R _31163_ (.A(_13844_),
    .B(_13847_),
    .Y(_13848_));
 INVx1_ASAP7_75t_R _31164_ (.A(_00593_),
    .Y(_13849_));
 NAND2x1_ASAP7_75t_R _31165_ (.A(_13842_),
    .B(_00589_),
    .Y(_13850_));
 OA211x2_ASAP7_75t_R _31166_ (.A1(_13711_),
    .A2(_13849_),
    .B(_13850_),
    .C(_13313_),
    .Y(_13851_));
 INVx1_ASAP7_75t_R _31167_ (.A(_00591_),
    .Y(_13852_));
 NAND2x1_ASAP7_75t_R _31168_ (.A(_13842_),
    .B(_00587_),
    .Y(_13853_));
 OA211x2_ASAP7_75t_R _31169_ (.A1(_13711_),
    .A2(_13852_),
    .B(_13853_),
    .C(_13317_),
    .Y(_13854_));
 NOR2x1_ASAP7_75t_R _31170_ (.A(_13851_),
    .B(_13854_),
    .Y(_13855_));
 AND2x6_ASAP7_75t_R _31171_ (.A(_13353_),
    .B(_13407_),
    .Y(_13856_));
 AOI22x1_ASAP7_75t_R _31172_ (.A1(_13840_),
    .A2(_13848_),
    .B1(_13855_),
    .B2(_13856_),
    .Y(_13857_));
 OR2x6_ASAP7_75t_R _31173_ (.A(_13352_),
    .B(_13459_),
    .Y(_13858_));
 NAND2x1_ASAP7_75t_R _31174_ (.A(_13695_),
    .B(_13461_),
    .Y(_13859_));
 AND2x2_ASAP7_75t_R _31175_ (.A(_13356_),
    .B(_00588_),
    .Y(_13860_));
 AO21x1_ASAP7_75t_R _31176_ (.A1(_13331_),
    .A2(_00592_),
    .B(_13860_),
    .Y(_13861_));
 AND2x2_ASAP7_75t_R _31177_ (.A(_13356_),
    .B(_00590_),
    .Y(_13862_));
 AO21x1_ASAP7_75t_R _31178_ (.A1(_13331_),
    .A2(_00594_),
    .B(_13862_),
    .Y(_13863_));
 OR2x2_ASAP7_75t_R _31179_ (.A(_13363_),
    .B(_13304_),
    .Y(_13864_));
 OAI22x1_ASAP7_75t_R _31180_ (.A1(_13859_),
    .A2(_13861_),
    .B1(_13863_),
    .B2(_13864_),
    .Y(_13865_));
 AND2x2_ASAP7_75t_R _31181_ (.A(_13326_),
    .B(_13304_),
    .Y(_13866_));
 INVx1_ASAP7_75t_R _31182_ (.A(_00578_),
    .Y(_13867_));
 NAND2x1_ASAP7_75t_R _31183_ (.A(_13356_),
    .B(_00574_),
    .Y(_13868_));
 OA21x2_ASAP7_75t_R _31184_ (.A1(_13842_),
    .A2(_13867_),
    .B(_13868_),
    .Y(_13869_));
 INVx1_ASAP7_75t_R _31185_ (.A(_00576_),
    .Y(_13870_));
 NAND2x1_ASAP7_75t_R _31186_ (.A(_13356_),
    .B(_00572_),
    .Y(_13871_));
 OA21x2_ASAP7_75t_R _31187_ (.A1(_13842_),
    .A2(_13870_),
    .B(_13871_),
    .Y(_13872_));
 AO22x2_ASAP7_75t_R _31188_ (.A1(_13866_),
    .A2(_13869_),
    .B1(_13872_),
    .B2(_13801_),
    .Y(_13873_));
 OR3x1_ASAP7_75t_R _31189_ (.A(_13858_),
    .B(_13865_),
    .C(_13873_),
    .Y(_13874_));
 INVx2_ASAP7_75t_R _31190_ (.A(_00566_),
    .Y(_13875_));
 NAND2x1_ASAP7_75t_R _31191_ (.A(_13391_),
    .B(_01790_),
    .Y(_13876_));
 OA211x2_ASAP7_75t_R _31192_ (.A1(_13347_),
    .A2(_13875_),
    .B(_13876_),
    .C(_13344_),
    .Y(_13877_));
 INVx2_ASAP7_75t_R _31193_ (.A(_00565_),
    .Y(_13878_));
 AND3x1_ASAP7_75t_R _31194_ (.A(_13393_),
    .B(_13326_),
    .C(_13878_),
    .Y(_13879_));
 OA21x2_ASAP7_75t_R _31195_ (.A1(_13877_),
    .A2(_13879_),
    .B(_13388_),
    .Y(_13880_));
 INVx2_ASAP7_75t_R _31196_ (.A(_00581_),
    .Y(_13881_));
 NAND2x1_ASAP7_75t_R _31197_ (.A(_13391_),
    .B(_00579_),
    .Y(_13882_));
 OA211x2_ASAP7_75t_R _31198_ (.A1(_13347_),
    .A2(_13881_),
    .B(_13882_),
    .C(_13393_),
    .Y(_13883_));
 INVx2_ASAP7_75t_R _31199_ (.A(_00582_),
    .Y(_13884_));
 NAND2x1_ASAP7_75t_R _31200_ (.A(_13391_),
    .B(_00580_),
    .Y(_13885_));
 OA211x2_ASAP7_75t_R _31201_ (.A1(_13481_),
    .A2(_13884_),
    .B(_13885_),
    .C(_13344_),
    .Y(_13886_));
 OA21x2_ASAP7_75t_R _31202_ (.A1(_13883_),
    .A2(_13886_),
    .B(_13461_),
    .Y(_13887_));
 OR3x1_ASAP7_75t_R _31203_ (.A(_13389_),
    .B(_13880_),
    .C(_13887_),
    .Y(_13888_));
 NOR2x1_ASAP7_75t_R _31204_ (.A(_13352_),
    .B(_13304_),
    .Y(_13889_));
 NAND2x1_ASAP7_75t_R _31205_ (.A(_13479_),
    .B(_00584_),
    .Y(_13890_));
 NAND2x1_ASAP7_75t_R _31206_ (.A(_13313_),
    .B(_00586_),
    .Y(_13891_));
 INVx1_ASAP7_75t_R _31207_ (.A(_00585_),
    .Y(_13892_));
 NAND2x1_ASAP7_75t_R _31208_ (.A(_13517_),
    .B(_00583_),
    .Y(_13893_));
 OA21x2_ASAP7_75t_R _31209_ (.A1(_13481_),
    .A2(_13892_),
    .B(_13893_),
    .Y(_13894_));
 AND2x4_ASAP7_75t_R _31210_ (.A(_13393_),
    .B(_13460_),
    .Y(_13895_));
 AO32x2_ASAP7_75t_R _31211_ (.A1(_13889_),
    .A2(_13890_),
    .A3(_13891_),
    .B1(_13894_),
    .B2(_13895_),
    .Y(_13896_));
 INVx1_ASAP7_75t_R _31212_ (.A(_00570_),
    .Y(_13897_));
 NAND2x1_ASAP7_75t_R _31213_ (.A(_13338_),
    .B(_00568_),
    .Y(_13898_));
 OA21x2_ASAP7_75t_R _31214_ (.A1(_13402_),
    .A2(_13897_),
    .B(_13898_),
    .Y(_13899_));
 AND2x4_ASAP7_75t_R _31215_ (.A(_13345_),
    .B(_13304_),
    .Y(_13900_));
 INVx1_ASAP7_75t_R _31216_ (.A(_00569_),
    .Y(_13901_));
 NAND2x1_ASAP7_75t_R _31217_ (.A(_13517_),
    .B(_00567_),
    .Y(_13902_));
 AND2x2_ASAP7_75t_R _31218_ (.A(_13321_),
    .B(_13303_),
    .Y(_13903_));
 OA211x2_ASAP7_75t_R _31219_ (.A1(_13616_),
    .A2(_13901_),
    .B(_13902_),
    .C(_13903_),
    .Y(_13904_));
 AO21x2_ASAP7_75t_R _31220_ (.A1(_13899_),
    .A2(_13900_),
    .B(_13904_),
    .Y(_13905_));
 OR3x1_ASAP7_75t_R _31221_ (.A(_13513_),
    .B(_13896_),
    .C(_13905_),
    .Y(_13906_));
 AND4x1_ASAP7_75t_R _31222_ (.A(_13857_),
    .B(_13874_),
    .C(_13888_),
    .D(_13906_),
    .Y(_13907_));
 BUFx12f_ASAP7_75t_R _31223_ (.A(_13907_),
    .Y(_13908_));
 AOI22x1_ASAP7_75t_R _31224_ (.A1(_13838_),
    .A2(_13839_),
    .B1(_13908_),
    .B2(_13302_),
    .Y(_18585_));
 INVx4_ASAP7_75t_R _31225_ (.A(_18585_),
    .Y(_18583_));
 BUFx6f_ASAP7_75t_R _31226_ (.A(_01514_),
    .Y(_13909_));
 INVx2_ASAP7_75t_R _31227_ (.A(_13909_),
    .Y(_13910_));
 INVx2_ASAP7_75t_R _31228_ (.A(_00607_),
    .Y(_13911_));
 NAND2x1_ASAP7_75t_R _31229_ (.A(_13675_),
    .B(_00603_),
    .Y(_13912_));
 OA211x2_ASAP7_75t_R _31230_ (.A1(_13496_),
    .A2(_13911_),
    .B(_13912_),
    .C(_13327_),
    .Y(_13913_));
 INVx1_ASAP7_75t_R _31231_ (.A(_00605_),
    .Y(_13914_));
 NAND2x1_ASAP7_75t_R _31232_ (.A(_13675_),
    .B(_00601_),
    .Y(_13915_));
 OA211x2_ASAP7_75t_R _31233_ (.A1(_13712_),
    .A2(_13914_),
    .B(_13915_),
    .C(_13773_),
    .Y(_13916_));
 NOR2x1_ASAP7_75t_R _31234_ (.A(_13913_),
    .B(_13916_),
    .Y(_13917_));
 INVx1_ASAP7_75t_R _31235_ (.A(_00623_),
    .Y(_13918_));
 NAND2x1_ASAP7_75t_R _31236_ (.A(_13487_),
    .B(_00619_),
    .Y(_13919_));
 OA211x2_ASAP7_75t_R _31237_ (.A1(_13712_),
    .A2(_13918_),
    .B(_13919_),
    .C(_13314_),
    .Y(_13920_));
 INVx1_ASAP7_75t_R _31238_ (.A(_00621_),
    .Y(_13921_));
 NAND2x1_ASAP7_75t_R _31239_ (.A(_13487_),
    .B(_00617_),
    .Y(_13922_));
 OA211x2_ASAP7_75t_R _31240_ (.A1(_13712_),
    .A2(_13921_),
    .B(_13922_),
    .C(_13734_),
    .Y(_13923_));
 NOR2x1_ASAP7_75t_R _31241_ (.A(_13920_),
    .B(_13923_),
    .Y(_13924_));
 AOI22x1_ASAP7_75t_R _31242_ (.A1(_13840_),
    .A2(_13917_),
    .B1(_13924_),
    .B2(_13856_),
    .Y(_13925_));
 NAND2x1_ASAP7_75t_R _31243_ (.A(_13651_),
    .B(_00618_),
    .Y(_13926_));
 NAND2x1_ASAP7_75t_R _31244_ (.A(_13331_),
    .B(_00622_),
    .Y(_13927_));
 INVx1_ASAP7_75t_R _31245_ (.A(_00624_),
    .Y(_13928_));
 NAND2x1_ASAP7_75t_R _31246_ (.A(_13354_),
    .B(_00620_),
    .Y(_13929_));
 OA21x2_ASAP7_75t_R _31247_ (.A1(_13711_),
    .A2(_13928_),
    .B(_13929_),
    .Y(_13930_));
 AO32x2_ASAP7_75t_R _31248_ (.A1(_13797_),
    .A2(_13926_),
    .A3(_13927_),
    .B1(_13930_),
    .B2(_13805_),
    .Y(_13931_));
 AND2x2_ASAP7_75t_R _31249_ (.A(_13334_),
    .B(_00604_),
    .Y(_13932_));
 AO21x1_ASAP7_75t_R _31250_ (.A1(_13332_),
    .A2(_00608_),
    .B(_13932_),
    .Y(_13933_));
 AND2x2_ASAP7_75t_R _31251_ (.A(_13334_),
    .B(_00602_),
    .Y(_13934_));
 AO21x1_ASAP7_75t_R _31252_ (.A1(_13332_),
    .A2(_00606_),
    .B(_13934_),
    .Y(_13935_));
 BUFx6f_ASAP7_75t_R _31253_ (.A(_13378_),
    .Y(_13936_));
 NAND2x1_ASAP7_75t_R _31254_ (.A(_13936_),
    .B(_13305_),
    .Y(_13937_));
 OAI22x1_ASAP7_75t_R _31255_ (.A1(_13809_),
    .A2(_13933_),
    .B1(_13935_),
    .B2(_13937_),
    .Y(_13938_));
 OR3x1_ASAP7_75t_R _31256_ (.A(_13858_),
    .B(_13931_),
    .C(_13938_),
    .Y(_13939_));
 AND2x2_ASAP7_75t_R _31257_ (.A(_13479_),
    .B(_01789_),
    .Y(_13940_));
 AO211x2_ASAP7_75t_R _31258_ (.A1(_13327_),
    .A2(_00596_),
    .B(_13940_),
    .C(_13673_),
    .Y(_13941_));
 OR3x1_ASAP7_75t_R _31259_ (.A(_13346_),
    .B(_13753_),
    .C(_00595_),
    .Y(_13942_));
 AO21x2_ASAP7_75t_R _31260_ (.A1(_13941_),
    .A2(_13942_),
    .B(_13764_),
    .Y(_13943_));
 INVx1_ASAP7_75t_R _31261_ (.A(_00611_),
    .Y(_13944_));
 NAND2x1_ASAP7_75t_R _31262_ (.A(_13339_),
    .B(_00609_),
    .Y(_13945_));
 OA211x2_ASAP7_75t_R _31263_ (.A1(_13773_),
    .A2(_13944_),
    .B(_13945_),
    .C(_13673_),
    .Y(_13946_));
 INVx2_ASAP7_75t_R _31264_ (.A(_00612_),
    .Y(_13947_));
 NAND2x1_ASAP7_75t_R _31265_ (.A(_13748_),
    .B(_00610_),
    .Y(_13948_));
 OA211x2_ASAP7_75t_R _31266_ (.A1(_13746_),
    .A2(_13947_),
    .B(_13948_),
    .C(_13750_),
    .Y(_13949_));
 OAI21x1_ASAP7_75t_R _31267_ (.A1(_13946_),
    .A2(_13949_),
    .B(_13764_),
    .Y(_13950_));
 NAND3x1_ASAP7_75t_R _31268_ (.A(_13310_),
    .B(_13943_),
    .C(_13950_),
    .Y(_13951_));
 INVx1_ASAP7_75t_R _31269_ (.A(_00599_),
    .Y(_13952_));
 NAND2x1_ASAP7_75t_R _31270_ (.A(_13725_),
    .B(_00597_),
    .Y(_13953_));
 OA21x2_ASAP7_75t_R _31271_ (.A1(_13936_),
    .A2(_13952_),
    .B(_13953_),
    .Y(_13954_));
 INVx2_ASAP7_75t_R _31272_ (.A(_00615_),
    .Y(_13955_));
 NAND2x1_ASAP7_75t_R _31273_ (.A(_13701_),
    .B(_00613_),
    .Y(_13956_));
 OA211x2_ASAP7_75t_R _31274_ (.A1(_13734_),
    .A2(_13955_),
    .B(_13956_),
    .C(_13461_),
    .Y(_13957_));
 AOI211x1_ASAP7_75t_R _31275_ (.A1(_13306_),
    .A2(_13954_),
    .B(_13957_),
    .C(_13434_),
    .Y(_13958_));
 INVx1_ASAP7_75t_R _31276_ (.A(_00600_),
    .Y(_13959_));
 NAND2x1_ASAP7_75t_R _31277_ (.A(_13725_),
    .B(_00598_),
    .Y(_13960_));
 OA21x2_ASAP7_75t_R _31278_ (.A1(_13936_),
    .A2(_13959_),
    .B(_13960_),
    .Y(_13961_));
 INVx2_ASAP7_75t_R _31279_ (.A(_00616_),
    .Y(_13962_));
 NAND2x1_ASAP7_75t_R _31280_ (.A(_13701_),
    .B(_00614_),
    .Y(_13963_));
 OA211x2_ASAP7_75t_R _31281_ (.A1(_13734_),
    .A2(_13962_),
    .B(_13963_),
    .C(_13461_),
    .Y(_13964_));
 AOI211x1_ASAP7_75t_R _31282_ (.A1(_13306_),
    .A2(_13961_),
    .B(_13964_),
    .C(_13323_),
    .Y(_13965_));
 OAI21x1_ASAP7_75t_R _31283_ (.A1(_13958_),
    .A2(_13965_),
    .B(_13694_),
    .Y(_13966_));
 AND4x1_ASAP7_75t_R _31284_ (.A(_13925_),
    .B(_13939_),
    .C(_13951_),
    .D(_13966_),
    .Y(_13967_));
 BUFx12f_ASAP7_75t_R _31285_ (.A(_13967_),
    .Y(_13968_));
 BUFx12f_ASAP7_75t_R _31286_ (.A(_13302_),
    .Y(_13969_));
 AOI22x1_ASAP7_75t_R _31287_ (.A1(_13910_),
    .A2(_13839_),
    .B1(_13968_),
    .B2(_13969_),
    .Y(_18590_));
 INVx2_ASAP7_75t_R _31288_ (.A(_18590_),
    .Y(_18588_));
 INVx2_ASAP7_75t_R _31289_ (.A(_01513_),
    .Y(_13970_));
 INVx2_ASAP7_75t_R _31290_ (.A(_00650_),
    .Y(_13971_));
 NAND2x1_ASAP7_75t_R _31291_ (.A(_13738_),
    .B(_00648_),
    .Y(_13972_));
 OA21x2_ASAP7_75t_R _31292_ (.A1(_13340_),
    .A2(_13971_),
    .B(_13972_),
    .Y(_13973_));
 INVx1_ASAP7_75t_R _31293_ (.A(_00651_),
    .Y(_13974_));
 NOR2x1_ASAP7_75t_R _31294_ (.A(_13340_),
    .B(_00653_),
    .Y(_13975_));
 AO21x1_ASAP7_75t_R _31295_ (.A1(_13813_),
    .A2(_13974_),
    .B(_13975_),
    .Y(_13976_));
 INVx2_ASAP7_75t_R _31296_ (.A(_00649_),
    .Y(_13977_));
 NAND2x1_ASAP7_75t_R _31297_ (.A(_13734_),
    .B(_00647_),
    .Y(_13978_));
 OA211x2_ASAP7_75t_R _31298_ (.A1(_13340_),
    .A2(_13977_),
    .B(_13646_),
    .C(_13978_),
    .Y(_13979_));
 AOI221x1_ASAP7_75t_R _31299_ (.A1(_13641_),
    .A2(_13973_),
    .B1(_13976_),
    .B2(_13632_),
    .C(_13979_),
    .Y(_13980_));
 INVx1_ASAP7_75t_R _31300_ (.A(_00654_),
    .Y(_13981_));
 NAND2x1_ASAP7_75t_R _31301_ (.A(_13936_),
    .B(_00652_),
    .Y(_13982_));
 OA211x2_ASAP7_75t_R _31302_ (.A1(_13813_),
    .A2(_13981_),
    .B(_13637_),
    .C(_13982_),
    .Y(_13983_));
 NOR2x1_ASAP7_75t_R _31303_ (.A(_13365_),
    .B(_13983_),
    .Y(_13984_));
 INVx2_ASAP7_75t_R _31304_ (.A(_00642_),
    .Y(_13985_));
 NAND2x1_ASAP7_75t_R _31305_ (.A(_13936_),
    .B(_00640_),
    .Y(_13986_));
 OA211x2_ASAP7_75t_R _31306_ (.A1(_13340_),
    .A2(_13985_),
    .B(_13986_),
    .C(_13434_),
    .Y(_13987_));
 INVx1_ASAP7_75t_R _31307_ (.A(_00641_),
    .Y(_13988_));
 NAND2x1_ASAP7_75t_R _31308_ (.A(_13738_),
    .B(_00639_),
    .Y(_13989_));
 OA211x2_ASAP7_75t_R _31309_ (.A1(_13813_),
    .A2(_13988_),
    .B(_13989_),
    .C(_13323_),
    .Y(_13990_));
 NOR2x1_ASAP7_75t_R _31310_ (.A(_13987_),
    .B(_13990_),
    .Y(_13991_));
 AND2x2_ASAP7_75t_R _31311_ (.A(_13753_),
    .B(_01788_),
    .Y(_13992_));
 AO21x1_ASAP7_75t_R _31312_ (.A1(_13328_),
    .A2(_00626_),
    .B(_13992_),
    .Y(_13993_));
 OA221x2_ASAP7_75t_R _31313_ (.A1(_00625_),
    .A2(_13670_),
    .B1(_13993_),
    .B2(_13323_),
    .C(_13484_),
    .Y(_13994_));
 AOI221x1_ASAP7_75t_R _31314_ (.A1(_13980_),
    .A2(_13984_),
    .B1(_13991_),
    .B2(_13666_),
    .C(_13994_),
    .Y(_13995_));
 INVx1_ASAP7_75t_R _31315_ (.A(_00638_),
    .Y(_13996_));
 NAND2x1_ASAP7_75t_R _31316_ (.A(_13675_),
    .B(_00634_),
    .Y(_13997_));
 OA211x2_ASAP7_75t_R _31317_ (.A1(_13496_),
    .A2(_13996_),
    .B(_13997_),
    .C(_13314_),
    .Y(_13998_));
 INVx1_ASAP7_75t_R _31318_ (.A(_00636_),
    .Y(_13999_));
 NAND2x1_ASAP7_75t_R _31319_ (.A(_13675_),
    .B(_00632_),
    .Y(_14000_));
 OA211x2_ASAP7_75t_R _31320_ (.A1(_13496_),
    .A2(_13999_),
    .B(_14000_),
    .C(_13773_),
    .Y(_14001_));
 OR3x1_ASAP7_75t_R _31321_ (.A(_13417_),
    .B(_13998_),
    .C(_14001_),
    .Y(_14002_));
 INVx1_ASAP7_75t_R _31322_ (.A(_00637_),
    .Y(_14003_));
 NAND2x1_ASAP7_75t_R _31323_ (.A(_13675_),
    .B(_00633_),
    .Y(_14004_));
 OA211x2_ASAP7_75t_R _31324_ (.A1(_13496_),
    .A2(_14003_),
    .B(_14004_),
    .C(_13327_),
    .Y(_14005_));
 INVx1_ASAP7_75t_R _31325_ (.A(_00635_),
    .Y(_14006_));
 NAND2x1_ASAP7_75t_R _31326_ (.A(_13675_),
    .B(_00631_),
    .Y(_14007_));
 OA211x2_ASAP7_75t_R _31327_ (.A1(_13496_),
    .A2(_14006_),
    .B(_14007_),
    .C(_13773_),
    .Y(_14008_));
 OR3x1_ASAP7_75t_R _31328_ (.A(_13544_),
    .B(_14005_),
    .C(_14008_),
    .Y(_14009_));
 INVx2_ASAP7_75t_R _31329_ (.A(_00629_),
    .Y(_14010_));
 NAND2x1_ASAP7_75t_R _31330_ (.A(_13695_),
    .B(_00627_),
    .Y(_14011_));
 OA211x2_ASAP7_75t_R _31331_ (.A1(_13746_),
    .A2(_14010_),
    .B(_14011_),
    .C(_13673_),
    .Y(_14012_));
 INVx2_ASAP7_75t_R _31332_ (.A(_00630_),
    .Y(_14013_));
 NAND2x1_ASAP7_75t_R _31333_ (.A(_13695_),
    .B(_00628_),
    .Y(_14014_));
 OA211x2_ASAP7_75t_R _31334_ (.A1(_13746_),
    .A2(_14013_),
    .B(_14014_),
    .C(_13750_),
    .Y(_14015_));
 OR3x1_ASAP7_75t_R _31335_ (.A(_13375_),
    .B(_14012_),
    .C(_14015_),
    .Y(_14016_));
 INVx2_ASAP7_75t_R _31336_ (.A(_00646_),
    .Y(_14017_));
 NAND2x1_ASAP7_75t_R _31337_ (.A(_13748_),
    .B(_00644_),
    .Y(_14018_));
 OA211x2_ASAP7_75t_R _31338_ (.A1(_13746_),
    .A2(_14017_),
    .B(_14018_),
    .C(_13750_),
    .Y(_14019_));
 INVx2_ASAP7_75t_R _31339_ (.A(_00645_),
    .Y(_14020_));
 NAND2x1_ASAP7_75t_R _31340_ (.A(_13748_),
    .B(_00643_),
    .Y(_14021_));
 OA211x2_ASAP7_75t_R _31341_ (.A1(_13746_),
    .A2(_14020_),
    .B(_14021_),
    .C(_13673_),
    .Y(_14022_));
 OR3x1_ASAP7_75t_R _31342_ (.A(_13386_),
    .B(_14019_),
    .C(_14022_),
    .Y(_14023_));
 AND4x1_ASAP7_75t_R _31343_ (.A(_14002_),
    .B(_14009_),
    .C(_14016_),
    .D(_14023_),
    .Y(_14024_));
 AND3x4_ASAP7_75t_R _31344_ (.A(_13302_),
    .B(_13995_),
    .C(_14024_),
    .Y(_14025_));
 AO21x1_ASAP7_75t_R _31345_ (.A1(_13970_),
    .A2(_13839_),
    .B(_14025_),
    .Y(_14026_));
 BUFx3_ASAP7_75t_R _31346_ (.A(_14026_),
    .Y(_18593_));
 INVx1_ASAP7_75t_R _31347_ (.A(_18593_),
    .Y(_18595_));
 INVx2_ASAP7_75t_R _31348_ (.A(_01512_),
    .Y(_14027_));
 AND2x4_ASAP7_75t_R _31349_ (.A(_13332_),
    .B(_13374_),
    .Y(_14028_));
 INVx2_ASAP7_75t_R _31350_ (.A(_00660_),
    .Y(_14029_));
 NAND2x1_ASAP7_75t_R _31351_ (.A(_13518_),
    .B(_00658_),
    .Y(_14030_));
 OA21x2_ASAP7_75t_R _31352_ (.A1(_13701_),
    .A2(_14029_),
    .B(_14030_),
    .Y(_14031_));
 INVx2_ASAP7_75t_R _31353_ (.A(_00659_),
    .Y(_14032_));
 NAND2x1_ASAP7_75t_R _31354_ (.A(_13363_),
    .B(_00657_),
    .Y(_14033_));
 OA211x2_ASAP7_75t_R _31355_ (.A1(_13748_),
    .A2(_14032_),
    .B(_14033_),
    .C(_13352_),
    .Y(_14034_));
 AO21x1_ASAP7_75t_R _31356_ (.A1(_13750_),
    .A2(_14031_),
    .B(_14034_),
    .Y(_14035_));
 INVx2_ASAP7_75t_R _31357_ (.A(_00676_),
    .Y(_14036_));
 NAND2x1_ASAP7_75t_R _31358_ (.A(_13317_),
    .B(_00674_),
    .Y(_14037_));
 OA21x2_ASAP7_75t_R _31359_ (.A1(_13701_),
    .A2(_14036_),
    .B(_14037_),
    .Y(_14038_));
 INVx2_ASAP7_75t_R _31360_ (.A(_00675_),
    .Y(_14039_));
 NAND2x1_ASAP7_75t_R _31361_ (.A(_13479_),
    .B(_00673_),
    .Y(_14040_));
 OA211x2_ASAP7_75t_R _31362_ (.A1(_13695_),
    .A2(_14039_),
    .B(_14040_),
    .C(_13352_),
    .Y(_14041_));
 AO21x2_ASAP7_75t_R _31363_ (.A1(_13434_),
    .A2(_14038_),
    .B(_14041_),
    .Y(_14042_));
 INVx1_ASAP7_75t_R _31364_ (.A(_13386_),
    .Y(_14043_));
 AO22x1_ASAP7_75t_R _31365_ (.A1(_14028_),
    .A2(_14035_),
    .B1(_14042_),
    .B2(_14043_),
    .Y(_14044_));
 AND2x2_ASAP7_75t_R _31366_ (.A(_13363_),
    .B(_01787_),
    .Y(_14045_));
 AO21x1_ASAP7_75t_R _31367_ (.A1(_13327_),
    .A2(_00656_),
    .B(_14045_),
    .Y(_14046_));
 OR3x1_ASAP7_75t_R _31368_ (.A(_13369_),
    .B(_13748_),
    .C(_00655_),
    .Y(_14047_));
 OA211x2_ASAP7_75t_R _31369_ (.A1(_13353_),
    .A2(_14046_),
    .B(_14047_),
    .C(_13305_),
    .Y(_14048_));
 INVx1_ASAP7_75t_R _31370_ (.A(_00669_),
    .Y(_14049_));
 NOR2x1_ASAP7_75t_R _31371_ (.A(_13748_),
    .B(_00671_),
    .Y(_14050_));
 AO21x1_ASAP7_75t_R _31372_ (.A1(_13753_),
    .A2(_14049_),
    .B(_14050_),
    .Y(_14051_));
 INVx2_ASAP7_75t_R _31373_ (.A(_00672_),
    .Y(_14052_));
 NAND2x1_ASAP7_75t_R _31374_ (.A(_13518_),
    .B(_00670_),
    .Y(_14053_));
 OA211x2_ASAP7_75t_R _31375_ (.A1(_13725_),
    .A2(_14052_),
    .B(_14053_),
    .C(_13346_),
    .Y(_14054_));
 AOI211x1_ASAP7_75t_R _31376_ (.A1(_13323_),
    .A2(_14051_),
    .B(_14054_),
    .C(_13305_),
    .Y(_14055_));
 NOR3x1_ASAP7_75t_R _31377_ (.A(_13389_),
    .B(_14048_),
    .C(_14055_),
    .Y(_14056_));
 INVx1_ASAP7_75t_R _31378_ (.A(_00661_),
    .Y(_14057_));
 NOR2x1_ASAP7_75t_R _31379_ (.A(_13334_),
    .B(_00665_),
    .Y(_14058_));
 AO21x1_ASAP7_75t_R _31380_ (.A1(_13487_),
    .A2(_14057_),
    .B(_14058_),
    .Y(_14059_));
 INVx2_ASAP7_75t_R _31381_ (.A(_00667_),
    .Y(_14060_));
 NAND2x1_ASAP7_75t_R _31382_ (.A(_13842_),
    .B(_00663_),
    .Y(_14061_));
 OA211x2_ASAP7_75t_R _31383_ (.A1(_13711_),
    .A2(_14060_),
    .B(_14061_),
    .C(_13313_),
    .Y(_14062_));
 AO21x2_ASAP7_75t_R _31384_ (.A1(_13738_),
    .A2(_14059_),
    .B(_14062_),
    .Y(_14063_));
 INVx2_ASAP7_75t_R _31385_ (.A(_00677_),
    .Y(_14064_));
 NOR2x1_ASAP7_75t_R _31386_ (.A(_13334_),
    .B(_00681_),
    .Y(_14065_));
 AO21x1_ASAP7_75t_R _31387_ (.A1(_13487_),
    .A2(_14064_),
    .B(_14065_),
    .Y(_14066_));
 INVx1_ASAP7_75t_R _31388_ (.A(_00683_),
    .Y(_14067_));
 NAND2x1_ASAP7_75t_R _31389_ (.A(_13842_),
    .B(_00679_),
    .Y(_14068_));
 OA211x2_ASAP7_75t_R _31390_ (.A1(_13711_),
    .A2(_14067_),
    .B(_14068_),
    .C(_13313_),
    .Y(_14069_));
 AO21x2_ASAP7_75t_R _31391_ (.A1(_13738_),
    .A2(_14066_),
    .B(_14069_),
    .Y(_14070_));
 AO22x1_ASAP7_75t_R _31392_ (.A1(_13840_),
    .A2(_14063_),
    .B1(_14070_),
    .B2(_13856_),
    .Y(_14071_));
 INVx2_ASAP7_75t_R _31393_ (.A(_00682_),
    .Y(_14072_));
 NAND2x1_ASAP7_75t_R _31394_ (.A(_13304_),
    .B(_00666_),
    .Y(_14073_));
 OA211x2_ASAP7_75t_R _31395_ (.A1(_13388_),
    .A2(_14072_),
    .B(_14073_),
    .C(_13331_),
    .Y(_14074_));
 INVx2_ASAP7_75t_R _31396_ (.A(_00678_),
    .Y(_14075_));
 NAND2x1_ASAP7_75t_R _31397_ (.A(_13304_),
    .B(_00662_),
    .Y(_14076_));
 OA211x2_ASAP7_75t_R _31398_ (.A1(_13388_),
    .A2(_14075_),
    .B(_14076_),
    .C(_13651_),
    .Y(_14077_));
 NOR2x1_ASAP7_75t_R _31399_ (.A(_14074_),
    .B(_14077_),
    .Y(_14078_));
 INVx2_ASAP7_75t_R _31400_ (.A(_00684_),
    .Y(_14079_));
 NAND2x1_ASAP7_75t_R _31401_ (.A(_13304_),
    .B(_00668_),
    .Y(_14080_));
 OA211x2_ASAP7_75t_R _31402_ (.A1(_13388_),
    .A2(_14079_),
    .B(_14080_),
    .C(_13332_),
    .Y(_14081_));
 INVx2_ASAP7_75t_R _31403_ (.A(_00680_),
    .Y(_14082_));
 NAND2x1_ASAP7_75t_R _31404_ (.A(_13388_),
    .B(_00664_),
    .Y(_14083_));
 OA211x2_ASAP7_75t_R _31405_ (.A1(_13388_),
    .A2(_14082_),
    .B(_14083_),
    .C(_13651_),
    .Y(_14084_));
 NOR2x1_ASAP7_75t_R _31406_ (.A(_14081_),
    .B(_14084_),
    .Y(_14085_));
 OR3x1_ASAP7_75t_R _31407_ (.A(_13353_),
    .B(_13340_),
    .C(_13459_),
    .Y(_14086_));
 OAI22x1_ASAP7_75t_R _31408_ (.A1(_13716_),
    .A2(_14078_),
    .B1(_14085_),
    .B2(_14086_),
    .Y(_14087_));
 OR4x1_ASAP7_75t_R _31409_ (.A(_14044_),
    .B(_14056_),
    .C(_14071_),
    .D(_14087_),
    .Y(_14088_));
 BUFx12f_ASAP7_75t_R _31410_ (.A(_14088_),
    .Y(_14089_));
 BUFx12f_ASAP7_75t_R _31411_ (.A(_13969_),
    .Y(_14090_));
 AOI22x1_ASAP7_75t_R _31412_ (.A1(_14027_),
    .A2(_13839_),
    .B1(_14089_),
    .B2(_14090_),
    .Y(_18600_));
 INVx1_ASAP7_75t_R _31413_ (.A(_18600_),
    .Y(_18598_));
 AND2x4_ASAP7_75t_R _31414_ (.A(_00344_),
    .B(_00341_),
    .Y(_14091_));
 AND3x4_ASAP7_75t_R _31415_ (.A(_13123_),
    .B(_13163_),
    .C(_14091_),
    .Y(_14092_));
 AND2x4_ASAP7_75t_R _31416_ (.A(_13094_),
    .B(_14092_),
    .Y(_14093_));
 AND2x6_ASAP7_75t_R _31417_ (.A(_13685_),
    .B(_13602_),
    .Y(_14094_));
 AND4x1_ASAP7_75t_R _31418_ (.A(_13287_),
    .B(_00339_),
    .C(_13455_),
    .D(_01506_),
    .Y(_14095_));
 AND3x1_ASAP7_75t_R _31419_ (.A(_14093_),
    .B(_14094_),
    .C(_14095_),
    .Y(_14096_));
 AND3x4_ASAP7_75t_R _31420_ (.A(_13837_),
    .B(_13909_),
    .C(_13831_),
    .Y(_14097_));
 BUFx12f_ASAP7_75t_R _31421_ (.A(_14097_),
    .Y(_14098_));
 BUFx12f_ASAP7_75t_R _31422_ (.A(_00412_),
    .Y(_14099_));
 AND3x1_ASAP7_75t_R _31423_ (.A(_14099_),
    .B(_01512_),
    .C(_01513_),
    .Y(_14100_));
 BUFx6f_ASAP7_75t_R _31424_ (.A(_14100_),
    .Y(_14101_));
 AND5x2_ASAP7_75t_R _31425_ (.A(_13378_),
    .B(_13354_),
    .C(_13459_),
    .D(_13304_),
    .E(_01510_),
    .Y(_14102_));
 AND3x4_ASAP7_75t_R _31426_ (.A(_14098_),
    .B(_14101_),
    .C(_14102_),
    .Y(_14103_));
 NOR2x1_ASAP7_75t_R _31427_ (.A(_01510_),
    .B(_13831_),
    .Y(_14104_));
 AND5x2_ASAP7_75t_R _31428_ (.A(_13460_),
    .B(_14099_),
    .C(_13837_),
    .D(_13910_),
    .E(_14104_),
    .Y(_14105_));
 AND4x1_ASAP7_75t_R _31429_ (.A(_13303_),
    .B(_14099_),
    .C(_01510_),
    .D(_14098_),
    .Y(_14106_));
 NOR2x2_ASAP7_75t_R _31430_ (.A(_01512_),
    .B(_01513_),
    .Y(_14107_));
 AND4x1_ASAP7_75t_R _31431_ (.A(_13322_),
    .B(_13327_),
    .C(_13310_),
    .D(_14107_),
    .Y(_14108_));
 OA21x2_ASAP7_75t_R _31432_ (.A1(_14105_),
    .A2(_14106_),
    .B(_14108_),
    .Y(_14109_));
 AND5x2_ASAP7_75t_R _31433_ (.A(_01512_),
    .B(_13970_),
    .C(_13694_),
    .D(_13467_),
    .E(_14106_),
    .Y(_14110_));
 OR3x1_ASAP7_75t_R _31434_ (.A(_14103_),
    .B(_14109_),
    .C(_14110_),
    .Y(_14111_));
 BUFx6f_ASAP7_75t_R _31435_ (.A(_13227_),
    .Y(_14112_));
 AND3x1_ASAP7_75t_R _31436_ (.A(_14112_),
    .B(_13421_),
    .C(_13265_),
    .Y(_14113_));
 INVx1_ASAP7_75t_R _31437_ (.A(_14113_),
    .Y(_14114_));
 AO21x2_ASAP7_75t_R _31438_ (.A1(_14096_),
    .A2(_14111_),
    .B(_14114_),
    .Y(_14115_));
 INVx1_ASAP7_75t_R _31439_ (.A(_13421_),
    .Y(_14116_));
 BUFx6f_ASAP7_75t_R _31440_ (.A(_14116_),
    .Y(_14117_));
 OR2x6_ASAP7_75t_R _31441_ (.A(_14117_),
    .B(_13422_),
    .Y(_14118_));
 BUFx12f_ASAP7_75t_R _31442_ (.A(_14118_),
    .Y(_14119_));
 AND2x6_ASAP7_75t_R _31443_ (.A(_14119_),
    .B(_13265_),
    .Y(_14120_));
 INVx4_ASAP7_75t_R _31444_ (.A(_13227_),
    .Y(_14121_));
 BUFx6f_ASAP7_75t_R _31445_ (.A(_01510_),
    .Y(_14122_));
 OA211x2_ASAP7_75t_R _31446_ (.A1(_13261_),
    .A2(_14122_),
    .B(_14098_),
    .C(_14101_),
    .Y(_14123_));
 INVx2_ASAP7_75t_R _31447_ (.A(_13217_),
    .Y(_14124_));
 OR5x2_ASAP7_75t_R _31448_ (.A(_13280_),
    .B(_13230_),
    .C(_14124_),
    .D(_13285_),
    .E(_13225_),
    .Y(_14125_));
 OR4x1_ASAP7_75t_R _31449_ (.A(_14121_),
    .B(_13421_),
    .C(_14123_),
    .D(_14125_),
    .Y(_14126_));
 AOI21x1_ASAP7_75t_R _31450_ (.A1(_13276_),
    .A2(_13278_),
    .B(_13242_),
    .Y(_14127_));
 AND2x2_ASAP7_75t_R _31451_ (.A(_13246_),
    .B(_13247_),
    .Y(_14128_));
 OA21x2_ASAP7_75t_R _31452_ (.A1(_14128_),
    .A2(_13282_),
    .B(_13277_),
    .Y(_14129_));
 AND3x1_ASAP7_75t_R _31453_ (.A(_01540_),
    .B(_13240_),
    .C(_13290_),
    .Y(_14130_));
 NAND2x1_ASAP7_75t_R _31454_ (.A(_13263_),
    .B(_13240_),
    .Y(_14131_));
 AO21x1_ASAP7_75t_R _31455_ (.A1(_13226_),
    .A2(_13421_),
    .B(_13217_),
    .Y(_14132_));
 OA21x2_ASAP7_75t_R _31456_ (.A1(_13261_),
    .A2(_13227_),
    .B(_14132_),
    .Y(_14133_));
 NAND2x1_ASAP7_75t_R _31457_ (.A(_13277_),
    .B(_13218_),
    .Y(_14134_));
 OR3x2_ASAP7_75t_R _31458_ (.A(_13276_),
    .B(_13285_),
    .C(_14134_),
    .Y(_14135_));
 AND2x2_ASAP7_75t_R _31459_ (.A(_13227_),
    .B(_13242_),
    .Y(_14136_));
 NOR2x1_ASAP7_75t_R _31460_ (.A(_13227_),
    .B(_13421_),
    .Y(_14137_));
 NOR2x1_ASAP7_75t_R _31461_ (.A(_13262_),
    .B(_14137_),
    .Y(_14138_));
 OA33x2_ASAP7_75t_R _31462_ (.A1(_13441_),
    .A2(_14131_),
    .A3(_14133_),
    .B1(_14135_),
    .B2(_14136_),
    .B3(_14138_),
    .Y(_14139_));
 OA211x2_ASAP7_75t_R _31463_ (.A1(_14127_),
    .A2(_14129_),
    .B(_14130_),
    .C(_14139_),
    .Y(_14140_));
 AND3x4_ASAP7_75t_R _31464_ (.A(_14120_),
    .B(_14126_),
    .C(_14140_),
    .Y(_14141_));
 NAND2x2_ASAP7_75t_R _31465_ (.A(_14115_),
    .B(_14141_),
    .Y(_14142_));
 BUFx6f_ASAP7_75t_R _31466_ (.A(_14142_),
    .Y(_14143_));
 BUFx6f_ASAP7_75t_R _31467_ (.A(_14143_),
    .Y(_14144_));
 NOR2x1_ASAP7_75t_R _31468_ (.A(_18600_),
    .B(_14144_),
    .Y(_18081_));
 INVx1_ASAP7_75t_R _31469_ (.A(_00710_),
    .Y(_14145_));
 NAND2x1_ASAP7_75t_R _31470_ (.A(_13701_),
    .B(_00708_),
    .Y(_14146_));
 OA211x2_ASAP7_75t_R _31471_ (.A1(_13936_),
    .A2(_14145_),
    .B(_14146_),
    .C(_13750_),
    .Y(_14147_));
 INVx1_ASAP7_75t_R _31472_ (.A(_00709_),
    .Y(_14148_));
 NAND2x1_ASAP7_75t_R _31473_ (.A(_13701_),
    .B(_00707_),
    .Y(_14149_));
 OA211x2_ASAP7_75t_R _31474_ (.A1(_13936_),
    .A2(_14148_),
    .B(_14149_),
    .C(_13353_),
    .Y(_14150_));
 OA21x2_ASAP7_75t_R _31475_ (.A1(_14147_),
    .A2(_14150_),
    .B(_13688_),
    .Y(_14151_));
 INVx2_ASAP7_75t_R _31476_ (.A(_00706_),
    .Y(_14152_));
 NAND2x1_ASAP7_75t_R _31477_ (.A(_13348_),
    .B(_00704_),
    .Y(_14153_));
 OA211x2_ASAP7_75t_R _31478_ (.A1(_13936_),
    .A2(_14152_),
    .B(_14153_),
    .C(_13750_),
    .Y(_14154_));
 INVx1_ASAP7_75t_R _31479_ (.A(_00705_),
    .Y(_14155_));
 NAND2x1_ASAP7_75t_R _31480_ (.A(_13701_),
    .B(_00703_),
    .Y(_14156_));
 OA211x2_ASAP7_75t_R _31481_ (.A1(_13936_),
    .A2(_14155_),
    .B(_14156_),
    .C(_13353_),
    .Y(_14157_));
 OA21x2_ASAP7_75t_R _31482_ (.A1(_14154_),
    .A2(_14157_),
    .B(_13694_),
    .Y(_14158_));
 AO21x2_ASAP7_75t_R _31483_ (.A1(_13814_),
    .A2(_14151_),
    .B(_14158_),
    .Y(_14159_));
 INVx1_ASAP7_75t_R _31484_ (.A(_00714_),
    .Y(_14160_));
 NAND2x1_ASAP7_75t_R _31485_ (.A(_13339_),
    .B(_00712_),
    .Y(_14161_));
 OA211x2_ASAP7_75t_R _31486_ (.A1(_13753_),
    .A2(_14160_),
    .B(_14161_),
    .C(_13346_),
    .Y(_14162_));
 INVx2_ASAP7_75t_R _31487_ (.A(_00713_),
    .Y(_14163_));
 NAND2x1_ASAP7_75t_R _31488_ (.A(_13339_),
    .B(_00711_),
    .Y(_14164_));
 OA211x2_ASAP7_75t_R _31489_ (.A1(_13753_),
    .A2(_14163_),
    .B(_14164_),
    .C(_13322_),
    .Y(_14165_));
 OA211x2_ASAP7_75t_R _31490_ (.A1(_14162_),
    .A2(_14165_),
    .B(_13669_),
    .C(_13407_),
    .Y(_14166_));
 INVx1_ASAP7_75t_R _31491_ (.A(_00697_),
    .Y(_14167_));
 NAND2x1_ASAP7_75t_R _31492_ (.A(_13675_),
    .B(_00693_),
    .Y(_14168_));
 OA211x2_ASAP7_75t_R _31493_ (.A1(_13496_),
    .A2(_14167_),
    .B(_14168_),
    .C(_13327_),
    .Y(_14169_));
 INVx1_ASAP7_75t_R _31494_ (.A(_00695_),
    .Y(_14170_));
 NAND2x1_ASAP7_75t_R _31495_ (.A(_13675_),
    .B(_00691_),
    .Y(_14171_));
 OA211x2_ASAP7_75t_R _31496_ (.A1(_13496_),
    .A2(_14170_),
    .B(_14171_),
    .C(_13753_),
    .Y(_14172_));
 OA21x2_ASAP7_75t_R _31497_ (.A1(_14169_),
    .A2(_14172_),
    .B(_13840_),
    .Y(_14173_));
 INVx2_ASAP7_75t_R _31498_ (.A(_00690_),
    .Y(_14174_));
 NAND2x1_ASAP7_75t_R _31499_ (.A(_13748_),
    .B(_00688_),
    .Y(_14175_));
 OA211x2_ASAP7_75t_R _31500_ (.A1(_13746_),
    .A2(_14174_),
    .B(_14175_),
    .C(_13346_),
    .Y(_14176_));
 INVx2_ASAP7_75t_R _31501_ (.A(_00689_),
    .Y(_14177_));
 NAND2x1_ASAP7_75t_R _31502_ (.A(_13748_),
    .B(_00687_),
    .Y(_14178_));
 OA211x2_ASAP7_75t_R _31503_ (.A1(_13773_),
    .A2(_14177_),
    .B(_14178_),
    .C(_13673_),
    .Y(_14179_));
 OA21x2_ASAP7_75t_R _31504_ (.A1(_14176_),
    .A2(_14179_),
    .B(_14028_),
    .Y(_14180_));
 INVx2_ASAP7_75t_R _31505_ (.A(_00698_),
    .Y(_14181_));
 NAND2x1_ASAP7_75t_R _31506_ (.A(_13711_),
    .B(_00694_),
    .Y(_14182_));
 OA211x2_ASAP7_75t_R _31507_ (.A1(_13651_),
    .A2(_14181_),
    .B(_14182_),
    .C(_13327_),
    .Y(_14183_));
 INVx1_ASAP7_75t_R _31508_ (.A(_00696_),
    .Y(_14184_));
 NAND2x1_ASAP7_75t_R _31509_ (.A(_13711_),
    .B(_00692_),
    .Y(_14185_));
 OA211x2_ASAP7_75t_R _31510_ (.A1(_13651_),
    .A2(_14184_),
    .B(_14185_),
    .C(_13348_),
    .Y(_14186_));
 OA211x2_ASAP7_75t_R _31511_ (.A1(_14183_),
    .A2(_14186_),
    .B(_13305_),
    .C(_13416_),
    .Y(_14187_));
 OR4x1_ASAP7_75t_R _31512_ (.A(_14166_),
    .B(_14173_),
    .C(_14180_),
    .D(_14187_),
    .Y(_14188_));
 AND2x2_ASAP7_75t_R _31513_ (.A(_13773_),
    .B(_01786_),
    .Y(_14189_));
 AO21x1_ASAP7_75t_R _31514_ (.A1(_13328_),
    .A2(_00686_),
    .B(_14189_),
    .Y(_14190_));
 BUFx12f_ASAP7_75t_R _31515_ (.A(_13323_),
    .Y(_14191_));
 OAI22x1_ASAP7_75t_R _31516_ (.A1(_00685_),
    .A2(_13670_),
    .B1(_14190_),
    .B2(_14191_),
    .Y(_14192_));
 INVx2_ASAP7_75t_R _31517_ (.A(_00702_),
    .Y(_14193_));
 NAND2x1_ASAP7_75t_R _31518_ (.A(_13695_),
    .B(_00700_),
    .Y(_14194_));
 OA211x2_ASAP7_75t_R _31519_ (.A1(_13734_),
    .A2(_14193_),
    .B(_14194_),
    .C(_13750_),
    .Y(_14195_));
 INVx1_ASAP7_75t_R _31520_ (.A(_00701_),
    .Y(_14196_));
 NAND2x1_ASAP7_75t_R _31521_ (.A(_13695_),
    .B(_00699_),
    .Y(_14197_));
 OA211x2_ASAP7_75t_R _31522_ (.A1(_13734_),
    .A2(_14196_),
    .B(_14197_),
    .C(_13673_),
    .Y(_14198_));
 OR3x2_ASAP7_75t_R _31523_ (.A(_13306_),
    .B(_14195_),
    .C(_14198_),
    .Y(_14199_));
 OA211x2_ASAP7_75t_R _31524_ (.A1(_13764_),
    .A2(_14192_),
    .B(_14199_),
    .C(_13310_),
    .Y(_14200_));
 AO211x2_ASAP7_75t_R _31525_ (.A1(_13764_),
    .A2(_14159_),
    .B(_14188_),
    .C(_14200_),
    .Y(_14201_));
 INVx3_ASAP7_75t_R _31526_ (.A(_01510_),
    .Y(_14202_));
 AO32x1_ASAP7_75t_R _31527_ (.A1(_13260_),
    .A2(_13300_),
    .A3(_14201_),
    .B1(_13839_),
    .B2(_14202_),
    .Y(_14203_));
 BUFx3_ASAP7_75t_R _31528_ (.A(_14203_),
    .Y(_18603_));
 INVx1_ASAP7_75t_R _31529_ (.A(_18603_),
    .Y(_18605_));
 INVx1_ASAP7_75t_R _31530_ (.A(_00733_),
    .Y(_14204_));
 NOR2x1_ASAP7_75t_R _31531_ (.A(_13347_),
    .B(_00735_),
    .Y(_14205_));
 AO21x1_ASAP7_75t_R _31532_ (.A1(_13518_),
    .A2(_14204_),
    .B(_14205_),
    .Y(_14206_));
 INVx2_ASAP7_75t_R _31533_ (.A(_00736_),
    .Y(_14207_));
 NAND2x1_ASAP7_75t_R _31534_ (.A(_13316_),
    .B(_00734_),
    .Y(_14208_));
 OA211x2_ASAP7_75t_R _31535_ (.A1(_13402_),
    .A2(_14207_),
    .B(_14208_),
    .C(_13345_),
    .Y(_14209_));
 AO21x1_ASAP7_75t_R _31536_ (.A1(_13673_),
    .A2(_14206_),
    .B(_14209_),
    .Y(_14210_));
 INVx1_ASAP7_75t_R _31537_ (.A(_00720_),
    .Y(_14211_));
 NAND2x1_ASAP7_75t_R _31538_ (.A(_13517_),
    .B(_00718_),
    .Y(_14212_));
 OA211x2_ASAP7_75t_R _31539_ (.A1(_13616_),
    .A2(_14211_),
    .B(_14212_),
    .C(_13345_),
    .Y(_14213_));
 INVx1_ASAP7_75t_R _31540_ (.A(_00719_),
    .Y(_14214_));
 NAND2x1_ASAP7_75t_R _31541_ (.A(_13517_),
    .B(_00717_),
    .Y(_14215_));
 OA211x2_ASAP7_75t_R _31542_ (.A1(_13616_),
    .A2(_14214_),
    .B(_14215_),
    .C(_13393_),
    .Y(_14216_));
 OR3x1_ASAP7_75t_R _31543_ (.A(_13375_),
    .B(_14213_),
    .C(_14216_),
    .Y(_14217_));
 OA21x2_ASAP7_75t_R _31544_ (.A1(_13386_),
    .A2(_14210_),
    .B(_14217_),
    .Y(_14218_));
 AND2x2_ASAP7_75t_R _31545_ (.A(_13338_),
    .B(_01785_),
    .Y(_14219_));
 AO21x1_ASAP7_75t_R _31546_ (.A1(_13313_),
    .A2(_00716_),
    .B(_14219_),
    .Y(_14220_));
 OAI22x1_ASAP7_75t_R _31547_ (.A1(_00715_),
    .A2(_13670_),
    .B1(_14220_),
    .B2(_13353_),
    .Y(_14221_));
 INVx2_ASAP7_75t_R _31548_ (.A(_00732_),
    .Y(_14222_));
 NAND2x1_ASAP7_75t_R _31549_ (.A(net1977),
    .B(_00730_),
    .Y(_14223_));
 OA211x2_ASAP7_75t_R _31550_ (.A1(_13498_),
    .A2(_14222_),
    .B(_14223_),
    .C(_13344_),
    .Y(_14224_));
 INVx2_ASAP7_75t_R _31551_ (.A(_00731_),
    .Y(_14225_));
 NAND2x1_ASAP7_75t_R _31552_ (.A(net1977),
    .B(_00729_),
    .Y(_14226_));
 OA211x2_ASAP7_75t_R _31553_ (.A1(_13498_),
    .A2(_14225_),
    .B(_14226_),
    .C(_13321_),
    .Y(_14227_));
 OR4x1_ASAP7_75t_R _31554_ (.A(_13388_),
    .B(_13389_),
    .C(_14224_),
    .D(_14227_),
    .Y(_14228_));
 OA21x2_ASAP7_75t_R _31555_ (.A1(_13485_),
    .A2(_14221_),
    .B(_14228_),
    .Y(_14229_));
 INVx2_ASAP7_75t_R _31556_ (.A(_00728_),
    .Y(_14230_));
 NAND2x1_ASAP7_75t_R _31557_ (.A(_13338_),
    .B(_00726_),
    .Y(_14231_));
 OA211x2_ASAP7_75t_R _31558_ (.A1(_13378_),
    .A2(_14230_),
    .B(_13637_),
    .C(_14231_),
    .Y(_14232_));
 INVx1_ASAP7_75t_R _31559_ (.A(_00725_),
    .Y(_14233_));
 NOR2x1_ASAP7_75t_R _31560_ (.A(_13391_),
    .B(_00727_),
    .Y(_14234_));
 AO21x1_ASAP7_75t_R _31561_ (.A1(_13481_),
    .A2(_14233_),
    .B(_14234_),
    .Y(_14235_));
 INVx1_ASAP7_75t_R _31562_ (.A(_00723_),
    .Y(_14236_));
 NAND2x1_ASAP7_75t_R _31563_ (.A(_13362_),
    .B(_00721_),
    .Y(_14237_));
 OA211x2_ASAP7_75t_R _31564_ (.A1(_13316_),
    .A2(_14236_),
    .B(_13646_),
    .C(_14237_),
    .Y(_14238_));
 AO21x1_ASAP7_75t_R _31565_ (.A1(_13632_),
    .A2(_14235_),
    .B(_14238_),
    .Y(_14239_));
 INVx1_ASAP7_75t_R _31566_ (.A(_00724_),
    .Y(_14240_));
 NAND2x1_ASAP7_75t_R _31567_ (.A(_13498_),
    .B(_00722_),
    .Y(_14241_));
 OA211x2_ASAP7_75t_R _31568_ (.A1(_13378_),
    .A2(_14240_),
    .B(_13641_),
    .C(_14241_),
    .Y(_14242_));
 OR5x1_ASAP7_75t_R _31569_ (.A(_13459_),
    .B(_13461_),
    .C(_14232_),
    .D(_14239_),
    .E(_14242_),
    .Y(_14243_));
 INVx2_ASAP7_75t_R _31570_ (.A(_00743_),
    .Y(_14244_));
 NAND2x1_ASAP7_75t_R _31571_ (.A(_13333_),
    .B(_00739_),
    .Y(_14245_));
 OA211x2_ASAP7_75t_R _31572_ (.A1(_13842_),
    .A2(_14244_),
    .B(_14245_),
    .C(_13326_),
    .Y(_14246_));
 INVx1_ASAP7_75t_R _31573_ (.A(_00741_),
    .Y(_14247_));
 NAND2x1_ASAP7_75t_R _31574_ (.A(_13333_),
    .B(_00737_),
    .Y(_14248_));
 OA211x2_ASAP7_75t_R _31575_ (.A1(_13400_),
    .A2(_14247_),
    .B(_14248_),
    .C(_13481_),
    .Y(_14249_));
 OR3x1_ASAP7_75t_R _31576_ (.A(_13346_),
    .B(_14246_),
    .C(_14249_),
    .Y(_14250_));
 INVx1_ASAP7_75t_R _31577_ (.A(_00744_),
    .Y(_14251_));
 NAND2x1_ASAP7_75t_R _31578_ (.A(_13333_),
    .B(_00740_),
    .Y(_14252_));
 OA211x2_ASAP7_75t_R _31579_ (.A1(_13842_),
    .A2(_14251_),
    .B(_14252_),
    .C(_13326_),
    .Y(_14253_));
 INVx1_ASAP7_75t_R _31580_ (.A(_00742_),
    .Y(_14254_));
 NAND2x1_ASAP7_75t_R _31581_ (.A(_13333_),
    .B(_00738_),
    .Y(_14255_));
 OA211x2_ASAP7_75t_R _31582_ (.A1(_13400_),
    .A2(_14254_),
    .B(_14255_),
    .C(_13481_),
    .Y(_14256_));
 OR3x1_ASAP7_75t_R _31583_ (.A(_13322_),
    .B(_14253_),
    .C(_14256_),
    .Y(_14257_));
 AO21x1_ASAP7_75t_R _31584_ (.A1(_14250_),
    .A2(_14257_),
    .B(_13365_),
    .Y(_14258_));
 AND4x1_ASAP7_75t_R _31585_ (.A(_14218_),
    .B(_14229_),
    .C(_14243_),
    .D(_14258_),
    .Y(_14259_));
 BUFx12f_ASAP7_75t_R _31586_ (.A(_14259_),
    .Y(_14260_));
 OR2x6_ASAP7_75t_R _31587_ (.A(_13763_),
    .B(_14260_),
    .Y(_14261_));
 NAND3x1_ASAP7_75t_R _31588_ (.A(_13259_),
    .B(_13427_),
    .C(_13438_),
    .Y(_14262_));
 AOI21x1_ASAP7_75t_R _31589_ (.A1(_13426_),
    .A2(_13429_),
    .B(_13272_),
    .Y(_14263_));
 NAND3x1_ASAP7_75t_R _31590_ (.A(_13434_),
    .B(_13440_),
    .C(_13443_),
    .Y(_14264_));
 NAND2x1_ASAP7_75t_R _31591_ (.A(_13248_),
    .B(_13240_),
    .Y(_14265_));
 OR3x1_ASAP7_75t_R _31592_ (.A(_13430_),
    .B(_13236_),
    .C(_14265_),
    .Y(_14266_));
 AND4x1_ASAP7_75t_R _31593_ (.A(_13277_),
    .B(_13220_),
    .C(_13263_),
    .D(_13440_),
    .Y(_14267_));
 AO211x2_ASAP7_75t_R _31594_ (.A1(_13296_),
    .A2(_13437_),
    .B(_14267_),
    .C(_14099_),
    .Y(_14268_));
 AO221x1_ASAP7_75t_R _31595_ (.A1(_13440_),
    .A2(_13443_),
    .B1(_14266_),
    .B2(_14268_),
    .C(_13272_),
    .Y(_14269_));
 OA31x2_ASAP7_75t_R _31596_ (.A1(_14262_),
    .A2(_14263_),
    .A3(_14264_),
    .B1(_14269_),
    .Y(_14270_));
 NAND2x1_ASAP7_75t_R _31597_ (.A(_13763_),
    .B(_14270_),
    .Y(_14271_));
 NAND2x2_ASAP7_75t_R _31598_ (.A(_14261_),
    .B(_14271_),
    .Y(_18610_));
 INVx4_ASAP7_75t_R _31599_ (.A(_18610_),
    .Y(_18608_));
 BUFx6f_ASAP7_75t_R _31600_ (.A(_13421_),
    .Y(_14272_));
 BUFx6f_ASAP7_75t_R _31601_ (.A(_14272_),
    .Y(_14273_));
 BUFx12f_ASAP7_75t_R _31602_ (.A(_14121_),
    .Y(_14274_));
 OR5x2_ASAP7_75t_R _31603_ (.A(_13280_),
    .B(_13230_),
    .C(_14124_),
    .D(_13285_),
    .E(_13223_),
    .Y(_14275_));
 AO21x1_ASAP7_75t_R _31604_ (.A1(_14274_),
    .A2(_14093_),
    .B(_14275_),
    .Y(_14276_));
 OR2x6_ASAP7_75t_R _31605_ (.A(_14273_),
    .B(_14276_),
    .Y(_18075_));
 INVx1_ASAP7_75t_R _31606_ (.A(_18075_),
    .Y(_18076_));
 BUFx12f_ASAP7_75t_R _31607_ (.A(_13188_),
    .Y(_14277_));
 BUFx12f_ASAP7_75t_R _31608_ (.A(_14277_),
    .Y(_14278_));
 NAND2x1_ASAP7_75t_R _31609_ (.A(_14278_),
    .B(_14092_),
    .Y(_14279_));
 AND3x4_ASAP7_75t_R _31610_ (.A(_14274_),
    .B(_13265_),
    .C(_14279_),
    .Y(_14280_));
 BUFx6f_ASAP7_75t_R _31611_ (.A(_14280_),
    .Y(_18074_));
 INVx1_ASAP7_75t_R _31612_ (.A(_18074_),
    .Y(_18078_));
 BUFx12f_ASAP7_75t_R _31613_ (.A(_13081_),
    .Y(_14281_));
 BUFx12f_ASAP7_75t_R _31614_ (.A(_13084_),
    .Y(_14282_));
 BUFx12f_ASAP7_75t_R _31615_ (.A(_14282_),
    .Y(_14283_));
 BUFx12f_ASAP7_75t_R _31616_ (.A(_13101_),
    .Y(_14284_));
 BUFx12f_ASAP7_75t_R _31617_ (.A(_13091_),
    .Y(_14285_));
 BUFx6f_ASAP7_75t_R _31618_ (.A(_14285_),
    .Y(_14286_));
 AND2x2_ASAP7_75t_R _31619_ (.A(_13193_),
    .B(_01785_),
    .Y(_14287_));
 AO21x1_ASAP7_75t_R _31620_ (.A1(_14286_),
    .A2(_00716_),
    .B(_14287_),
    .Y(_14288_));
 BUFx12f_ASAP7_75t_R _31621_ (.A(_13089_),
    .Y(_14289_));
 OAI22x1_ASAP7_75t_R _31622_ (.A1(_00715_),
    .A2(_14284_),
    .B1(_14288_),
    .B2(_14289_),
    .Y(_14290_));
 BUFx12f_ASAP7_75t_R _31623_ (.A(_13152_),
    .Y(_14291_));
 BUFx12f_ASAP7_75t_R _31624_ (.A(_13109_),
    .Y(_14292_));
 BUFx12f_ASAP7_75t_R _31625_ (.A(_14292_),
    .Y(_14293_));
 NAND2x1_ASAP7_75t_R _31626_ (.A(_14277_),
    .B(_00722_),
    .Y(_14294_));
 BUFx12f_ASAP7_75t_R _31627_ (.A(_13113_),
    .Y(_14295_));
 BUFx6f_ASAP7_75t_R _31628_ (.A(_14295_),
    .Y(_14296_));
 OA211x2_ASAP7_75t_R _31629_ (.A1(_14293_),
    .A2(_14240_),
    .B(_14294_),
    .C(_14296_),
    .Y(_14297_));
 BUFx12f_ASAP7_75t_R _31630_ (.A(_13095_),
    .Y(_14298_));
 BUFx6f_ASAP7_75t_R _31631_ (.A(_14298_),
    .Y(_14299_));
 BUFx12f_ASAP7_75t_R _31632_ (.A(_13135_),
    .Y(_14300_));
 BUFx12f_ASAP7_75t_R _31633_ (.A(_14300_),
    .Y(_14301_));
 NAND2x1_ASAP7_75t_R _31634_ (.A(_14301_),
    .B(_00721_),
    .Y(_14302_));
 OA211x2_ASAP7_75t_R _31635_ (.A1(_14299_),
    .A2(_14236_),
    .B(_14302_),
    .C(_13149_),
    .Y(_14303_));
 OR3x1_ASAP7_75t_R _31636_ (.A(_14291_),
    .B(_14297_),
    .C(_14303_),
    .Y(_14304_));
 BUFx12f_ASAP7_75t_R _31637_ (.A(_13124_),
    .Y(_14305_));
 OA211x2_ASAP7_75t_R _31638_ (.A1(_14283_),
    .A2(_14290_),
    .B(_14304_),
    .C(_14305_),
    .Y(_14306_));
 BUFx12f_ASAP7_75t_R _31639_ (.A(_13128_),
    .Y(_14307_));
 BUFx12f_ASAP7_75t_R _31640_ (.A(_13084_),
    .Y(_14308_));
 BUFx12f_ASAP7_75t_R _31641_ (.A(_14308_),
    .Y(_14309_));
 BUFx12f_ASAP7_75t_R _31642_ (.A(_13188_),
    .Y(_14310_));
 BUFx6f_ASAP7_75t_R _31643_ (.A(_14310_),
    .Y(_14311_));
 BUFx12f_ASAP7_75t_R _31644_ (.A(_13096_),
    .Y(_14312_));
 NAND2x1_ASAP7_75t_R _31645_ (.A(_14312_),
    .B(_00718_),
    .Y(_14313_));
 BUFx12f_ASAP7_75t_R _31646_ (.A(_13113_),
    .Y(_14314_));
 BUFx6f_ASAP7_75t_R _31647_ (.A(_14314_),
    .Y(_14315_));
 OA211x2_ASAP7_75t_R _31648_ (.A1(_14311_),
    .A2(_14211_),
    .B(_14313_),
    .C(_14315_),
    .Y(_14316_));
 BUFx12f_ASAP7_75t_R _31649_ (.A(_13109_),
    .Y(_14317_));
 BUFx6f_ASAP7_75t_R _31650_ (.A(_14317_),
    .Y(_14318_));
 BUFx12f_ASAP7_75t_R _31651_ (.A(_13135_),
    .Y(_14319_));
 BUFx12f_ASAP7_75t_R _31652_ (.A(_14319_),
    .Y(_14320_));
 NAND2x1_ASAP7_75t_R _31653_ (.A(_14320_),
    .B(_00717_),
    .Y(_14321_));
 BUFx6f_ASAP7_75t_R _31654_ (.A(_13087_),
    .Y(_14322_));
 BUFx6f_ASAP7_75t_R _31655_ (.A(_14322_),
    .Y(_14323_));
 OA211x2_ASAP7_75t_R _31656_ (.A1(_14318_),
    .A2(_14214_),
    .B(_14321_),
    .C(_14323_),
    .Y(_14324_));
 OR3x1_ASAP7_75t_R _31657_ (.A(_14309_),
    .B(_14316_),
    .C(_14324_),
    .Y(_14325_));
 BUFx12f_ASAP7_75t_R _31658_ (.A(_13104_),
    .Y(_14326_));
 BUFx12f_ASAP7_75t_R _31659_ (.A(_14326_),
    .Y(_14327_));
 NAND2x1_ASAP7_75t_R _31660_ (.A(_14312_),
    .B(_00726_),
    .Y(_14328_));
 BUFx6f_ASAP7_75t_R _31661_ (.A(_14314_),
    .Y(_14329_));
 OA211x2_ASAP7_75t_R _31662_ (.A1(_14318_),
    .A2(_14230_),
    .B(_14328_),
    .C(_14329_),
    .Y(_14330_));
 BUFx6f_ASAP7_75t_R _31663_ (.A(_13211_),
    .Y(_14331_));
 INVx1_ASAP7_75t_R _31664_ (.A(_00727_),
    .Y(_14332_));
 BUFx12f_ASAP7_75t_R _31665_ (.A(_14319_),
    .Y(_14333_));
 NAND2x1_ASAP7_75t_R _31666_ (.A(_14333_),
    .B(_00725_),
    .Y(_14334_));
 OA211x2_ASAP7_75t_R _31667_ (.A1(_14331_),
    .A2(_14332_),
    .B(_14334_),
    .C(_14323_),
    .Y(_14335_));
 OR3x1_ASAP7_75t_R _31668_ (.A(_14327_),
    .B(_14330_),
    .C(_14335_),
    .Y(_14336_));
 AND3x4_ASAP7_75t_R _31669_ (.A(_14307_),
    .B(_14325_),
    .C(_14336_),
    .Y(_14337_));
 OR3x2_ASAP7_75t_R _31670_ (.A(_14281_),
    .B(_14306_),
    .C(_14337_),
    .Y(_14338_));
 BUFx12f_ASAP7_75t_R _31671_ (.A(_13163_),
    .Y(_14339_));
 BUFx12f_ASAP7_75t_R _31672_ (.A(_13128_),
    .Y(_14340_));
 NAND2x1_ASAP7_75t_R _31673_ (.A(_14312_),
    .B(_00734_),
    .Y(_14341_));
 OA211x2_ASAP7_75t_R _31674_ (.A1(_14311_),
    .A2(_14207_),
    .B(_14341_),
    .C(_14315_),
    .Y(_14342_));
 INVx1_ASAP7_75t_R _31675_ (.A(_00735_),
    .Y(_14343_));
 NAND2x1_ASAP7_75t_R _31676_ (.A(_14320_),
    .B(_00733_),
    .Y(_14344_));
 OA211x2_ASAP7_75t_R _31677_ (.A1(_14318_),
    .A2(_14343_),
    .B(_14344_),
    .C(_14323_),
    .Y(_14345_));
 OR3x1_ASAP7_75t_R _31678_ (.A(_14309_),
    .B(_14342_),
    .C(_14345_),
    .Y(_14346_));
 NAND2x1_ASAP7_75t_R _31679_ (.A(_14312_),
    .B(_00742_),
    .Y(_14347_));
 OA211x2_ASAP7_75t_R _31680_ (.A1(_14318_),
    .A2(_14251_),
    .B(_14347_),
    .C(_14329_),
    .Y(_14348_));
 NAND2x1_ASAP7_75t_R _31681_ (.A(_14333_),
    .B(_00741_),
    .Y(_14349_));
 OA211x2_ASAP7_75t_R _31682_ (.A1(_14331_),
    .A2(_14244_),
    .B(_14349_),
    .C(_14323_),
    .Y(_14350_));
 OR3x1_ASAP7_75t_R _31683_ (.A(_14327_),
    .B(_14348_),
    .C(_14350_),
    .Y(_14351_));
 AND3x1_ASAP7_75t_R _31684_ (.A(_14340_),
    .B(_14346_),
    .C(_14351_),
    .Y(_14352_));
 BUFx12f_ASAP7_75t_R _31685_ (.A(_13104_),
    .Y(_14353_));
 BUFx12f_ASAP7_75t_R _31686_ (.A(_14353_),
    .Y(_14354_));
 INVx1_ASAP7_75t_R _31687_ (.A(_00737_),
    .Y(_14355_));
 NOR2x1_ASAP7_75t_R _31688_ (.A(_13143_),
    .B(_00739_),
    .Y(_14356_));
 AO21x1_ASAP7_75t_R _31689_ (.A1(_14278_),
    .A2(_14355_),
    .B(_14356_),
    .Y(_14357_));
 BUFx6f_ASAP7_75t_R _31690_ (.A(_14310_),
    .Y(_14358_));
 INVx1_ASAP7_75t_R _31691_ (.A(_00740_),
    .Y(_14359_));
 BUFx12f_ASAP7_75t_R _31692_ (.A(_14319_),
    .Y(_14360_));
 NAND2x1_ASAP7_75t_R _31693_ (.A(_14360_),
    .B(_00738_),
    .Y(_14361_));
 BUFx6f_ASAP7_75t_R _31694_ (.A(_13113_),
    .Y(_14362_));
 BUFx12f_ASAP7_75t_R _31695_ (.A(_14362_),
    .Y(_14363_));
 OA211x2_ASAP7_75t_R _31696_ (.A1(_14358_),
    .A2(_14359_),
    .B(_14361_),
    .C(_14363_),
    .Y(_14364_));
 AO21x1_ASAP7_75t_R _31697_ (.A1(_13090_),
    .A2(_14357_),
    .B(_14364_),
    .Y(_14365_));
 BUFx12f_ASAP7_75t_R _31698_ (.A(_13106_),
    .Y(_14366_));
 BUFx12f_ASAP7_75t_R _31699_ (.A(_13188_),
    .Y(_14367_));
 NAND2x1_ASAP7_75t_R _31700_ (.A(_14367_),
    .B(_00730_),
    .Y(_14368_));
 BUFx12f_ASAP7_75t_R _31701_ (.A(_14295_),
    .Y(_14369_));
 OA211x2_ASAP7_75t_R _31702_ (.A1(_14366_),
    .A2(_14222_),
    .B(_14368_),
    .C(_14369_),
    .Y(_14370_));
 NAND2x1_ASAP7_75t_R _31703_ (.A(_14367_),
    .B(_00729_),
    .Y(_14371_));
 BUFx12f_ASAP7_75t_R _31704_ (.A(_13148_),
    .Y(_14372_));
 OA211x2_ASAP7_75t_R _31705_ (.A1(_14366_),
    .A2(_14225_),
    .B(_14371_),
    .C(_14372_),
    .Y(_14373_));
 OR3x1_ASAP7_75t_R _31706_ (.A(_14282_),
    .B(_14370_),
    .C(_14373_),
    .Y(_14374_));
 OA211x2_ASAP7_75t_R _31707_ (.A1(_14354_),
    .A2(_14365_),
    .B(_14374_),
    .C(_14305_),
    .Y(_14375_));
 OR3x2_ASAP7_75t_R _31708_ (.A(_14339_),
    .B(_14352_),
    .C(_14375_),
    .Y(_14376_));
 BUFx6f_ASAP7_75t_R _31709_ (.A(_13267_),
    .Y(_14377_));
 AO21x2_ASAP7_75t_R _31710_ (.A1(_14338_),
    .A2(_14376_),
    .B(_14377_),
    .Y(_14378_));
 BUFx6f_ASAP7_75t_R _31711_ (.A(_01504_),
    .Y(_14379_));
 AO211x2_ASAP7_75t_R _31712_ (.A1(_13279_),
    .A2(_13284_),
    .B(_13286_),
    .C(_13291_),
    .Y(_14380_));
 BUFx6f_ASAP7_75t_R _31713_ (.A(_14380_),
    .Y(_14381_));
 BUFx12f_ASAP7_75t_R _31714_ (.A(_14381_),
    .Y(_14382_));
 AOI21x1_ASAP7_75t_R _31715_ (.A1(_13252_),
    .A2(_13266_),
    .B(_13272_),
    .Y(_14383_));
 BUFx12f_ASAP7_75t_R _31716_ (.A(_14383_),
    .Y(_14384_));
 BUFx6f_ASAP7_75t_R _31717_ (.A(_14384_),
    .Y(_14385_));
 AND2x2_ASAP7_75t_R _31718_ (.A(_01475_),
    .B(_14381_),
    .Y(_14386_));
 OAI22x1_ASAP7_75t_R _31719_ (.A1(_14379_),
    .A2(_14382_),
    .B1(_14385_),
    .B2(_14386_),
    .Y(_14387_));
 AND2x6_ASAP7_75t_R _31720_ (.A(_14378_),
    .B(_14387_),
    .Y(_18607_));
 INVx2_ASAP7_75t_R _31721_ (.A(_18607_),
    .Y(_18609_));
 NAND2x2_ASAP7_75t_R _31722_ (.A(_14119_),
    .B(_13265_),
    .Y(_14388_));
 OR3x1_ASAP7_75t_R _31723_ (.A(_14289_),
    .B(_13292_),
    .C(_14388_),
    .Y(_14389_));
 AOI22x1_ASAP7_75t_R _31724_ (.A1(_01477_),
    .A2(_13272_),
    .B1(_14384_),
    .B2(_14389_),
    .Y(_14390_));
 BUFx12f_ASAP7_75t_R _31725_ (.A(_13135_),
    .Y(_14391_));
 AND2x2_ASAP7_75t_R _31726_ (.A(_14391_),
    .B(_01796_),
    .Y(_14392_));
 AO21x1_ASAP7_75t_R _31727_ (.A1(_14285_),
    .A2(_00382_),
    .B(_14392_),
    .Y(_14393_));
 OAI22x1_ASAP7_75t_R _31728_ (.A1(_00381_),
    .A2(_13101_),
    .B1(_14393_),
    .B2(_13089_),
    .Y(_14394_));
 INVx1_ASAP7_75t_R _31729_ (.A(_00390_),
    .Y(_14395_));
 NAND2x1_ASAP7_75t_R _31730_ (.A(_13188_),
    .B(_00388_),
    .Y(_14396_));
 OA211x2_ASAP7_75t_R _31731_ (.A1(_13205_),
    .A2(_14395_),
    .B(_14396_),
    .C(_13114_),
    .Y(_14397_));
 INVx1_ASAP7_75t_R _31732_ (.A(_00389_),
    .Y(_14398_));
 NAND2x1_ASAP7_75t_R _31733_ (.A(_13109_),
    .B(_00387_),
    .Y(_14399_));
 OA211x2_ASAP7_75t_R _31734_ (.A1(_13205_),
    .A2(_14398_),
    .B(_14399_),
    .C(_13100_),
    .Y(_14400_));
 OR3x1_ASAP7_75t_R _31735_ (.A(_13104_),
    .B(_14397_),
    .C(_14400_),
    .Y(_14401_));
 OA211x2_ASAP7_75t_R _31736_ (.A1(_13085_),
    .A2(_14394_),
    .B(_14401_),
    .C(_13124_),
    .Y(_14402_));
 BUFx12f_ASAP7_75t_R _31737_ (.A(_13095_),
    .Y(_14403_));
 NAND2x1_ASAP7_75t_R _31738_ (.A(_13199_),
    .B(_00384_),
    .Y(_14404_));
 OA211x2_ASAP7_75t_R _31739_ (.A1(_14403_),
    .A2(_13367_),
    .B(_14404_),
    .C(_14295_),
    .Y(_14405_));
 NAND2x1_ASAP7_75t_R _31740_ (.A(_13145_),
    .B(_00383_),
    .Y(_14406_));
 OA211x2_ASAP7_75t_R _31741_ (.A1(_13132_),
    .A2(_13371_),
    .B(_14406_),
    .C(_13148_),
    .Y(_14407_));
 OR3x1_ASAP7_75t_R _31742_ (.A(_13130_),
    .B(_14405_),
    .C(_14407_),
    .Y(_14408_));
 NAND2x1_ASAP7_75t_R _31743_ (.A(_14300_),
    .B(_00392_),
    .Y(_14409_));
 OA211x2_ASAP7_75t_R _31744_ (.A1(_14403_),
    .A2(_13410_),
    .B(_14409_),
    .C(_14295_),
    .Y(_14410_));
 INVx1_ASAP7_75t_R _31745_ (.A(_00393_),
    .Y(_14411_));
 NAND2x1_ASAP7_75t_R _31746_ (.A(_13145_),
    .B(_00391_),
    .Y(_14412_));
 OA211x2_ASAP7_75t_R _31747_ (.A1(_13132_),
    .A2(_14411_),
    .B(_14412_),
    .C(_13148_),
    .Y(_14413_));
 OR3x1_ASAP7_75t_R _31748_ (.A(_13152_),
    .B(_14410_),
    .C(_14413_),
    .Y(_14414_));
 AND3x1_ASAP7_75t_R _31749_ (.A(_13128_),
    .B(_14408_),
    .C(_14414_),
    .Y(_14415_));
 OR3x2_ASAP7_75t_R _31750_ (.A(_13081_),
    .B(_14402_),
    .C(_14415_),
    .Y(_14416_));
 NAND2x1_ASAP7_75t_R _31751_ (.A(_13199_),
    .B(_00400_),
    .Y(_14417_));
 OA211x2_ASAP7_75t_R _31752_ (.A1(_14298_),
    .A2(_13379_),
    .B(_14417_),
    .C(_13139_),
    .Y(_14418_));
 NAND2x1_ASAP7_75t_R _31753_ (.A(_14300_),
    .B(_00399_),
    .Y(_14419_));
 OA211x2_ASAP7_75t_R _31754_ (.A1(_14403_),
    .A2(_13382_),
    .B(_14419_),
    .C(_13173_),
    .Y(_14420_));
 OR3x1_ASAP7_75t_R _31755_ (.A(_13130_),
    .B(_14418_),
    .C(_14420_),
    .Y(_14421_));
 NAND2x1_ASAP7_75t_R _31756_ (.A(_13199_),
    .B(_00408_),
    .Y(_14422_));
 OA211x2_ASAP7_75t_R _31757_ (.A1(_14403_),
    .A2(_13355_),
    .B(_14422_),
    .C(_14295_),
    .Y(_14423_));
 NAND2x1_ASAP7_75t_R _31758_ (.A(_14300_),
    .B(_00407_),
    .Y(_14424_));
 OA211x2_ASAP7_75t_R _31759_ (.A1(_14403_),
    .A2(_13404_),
    .B(_14424_),
    .C(_13148_),
    .Y(_14425_));
 OR3x1_ASAP7_75t_R _31760_ (.A(_13152_),
    .B(_14423_),
    .C(_14425_),
    .Y(_14426_));
 AND3x1_ASAP7_75t_R _31761_ (.A(_13128_),
    .B(_14421_),
    .C(_14426_),
    .Y(_14427_));
 BUFx12f_ASAP7_75t_R _31762_ (.A(_13124_),
    .Y(_14428_));
 NAND2x1_ASAP7_75t_R _31763_ (.A(_14300_),
    .B(_00396_),
    .Y(_14429_));
 OA211x2_ASAP7_75t_R _31764_ (.A1(_14403_),
    .A2(_13395_),
    .B(_14429_),
    .C(_14295_),
    .Y(_14430_));
 NAND2x1_ASAP7_75t_R _31765_ (.A(_13145_),
    .B(_00395_),
    .Y(_14431_));
 OA211x2_ASAP7_75t_R _31766_ (.A1(_13132_),
    .A2(_13390_),
    .B(_14431_),
    .C(_13148_),
    .Y(_14432_));
 OR3x1_ASAP7_75t_R _31767_ (.A(_13084_),
    .B(_14430_),
    .C(_14432_),
    .Y(_14433_));
 INVx1_ASAP7_75t_R _31768_ (.A(_00406_),
    .Y(_14434_));
 NAND2x1_ASAP7_75t_R _31769_ (.A(_13145_),
    .B(_00404_),
    .Y(_14435_));
 OA211x2_ASAP7_75t_R _31770_ (.A1(_13132_),
    .A2(_14434_),
    .B(_14435_),
    .C(_14295_),
    .Y(_14436_));
 BUFx12f_ASAP7_75t_R _31771_ (.A(_13095_),
    .Y(_14437_));
 INVx1_ASAP7_75t_R _31772_ (.A(_00405_),
    .Y(_14438_));
 NAND2x1_ASAP7_75t_R _31773_ (.A(_13145_),
    .B(_00403_),
    .Y(_14439_));
 OA211x2_ASAP7_75t_R _31774_ (.A1(_14437_),
    .A2(_14438_),
    .B(_14439_),
    .C(_13148_),
    .Y(_14440_));
 OR3x1_ASAP7_75t_R _31775_ (.A(_13152_),
    .B(_14436_),
    .C(_14440_),
    .Y(_14441_));
 AND3x1_ASAP7_75t_R _31776_ (.A(_14428_),
    .B(_14433_),
    .C(_14441_),
    .Y(_14442_));
 OR3x2_ASAP7_75t_R _31777_ (.A(_13163_),
    .B(_14427_),
    .C(_14442_),
    .Y(_14443_));
 AO21x2_ASAP7_75t_R _31778_ (.A1(_14416_),
    .A2(_14443_),
    .B(_13267_),
    .Y(_14444_));
 AND2x6_ASAP7_75t_R _31779_ (.A(_14390_),
    .B(_14444_),
    .Y(_18554_));
 INVx2_ASAP7_75t_R _31780_ (.A(_18554_),
    .Y(_18556_));
 INVx1_ASAP7_75t_R _31781_ (.A(_01496_),
    .Y(\cs_registers_i.pc_id_i[1] ));
 AND3x1_ASAP7_75t_R _31782_ (.A(_13252_),
    .B(_13259_),
    .C(_13266_),
    .Y(_14445_));
 BUFx6f_ASAP7_75t_R _31783_ (.A(_14445_),
    .Y(_14446_));
 BUFx12f_ASAP7_75t_R _31784_ (.A(_13081_),
    .Y(_14447_));
 BUFx12f_ASAP7_75t_R _31785_ (.A(_14308_),
    .Y(_14448_));
 AND2x4_ASAP7_75t_R _31786_ (.A(_13087_),
    .B(_13091_),
    .Y(_14449_));
 BUFx12f_ASAP7_75t_R _31787_ (.A(_13145_),
    .Y(_14450_));
 NAND2x1_ASAP7_75t_R _31788_ (.A(_14450_),
    .B(_01795_),
    .Y(_14451_));
 OA211x2_ASAP7_75t_R _31789_ (.A1(_14366_),
    .A2(_13480_),
    .B(_14451_),
    .C(_14369_),
    .Y(_14452_));
 AO21x1_ASAP7_75t_R _31790_ (.A1(_13478_),
    .A2(_14449_),
    .B(_14452_),
    .Y(_14453_));
 BUFx12f_ASAP7_75t_R _31791_ (.A(_13104_),
    .Y(_14454_));
 BUFx12f_ASAP7_75t_R _31792_ (.A(_13136_),
    .Y(_14455_));
 INVx1_ASAP7_75t_R _31793_ (.A(_00423_),
    .Y(_14456_));
 NAND2x1_ASAP7_75t_R _31794_ (.A(_13142_),
    .B(_00421_),
    .Y(_14457_));
 BUFx12f_ASAP7_75t_R _31795_ (.A(_13114_),
    .Y(_14458_));
 OA211x2_ASAP7_75t_R _31796_ (.A1(_14455_),
    .A2(_14456_),
    .B(_14457_),
    .C(_14458_),
    .Y(_14459_));
 BUFx12f_ASAP7_75t_R _31797_ (.A(_13135_),
    .Y(_14460_));
 BUFx12f_ASAP7_75t_R _31798_ (.A(_14460_),
    .Y(_14461_));
 NAND2x1_ASAP7_75t_R _31799_ (.A(_14292_),
    .B(_00420_),
    .Y(_14462_));
 BUFx6f_ASAP7_75t_R _31800_ (.A(_13100_),
    .Y(_14463_));
 OA211x2_ASAP7_75t_R _31801_ (.A1(_14461_),
    .A2(_13473_),
    .B(_14462_),
    .C(_14463_),
    .Y(_14464_));
 OR3x1_ASAP7_75t_R _31802_ (.A(_14454_),
    .B(_14459_),
    .C(_14464_),
    .Y(_14465_));
 BUFx12f_ASAP7_75t_R _31803_ (.A(_13124_),
    .Y(_14466_));
 OA211x2_ASAP7_75t_R _31804_ (.A1(_14448_),
    .A2(_14453_),
    .B(_14465_),
    .C(_14466_),
    .Y(_14467_));
 BUFx12f_ASAP7_75t_R _31805_ (.A(_13128_),
    .Y(_14468_));
 BUFx12f_ASAP7_75t_R _31806_ (.A(_13084_),
    .Y(_14469_));
 BUFx12f_ASAP7_75t_R _31807_ (.A(_13188_),
    .Y(_14470_));
 NAND2x1_ASAP7_75t_R _31808_ (.A(_14470_),
    .B(_00417_),
    .Y(_14471_));
 BUFx12f_ASAP7_75t_R _31809_ (.A(_13114_),
    .Y(_14472_));
 OA211x2_ASAP7_75t_R _31810_ (.A1(_13193_),
    .A2(_13497_),
    .B(_14471_),
    .C(_14472_),
    .Y(_14473_));
 BUFx12f_ASAP7_75t_R _31811_ (.A(_13192_),
    .Y(_14474_));
 NAND2x1_ASAP7_75t_R _31812_ (.A(_14310_),
    .B(_00416_),
    .Y(_14475_));
 BUFx12f_ASAP7_75t_R _31813_ (.A(_13100_),
    .Y(_14476_));
 OA211x2_ASAP7_75t_R _31814_ (.A1(_14474_),
    .A2(_13501_),
    .B(_14475_),
    .C(_14476_),
    .Y(_14477_));
 OR3x1_ASAP7_75t_R _31815_ (.A(_14469_),
    .B(_14473_),
    .C(_14477_),
    .Y(_14478_));
 NAND2x1_ASAP7_75t_R _31816_ (.A(_14470_),
    .B(_00425_),
    .Y(_14479_));
 OA211x2_ASAP7_75t_R _31817_ (.A1(_13193_),
    .A2(_13462_),
    .B(_14479_),
    .C(_14472_),
    .Y(_14480_));
 INVx1_ASAP7_75t_R _31818_ (.A(_00426_),
    .Y(_14481_));
 NAND2x1_ASAP7_75t_R _31819_ (.A(_14317_),
    .B(_00424_),
    .Y(_14482_));
 OA211x2_ASAP7_75t_R _31820_ (.A1(_14474_),
    .A2(_14481_),
    .B(_14482_),
    .C(_14476_),
    .Y(_14483_));
 OR3x1_ASAP7_75t_R _31821_ (.A(_13105_),
    .B(_14480_),
    .C(_14483_),
    .Y(_14484_));
 AND3x1_ASAP7_75t_R _31822_ (.A(_14468_),
    .B(_14478_),
    .C(_14484_),
    .Y(_14485_));
 OR3x2_ASAP7_75t_R _31823_ (.A(_14447_),
    .B(_14467_),
    .C(_14485_),
    .Y(_14486_));
 BUFx12f_ASAP7_75t_R _31824_ (.A(_13163_),
    .Y(_14487_));
 BUFx12f_ASAP7_75t_R _31825_ (.A(_13128_),
    .Y(_14488_));
 BUFx12f_ASAP7_75t_R _31826_ (.A(_13084_),
    .Y(_14489_));
 BUFx12f_ASAP7_75t_R _31827_ (.A(_13095_),
    .Y(_14490_));
 BUFx12f_ASAP7_75t_R _31828_ (.A(_14490_),
    .Y(_14491_));
 BUFx12f_ASAP7_75t_R _31829_ (.A(_13199_),
    .Y(_14492_));
 NAND2x1_ASAP7_75t_R _31830_ (.A(_14492_),
    .B(_00433_),
    .Y(_14493_));
 BUFx12f_ASAP7_75t_R _31831_ (.A(_13114_),
    .Y(_14494_));
 OA211x2_ASAP7_75t_R _31832_ (.A1(_14491_),
    .A2(_13514_),
    .B(_14493_),
    .C(_14494_),
    .Y(_14495_));
 BUFx12f_ASAP7_75t_R _31833_ (.A(_14437_),
    .Y(_14496_));
 NAND2x1_ASAP7_75t_R _31834_ (.A(_13189_),
    .B(_00432_),
    .Y(_14497_));
 BUFx12f_ASAP7_75t_R _31835_ (.A(_13100_),
    .Y(_14498_));
 OA211x2_ASAP7_75t_R _31836_ (.A1(_14496_),
    .A2(_13519_),
    .B(_14497_),
    .C(_14498_),
    .Y(_14499_));
 OR3x1_ASAP7_75t_R _31837_ (.A(_14489_),
    .B(_14495_),
    .C(_14499_),
    .Y(_14500_));
 BUFx12f_ASAP7_75t_R _31838_ (.A(_14437_),
    .Y(_14501_));
 BUFx12f_ASAP7_75t_R _31839_ (.A(_14300_),
    .Y(_14502_));
 NAND2x1_ASAP7_75t_R _31840_ (.A(_14502_),
    .B(_00441_),
    .Y(_14503_));
 BUFx12f_ASAP7_75t_R _31841_ (.A(_13114_),
    .Y(_14504_));
 OA211x2_ASAP7_75t_R _31842_ (.A1(_14501_),
    .A2(_13491_),
    .B(_14503_),
    .C(_14504_),
    .Y(_14505_));
 BUFx12f_ASAP7_75t_R _31843_ (.A(_14437_),
    .Y(_14506_));
 BUFx12f_ASAP7_75t_R _31844_ (.A(_13188_),
    .Y(_14507_));
 NAND2x1_ASAP7_75t_R _31845_ (.A(_14507_),
    .B(_00440_),
    .Y(_14508_));
 BUFx12f_ASAP7_75t_R _31846_ (.A(_13100_),
    .Y(_14509_));
 OA211x2_ASAP7_75t_R _31847_ (.A1(_14506_),
    .A2(_13488_),
    .B(_14508_),
    .C(_14509_),
    .Y(_14510_));
 OR3x1_ASAP7_75t_R _31848_ (.A(_14353_),
    .B(_14505_),
    .C(_14510_),
    .Y(_14511_));
 AND3x1_ASAP7_75t_R _31849_ (.A(_14488_),
    .B(_14500_),
    .C(_14511_),
    .Y(_14512_));
 NAND2x1_ASAP7_75t_R _31850_ (.A(_13189_),
    .B(_00429_),
    .Y(_14513_));
 OA211x2_ASAP7_75t_R _31851_ (.A1(_14496_),
    .A2(_13505_),
    .B(_14513_),
    .C(_14504_),
    .Y(_14514_));
 BUFx12f_ASAP7_75t_R _31852_ (.A(_13095_),
    .Y(_14515_));
 BUFx12f_ASAP7_75t_R _31853_ (.A(_14515_),
    .Y(_14516_));
 BUFx12f_ASAP7_75t_R _31854_ (.A(_13145_),
    .Y(_14517_));
 NAND2x1_ASAP7_75t_R _31855_ (.A(_14517_),
    .B(_00428_),
    .Y(_14518_));
 OA211x2_ASAP7_75t_R _31856_ (.A1(_14516_),
    .A2(_13508_),
    .B(_14518_),
    .C(_14509_),
    .Y(_14519_));
 OR3x1_ASAP7_75t_R _31857_ (.A(_14469_),
    .B(_14514_),
    .C(_14519_),
    .Y(_14520_));
 NAND2x1_ASAP7_75t_R _31858_ (.A(_14507_),
    .B(_00437_),
    .Y(_14521_));
 OA211x2_ASAP7_75t_R _31859_ (.A1(_14506_),
    .A2(_13523_),
    .B(_14521_),
    .C(_14504_),
    .Y(_14522_));
 NAND2x1_ASAP7_75t_R _31860_ (.A(_14517_),
    .B(_00436_),
    .Y(_14523_));
 OA211x2_ASAP7_75t_R _31861_ (.A1(_14516_),
    .A2(_13526_),
    .B(_14523_),
    .C(_14509_),
    .Y(_14524_));
 OR3x1_ASAP7_75t_R _31862_ (.A(_14353_),
    .B(_14522_),
    .C(_14524_),
    .Y(_14525_));
 AND3x1_ASAP7_75t_R _31863_ (.A(_14305_),
    .B(_14520_),
    .C(_14525_),
    .Y(_14526_));
 OR3x2_ASAP7_75t_R _31864_ (.A(_14487_),
    .B(_14512_),
    .C(_14526_),
    .Y(_14527_));
 NAND2x2_ASAP7_75t_R _31865_ (.A(_14486_),
    .B(_14527_),
    .Y(_14528_));
 OR3x1_ASAP7_75t_R _31866_ (.A(_14278_),
    .B(_13228_),
    .C(_14275_),
    .Y(_14529_));
 OA22x2_ASAP7_75t_R _31867_ (.A1(_01466_),
    .A2(_13260_),
    .B1(_14380_),
    .B2(_01496_),
    .Y(_14530_));
 OA211x2_ASAP7_75t_R _31868_ (.A1(_13273_),
    .A2(_14529_),
    .B(_14530_),
    .C(_13267_),
    .Y(_14531_));
 AOI21x1_ASAP7_75t_R _31869_ (.A1(_14446_),
    .A2(_14528_),
    .B(_14531_),
    .Y(_18558_));
 INVx3_ASAP7_75t_R _31870_ (.A(_18558_),
    .Y(_18560_));
 INVx1_ASAP7_75t_R _31871_ (.A(_02178_),
    .Y(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ));
 INVx1_ASAP7_75t_R _31872_ (.A(_02115_),
    .Y(\cs_registers_i.mhpmcounter[1857] ));
 OR3x2_ASAP7_75t_R _31873_ (.A(_13261_),
    .B(_14122_),
    .C(_14116_),
    .Y(_14532_));
 BUFx12f_ASAP7_75t_R _31874_ (.A(_13287_),
    .Y(_14533_));
 BUFx12f_ASAP7_75t_R _31875_ (.A(_14533_),
    .Y(_14534_));
 OR3x1_ASAP7_75t_R _31876_ (.A(_14534_),
    .B(_14202_),
    .C(_14273_),
    .Y(_14535_));
 AOI21x1_ASAP7_75t_R _31877_ (.A1(_14532_),
    .A2(_14535_),
    .B(_14274_),
    .Y(_14536_));
 AND3x1_ASAP7_75t_R _31878_ (.A(_14274_),
    .B(_14122_),
    .C(_14273_),
    .Y(_14537_));
 AND2x4_ASAP7_75t_R _31879_ (.A(_14098_),
    .B(_14101_),
    .Y(_14538_));
 AND5x2_ASAP7_75t_R _31880_ (.A(_13277_),
    .B(_13243_),
    .C(_13220_),
    .D(_13248_),
    .E(_13240_),
    .Y(_14539_));
 OA211x2_ASAP7_75t_R _31881_ (.A1(_14536_),
    .A2(_14537_),
    .B(_14538_),
    .C(_14539_),
    .Y(_14540_));
 BUFx12f_ASAP7_75t_R _31882_ (.A(_13262_),
    .Y(_14541_));
 AND2x4_ASAP7_75t_R _31883_ (.A(_13234_),
    .B(_13235_),
    .Y(_14542_));
 AND4x1_ASAP7_75t_R _31884_ (.A(_13280_),
    .B(_13248_),
    .C(_13240_),
    .D(_13264_),
    .Y(_14543_));
 AND2x6_ASAP7_75t_R _31885_ (.A(_14542_),
    .B(_14543_),
    .Y(_14544_));
 AND2x2_ASAP7_75t_R _31886_ (.A(_13222_),
    .B(_13242_),
    .Y(_14545_));
 AND5x2_ASAP7_75t_R _31887_ (.A(_13220_),
    .B(_13263_),
    .C(_13217_),
    .D(_13240_),
    .E(_14545_),
    .Y(_14546_));
 AND4x1_ASAP7_75t_R _31888_ (.A(_14099_),
    .B(_01512_),
    .C(_01513_),
    .D(_13909_),
    .Y(_14547_));
 AND4x1_ASAP7_75t_R _31889_ (.A(_14122_),
    .B(_14117_),
    .C(_14546_),
    .D(_14547_),
    .Y(_14548_));
 OA22x2_ASAP7_75t_R _31890_ (.A1(_14541_),
    .A2(_14273_),
    .B1(_14544_),
    .B2(_14548_),
    .Y(_14549_));
 AND3x1_ASAP7_75t_R _31891_ (.A(_14274_),
    .B(_14273_),
    .C(_14546_),
    .Y(_14550_));
 AO21x1_ASAP7_75t_R _31892_ (.A1(_14112_),
    .A2(_14549_),
    .B(_14550_),
    .Y(_14551_));
 NOR2x1_ASAP7_75t_R _31893_ (.A(_14540_),
    .B(_14551_),
    .Y(_18001_));
 INVx1_ASAP7_75t_R _31894_ (.A(_18001_),
    .Y(_18002_));
 NOR2x1_ASAP7_75t_R _31895_ (.A(_14272_),
    .B(_13422_),
    .Y(_14552_));
 AO21x1_ASAP7_75t_R _31896_ (.A1(_14541_),
    .A2(_14272_),
    .B(_14552_),
    .Y(_14553_));
 AND3x1_ASAP7_75t_R _31897_ (.A(_14122_),
    .B(_13831_),
    .C(_14553_),
    .Y(_14554_));
 NAND2x1_ASAP7_75t_R _31898_ (.A(_14098_),
    .B(_14101_),
    .Y(_14555_));
 NAND2x1_ASAP7_75t_R _31899_ (.A(_14122_),
    .B(_14117_),
    .Y(_14556_));
 OR4x1_ASAP7_75t_R _31900_ (.A(_13287_),
    .B(_13227_),
    .C(_14555_),
    .D(_14556_),
    .Y(_14557_));
 AO21x1_ASAP7_75t_R _31901_ (.A1(_13287_),
    .A2(_14202_),
    .B(_13421_),
    .Y(_14558_));
 NAND3x1_ASAP7_75t_R _31902_ (.A(_13227_),
    .B(_14098_),
    .C(_14101_),
    .Y(_14559_));
 AOI21x1_ASAP7_75t_R _31903_ (.A1(_14532_),
    .A2(_14558_),
    .B(_14559_),
    .Y(_14560_));
 AND3x1_ASAP7_75t_R _31904_ (.A(_13837_),
    .B(_01510_),
    .C(_13909_),
    .Y(_14561_));
 AND2x4_ASAP7_75t_R _31905_ (.A(_14101_),
    .B(_14561_),
    .Y(_14562_));
 OA21x2_ASAP7_75t_R _31906_ (.A1(_13832_),
    .A2(_14272_),
    .B(_14562_),
    .Y(_14563_));
 NOR2x1_ASAP7_75t_R _31907_ (.A(_14560_),
    .B(_14563_),
    .Y(_14564_));
 AO221x1_ASAP7_75t_R _31908_ (.A1(_14547_),
    .A2(_14554_),
    .B1(_14557_),
    .B2(_14564_),
    .C(_13838_),
    .Y(_14565_));
 NAND2x1_ASAP7_75t_R _31909_ (.A(_14542_),
    .B(_14543_),
    .Y(_14566_));
 OR3x1_ASAP7_75t_R _31910_ (.A(_14534_),
    .B(_14125_),
    .C(_14547_),
    .Y(_14567_));
 OAI21x1_ASAP7_75t_R _31911_ (.A1(_14117_),
    .A2(_14566_),
    .B(_14567_),
    .Y(_14568_));
 AO21x1_ASAP7_75t_R _31912_ (.A1(_14273_),
    .A2(_14546_),
    .B(_14534_),
    .Y(_14569_));
 AO221x1_ASAP7_75t_R _31913_ (.A1(_14117_),
    .A2(_14546_),
    .B1(_14544_),
    .B2(_14274_),
    .C(_14541_),
    .Y(_14570_));
 AND2x2_ASAP7_75t_R _31914_ (.A(_13277_),
    .B(_13282_),
    .Y(_14571_));
 OA21x2_ASAP7_75t_R _31915_ (.A1(_13263_),
    .A2(_14124_),
    .B(_13264_),
    .Y(_14572_));
 AND2x2_ASAP7_75t_R _31916_ (.A(_13246_),
    .B(_14545_),
    .Y(_14573_));
 OA21x2_ASAP7_75t_R _31917_ (.A1(_14572_),
    .A2(_14573_),
    .B(_13280_),
    .Y(_14574_));
 AND2x2_ASAP7_75t_R _31918_ (.A(_13240_),
    .B(_13290_),
    .Y(_14575_));
 OAI21x1_ASAP7_75t_R _31919_ (.A1(_14571_),
    .A2(_14574_),
    .B(_14575_),
    .Y(_14576_));
 AO21x1_ASAP7_75t_R _31920_ (.A1(_14569_),
    .A2(_14570_),
    .B(_14576_),
    .Y(_14577_));
 AO221x1_ASAP7_75t_R _31921_ (.A1(_14137_),
    .A2(_14544_),
    .B1(_14568_),
    .B2(_14112_),
    .C(_14577_),
    .Y(_14578_));
 AO21x2_ASAP7_75t_R _31922_ (.A1(_14539_),
    .A2(_14565_),
    .B(_14578_),
    .Y(_18000_));
 INVx1_ASAP7_75t_R _31923_ (.A(_18000_),
    .Y(_18004_));
 NOR2x1_ASAP7_75t_R _31924_ (.A(_00751_),
    .B(_14544_),
    .Y(_14579_));
 OA21x2_ASAP7_75t_R _31925_ (.A1(_14571_),
    .A2(_14574_),
    .B(_14575_),
    .Y(_14580_));
 OR5x2_ASAP7_75t_R _31926_ (.A(_13244_),
    .B(_13242_),
    .C(_13218_),
    .D(_13276_),
    .E(_13285_),
    .Y(_14581_));
 AND3x1_ASAP7_75t_R _31927_ (.A(_14121_),
    .B(_01510_),
    .C(_14116_),
    .Y(_14582_));
 AND3x1_ASAP7_75t_R _31928_ (.A(_13262_),
    .B(_14538_),
    .C(_14582_),
    .Y(_14583_));
 AO21x1_ASAP7_75t_R _31929_ (.A1(_13287_),
    .A2(_14121_),
    .B(_14117_),
    .Y(_14584_));
 NAND2x1_ASAP7_75t_R _31930_ (.A(_14101_),
    .B(_14561_),
    .Y(_14585_));
 AOI21x1_ASAP7_75t_R _31931_ (.A1(_13831_),
    .A2(_14584_),
    .B(_14585_),
    .Y(_14586_));
 OR4x1_ASAP7_75t_R _31932_ (.A(_14560_),
    .B(_14581_),
    .C(_14583_),
    .D(_14586_),
    .Y(_14587_));
 NAND2x2_ASAP7_75t_R _31933_ (.A(_13287_),
    .B(_14121_),
    .Y(_14588_));
 OR4x1_ASAP7_75t_R _31934_ (.A(_13226_),
    .B(_14121_),
    .C(_13421_),
    .D(_14547_),
    .Y(_14589_));
 AO21x2_ASAP7_75t_R _31935_ (.A1(_14588_),
    .A2(_14589_),
    .B(_14125_),
    .Y(_14590_));
 NAND2x2_ASAP7_75t_R _31936_ (.A(_13234_),
    .B(_13235_),
    .Y(_14591_));
 OR4x1_ASAP7_75t_R _31937_ (.A(_13220_),
    .B(_13276_),
    .C(_13285_),
    .D(_13223_),
    .Y(_14592_));
 OR3x1_ASAP7_75t_R _31938_ (.A(_14112_),
    .B(_14591_),
    .C(_14592_),
    .Y(_14593_));
 NAND2x1_ASAP7_75t_R _31939_ (.A(_14546_),
    .B(_14137_),
    .Y(_14594_));
 XOR2x2_ASAP7_75t_R _31940_ (.A(_13226_),
    .B(_13421_),
    .Y(_14595_));
 OR3x1_ASAP7_75t_R _31941_ (.A(_14591_),
    .B(_14592_),
    .C(_14595_),
    .Y(_14596_));
 OR5x1_ASAP7_75t_R _31942_ (.A(_13287_),
    .B(_14112_),
    .C(_14555_),
    .D(_14581_),
    .E(_14556_),
    .Y(_14597_));
 AND5x1_ASAP7_75t_R _31943_ (.A(_14590_),
    .B(_14593_),
    .C(_14594_),
    .D(_14596_),
    .E(_14597_),
    .Y(_14598_));
 AO32x2_ASAP7_75t_R _31944_ (.A1(_13909_),
    .A2(_14101_),
    .A3(_14546_),
    .B1(_14539_),
    .B2(_14123_),
    .Y(_14599_));
 AND3x1_ASAP7_75t_R _31945_ (.A(_13287_),
    .B(_13234_),
    .C(_13235_),
    .Y(_14600_));
 AO22x2_ASAP7_75t_R _31946_ (.A1(_13287_),
    .A2(_14546_),
    .B1(_14543_),
    .B2(_14600_),
    .Y(_14601_));
 AND2x6_ASAP7_75t_R _31947_ (.A(_14112_),
    .B(_14117_),
    .Y(_14602_));
 OAI21x1_ASAP7_75t_R _31948_ (.A1(_14599_),
    .A2(_14601_),
    .B(_14602_),
    .Y(_14603_));
 AND4x1_ASAP7_75t_R _31949_ (.A(_14580_),
    .B(_14587_),
    .C(_14598_),
    .D(_14603_),
    .Y(_14604_));
 AND3x4_ASAP7_75t_R _31950_ (.A(_14542_),
    .B(_14588_),
    .C(_14543_),
    .Y(_14605_));
 INVx1_ASAP7_75t_R _31951_ (.A(_02221_),
    .Y(_14606_));
 AO21x1_ASAP7_75t_R _31952_ (.A1(_14532_),
    .A2(_14558_),
    .B(_14559_),
    .Y(_14607_));
 AO21x1_ASAP7_75t_R _31953_ (.A1(_13831_),
    .A2(_14584_),
    .B(_14585_),
    .Y(_14608_));
 AND4x1_ASAP7_75t_R _31954_ (.A(_14607_),
    .B(_14539_),
    .C(_14557_),
    .D(_14608_),
    .Y(_14609_));
 AOI21x1_ASAP7_75t_R _31955_ (.A1(_14588_),
    .A2(_14589_),
    .B(_14125_),
    .Y(_14610_));
 AO32x1_ASAP7_75t_R _31956_ (.A1(_14121_),
    .A2(_14542_),
    .A3(_14543_),
    .B1(_14137_),
    .B2(_14546_),
    .Y(_14611_));
 NOR3x1_ASAP7_75t_R _31957_ (.A(_14591_),
    .B(_14592_),
    .C(_14595_),
    .Y(_14612_));
 AND4x1_ASAP7_75t_R _31958_ (.A(_13262_),
    .B(_14538_),
    .C(_14539_),
    .D(_14582_),
    .Y(_14613_));
 OR4x1_ASAP7_75t_R _31959_ (.A(_14610_),
    .B(_14611_),
    .C(_14612_),
    .D(_14613_),
    .Y(_14614_));
 OA21x2_ASAP7_75t_R _31960_ (.A1(_14599_),
    .A2(_14601_),
    .B(_14602_),
    .Y(_14615_));
 OR5x1_ASAP7_75t_R _31961_ (.A(_14606_),
    .B(_14576_),
    .C(_14609_),
    .D(_14614_),
    .E(_14615_),
    .Y(_14616_));
 OAI21x1_ASAP7_75t_R _31962_ (.A1(_14588_),
    .A2(_14566_),
    .B(_14590_),
    .Y(_14617_));
 OA31x2_ASAP7_75t_R _31963_ (.A1(_14576_),
    .A2(_14609_),
    .A3(_14617_),
    .B1(_02220_),
    .Y(_14618_));
 AOI221x1_ASAP7_75t_R _31964_ (.A1(_14579_),
    .A2(_14604_),
    .B1(_14605_),
    .B2(_14616_),
    .C(_14618_),
    .Y(_14619_));
 OR3x2_ASAP7_75t_R _31965_ (.A(_13831_),
    .B(_14585_),
    .C(_14581_),
    .Y(_14620_));
 AND2x6_ASAP7_75t_R _31966_ (.A(_14619_),
    .B(_14620_),
    .Y(_14621_));
 BUFx6f_ASAP7_75t_R _31967_ (.A(_14621_),
    .Y(_16998_));
 AND3x4_ASAP7_75t_R _31968_ (.A(_13832_),
    .B(_14562_),
    .C(_14539_),
    .Y(_14622_));
 BUFx12f_ASAP7_75t_R _31969_ (.A(_14622_),
    .Y(_14623_));
 BUFx12f_ASAP7_75t_R _31970_ (.A(_14623_),
    .Y(_14624_));
 BUFx6f_ASAP7_75t_R _31971_ (.A(_14624_),
    .Y(_14625_));
 OR3x2_ASAP7_75t_R _31972_ (.A(_13831_),
    .B(_14585_),
    .C(_14581_),
    .Y(_14626_));
 BUFx6f_ASAP7_75t_R _31973_ (.A(_14626_),
    .Y(_14627_));
 AND2x6_ASAP7_75t_R _31974_ (.A(_01798_),
    .B(_02198_),
    .Y(_14628_));
 BUFx6f_ASAP7_75t_R _31975_ (.A(_14628_),
    .Y(_14629_));
 OR3x1_ASAP7_75t_R _31976_ (.A(_00062_),
    .B(_14627_),
    .C(_14629_),
    .Y(_14630_));
 OA21x2_ASAP7_75t_R _31977_ (.A1(_18556_),
    .A2(_14625_),
    .B(_14630_),
    .Y(_16997_));
 INVx1_ASAP7_75t_R _31978_ (.A(_16997_),
    .Y(_18008_));
 AO221x1_ASAP7_75t_R _31979_ (.A1(_14579_),
    .A2(_14604_),
    .B1(_14605_),
    .B2(_14616_),
    .C(_14618_),
    .Y(_14631_));
 BUFx6f_ASAP7_75t_R _31980_ (.A(_14631_),
    .Y(_14632_));
 BUFx6f_ASAP7_75t_R _31981_ (.A(_00752_),
    .Y(_14633_));
 BUFx12f_ASAP7_75t_R _31982_ (.A(_14633_),
    .Y(_14634_));
 AND2x6_ASAP7_75t_R _31983_ (.A(_14416_),
    .B(_14443_),
    .Y(_14635_));
 BUFx6f_ASAP7_75t_R _31984_ (.A(_00753_),
    .Y(_14636_));
 INVx1_ASAP7_75t_R _31985_ (.A(_00062_),
    .Y(_14637_));
 INVx1_ASAP7_75t_R _31986_ (.A(_01756_),
    .Y(_14638_));
 INVx3_ASAP7_75t_R _31987_ (.A(_00753_),
    .Y(_14639_));
 INVx5_ASAP7_75t_R _31988_ (.A(_14633_),
    .Y(_14640_));
 NAND2x2_ASAP7_75t_R _31989_ (.A(_01798_),
    .B(_02198_),
    .Y(_14641_));
 OR3x2_ASAP7_75t_R _31990_ (.A(_14639_),
    .B(_14640_),
    .C(_14641_),
    .Y(_14642_));
 OA222x2_ASAP7_75t_R _31991_ (.A1(_14636_),
    .A2(_14637_),
    .B1(_14638_),
    .B2(_14628_),
    .C1(_14642_),
    .C2(_13420_),
    .Y(_14643_));
 OAI21x1_ASAP7_75t_R _31992_ (.A1(_14634_),
    .A2(_14635_),
    .B(_14643_),
    .Y(_14644_));
 AO22x1_ASAP7_75t_R _31993_ (.A1(_18553_),
    .A2(_14632_),
    .B1(_14624_),
    .B2(_14644_),
    .Y(_14645_));
 AO21x1_ASAP7_75t_R _31994_ (.A1(_18555_),
    .A2(_14621_),
    .B(_14645_),
    .Y(_18007_));
 INVx1_ASAP7_75t_R _31995_ (.A(_18007_),
    .Y(_16996_));
 BUFx12f_ASAP7_75t_R _31996_ (.A(_14624_),
    .Y(_14646_));
 BUFx12f_ASAP7_75t_R _31997_ (.A(_14646_),
    .Y(_14647_));
 BUFx6f_ASAP7_75t_R _31998_ (.A(_14627_),
    .Y(_14648_));
 BUFx6f_ASAP7_75t_R _31999_ (.A(_14628_),
    .Y(_14649_));
 BUFx6f_ASAP7_75t_R _32000_ (.A(_14649_),
    .Y(_14650_));
 OR3x1_ASAP7_75t_R _32001_ (.A(_00097_),
    .B(_14648_),
    .C(_14650_),
    .Y(_14651_));
 OAI21x1_ASAP7_75t_R _32002_ (.A1(_18560_),
    .A2(_14647_),
    .B(_14651_),
    .Y(_18010_));
 XNOR2x1_ASAP7_75t_R _32003_ (.B(_00755_),
    .Y(\alu_adder_result_ex[1] ),
    .A(_00757_));
 INVx8_ASAP7_75t_R _32004_ (.A(\alu_adder_result_ex[1] ),
    .Y(_18712_));
 INVx2_ASAP7_75t_R _32005_ (.A(_00016_),
    .Y(\cs_registers_i.pc_id_i[2] ));
 BUFx12f_ASAP7_75t_R _32006_ (.A(_14314_),
    .Y(_14652_));
 BUFx12f_ASAP7_75t_R _32007_ (.A(_14300_),
    .Y(_14653_));
 NAND2x1_ASAP7_75t_R _32008_ (.A(_14653_),
    .B(_01794_),
    .Y(_14654_));
 NAND2x1_ASAP7_75t_R _32009_ (.A(_13091_),
    .B(_00446_),
    .Y(_14655_));
 AO32x1_ASAP7_75t_R _32010_ (.A1(_14652_),
    .A2(_14654_),
    .A3(_14655_),
    .B1(_13554_),
    .B2(_14449_),
    .Y(_14656_));
 INVx1_ASAP7_75t_R _32011_ (.A(_00454_),
    .Y(_14657_));
 NAND2x1_ASAP7_75t_R _32012_ (.A(_13188_),
    .B(_00452_),
    .Y(_14658_));
 OA211x2_ASAP7_75t_R _32013_ (.A1(_13192_),
    .A2(_14657_),
    .B(_14658_),
    .C(_14295_),
    .Y(_14659_));
 INVx1_ASAP7_75t_R _32014_ (.A(_00453_),
    .Y(_14660_));
 NAND2x1_ASAP7_75t_R _32015_ (.A(_13188_),
    .B(_00451_),
    .Y(_14661_));
 OA211x2_ASAP7_75t_R _32016_ (.A1(_13192_),
    .A2(_14660_),
    .B(_14661_),
    .C(_13148_),
    .Y(_14662_));
 OR3x1_ASAP7_75t_R _32017_ (.A(_13104_),
    .B(_14659_),
    .C(_14662_),
    .Y(_14663_));
 OA211x2_ASAP7_75t_R _32018_ (.A1(_14469_),
    .A2(_14656_),
    .B(_14663_),
    .C(_13124_),
    .Y(_14664_));
 NAND2x1_ASAP7_75t_R _32019_ (.A(_13136_),
    .B(_00448_),
    .Y(_14665_));
 OA211x2_ASAP7_75t_R _32020_ (.A1(_13196_),
    .A2(_13559_),
    .B(_14665_),
    .C(_14314_),
    .Y(_14666_));
 BUFx12f_ASAP7_75t_R _32021_ (.A(_13135_),
    .Y(_14667_));
 NAND2x1_ASAP7_75t_R _32022_ (.A(_14667_),
    .B(_00447_),
    .Y(_14668_));
 OA211x2_ASAP7_75t_R _32023_ (.A1(_13165_),
    .A2(_13556_),
    .B(_14668_),
    .C(_14322_),
    .Y(_14669_));
 OR3x2_ASAP7_75t_R _32024_ (.A(_13130_),
    .B(_14666_),
    .C(_14669_),
    .Y(_14670_));
 NAND2x1_ASAP7_75t_R _32025_ (.A(_14667_),
    .B(_00456_),
    .Y(_14671_));
 OA211x2_ASAP7_75t_R _32026_ (.A1(_13196_),
    .A2(_13567_),
    .B(_14671_),
    .C(_14314_),
    .Y(_14672_));
 NAND2x1_ASAP7_75t_R _32027_ (.A(_14667_),
    .B(_00455_),
    .Y(_14673_));
 OA211x2_ASAP7_75t_R _32028_ (.A1(_13165_),
    .A2(_13548_),
    .B(_14673_),
    .C(_14322_),
    .Y(_14674_));
 OR3x1_ASAP7_75t_R _32029_ (.A(_14326_),
    .B(_14672_),
    .C(_14674_),
    .Y(_14675_));
 AND3x1_ASAP7_75t_R _32030_ (.A(_13128_),
    .B(_14670_),
    .C(_14675_),
    .Y(_14676_));
 OR3x2_ASAP7_75t_R _32031_ (.A(_13081_),
    .B(_14664_),
    .C(_14676_),
    .Y(_14677_));
 BUFx12f_ASAP7_75t_R _32032_ (.A(_13109_),
    .Y(_14678_));
 NAND2x1_ASAP7_75t_R _32033_ (.A(_13136_),
    .B(_00464_),
    .Y(_14679_));
 OA211x2_ASAP7_75t_R _32034_ (.A1(_14678_),
    .A2(_13571_),
    .B(_14679_),
    .C(_14314_),
    .Y(_14680_));
 NAND2x1_ASAP7_75t_R _32035_ (.A(_13136_),
    .B(_00463_),
    .Y(_14681_));
 OA211x2_ASAP7_75t_R _32036_ (.A1(_13196_),
    .A2(_13574_),
    .B(_14681_),
    .C(_14322_),
    .Y(_14682_));
 OR3x1_ASAP7_75t_R _32037_ (.A(_13130_),
    .B(_14680_),
    .C(_14682_),
    .Y(_14683_));
 NAND2x1_ASAP7_75t_R _32038_ (.A(_13136_),
    .B(_00472_),
    .Y(_14684_));
 OA211x2_ASAP7_75t_R _32039_ (.A1(_14678_),
    .A2(_13588_),
    .B(_14684_),
    .C(_14314_),
    .Y(_14685_));
 NAND2x1_ASAP7_75t_R _32040_ (.A(_14667_),
    .B(_00471_),
    .Y(_14686_));
 OA211x2_ASAP7_75t_R _32041_ (.A1(_13196_),
    .A2(_13585_),
    .B(_14686_),
    .C(_14322_),
    .Y(_14687_));
 OR3x1_ASAP7_75t_R _32042_ (.A(_14326_),
    .B(_14685_),
    .C(_14687_),
    .Y(_14688_));
 AND3x1_ASAP7_75t_R _32043_ (.A(_13128_),
    .B(_14683_),
    .C(_14688_),
    .Y(_14689_));
 NAND2x1_ASAP7_75t_R _32044_ (.A(_13136_),
    .B(_00460_),
    .Y(_14690_));
 OA211x2_ASAP7_75t_R _32045_ (.A1(_13196_),
    .A2(_13578_),
    .B(_14690_),
    .C(_14314_),
    .Y(_14691_));
 NAND2x1_ASAP7_75t_R _32046_ (.A(_14667_),
    .B(_00459_),
    .Y(_14692_));
 OA211x2_ASAP7_75t_R _32047_ (.A1(_13165_),
    .A2(_13581_),
    .B(_14692_),
    .C(_14322_),
    .Y(_14693_));
 OR3x1_ASAP7_75t_R _32048_ (.A(_13130_),
    .B(_14691_),
    .C(_14693_),
    .Y(_14694_));
 NAND2x1_ASAP7_75t_R _32049_ (.A(_14667_),
    .B(_00468_),
    .Y(_14695_));
 OA211x2_ASAP7_75t_R _32050_ (.A1(_13196_),
    .A2(_13595_),
    .B(_14695_),
    .C(_14314_),
    .Y(_14696_));
 BUFx12f_ASAP7_75t_R _32051_ (.A(_13109_),
    .Y(_14697_));
 NAND2x1_ASAP7_75t_R _32052_ (.A(_14667_),
    .B(_00467_),
    .Y(_14698_));
 OA211x2_ASAP7_75t_R _32053_ (.A1(_14697_),
    .A2(_13592_),
    .B(_14698_),
    .C(_14322_),
    .Y(_14699_));
 OR3x1_ASAP7_75t_R _32054_ (.A(_14326_),
    .B(_14696_),
    .C(_14699_),
    .Y(_14700_));
 AND3x1_ASAP7_75t_R _32055_ (.A(_14428_),
    .B(_14694_),
    .C(_14700_),
    .Y(_14701_));
 OR3x2_ASAP7_75t_R _32056_ (.A(_13163_),
    .B(_14689_),
    .C(_14701_),
    .Y(_14702_));
 AND2x6_ASAP7_75t_R _32057_ (.A(_14677_),
    .B(_14702_),
    .Y(_14703_));
 AND3x1_ASAP7_75t_R _32058_ (.A(_14307_),
    .B(_14119_),
    .C(_13265_),
    .Y(_14704_));
 OAI22x1_ASAP7_75t_R _32059_ (.A1(_01455_),
    .A2(_13260_),
    .B1(_14380_),
    .B2(_00016_),
    .Y(_14705_));
 AO211x2_ASAP7_75t_R _32060_ (.A1(_14384_),
    .A2(_14704_),
    .B(_14705_),
    .C(_14446_),
    .Y(_14706_));
 OA21x2_ASAP7_75t_R _32061_ (.A1(_14377_),
    .A2(_14703_),
    .B(_14706_),
    .Y(_14707_));
 BUFx6f_ASAP7_75t_R _32062_ (.A(_14707_),
    .Y(_18562_));
 INVx2_ASAP7_75t_R _32063_ (.A(_18562_),
    .Y(_18564_));
 OR3x1_ASAP7_75t_R _32064_ (.A(_00100_),
    .B(_14648_),
    .C(_14650_),
    .Y(_14708_));
 OAI21x1_ASAP7_75t_R _32065_ (.A1(_14647_),
    .A2(_18564_),
    .B(_14708_),
    .Y(_18012_));
 BUFx6f_ASAP7_75t_R _32066_ (.A(_13267_),
    .Y(_14709_));
 BUFx12f_ASAP7_75t_R _32067_ (.A(_13120_),
    .Y(_14710_));
 BUFx12f_ASAP7_75t_R _32068_ (.A(_14678_),
    .Y(_14711_));
 NOR2x1_ASAP7_75t_R _32069_ (.A(_14312_),
    .B(_00487_),
    .Y(_14712_));
 AO21x1_ASAP7_75t_R _32070_ (.A1(_14711_),
    .A2(_13633_),
    .B(_14712_),
    .Y(_14713_));
 NAND2x1_ASAP7_75t_R _32071_ (.A(_14310_),
    .B(_00486_),
    .Y(_14714_));
 OA211x2_ASAP7_75t_R _32072_ (.A1(_14474_),
    .A2(_13636_),
    .B(_14714_),
    .C(_14472_),
    .Y(_14715_));
 AO21x1_ASAP7_75t_R _32073_ (.A1(_14710_),
    .A2(_14713_),
    .B(_14715_),
    .Y(_14716_));
 BUFx12f_ASAP7_75t_R _32074_ (.A(_14460_),
    .Y(_14717_));
 NAND2x1_ASAP7_75t_R _32075_ (.A(_14678_),
    .B(_00478_),
    .Y(_14718_));
 OA211x2_ASAP7_75t_R _32076_ (.A1(_14717_),
    .A2(_13676_),
    .B(_14718_),
    .C(_13115_),
    .Y(_14719_));
 NAND2x1_ASAP7_75t_R _32077_ (.A(_14678_),
    .B(_00477_),
    .Y(_14720_));
 OA211x2_ASAP7_75t_R _32078_ (.A1(_13097_),
    .A2(_13679_),
    .B(_14720_),
    .C(_13120_),
    .Y(_14721_));
 OR3x1_ASAP7_75t_R _32079_ (.A(_13085_),
    .B(_14719_),
    .C(_14721_),
    .Y(_14722_));
 OA21x2_ASAP7_75t_R _32080_ (.A1(_13186_),
    .A2(_14716_),
    .B(_14722_),
    .Y(_14723_));
 AND2x2_ASAP7_75t_R _32081_ (.A(_14470_),
    .B(_01793_),
    .Y(_14724_));
 AO21x1_ASAP7_75t_R _32082_ (.A1(_14285_),
    .A2(_00476_),
    .B(_14724_),
    .Y(_14725_));
 OAI22x1_ASAP7_75t_R _32083_ (.A1(_00475_),
    .A2(_13102_),
    .B1(_14725_),
    .B2(_13187_),
    .Y(_14726_));
 INVx1_ASAP7_75t_R _32084_ (.A(_00484_),
    .Y(_14727_));
 NAND2x1_ASAP7_75t_R _32085_ (.A(_14515_),
    .B(_00482_),
    .Y(_14728_));
 BUFx12f_ASAP7_75t_R _32086_ (.A(_13114_),
    .Y(_14729_));
 OA211x2_ASAP7_75t_R _32087_ (.A1(_14277_),
    .A2(_14727_),
    .B(_14728_),
    .C(_14729_),
    .Y(_14730_));
 NAND2x1_ASAP7_75t_R _32088_ (.A(_14515_),
    .B(_00481_),
    .Y(_14731_));
 BUFx12f_ASAP7_75t_R _32089_ (.A(_13100_),
    .Y(_14732_));
 OA211x2_ASAP7_75t_R _32090_ (.A1(_14301_),
    .A2(_13645_),
    .B(_14731_),
    .C(_14732_),
    .Y(_14733_));
 OR3x1_ASAP7_75t_R _32091_ (.A(_13185_),
    .B(_14730_),
    .C(_14733_),
    .Y(_14734_));
 OA211x2_ASAP7_75t_R _32092_ (.A1(_14448_),
    .A2(_14726_),
    .B(_14734_),
    .C(_14466_),
    .Y(_14735_));
 AO21x1_ASAP7_75t_R _32093_ (.A1(_14307_),
    .A2(_14723_),
    .B(_14735_),
    .Y(_14736_));
 BUFx12f_ASAP7_75t_R _32094_ (.A(_13084_),
    .Y(_14737_));
 BUFx12f_ASAP7_75t_R _32095_ (.A(_14667_),
    .Y(_14738_));
 NAND2x1_ASAP7_75t_R _32096_ (.A(_14490_),
    .B(_00494_),
    .Y(_14739_));
 BUFx12f_ASAP7_75t_R _32097_ (.A(_13114_),
    .Y(_14740_));
 OA211x2_ASAP7_75t_R _32098_ (.A1(_14738_),
    .A2(_13627_),
    .B(_14739_),
    .C(_14740_),
    .Y(_14741_));
 NAND2x1_ASAP7_75t_R _32099_ (.A(_14490_),
    .B(_00493_),
    .Y(_14742_));
 BUFx12f_ASAP7_75t_R _32100_ (.A(_13100_),
    .Y(_14743_));
 OA211x2_ASAP7_75t_R _32101_ (.A1(_14653_),
    .A2(_13620_),
    .B(_14742_),
    .C(_14743_),
    .Y(_14744_));
 OR3x1_ASAP7_75t_R _32102_ (.A(_14737_),
    .B(_14741_),
    .C(_14744_),
    .Y(_14745_));
 NAND2x1_ASAP7_75t_R _32103_ (.A(_14490_),
    .B(_00502_),
    .Y(_14746_));
 OA211x2_ASAP7_75t_R _32104_ (.A1(_13200_),
    .A2(_13624_),
    .B(_14746_),
    .C(_14740_),
    .Y(_14747_));
 NAND2x1_ASAP7_75t_R _32105_ (.A(_13192_),
    .B(_00501_),
    .Y(_14748_));
 OA211x2_ASAP7_75t_R _32106_ (.A1(_14653_),
    .A2(_13617_),
    .B(_14748_),
    .C(_14743_),
    .Y(_14749_));
 OR3x1_ASAP7_75t_R _32107_ (.A(_14454_),
    .B(_14747_),
    .C(_14749_),
    .Y(_14750_));
 AND3x1_ASAP7_75t_R _32108_ (.A(_14468_),
    .B(_14745_),
    .C(_14750_),
    .Y(_14751_));
 BUFx12f_ASAP7_75t_R _32109_ (.A(_13199_),
    .Y(_14752_));
 NOR2x1_ASAP7_75t_R _32110_ (.A(_14752_),
    .B(_00499_),
    .Y(_14753_));
 AO21x1_ASAP7_75t_R _32111_ (.A1(_14474_),
    .A2(_13653_),
    .B(_14753_),
    .Y(_14754_));
 BUFx12f_ASAP7_75t_R _32112_ (.A(_13135_),
    .Y(_14755_));
 BUFx12f_ASAP7_75t_R _32113_ (.A(_14755_),
    .Y(_14756_));
 NAND2x1_ASAP7_75t_R _32114_ (.A(_13132_),
    .B(_00498_),
    .Y(_14757_));
 OA211x2_ASAP7_75t_R _32115_ (.A1(_14756_),
    .A2(_13656_),
    .B(_14757_),
    .C(_14458_),
    .Y(_14758_));
 AO21x1_ASAP7_75t_R _32116_ (.A1(_14710_),
    .A2(_14754_),
    .B(_14758_),
    .Y(_14759_));
 BUFx12f_ASAP7_75t_R _32117_ (.A(_13135_),
    .Y(_14760_));
 NAND2x1_ASAP7_75t_R _32118_ (.A(_14760_),
    .B(_00490_),
    .Y(_14761_));
 BUFx12f_ASAP7_75t_R _32119_ (.A(_13114_),
    .Y(_14762_));
 OA211x2_ASAP7_75t_R _32120_ (.A1(_14470_),
    .A2(_13660_),
    .B(_14761_),
    .C(_14762_),
    .Y(_14763_));
 NAND2x1_ASAP7_75t_R _32121_ (.A(_14760_),
    .B(_00489_),
    .Y(_14764_));
 BUFx12f_ASAP7_75t_R _32122_ (.A(_13087_),
    .Y(_14765_));
 OA211x2_ASAP7_75t_R _32123_ (.A1(_14310_),
    .A2(_13663_),
    .B(_14764_),
    .C(_14765_),
    .Y(_14766_));
 OR3x1_ASAP7_75t_R _32124_ (.A(_14308_),
    .B(_14763_),
    .C(_14766_),
    .Y(_14767_));
 OA211x2_ASAP7_75t_R _32125_ (.A1(_13186_),
    .A2(_14759_),
    .B(_14767_),
    .C(_14428_),
    .Y(_14768_));
 OR3x1_ASAP7_75t_R _32126_ (.A(_14487_),
    .B(_14751_),
    .C(_14768_),
    .Y(_14769_));
 OA21x2_ASAP7_75t_R _32127_ (.A1(_14281_),
    .A2(_14736_),
    .B(_14769_),
    .Y(_14770_));
 AND3x1_ASAP7_75t_R _32128_ (.A(_14283_),
    .B(_14119_),
    .C(_13265_),
    .Y(_14771_));
 BUFx6f_ASAP7_75t_R _32129_ (.A(_14380_),
    .Y(_14772_));
 BUFx6f_ASAP7_75t_R _32130_ (.A(_00018_),
    .Y(_14773_));
 OAI22x1_ASAP7_75t_R _32131_ (.A1(_01452_),
    .A2(_13260_),
    .B1(_14772_),
    .B2(_14773_),
    .Y(_14774_));
 AO211x2_ASAP7_75t_R _32132_ (.A1(_14384_),
    .A2(_14771_),
    .B(_14774_),
    .C(_14446_),
    .Y(_14775_));
 OA21x2_ASAP7_75t_R _32133_ (.A1(_14709_),
    .A2(_14770_),
    .B(_14775_),
    .Y(_14776_));
 BUFx6f_ASAP7_75t_R _32134_ (.A(_14776_),
    .Y(_18567_));
 INVx3_ASAP7_75t_R _32135_ (.A(_18567_),
    .Y(_18569_));
 OR3x1_ASAP7_75t_R _32136_ (.A(_00104_),
    .B(_14648_),
    .C(_14650_),
    .Y(_14777_));
 OAI21x1_ASAP7_75t_R _32137_ (.A1(_14647_),
    .A2(_18569_),
    .B(_14777_),
    .Y(_18014_));
 BUFx12f_ASAP7_75t_R _32138_ (.A(_14428_),
    .Y(_14778_));
 AND2x2_ASAP7_75t_R _32139_ (.A(_14317_),
    .B(_01792_),
    .Y(_14779_));
 AO21x1_ASAP7_75t_R _32140_ (.A1(_14285_),
    .A2(_00506_),
    .B(_14779_),
    .Y(_14780_));
 OAI22x1_ASAP7_75t_R _32141_ (.A1(_00505_),
    .A2(_13101_),
    .B1(_14780_),
    .B2(_14710_),
    .Y(_14781_));
 BUFx12f_ASAP7_75t_R _32142_ (.A(_14460_),
    .Y(_14782_));
 INVx1_ASAP7_75t_R _32143_ (.A(_00514_),
    .Y(_14783_));
 NAND2x1_ASAP7_75t_R _32144_ (.A(_14437_),
    .B(_00512_),
    .Y(_14784_));
 OA211x2_ASAP7_75t_R _32145_ (.A1(_14782_),
    .A2(_14783_),
    .B(_14784_),
    .C(_14458_),
    .Y(_14785_));
 INVx1_ASAP7_75t_R _32146_ (.A(_00513_),
    .Y(_14786_));
 NAND2x1_ASAP7_75t_R _32147_ (.A(_14490_),
    .B(_00511_),
    .Y(_14787_));
 OA211x2_ASAP7_75t_R _32148_ (.A1(_14738_),
    .A2(_14786_),
    .B(_14787_),
    .C(_14743_),
    .Y(_14788_));
 OR3x1_ASAP7_75t_R _32149_ (.A(_14454_),
    .B(_14785_),
    .C(_14788_),
    .Y(_14789_));
 OA21x2_ASAP7_75t_R _32150_ (.A1(_14448_),
    .A2(_14781_),
    .B(_14789_),
    .Y(_14790_));
 INVx1_ASAP7_75t_R _32151_ (.A(_00510_),
    .Y(_14791_));
 NAND2x1_ASAP7_75t_R _32152_ (.A(_13106_),
    .B(_00508_),
    .Y(_14792_));
 OA211x2_ASAP7_75t_R _32153_ (.A1(_13146_),
    .A2(_14791_),
    .B(_14792_),
    .C(_14740_),
    .Y(_14793_));
 BUFx12f_ASAP7_75t_R _32154_ (.A(_13145_),
    .Y(_14794_));
 INVx1_ASAP7_75t_R _32155_ (.A(_00509_),
    .Y(_14795_));
 NAND2x1_ASAP7_75t_R _32156_ (.A(_13106_),
    .B(_00507_),
    .Y(_14796_));
 OA211x2_ASAP7_75t_R _32157_ (.A1(_14794_),
    .A2(_14795_),
    .B(_14796_),
    .C(_14732_),
    .Y(_14797_));
 OR3x1_ASAP7_75t_R _32158_ (.A(_14737_),
    .B(_14793_),
    .C(_14797_),
    .Y(_14798_));
 INVx1_ASAP7_75t_R _32159_ (.A(_00518_),
    .Y(_14799_));
 NAND2x1_ASAP7_75t_R _32160_ (.A(_13106_),
    .B(_00516_),
    .Y(_14800_));
 OA211x2_ASAP7_75t_R _32161_ (.A1(_13146_),
    .A2(_14799_),
    .B(_14800_),
    .C(_14740_),
    .Y(_14801_));
 NAND2x1_ASAP7_75t_R _32162_ (.A(_13106_),
    .B(_00515_),
    .Y(_14802_));
 OA211x2_ASAP7_75t_R _32163_ (.A1(_14794_),
    .A2(_13703_),
    .B(_14802_),
    .C(_14732_),
    .Y(_14803_));
 OR3x1_ASAP7_75t_R _32164_ (.A(_13185_),
    .B(_14801_),
    .C(_14803_),
    .Y(_14804_));
 AND3x1_ASAP7_75t_R _32165_ (.A(_14468_),
    .B(_14798_),
    .C(_14804_),
    .Y(_14805_));
 AO21x1_ASAP7_75t_R _32166_ (.A1(_14778_),
    .A2(_14790_),
    .B(_14805_),
    .Y(_14806_));
 BUFx12f_ASAP7_75t_R _32167_ (.A(_13128_),
    .Y(_14807_));
 BUFx12f_ASAP7_75t_R _32168_ (.A(_14755_),
    .Y(_14808_));
 INVx1_ASAP7_75t_R _32169_ (.A(_00526_),
    .Y(_14809_));
 NAND2x1_ASAP7_75t_R _32170_ (.A(_13205_),
    .B(_00524_),
    .Y(_14810_));
 OA211x2_ASAP7_75t_R _32171_ (.A1(_14808_),
    .A2(_14809_),
    .B(_14810_),
    .C(_14729_),
    .Y(_14811_));
 NAND2x1_ASAP7_75t_R _32172_ (.A(_13096_),
    .B(_00523_),
    .Y(_14812_));
 OA211x2_ASAP7_75t_R _32173_ (.A1(_14492_),
    .A2(_13729_),
    .B(_14812_),
    .C(_14765_),
    .Y(_14813_));
 OR3x1_ASAP7_75t_R _32174_ (.A(_14737_),
    .B(_14811_),
    .C(_14813_),
    .Y(_14814_));
 BUFx12f_ASAP7_75t_R _32175_ (.A(_13199_),
    .Y(_14815_));
 NAND2x1_ASAP7_75t_R _32176_ (.A(_13096_),
    .B(_00532_),
    .Y(_14816_));
 OA211x2_ASAP7_75t_R _32177_ (.A1(_14815_),
    .A2(_13739_),
    .B(_14816_),
    .C(_14729_),
    .Y(_14817_));
 INVx1_ASAP7_75t_R _32178_ (.A(_00533_),
    .Y(_14818_));
 NAND2x1_ASAP7_75t_R _32179_ (.A(_13096_),
    .B(_00531_),
    .Y(_14819_));
 OA211x2_ASAP7_75t_R _32180_ (.A1(_14502_),
    .A2(_14818_),
    .B(_14819_),
    .C(_14765_),
    .Y(_14820_));
 OR3x1_ASAP7_75t_R _32181_ (.A(_13185_),
    .B(_14817_),
    .C(_14820_),
    .Y(_14821_));
 AND3x1_ASAP7_75t_R _32182_ (.A(_14807_),
    .B(_14814_),
    .C(_14821_),
    .Y(_14822_));
 NOR2x1_ASAP7_75t_R _32183_ (.A(_14678_),
    .B(_00529_),
    .Y(_14823_));
 AO21x1_ASAP7_75t_R _32184_ (.A1(_14455_),
    .A2(_13743_),
    .B(_14823_),
    .Y(_14824_));
 NAND2x1_ASAP7_75t_R _32185_ (.A(_13205_),
    .B(_00528_),
    .Y(_14825_));
 OA211x2_ASAP7_75t_R _32186_ (.A1(_14367_),
    .A2(_13747_),
    .B(_14825_),
    .C(_14729_),
    .Y(_14826_));
 AO21x1_ASAP7_75t_R _32187_ (.A1(_13089_),
    .A2(_14824_),
    .B(_14826_),
    .Y(_14827_));
 NAND2x1_ASAP7_75t_R _32188_ (.A(_14667_),
    .B(_00520_),
    .Y(_14828_));
 OA211x2_ASAP7_75t_R _32189_ (.A1(_14697_),
    .A2(_13754_),
    .B(_14828_),
    .C(_14314_),
    .Y(_14829_));
 NAND2x1_ASAP7_75t_R _32190_ (.A(_14755_),
    .B(_00519_),
    .Y(_14830_));
 OA211x2_ASAP7_75t_R _32191_ (.A1(_13142_),
    .A2(_13757_),
    .B(_14830_),
    .C(_13173_),
    .Y(_14831_));
 OR3x1_ASAP7_75t_R _32192_ (.A(_13130_),
    .B(_14829_),
    .C(_14831_),
    .Y(_14832_));
 OA211x2_ASAP7_75t_R _32193_ (.A1(_13153_),
    .A2(_14827_),
    .B(_14832_),
    .C(_14428_),
    .Y(_14833_));
 OR3x1_ASAP7_75t_R _32194_ (.A(_14487_),
    .B(_14822_),
    .C(_14833_),
    .Y(_14834_));
 OA21x2_ASAP7_75t_R _32195_ (.A1(_14281_),
    .A2(_14806_),
    .B(_14834_),
    .Y(_14835_));
 AND3x1_ASAP7_75t_R _32196_ (.A(_14447_),
    .B(_14119_),
    .C(_13265_),
    .Y(_14836_));
 BUFx6f_ASAP7_75t_R _32197_ (.A(_01483_),
    .Y(_14837_));
 OAI22x1_ASAP7_75t_R _32198_ (.A1(_01451_),
    .A2(_13260_),
    .B1(_14380_),
    .B2(_14837_),
    .Y(_14838_));
 AO211x2_ASAP7_75t_R _32199_ (.A1(_14383_),
    .A2(_14836_),
    .B(_14838_),
    .C(_14446_),
    .Y(_14839_));
 OA21x2_ASAP7_75t_R _32200_ (.A1(_14377_),
    .A2(_14835_),
    .B(_14839_),
    .Y(_14840_));
 BUFx6f_ASAP7_75t_R _32201_ (.A(_14840_),
    .Y(_18572_));
 INVx3_ASAP7_75t_R _32202_ (.A(_18572_),
    .Y(_18574_));
 OR3x1_ASAP7_75t_R _32203_ (.A(_00109_),
    .B(_14648_),
    .C(_14650_),
    .Y(_14841_));
 OAI21x1_ASAP7_75t_R _32204_ (.A1(_14647_),
    .A2(_18574_),
    .B(_14841_),
    .Y(_18016_));
 AND2x2_ASAP7_75t_R _32205_ (.A(_14717_),
    .B(_01791_),
    .Y(_14842_));
 AO21x1_ASAP7_75t_R _32206_ (.A1(_13092_),
    .A2(_00536_),
    .B(_14842_),
    .Y(_14843_));
 OAI22x1_ASAP7_75t_R _32207_ (.A1(_00535_),
    .A2(_14284_),
    .B1(_14843_),
    .B2(_13090_),
    .Y(_14844_));
 INVx1_ASAP7_75t_R _32208_ (.A(_00544_),
    .Y(_14845_));
 NAND2x1_ASAP7_75t_R _32209_ (.A(_14517_),
    .B(_00542_),
    .Y(_14846_));
 OA211x2_ASAP7_75t_R _32210_ (.A1(_13193_),
    .A2(_14845_),
    .B(_14846_),
    .C(_14472_),
    .Y(_14847_));
 INVx1_ASAP7_75t_R _32211_ (.A(_00543_),
    .Y(_14848_));
 NAND2x1_ASAP7_75t_R _32212_ (.A(_14470_),
    .B(_00541_),
    .Y(_14849_));
 OA211x2_ASAP7_75t_R _32213_ (.A1(_14474_),
    .A2(_14848_),
    .B(_14849_),
    .C(_14476_),
    .Y(_14850_));
 OR3x1_ASAP7_75t_R _32214_ (.A(_14353_),
    .B(_14847_),
    .C(_14850_),
    .Y(_14851_));
 BUFx12f_ASAP7_75t_R _32215_ (.A(_13124_),
    .Y(_14852_));
 OA211x2_ASAP7_75t_R _32216_ (.A1(_13086_),
    .A2(_14844_),
    .B(_14851_),
    .C(_14852_),
    .Y(_14853_));
 BUFx6f_ASAP7_75t_R _32217_ (.A(_14678_),
    .Y(_14854_));
 NAND2x1_ASAP7_75t_R _32218_ (.A(_14653_),
    .B(_00538_),
    .Y(_14855_));
 BUFx12f_ASAP7_75t_R _32219_ (.A(_13139_),
    .Y(_14856_));
 OA211x2_ASAP7_75t_R _32220_ (.A1(_14854_),
    .A2(_13770_),
    .B(_14855_),
    .C(_14856_),
    .Y(_14857_));
 BUFx12f_ASAP7_75t_R _32221_ (.A(_13136_),
    .Y(_14858_));
 NAND2x1_ASAP7_75t_R _32222_ (.A(_14858_),
    .B(_00537_),
    .Y(_14859_));
 OA211x2_ASAP7_75t_R _32223_ (.A1(_13166_),
    .A2(_13774_),
    .B(_14859_),
    .C(_13174_),
    .Y(_14860_));
 OR3x1_ASAP7_75t_R _32224_ (.A(_13131_),
    .B(_14857_),
    .C(_14860_),
    .Y(_14861_));
 INVx1_ASAP7_75t_R _32225_ (.A(_00548_),
    .Y(_14862_));
 NAND2x1_ASAP7_75t_R _32226_ (.A(_14858_),
    .B(_00546_),
    .Y(_14863_));
 OA211x2_ASAP7_75t_R _32227_ (.A1(_14854_),
    .A2(_14862_),
    .B(_14863_),
    .C(_14856_),
    .Y(_14864_));
 NAND2x1_ASAP7_75t_R _32228_ (.A(_14858_),
    .B(_00545_),
    .Y(_14865_));
 OA211x2_ASAP7_75t_R _32229_ (.A1(_13166_),
    .A2(_13822_),
    .B(_14865_),
    .C(_13174_),
    .Y(_14866_));
 OR3x1_ASAP7_75t_R _32230_ (.A(_13153_),
    .B(_14864_),
    .C(_14866_),
    .Y(_14867_));
 AND3x1_ASAP7_75t_R _32231_ (.A(_13129_),
    .B(_14861_),
    .C(_14867_),
    .Y(_14868_));
 OR3x2_ASAP7_75t_R _32232_ (.A(_13082_),
    .B(_14853_),
    .C(_14868_),
    .Y(_14869_));
 NAND2x1_ASAP7_75t_R _32233_ (.A(_14653_),
    .B(_00554_),
    .Y(_14870_));
 OA211x2_ASAP7_75t_R _32234_ (.A1(_14854_),
    .A2(_13781_),
    .B(_14870_),
    .C(_14856_),
    .Y(_14871_));
 INVx1_ASAP7_75t_R _32235_ (.A(_00555_),
    .Y(_14872_));
 NAND2x1_ASAP7_75t_R _32236_ (.A(_14858_),
    .B(_00553_),
    .Y(_14873_));
 BUFx12f_ASAP7_75t_R _32237_ (.A(_13173_),
    .Y(_14874_));
 OA211x2_ASAP7_75t_R _32238_ (.A1(_14854_),
    .A2(_14872_),
    .B(_14873_),
    .C(_14874_),
    .Y(_14875_));
 OR3x1_ASAP7_75t_R _32239_ (.A(_13131_),
    .B(_14871_),
    .C(_14875_),
    .Y(_14876_));
 BUFx12f_ASAP7_75t_R _32240_ (.A(_13152_),
    .Y(_14877_));
 NAND2x1_ASAP7_75t_R _32241_ (.A(_14653_),
    .B(_00562_),
    .Y(_14878_));
 OA211x2_ASAP7_75t_R _32242_ (.A1(_14854_),
    .A2(_13804_),
    .B(_14878_),
    .C(_14856_),
    .Y(_14879_));
 NAND2x1_ASAP7_75t_R _32243_ (.A(_14858_),
    .B(_00561_),
    .Y(_14880_));
 OA211x2_ASAP7_75t_R _32244_ (.A1(_13166_),
    .A2(_13818_),
    .B(_14880_),
    .C(_14874_),
    .Y(_14881_));
 OR3x1_ASAP7_75t_R _32245_ (.A(_14877_),
    .B(_14879_),
    .C(_14881_),
    .Y(_14882_));
 AND3x1_ASAP7_75t_R _32246_ (.A(_13129_),
    .B(_14876_),
    .C(_14882_),
    .Y(_14883_));
 NOR2x1_ASAP7_75t_R _32247_ (.A(_14491_),
    .B(_00559_),
    .Y(_14884_));
 AO21x1_ASAP7_75t_R _32248_ (.A1(_13190_),
    .A2(_13815_),
    .B(_14884_),
    .Y(_14885_));
 BUFx6f_ASAP7_75t_R _32249_ (.A(_13211_),
    .Y(_14886_));
 INVx1_ASAP7_75t_R _32250_ (.A(_00560_),
    .Y(_14887_));
 BUFx12f_ASAP7_75t_R _32251_ (.A(_13136_),
    .Y(_14888_));
 NAND2x1_ASAP7_75t_R _32252_ (.A(_14888_),
    .B(_00558_),
    .Y(_14889_));
 OA211x2_ASAP7_75t_R _32253_ (.A1(_14886_),
    .A2(_14887_),
    .B(_14889_),
    .C(_14652_),
    .Y(_14890_));
 AO21x1_ASAP7_75t_R _32254_ (.A1(_13187_),
    .A2(_14885_),
    .B(_14890_),
    .Y(_14891_));
 NAND2x1_ASAP7_75t_R _32255_ (.A(_14310_),
    .B(_00550_),
    .Y(_14892_));
 OA211x2_ASAP7_75t_R _32256_ (.A1(_14474_),
    .A2(_13789_),
    .B(_14892_),
    .C(_13115_),
    .Y(_14893_));
 NAND2x1_ASAP7_75t_R _32257_ (.A(_14317_),
    .B(_00549_),
    .Y(_14894_));
 OA211x2_ASAP7_75t_R _32258_ (.A1(_13107_),
    .A2(_13792_),
    .B(_14894_),
    .C(_14476_),
    .Y(_14895_));
 OR3x1_ASAP7_75t_R _32259_ (.A(_14469_),
    .B(_14893_),
    .C(_14895_),
    .Y(_14896_));
 OA211x2_ASAP7_75t_R _32260_ (.A1(_13186_),
    .A2(_14891_),
    .B(_14896_),
    .C(_13125_),
    .Y(_14897_));
 OR3x2_ASAP7_75t_R _32261_ (.A(_13164_),
    .B(_14883_),
    .C(_14897_),
    .Y(_14898_));
 AO21x2_ASAP7_75t_R _32262_ (.A1(_14869_),
    .A2(_14898_),
    .B(_14377_),
    .Y(_14899_));
 BUFx6f_ASAP7_75t_R _32263_ (.A(_01482_),
    .Y(_14900_));
 AND2x2_ASAP7_75t_R _32264_ (.A(_01450_),
    .B(_14381_),
    .Y(_14901_));
 OAI22x1_ASAP7_75t_R _32265_ (.A1(_14900_),
    .A2(_14382_),
    .B1(_14385_),
    .B2(_14901_),
    .Y(_14902_));
 NAND2x2_ASAP7_75t_R _32266_ (.A(_14899_),
    .B(_14902_),
    .Y(_18579_));
 INVx1_ASAP7_75t_R _32267_ (.A(_18579_),
    .Y(_18577_));
 BUFx6f_ASAP7_75t_R _32268_ (.A(_14627_),
    .Y(_14903_));
 INVx1_ASAP7_75t_R _32269_ (.A(_00114_),
    .Y(_14904_));
 BUFx6f_ASAP7_75t_R _32270_ (.A(_14641_),
    .Y(_14905_));
 BUFx6f_ASAP7_75t_R _32271_ (.A(_14905_),
    .Y(_14906_));
 BUFx6f_ASAP7_75t_R _32272_ (.A(_14906_),
    .Y(_14907_));
 AND3x1_ASAP7_75t_R _32273_ (.A(_14904_),
    .B(_14625_),
    .C(_14907_),
    .Y(_14908_));
 AO21x1_ASAP7_75t_R _32274_ (.A1(_14903_),
    .A2(_18577_),
    .B(_14908_),
    .Y(_18018_));
 NAND2x1_ASAP7_75t_R _32275_ (.A(_14794_),
    .B(_01790_),
    .Y(_14909_));
 OA211x2_ASAP7_75t_R _32276_ (.A1(_14293_),
    .A2(_13875_),
    .B(_14909_),
    .C(_14296_),
    .Y(_14910_));
 AO21x1_ASAP7_75t_R _32277_ (.A1(_13878_),
    .A2(_14449_),
    .B(_14910_),
    .Y(_14911_));
 INVx1_ASAP7_75t_R _32278_ (.A(_00574_),
    .Y(_14912_));
 NAND2x1_ASAP7_75t_R _32279_ (.A(_13196_),
    .B(_00572_),
    .Y(_14913_));
 BUFx12f_ASAP7_75t_R _32280_ (.A(_13114_),
    .Y(_14914_));
 OA211x2_ASAP7_75t_R _32281_ (.A1(_13097_),
    .A2(_14912_),
    .B(_14913_),
    .C(_14914_),
    .Y(_14915_));
 INVx1_ASAP7_75t_R _32282_ (.A(_00573_),
    .Y(_14916_));
 NAND2x1_ASAP7_75t_R _32283_ (.A(_13165_),
    .B(_00571_),
    .Y(_14917_));
 OA211x2_ASAP7_75t_R _32284_ (.A1(_13097_),
    .A2(_14916_),
    .B(_14917_),
    .C(_13120_),
    .Y(_14918_));
 OR3x1_ASAP7_75t_R _32285_ (.A(_13105_),
    .B(_14915_),
    .C(_14918_),
    .Y(_14919_));
 OA211x2_ASAP7_75t_R _32286_ (.A1(_13086_),
    .A2(_14911_),
    .B(_14919_),
    .C(_13125_),
    .Y(_14920_));
 BUFx12f_ASAP7_75t_R _32287_ (.A(_13132_),
    .Y(_14921_));
 NAND2x1_ASAP7_75t_R _32288_ (.A(_14752_),
    .B(_00568_),
    .Y(_14922_));
 BUFx12f_ASAP7_75t_R _32289_ (.A(_14295_),
    .Y(_14923_));
 OA211x2_ASAP7_75t_R _32290_ (.A1(_14921_),
    .A2(_13897_),
    .B(_14922_),
    .C(_14923_),
    .Y(_14924_));
 NAND2x1_ASAP7_75t_R _32291_ (.A(_14815_),
    .B(_00567_),
    .Y(_14925_));
 BUFx12f_ASAP7_75t_R _32292_ (.A(_13100_),
    .Y(_14926_));
 OA211x2_ASAP7_75t_R _32293_ (.A1(_14491_),
    .A2(_13901_),
    .B(_14925_),
    .C(_14926_),
    .Y(_14927_));
 OR3x1_ASAP7_75t_R _32294_ (.A(_14489_),
    .B(_14924_),
    .C(_14927_),
    .Y(_14928_));
 BUFx12f_ASAP7_75t_R _32295_ (.A(_13104_),
    .Y(_14929_));
 NAND2x1_ASAP7_75t_R _32296_ (.A(_14808_),
    .B(_00576_),
    .Y(_14930_));
 OA211x2_ASAP7_75t_R _32297_ (.A1(_14921_),
    .A2(_13867_),
    .B(_14930_),
    .C(_14494_),
    .Y(_14931_));
 NAND2x1_ASAP7_75t_R _32298_ (.A(_14502_),
    .B(_00575_),
    .Y(_14932_));
 OA211x2_ASAP7_75t_R _32299_ (.A1(_14501_),
    .A2(_13841_),
    .B(_14932_),
    .C(_14498_),
    .Y(_14933_));
 OR3x1_ASAP7_75t_R _32300_ (.A(_14929_),
    .B(_14931_),
    .C(_14933_),
    .Y(_14934_));
 AND3x1_ASAP7_75t_R _32301_ (.A(_14488_),
    .B(_14928_),
    .C(_14934_),
    .Y(_14935_));
 OR3x2_ASAP7_75t_R _32302_ (.A(_13082_),
    .B(_14920_),
    .C(_14935_),
    .Y(_14936_));
 INVx1_ASAP7_75t_R _32303_ (.A(_00586_),
    .Y(_14937_));
 NAND2x1_ASAP7_75t_R _32304_ (.A(_14752_),
    .B(_00584_),
    .Y(_14938_));
 OA211x2_ASAP7_75t_R _32305_ (.A1(_14921_),
    .A2(_14937_),
    .B(_14938_),
    .C(_14923_),
    .Y(_14939_));
 NAND2x1_ASAP7_75t_R _32306_ (.A(_14492_),
    .B(_00583_),
    .Y(_14940_));
 OA211x2_ASAP7_75t_R _32307_ (.A1(_14491_),
    .A2(_13892_),
    .B(_14940_),
    .C(_14926_),
    .Y(_14941_));
 OR3x1_ASAP7_75t_R _32308_ (.A(_14489_),
    .B(_14939_),
    .C(_14941_),
    .Y(_14942_));
 BUFx12f_ASAP7_75t_R _32309_ (.A(_14437_),
    .Y(_14943_));
 INVx1_ASAP7_75t_R _32310_ (.A(_00594_),
    .Y(_14944_));
 NAND2x1_ASAP7_75t_R _32311_ (.A(_14808_),
    .B(_00592_),
    .Y(_14945_));
 OA211x2_ASAP7_75t_R _32312_ (.A1(_14943_),
    .A2(_14944_),
    .B(_14945_),
    .C(_14494_),
    .Y(_14946_));
 NAND2x1_ASAP7_75t_R _32313_ (.A(_14502_),
    .B(_00591_),
    .Y(_14947_));
 OA211x2_ASAP7_75t_R _32314_ (.A1(_14501_),
    .A2(_13849_),
    .B(_14947_),
    .C(_14498_),
    .Y(_14948_));
 OR3x1_ASAP7_75t_R _32315_ (.A(_14929_),
    .B(_14946_),
    .C(_14948_),
    .Y(_14949_));
 AND3x1_ASAP7_75t_R _32316_ (.A(_14488_),
    .B(_14942_),
    .C(_14949_),
    .Y(_14950_));
 NAND2x1_ASAP7_75t_R _32317_ (.A(_14492_),
    .B(_00580_),
    .Y(_14951_));
 OA211x2_ASAP7_75t_R _32318_ (.A1(_14491_),
    .A2(_13884_),
    .B(_14951_),
    .C(_14504_),
    .Y(_14952_));
 NAND2x1_ASAP7_75t_R _32319_ (.A(_13189_),
    .B(_00579_),
    .Y(_14953_));
 OA211x2_ASAP7_75t_R _32320_ (.A1(_14506_),
    .A2(_13881_),
    .B(_14953_),
    .C(_14498_),
    .Y(_14954_));
 OR3x1_ASAP7_75t_R _32321_ (.A(_14489_),
    .B(_14952_),
    .C(_14954_),
    .Y(_14955_));
 INVx1_ASAP7_75t_R _32322_ (.A(_00590_),
    .Y(_14956_));
 NAND2x1_ASAP7_75t_R _32323_ (.A(_14502_),
    .B(_00588_),
    .Y(_14957_));
 OA211x2_ASAP7_75t_R _32324_ (.A1(_14501_),
    .A2(_14956_),
    .B(_14957_),
    .C(_14504_),
    .Y(_14958_));
 INVx1_ASAP7_75t_R _32325_ (.A(_00589_),
    .Y(_14959_));
 NAND2x1_ASAP7_75t_R _32326_ (.A(_14507_),
    .B(_00587_),
    .Y(_14960_));
 OA211x2_ASAP7_75t_R _32327_ (.A1(_14506_),
    .A2(_14959_),
    .B(_14960_),
    .C(_14509_),
    .Y(_14961_));
 OR3x1_ASAP7_75t_R _32328_ (.A(_14353_),
    .B(_14958_),
    .C(_14961_),
    .Y(_14962_));
 AND3x1_ASAP7_75t_R _32329_ (.A(_14305_),
    .B(_14955_),
    .C(_14962_),
    .Y(_14963_));
 OR3x2_ASAP7_75t_R _32330_ (.A(_14487_),
    .B(_14950_),
    .C(_14963_),
    .Y(_14964_));
 AO21x2_ASAP7_75t_R _32331_ (.A1(_14936_),
    .A2(_14964_),
    .B(_13267_),
    .Y(_14965_));
 BUFx6f_ASAP7_75t_R _32332_ (.A(_01481_),
    .Y(_14966_));
 BUFx12f_ASAP7_75t_R _32333_ (.A(_14772_),
    .Y(_14967_));
 BUFx6f_ASAP7_75t_R _32334_ (.A(_14383_),
    .Y(_14968_));
 AND2x2_ASAP7_75t_R _32335_ (.A(_01449_),
    .B(_14772_),
    .Y(_14969_));
 OAI22x1_ASAP7_75t_R _32336_ (.A1(_14966_),
    .A2(_14967_),
    .B1(_14968_),
    .B2(_14969_),
    .Y(_14970_));
 NAND2x2_ASAP7_75t_R _32337_ (.A(_14965_),
    .B(_14970_),
    .Y(_18584_));
 INVx2_ASAP7_75t_R _32338_ (.A(_18584_),
    .Y(_18582_));
 INVx1_ASAP7_75t_R _32339_ (.A(_00121_),
    .Y(_14971_));
 AND3x1_ASAP7_75t_R _32340_ (.A(_14971_),
    .B(_14625_),
    .C(_14907_),
    .Y(_14972_));
 AO21x1_ASAP7_75t_R _32341_ (.A1(_14903_),
    .A2(_18582_),
    .B(_14972_),
    .Y(_18020_));
 AND2x2_ASAP7_75t_R _32342_ (.A(_14333_),
    .B(_01789_),
    .Y(_14973_));
 AO21x1_ASAP7_75t_R _32343_ (.A1(_13092_),
    .A2(_00596_),
    .B(_14973_),
    .Y(_14974_));
 BUFx12f_ASAP7_75t_R _32344_ (.A(_13089_),
    .Y(_14975_));
 OAI22x1_ASAP7_75t_R _32345_ (.A1(_00595_),
    .A2(_13102_),
    .B1(_14974_),
    .B2(_14975_),
    .Y(_14976_));
 INVx1_ASAP7_75t_R _32346_ (.A(_00604_),
    .Y(_14977_));
 NAND2x1_ASAP7_75t_R _32347_ (.A(_13196_),
    .B(_00602_),
    .Y(_14978_));
 OA211x2_ASAP7_75t_R _32348_ (.A1(_13097_),
    .A2(_14977_),
    .B(_14978_),
    .C(_14914_),
    .Y(_14979_));
 INVx1_ASAP7_75t_R _32349_ (.A(_00603_),
    .Y(_14980_));
 NAND2x1_ASAP7_75t_R _32350_ (.A(_13165_),
    .B(_00601_),
    .Y(_14981_));
 OA211x2_ASAP7_75t_R _32351_ (.A1(_13097_),
    .A2(_14980_),
    .B(_14981_),
    .C(_13120_),
    .Y(_14982_));
 OR3x1_ASAP7_75t_R _32352_ (.A(_13105_),
    .B(_14979_),
    .C(_14982_),
    .Y(_14983_));
 OA211x2_ASAP7_75t_R _32353_ (.A1(_13086_),
    .A2(_14976_),
    .B(_14983_),
    .C(_13125_),
    .Y(_14984_));
 BUFx12f_ASAP7_75t_R _32354_ (.A(_13132_),
    .Y(_14985_));
 NAND2x1_ASAP7_75t_R _32355_ (.A(_14752_),
    .B(_00598_),
    .Y(_14986_));
 OA211x2_ASAP7_75t_R _32356_ (.A1(_14985_),
    .A2(_13959_),
    .B(_14986_),
    .C(_14923_),
    .Y(_14987_));
 NAND2x1_ASAP7_75t_R _32357_ (.A(_14815_),
    .B(_00597_),
    .Y(_14988_));
 OA211x2_ASAP7_75t_R _32358_ (.A1(_14943_),
    .A2(_13952_),
    .B(_14988_),
    .C(_14926_),
    .Y(_14989_));
 OR3x1_ASAP7_75t_R _32359_ (.A(_14282_),
    .B(_14987_),
    .C(_14989_),
    .Y(_14990_));
 INVx1_ASAP7_75t_R _32360_ (.A(_00608_),
    .Y(_14991_));
 NAND2x1_ASAP7_75t_R _32361_ (.A(_14752_),
    .B(_00606_),
    .Y(_14992_));
 OA211x2_ASAP7_75t_R _32362_ (.A1(_14921_),
    .A2(_14991_),
    .B(_14992_),
    .C(_14923_),
    .Y(_14993_));
 NAND2x1_ASAP7_75t_R _32363_ (.A(_14492_),
    .B(_00605_),
    .Y(_14994_));
 OA211x2_ASAP7_75t_R _32364_ (.A1(_14491_),
    .A2(_13911_),
    .B(_14994_),
    .C(_14926_),
    .Y(_14995_));
 OR3x1_ASAP7_75t_R _32365_ (.A(_14929_),
    .B(_14993_),
    .C(_14995_),
    .Y(_14996_));
 AND3x1_ASAP7_75t_R _32366_ (.A(_14488_),
    .B(_14990_),
    .C(_14996_),
    .Y(_14997_));
 OR3x2_ASAP7_75t_R _32367_ (.A(_13082_),
    .B(_14984_),
    .C(_14997_),
    .Y(_14998_));
 NAND2x1_ASAP7_75t_R _32368_ (.A(_14450_),
    .B(_00614_),
    .Y(_14999_));
 OA211x2_ASAP7_75t_R _32369_ (.A1(_14985_),
    .A2(_13962_),
    .B(_14999_),
    .C(_14369_),
    .Y(_15000_));
 NAND2x1_ASAP7_75t_R _32370_ (.A(_14752_),
    .B(_00613_),
    .Y(_15001_));
 OA211x2_ASAP7_75t_R _32371_ (.A1(_14921_),
    .A2(_13955_),
    .B(_15001_),
    .C(_14372_),
    .Y(_15002_));
 OR3x1_ASAP7_75t_R _32372_ (.A(_14282_),
    .B(_15000_),
    .C(_15002_),
    .Y(_15003_));
 NAND2x1_ASAP7_75t_R _32373_ (.A(_14450_),
    .B(_00622_),
    .Y(_15004_));
 OA211x2_ASAP7_75t_R _32374_ (.A1(_14985_),
    .A2(_13928_),
    .B(_15004_),
    .C(_14369_),
    .Y(_15005_));
 NAND2x1_ASAP7_75t_R _32375_ (.A(_14808_),
    .B(_00621_),
    .Y(_15006_));
 OA211x2_ASAP7_75t_R _32376_ (.A1(_14943_),
    .A2(_13918_),
    .B(_15006_),
    .C(_14372_),
    .Y(_15007_));
 OR3x1_ASAP7_75t_R _32377_ (.A(_14291_),
    .B(_15005_),
    .C(_15007_),
    .Y(_15008_));
 AND3x1_ASAP7_75t_R _32378_ (.A(_14488_),
    .B(_15003_),
    .C(_15008_),
    .Y(_15009_));
 NAND2x1_ASAP7_75t_R _32379_ (.A(_14808_),
    .B(_00610_),
    .Y(_15010_));
 OA211x2_ASAP7_75t_R _32380_ (.A1(_14921_),
    .A2(_13947_),
    .B(_15010_),
    .C(_14923_),
    .Y(_15011_));
 NAND2x1_ASAP7_75t_R _32381_ (.A(_14492_),
    .B(_00609_),
    .Y(_15012_));
 OA211x2_ASAP7_75t_R _32382_ (.A1(_14501_),
    .A2(_13944_),
    .B(_15012_),
    .C(_14926_),
    .Y(_15013_));
 OR3x1_ASAP7_75t_R _32383_ (.A(_14489_),
    .B(_15011_),
    .C(_15013_),
    .Y(_15014_));
 INVx1_ASAP7_75t_R _32384_ (.A(_00620_),
    .Y(_15015_));
 NAND2x1_ASAP7_75t_R _32385_ (.A(_14815_),
    .B(_00618_),
    .Y(_15016_));
 OA211x2_ASAP7_75t_R _32386_ (.A1(_14943_),
    .A2(_15015_),
    .B(_15016_),
    .C(_14494_),
    .Y(_15017_));
 INVx1_ASAP7_75t_R _32387_ (.A(_00619_),
    .Y(_15018_));
 NAND2x1_ASAP7_75t_R _32388_ (.A(_14502_),
    .B(_00617_),
    .Y(_15019_));
 OA211x2_ASAP7_75t_R _32389_ (.A1(_14496_),
    .A2(_15018_),
    .B(_15019_),
    .C(_14498_),
    .Y(_15020_));
 OR3x1_ASAP7_75t_R _32390_ (.A(_14929_),
    .B(_15017_),
    .C(_15020_),
    .Y(_15021_));
 AND3x1_ASAP7_75t_R _32391_ (.A(_14305_),
    .B(_15014_),
    .C(_15021_),
    .Y(_15022_));
 OR3x2_ASAP7_75t_R _32392_ (.A(_14487_),
    .B(_15009_),
    .C(_15022_),
    .Y(_15023_));
 AO21x2_ASAP7_75t_R _32393_ (.A1(_14998_),
    .A2(_15023_),
    .B(_13267_),
    .Y(_15024_));
 AND2x2_ASAP7_75t_R _32394_ (.A(_01448_),
    .B(_14381_),
    .Y(_15025_));
 OAI22x1_ASAP7_75t_R _32395_ (.A1(_01480_),
    .A2(_14967_),
    .B1(_14968_),
    .B2(_15025_),
    .Y(_15026_));
 AND2x6_ASAP7_75t_R _32396_ (.A(_15024_),
    .B(_15026_),
    .Y(_18587_));
 INVx2_ASAP7_75t_R _32397_ (.A(_18587_),
    .Y(_18589_));
 INVx2_ASAP7_75t_R _32398_ (.A(_00128_),
    .Y(_15027_));
 AND3x1_ASAP7_75t_R _32399_ (.A(_15027_),
    .B(_14625_),
    .C(_14907_),
    .Y(_15028_));
 AO21x1_ASAP7_75t_R _32400_ (.A1(_14903_),
    .A2(_18587_),
    .B(_15028_),
    .Y(_18022_));
 BUFx3_ASAP7_75t_R _32401_ (.A(_00765_),
    .Y(_15029_));
 AO21x1_ASAP7_75t_R _32402_ (.A1(_15029_),
    .A2(_00768_),
    .B(_00767_),
    .Y(_15030_));
 AND2x4_ASAP7_75t_R _32403_ (.A(_00770_),
    .B(_15030_),
    .Y(_15031_));
 INVx1_ASAP7_75t_R _32404_ (.A(_00757_),
    .Y(_15032_));
 OA21x2_ASAP7_75t_R _32405_ (.A1(_15032_),
    .A2(_00755_),
    .B(_00762_),
    .Y(_15033_));
 OR2x6_ASAP7_75t_R _32406_ (.A(_00761_),
    .B(_00763_),
    .Y(_15034_));
 OA21x2_ASAP7_75t_R _32407_ (.A1(_00764_),
    .A2(_00763_),
    .B(_00766_),
    .Y(_15035_));
 AND3x1_ASAP7_75t_R _32408_ (.A(_00768_),
    .B(_00770_),
    .C(_15035_),
    .Y(_15036_));
 OA21x2_ASAP7_75t_R _32409_ (.A1(_15033_),
    .A2(_15034_),
    .B(_15036_),
    .Y(_15037_));
 OR3x1_ASAP7_75t_R _32410_ (.A(_00769_),
    .B(_15031_),
    .C(_15037_),
    .Y(_15038_));
 AND2x2_ASAP7_75t_R _32411_ (.A(_00772_),
    .B(_15038_),
    .Y(_15039_));
 XNOR2x1_ASAP7_75t_R _32412_ (.B(_15039_),
    .Y(_15040_),
    .A(_00771_));
 INVx3_ASAP7_75t_R _32413_ (.A(_15040_),
    .Y(\alu_adder_result_ex[7] ));
 OA21x2_ASAP7_75t_R _32414_ (.A1(_15029_),
    .A2(_15035_),
    .B(_00768_),
    .Y(_15041_));
 OA21x2_ASAP7_75t_R _32415_ (.A1(_00755_),
    .A2(_00756_),
    .B(_00762_),
    .Y(_15042_));
 OA211x2_ASAP7_75t_R _32416_ (.A1(_00767_),
    .A2(_15041_),
    .B(_15042_),
    .C(_00770_),
    .Y(_15043_));
 OR2x6_ASAP7_75t_R _32417_ (.A(_00755_),
    .B(_00754_),
    .Y(_15044_));
 AO21x1_ASAP7_75t_R _32418_ (.A1(_15042_),
    .A2(_15044_),
    .B(_15034_),
    .Y(_15045_));
 AO21x1_ASAP7_75t_R _32419_ (.A1(_15035_),
    .A2(_15045_),
    .B(_15029_),
    .Y(_15046_));
 AO21x1_ASAP7_75t_R _32420_ (.A1(_00768_),
    .A2(_15046_),
    .B(_00767_),
    .Y(_15047_));
 AO32x1_ASAP7_75t_R _32421_ (.A1(net1953),
    .A2(_14626_),
    .A3(_15043_),
    .B1(_15047_),
    .B2(_00770_),
    .Y(_15048_));
 XOR2x1_ASAP7_75t_R _32422_ (.A(_00769_),
    .Y(\alu_adder_result_ex[6] ),
    .B(_15048_));
 AND2x2_ASAP7_75t_R _32423_ (.A(_14450_),
    .B(_01788_),
    .Y(_15049_));
 AO21x1_ASAP7_75t_R _32424_ (.A1(_13092_),
    .A2(_00626_),
    .B(_15049_),
    .Y(_15050_));
 OAI22x1_ASAP7_75t_R _32425_ (.A1(_00625_),
    .A2(_13102_),
    .B1(_15050_),
    .B2(_13187_),
    .Y(_15051_));
 BUFx12f_ASAP7_75t_R _32426_ (.A(_14460_),
    .Y(_15052_));
 INVx1_ASAP7_75t_R _32427_ (.A(_00634_),
    .Y(_15053_));
 NAND2x1_ASAP7_75t_R _32428_ (.A(_14292_),
    .B(_00632_),
    .Y(_15054_));
 OA211x2_ASAP7_75t_R _32429_ (.A1(_15052_),
    .A2(_15053_),
    .B(_15054_),
    .C(_14458_),
    .Y(_15055_));
 INVx1_ASAP7_75t_R _32430_ (.A(_00633_),
    .Y(_15056_));
 NAND2x1_ASAP7_75t_R _32431_ (.A(_14292_),
    .B(_00631_),
    .Y(_15057_));
 OA211x2_ASAP7_75t_R _32432_ (.A1(_14320_),
    .A2(_15056_),
    .B(_15057_),
    .C(_14743_),
    .Y(_15058_));
 OR3x1_ASAP7_75t_R _32433_ (.A(_14454_),
    .B(_15055_),
    .C(_15058_),
    .Y(_15059_));
 OA21x2_ASAP7_75t_R _32434_ (.A1(_14448_),
    .A2(_15051_),
    .B(_15059_),
    .Y(_15060_));
 BUFx12f_ASAP7_75t_R _32435_ (.A(_14667_),
    .Y(_15061_));
 NAND2x1_ASAP7_75t_R _32436_ (.A(_14437_),
    .B(_00628_),
    .Y(_15062_));
 OA211x2_ASAP7_75t_R _32437_ (.A1(_15061_),
    .A2(_14013_),
    .B(_15062_),
    .C(_14458_),
    .Y(_15063_));
 NAND2x1_ASAP7_75t_R _32438_ (.A(_14490_),
    .B(_00627_),
    .Y(_15064_));
 OA211x2_ASAP7_75t_R _32439_ (.A1(_13200_),
    .A2(_14010_),
    .B(_15064_),
    .C(_14743_),
    .Y(_15065_));
 OR3x1_ASAP7_75t_R _32440_ (.A(_14737_),
    .B(_15063_),
    .C(_15065_),
    .Y(_15066_));
 NAND2x1_ASAP7_75t_R _32441_ (.A(_14437_),
    .B(_00636_),
    .Y(_15067_));
 OA211x2_ASAP7_75t_R _32442_ (.A1(_14738_),
    .A2(_13996_),
    .B(_15067_),
    .C(_14740_),
    .Y(_15068_));
 NAND2x1_ASAP7_75t_R _32443_ (.A(_14490_),
    .B(_00635_),
    .Y(_15069_));
 OA211x2_ASAP7_75t_R _32444_ (.A1(_13200_),
    .A2(_14003_),
    .B(_15069_),
    .C(_14743_),
    .Y(_15070_));
 OR3x1_ASAP7_75t_R _32445_ (.A(_14454_),
    .B(_15068_),
    .C(_15070_),
    .Y(_15071_));
 AND3x1_ASAP7_75t_R _32446_ (.A(_14468_),
    .B(_15066_),
    .C(_15071_),
    .Y(_15072_));
 AO21x1_ASAP7_75t_R _32447_ (.A1(_14778_),
    .A2(_15060_),
    .B(_15072_),
    .Y(_15073_));
 NAND2x1_ASAP7_75t_R _32448_ (.A(_14515_),
    .B(_00644_),
    .Y(_15074_));
 OA211x2_ASAP7_75t_R _32449_ (.A1(_14794_),
    .A2(_14017_),
    .B(_15074_),
    .C(_14740_),
    .Y(_15075_));
 NAND2x1_ASAP7_75t_R _32450_ (.A(_14515_),
    .B(_00643_),
    .Y(_15076_));
 OA211x2_ASAP7_75t_R _32451_ (.A1(_14277_),
    .A2(_14020_),
    .B(_15076_),
    .C(_14732_),
    .Y(_15077_));
 OR3x1_ASAP7_75t_R _32452_ (.A(_14737_),
    .B(_15075_),
    .C(_15077_),
    .Y(_15078_));
 NAND2x1_ASAP7_75t_R _32453_ (.A(_14515_),
    .B(_00652_),
    .Y(_15079_));
 OA211x2_ASAP7_75t_R _32454_ (.A1(_14794_),
    .A2(_13981_),
    .B(_15079_),
    .C(_14729_),
    .Y(_15080_));
 INVx1_ASAP7_75t_R _32455_ (.A(_00653_),
    .Y(_15081_));
 NAND2x1_ASAP7_75t_R _32456_ (.A(_14515_),
    .B(_00651_),
    .Y(_15082_));
 OA211x2_ASAP7_75t_R _32457_ (.A1(_14301_),
    .A2(_15081_),
    .B(_15082_),
    .C(_14732_),
    .Y(_15083_));
 OR3x1_ASAP7_75t_R _32458_ (.A(_13185_),
    .B(_15080_),
    .C(_15083_),
    .Y(_15084_));
 AND3x1_ASAP7_75t_R _32459_ (.A(_14807_),
    .B(_15078_),
    .C(_15084_),
    .Y(_15085_));
 NAND2x1_ASAP7_75t_R _32460_ (.A(_14515_),
    .B(_00640_),
    .Y(_15086_));
 OA211x2_ASAP7_75t_R _32461_ (.A1(_14277_),
    .A2(_13985_),
    .B(_15086_),
    .C(_14729_),
    .Y(_15087_));
 NAND2x1_ASAP7_75t_R _32462_ (.A(_14515_),
    .B(_00639_),
    .Y(_15088_));
 OA211x2_ASAP7_75t_R _32463_ (.A1(_14301_),
    .A2(_13988_),
    .B(_15088_),
    .C(_14732_),
    .Y(_15089_));
 OR3x1_ASAP7_75t_R _32464_ (.A(_14737_),
    .B(_15087_),
    .C(_15089_),
    .Y(_15090_));
 NAND2x1_ASAP7_75t_R _32465_ (.A(_14515_),
    .B(_00648_),
    .Y(_15091_));
 OA211x2_ASAP7_75t_R _32466_ (.A1(_14277_),
    .A2(_13971_),
    .B(_15091_),
    .C(_14729_),
    .Y(_15092_));
 NAND2x1_ASAP7_75t_R _32467_ (.A(_13205_),
    .B(_00647_),
    .Y(_15093_));
 OA211x2_ASAP7_75t_R _32468_ (.A1(_14367_),
    .A2(_13977_),
    .B(_15093_),
    .C(_14732_),
    .Y(_15094_));
 OR3x1_ASAP7_75t_R _32469_ (.A(_13185_),
    .B(_15092_),
    .C(_15094_),
    .Y(_15095_));
 AND3x1_ASAP7_75t_R _32470_ (.A(_14466_),
    .B(_15090_),
    .C(_15095_),
    .Y(_15096_));
 OR3x2_ASAP7_75t_R _32471_ (.A(_14487_),
    .B(_15085_),
    .C(_15096_),
    .Y(_15097_));
 OA21x2_ASAP7_75t_R _32472_ (.A1(_14281_),
    .A2(_15073_),
    .B(_15097_),
    .Y(_15098_));
 BUFx6f_ASAP7_75t_R _32473_ (.A(_01479_),
    .Y(_15099_));
 BUFx6f_ASAP7_75t_R _32474_ (.A(_14380_),
    .Y(_15100_));
 AND2x2_ASAP7_75t_R _32475_ (.A(_01447_),
    .B(_14772_),
    .Y(_15101_));
 OAI22x1_ASAP7_75t_R _32476_ (.A1(_15099_),
    .A2(_15100_),
    .B1(_14384_),
    .B2(_15101_),
    .Y(_15102_));
 OA21x2_ASAP7_75t_R _32477_ (.A1(_13268_),
    .A2(_15098_),
    .B(_15102_),
    .Y(_15103_));
 BUFx6f_ASAP7_75t_R _32478_ (.A(_15103_),
    .Y(_18592_));
 INVx3_ASAP7_75t_R _32479_ (.A(_18592_),
    .Y(_18594_));
 BUFx6f_ASAP7_75t_R _32480_ (.A(_14627_),
    .Y(_15104_));
 OR3x1_ASAP7_75t_R _32481_ (.A(_00135_),
    .B(_15104_),
    .C(_14650_),
    .Y(_15105_));
 OAI21x1_ASAP7_75t_R _32482_ (.A1(_14647_),
    .A2(_18594_),
    .B(_15105_),
    .Y(_18024_));
 AND2x2_ASAP7_75t_R _32483_ (.A(_13206_),
    .B(_01787_),
    .Y(_15106_));
 AO21x1_ASAP7_75t_R _32484_ (.A1(_14286_),
    .A2(_00656_),
    .B(_15106_),
    .Y(_15107_));
 OAI22x1_ASAP7_75t_R _32485_ (.A1(_00655_),
    .A2(_14284_),
    .B1(_15107_),
    .B2(_14289_),
    .Y(_15108_));
 INVx1_ASAP7_75t_R _32486_ (.A(_00664_),
    .Y(_15109_));
 NAND2x1_ASAP7_75t_R _32487_ (.A(_14815_),
    .B(_00662_),
    .Y(_15110_));
 OA211x2_ASAP7_75t_R _32488_ (.A1(_14491_),
    .A2(_15109_),
    .B(_15110_),
    .C(_14494_),
    .Y(_15111_));
 INVx1_ASAP7_75t_R _32489_ (.A(_00663_),
    .Y(_15112_));
 NAND2x1_ASAP7_75t_R _32490_ (.A(_13189_),
    .B(_00661_),
    .Y(_15113_));
 OA211x2_ASAP7_75t_R _32491_ (.A1(_14496_),
    .A2(_15112_),
    .B(_15113_),
    .C(_14498_),
    .Y(_15114_));
 OR3x1_ASAP7_75t_R _32492_ (.A(_14929_),
    .B(_15111_),
    .C(_15114_),
    .Y(_15115_));
 OA211x2_ASAP7_75t_R _32493_ (.A1(_14283_),
    .A2(_15108_),
    .B(_15115_),
    .C(_14852_),
    .Y(_15116_));
 BUFx12f_ASAP7_75t_R _32494_ (.A(_13130_),
    .Y(_15117_));
 NAND2x1_ASAP7_75t_R _32495_ (.A(_15061_),
    .B(_00658_),
    .Y(_15118_));
 OA211x2_ASAP7_75t_R _32496_ (.A1(_14711_),
    .A2(_14029_),
    .B(_15118_),
    .C(_13202_),
    .Y(_15119_));
 BUFx12f_ASAP7_75t_R _32497_ (.A(_14678_),
    .Y(_15120_));
 NAND2x1_ASAP7_75t_R _32498_ (.A(_14738_),
    .B(_00657_),
    .Y(_15121_));
 BUFx6f_ASAP7_75t_R _32499_ (.A(_13173_),
    .Y(_15122_));
 OA211x2_ASAP7_75t_R _32500_ (.A1(_15120_),
    .A2(_14032_),
    .B(_15121_),
    .C(_15122_),
    .Y(_15123_));
 OR3x1_ASAP7_75t_R _32501_ (.A(_15117_),
    .B(_15119_),
    .C(_15123_),
    .Y(_15124_));
 INVx1_ASAP7_75t_R _32502_ (.A(_00668_),
    .Y(_15125_));
 NAND2x1_ASAP7_75t_R _32503_ (.A(_15061_),
    .B(_00666_),
    .Y(_15126_));
 OA211x2_ASAP7_75t_R _32504_ (.A1(_15120_),
    .A2(_15125_),
    .B(_15126_),
    .C(_13202_),
    .Y(_15127_));
 NAND2x1_ASAP7_75t_R _32505_ (.A(_14738_),
    .B(_00665_),
    .Y(_15128_));
 OA211x2_ASAP7_75t_R _32506_ (.A1(_13197_),
    .A2(_14060_),
    .B(_15128_),
    .C(_14874_),
    .Y(_15129_));
 OR3x1_ASAP7_75t_R _32507_ (.A(_14877_),
    .B(_15127_),
    .C(_15129_),
    .Y(_15130_));
 AND3x1_ASAP7_75t_R _32508_ (.A(_14340_),
    .B(_15124_),
    .C(_15130_),
    .Y(_15131_));
 OR3x2_ASAP7_75t_R _32509_ (.A(_13082_),
    .B(_15116_),
    .C(_15131_),
    .Y(_15132_));
 NAND2x1_ASAP7_75t_R _32510_ (.A(_14782_),
    .B(_00674_),
    .Y(_15133_));
 OA211x2_ASAP7_75t_R _32511_ (.A1(_14711_),
    .A2(_14036_),
    .B(_15133_),
    .C(_14652_),
    .Y(_15134_));
 NAND2x1_ASAP7_75t_R _32512_ (.A(_15061_),
    .B(_00673_),
    .Y(_15135_));
 OA211x2_ASAP7_75t_R _32513_ (.A1(_15120_),
    .A2(_14039_),
    .B(_15135_),
    .C(_15122_),
    .Y(_15136_));
 OR3x1_ASAP7_75t_R _32514_ (.A(_15117_),
    .B(_15134_),
    .C(_15136_),
    .Y(_15137_));
 NAND2x1_ASAP7_75t_R _32515_ (.A(_14782_),
    .B(_00682_),
    .Y(_15138_));
 OA211x2_ASAP7_75t_R _32516_ (.A1(_14711_),
    .A2(_14079_),
    .B(_15138_),
    .C(_13202_),
    .Y(_15139_));
 NAND2x1_ASAP7_75t_R _32517_ (.A(_14738_),
    .B(_00681_),
    .Y(_15140_));
 OA211x2_ASAP7_75t_R _32518_ (.A1(_15120_),
    .A2(_14067_),
    .B(_15140_),
    .C(_15122_),
    .Y(_15141_));
 OR3x1_ASAP7_75t_R _32519_ (.A(_14877_),
    .B(_15139_),
    .C(_15141_),
    .Y(_15142_));
 AND3x1_ASAP7_75t_R _32520_ (.A(_14340_),
    .B(_15137_),
    .C(_15142_),
    .Y(_15143_));
 NOR2x1_ASAP7_75t_R _32521_ (.A(_14366_),
    .B(_00679_),
    .Y(_15144_));
 AO21x1_ASAP7_75t_R _32522_ (.A1(_13190_),
    .A2(_14064_),
    .B(_15144_),
    .Y(_15145_));
 NAND2x1_ASAP7_75t_R _32523_ (.A(_14333_),
    .B(_00678_),
    .Y(_15146_));
 OA211x2_ASAP7_75t_R _32524_ (.A1(_14331_),
    .A2(_14082_),
    .B(_15146_),
    .C(_14329_),
    .Y(_15147_));
 AO21x1_ASAP7_75t_R _32525_ (.A1(_14975_),
    .A2(_15145_),
    .B(_15147_),
    .Y(_15148_));
 NAND2x1_ASAP7_75t_R _32526_ (.A(_14507_),
    .B(_00670_),
    .Y(_15149_));
 OA211x2_ASAP7_75t_R _32527_ (.A1(_14506_),
    .A2(_14052_),
    .B(_15149_),
    .C(_14472_),
    .Y(_15150_));
 INVx1_ASAP7_75t_R _32528_ (.A(_00671_),
    .Y(_15151_));
 NAND2x1_ASAP7_75t_R _32529_ (.A(_14517_),
    .B(_00669_),
    .Y(_15152_));
 OA211x2_ASAP7_75t_R _32530_ (.A1(_14516_),
    .A2(_15151_),
    .B(_15152_),
    .C(_14509_),
    .Y(_15153_));
 OR3x1_ASAP7_75t_R _32531_ (.A(_14469_),
    .B(_15150_),
    .C(_15153_),
    .Y(_15154_));
 OA211x2_ASAP7_75t_R _32532_ (.A1(_14354_),
    .A2(_15148_),
    .B(_15154_),
    .C(_14852_),
    .Y(_15155_));
 OR3x2_ASAP7_75t_R _32533_ (.A(_13164_),
    .B(_15143_),
    .C(_15155_),
    .Y(_15156_));
 AO21x2_ASAP7_75t_R _32534_ (.A1(_15132_),
    .A2(_15156_),
    .B(_13268_),
    .Y(_15157_));
 BUFx6f_ASAP7_75t_R _32535_ (.A(_01478_),
    .Y(_15158_));
 AND2x2_ASAP7_75t_R _32536_ (.A(_01446_),
    .B(_14381_),
    .Y(_15159_));
 OAI22x1_ASAP7_75t_R _32537_ (.A1(_15158_),
    .A2(_14382_),
    .B1(_14385_),
    .B2(_15159_),
    .Y(_15160_));
 NAND2x2_ASAP7_75t_R _32538_ (.A(_15157_),
    .B(_15160_),
    .Y(_18599_));
 INVx1_ASAP7_75t_R _32539_ (.A(_18599_),
    .Y(_18597_));
 OR3x1_ASAP7_75t_R _32540_ (.A(_00144_),
    .B(_15104_),
    .C(_14650_),
    .Y(_15161_));
 OAI21x1_ASAP7_75t_R _32541_ (.A1(_14647_),
    .A2(_18599_),
    .B(_15161_),
    .Y(_18026_));
 OR3x1_ASAP7_75t_R _32542_ (.A(_00769_),
    .B(_00771_),
    .C(net1948),
    .Y(_15162_));
 OA21x2_ASAP7_75t_R _32543_ (.A1(_00772_),
    .A2(_00771_),
    .B(_00774_),
    .Y(_15163_));
 OA21x2_ASAP7_75t_R _32544_ (.A1(net1948),
    .A2(_15163_),
    .B(_00776_),
    .Y(_15164_));
 OA31x2_ASAP7_75t_R _32545_ (.A1(_15031_),
    .A2(_15037_),
    .A3(_15162_),
    .B1(_15164_),
    .Y(_15165_));
 XNOR2x1_ASAP7_75t_R _32546_ (.B(_15165_),
    .Y(_15166_),
    .A(net1950));
 INVx3_ASAP7_75t_R _32547_ (.A(_15166_),
    .Y(\alu_adder_result_ex[9] ));
 OR2x6_ASAP7_75t_R _32548_ (.A(_00769_),
    .B(_00771_),
    .Y(_15167_));
 OA21x2_ASAP7_75t_R _32549_ (.A1(_15031_),
    .A2(_15167_),
    .B(_15163_),
    .Y(_15168_));
 BUFx6f_ASAP7_75t_R _32550_ (.A(_15168_),
    .Y(_15169_));
 OR2x6_ASAP7_75t_R _32551_ (.A(_15034_),
    .B(_15044_),
    .Y(_15170_));
 OA21x2_ASAP7_75t_R _32552_ (.A1(_00761_),
    .A2(_15042_),
    .B(_00764_),
    .Y(_15171_));
 OA22x2_ASAP7_75t_R _32553_ (.A1(_00763_),
    .A2(_15171_),
    .B1(_15170_),
    .B2(_14626_),
    .Y(_15172_));
 OA21x2_ASAP7_75t_R _32554_ (.A1(_00768_),
    .A2(_00767_),
    .B(_00770_),
    .Y(_15173_));
 OA211x2_ASAP7_75t_R _32555_ (.A1(_15167_),
    .A2(_15173_),
    .B(_00766_),
    .C(_15163_),
    .Y(_15174_));
 OA211x2_ASAP7_75t_R _32556_ (.A1(net1953),
    .A2(_15170_),
    .B(_15172_),
    .C(_15174_),
    .Y(_15175_));
 BUFx6f_ASAP7_75t_R _32557_ (.A(_15175_),
    .Y(_15176_));
 OAI21x1_ASAP7_75t_R _32558_ (.A1(_15169_),
    .A2(_15176_),
    .B(net1949),
    .Y(_15177_));
 OR3x2_ASAP7_75t_R _32559_ (.A(net1949),
    .B(_15169_),
    .C(_15176_),
    .Y(_15178_));
 NAND2x2_ASAP7_75t_R _32560_ (.A(_15177_),
    .B(_15178_),
    .Y(_15179_));
 INVx3_ASAP7_75t_R _32561_ (.A(_15179_),
    .Y(\alu_adder_result_ex[8] ));
 AND2x2_ASAP7_75t_R _32562_ (.A(_14516_),
    .B(_01786_),
    .Y(_15180_));
 AO21x1_ASAP7_75t_R _32563_ (.A1(_14286_),
    .A2(_00686_),
    .B(_15180_),
    .Y(_15181_));
 OAI22x1_ASAP7_75t_R _32564_ (.A1(_00685_),
    .A2(_14284_),
    .B1(_15181_),
    .B2(_14289_),
    .Y(_15182_));
 INVx1_ASAP7_75t_R _32565_ (.A(_00694_),
    .Y(_15183_));
 NAND2x1_ASAP7_75t_R _32566_ (.A(_14794_),
    .B(_00692_),
    .Y(_15184_));
 OA211x2_ASAP7_75t_R _32567_ (.A1(_14293_),
    .A2(_15183_),
    .B(_15184_),
    .C(_14296_),
    .Y(_15185_));
 INVx1_ASAP7_75t_R _32568_ (.A(_00693_),
    .Y(_15186_));
 NAND2x1_ASAP7_75t_R _32569_ (.A(_14301_),
    .B(_00691_),
    .Y(_15187_));
 OA211x2_ASAP7_75t_R _32570_ (.A1(_14299_),
    .A2(_15186_),
    .B(_15187_),
    .C(_13149_),
    .Y(_15188_));
 OR3x1_ASAP7_75t_R _32571_ (.A(_14291_),
    .B(_15185_),
    .C(_15188_),
    .Y(_15189_));
 OA211x2_ASAP7_75t_R _32572_ (.A1(_14283_),
    .A2(_15182_),
    .B(_15189_),
    .C(_14305_),
    .Y(_15190_));
 BUFx6f_ASAP7_75t_R _32573_ (.A(_14470_),
    .Y(_15191_));
 NAND2x1_ASAP7_75t_R _32574_ (.A(_15052_),
    .B(_00688_),
    .Y(_15192_));
 OA211x2_ASAP7_75t_R _32575_ (.A1(_15191_),
    .A2(_14174_),
    .B(_15192_),
    .C(_14315_),
    .Y(_15193_));
 NAND2x1_ASAP7_75t_R _32576_ (.A(_14320_),
    .B(_00687_),
    .Y(_15194_));
 BUFx6f_ASAP7_75t_R _32577_ (.A(_14322_),
    .Y(_15195_));
 OA211x2_ASAP7_75t_R _32578_ (.A1(_14318_),
    .A2(_14177_),
    .B(_15194_),
    .C(_15195_),
    .Y(_15196_));
 OR3x1_ASAP7_75t_R _32579_ (.A(_14309_),
    .B(_15193_),
    .C(_15196_),
    .Y(_15197_));
 NAND2x1_ASAP7_75t_R _32580_ (.A(_14312_),
    .B(_00696_),
    .Y(_15198_));
 OA211x2_ASAP7_75t_R _32581_ (.A1(_14311_),
    .A2(_14181_),
    .B(_15198_),
    .C(_14315_),
    .Y(_15199_));
 NAND2x1_ASAP7_75t_R _32582_ (.A(_14320_),
    .B(_00695_),
    .Y(_15200_));
 OA211x2_ASAP7_75t_R _32583_ (.A1(_14318_),
    .A2(_14167_),
    .B(_15200_),
    .C(_14323_),
    .Y(_15201_));
 OR3x1_ASAP7_75t_R _32584_ (.A(_14327_),
    .B(_15199_),
    .C(_15201_),
    .Y(_15202_));
 AND3x1_ASAP7_75t_R _32585_ (.A(_14307_),
    .B(_15197_),
    .C(_15202_),
    .Y(_15203_));
 OR3x2_ASAP7_75t_R _32586_ (.A(_14281_),
    .B(_15190_),
    .C(_15203_),
    .Y(_15204_));
 NAND2x1_ASAP7_75t_R _32587_ (.A(_15052_),
    .B(_00704_),
    .Y(_15205_));
 OA211x2_ASAP7_75t_R _32588_ (.A1(_14311_),
    .A2(_14152_),
    .B(_15205_),
    .C(_14315_),
    .Y(_15206_));
 NAND2x1_ASAP7_75t_R _32589_ (.A(_14320_),
    .B(_00703_),
    .Y(_15207_));
 OA211x2_ASAP7_75t_R _32590_ (.A1(_14318_),
    .A2(_14155_),
    .B(_15207_),
    .C(_15195_),
    .Y(_15208_));
 OR3x1_ASAP7_75t_R _32591_ (.A(_14309_),
    .B(_15206_),
    .C(_15208_),
    .Y(_15209_));
 NAND2x1_ASAP7_75t_R _32592_ (.A(_14312_),
    .B(_00712_),
    .Y(_15210_));
 OA211x2_ASAP7_75t_R _32593_ (.A1(_14311_),
    .A2(_14160_),
    .B(_15210_),
    .C(_14315_),
    .Y(_15211_));
 NAND2x1_ASAP7_75t_R _32594_ (.A(_14320_),
    .B(_00711_),
    .Y(_15212_));
 OA211x2_ASAP7_75t_R _32595_ (.A1(_14318_),
    .A2(_14163_),
    .B(_15212_),
    .C(_14323_),
    .Y(_15213_));
 OR3x1_ASAP7_75t_R _32596_ (.A(_14327_),
    .B(_15211_),
    .C(_15213_),
    .Y(_15214_));
 AND3x1_ASAP7_75t_R _32597_ (.A(_14307_),
    .B(_15209_),
    .C(_15214_),
    .Y(_15215_));
 NAND2x1_ASAP7_75t_R _32598_ (.A(_14320_),
    .B(_00700_),
    .Y(_15216_));
 OA211x2_ASAP7_75t_R _32599_ (.A1(_14318_),
    .A2(_14193_),
    .B(_15216_),
    .C(_14329_),
    .Y(_15217_));
 NAND2x1_ASAP7_75t_R _32600_ (.A(_14333_),
    .B(_00699_),
    .Y(_15218_));
 OA211x2_ASAP7_75t_R _32601_ (.A1(_14331_),
    .A2(_14196_),
    .B(_15218_),
    .C(_14323_),
    .Y(_15219_));
 OR3x1_ASAP7_75t_R _32602_ (.A(_14309_),
    .B(_15217_),
    .C(_15219_),
    .Y(_15220_));
 NAND2x1_ASAP7_75t_R _32603_ (.A(_14320_),
    .B(_00708_),
    .Y(_15221_));
 OA211x2_ASAP7_75t_R _32604_ (.A1(_14318_),
    .A2(_14145_),
    .B(_15221_),
    .C(_14329_),
    .Y(_15222_));
 NAND2x1_ASAP7_75t_R _32605_ (.A(_14333_),
    .B(_00707_),
    .Y(_15223_));
 OA211x2_ASAP7_75t_R _32606_ (.A1(_14331_),
    .A2(_14148_),
    .B(_15223_),
    .C(_14323_),
    .Y(_15224_));
 OR3x1_ASAP7_75t_R _32607_ (.A(_14327_),
    .B(_15222_),
    .C(_15224_),
    .Y(_15225_));
 AND3x1_ASAP7_75t_R _32608_ (.A(_14778_),
    .B(_15220_),
    .C(_15225_),
    .Y(_15226_));
 OR3x2_ASAP7_75t_R _32609_ (.A(_14339_),
    .B(_15215_),
    .C(_15226_),
    .Y(_15227_));
 AO21x2_ASAP7_75t_R _32610_ (.A1(_15204_),
    .A2(_15227_),
    .B(_14377_),
    .Y(_15228_));
 AND2x2_ASAP7_75t_R _32611_ (.A(_01476_),
    .B(_14381_),
    .Y(_15229_));
 OAI22x1_ASAP7_75t_R _32612_ (.A1(_00019_),
    .A2(_14382_),
    .B1(_14385_),
    .B2(_15229_),
    .Y(_15230_));
 AND2x4_ASAP7_75t_R _32613_ (.A(_15228_),
    .B(_15230_),
    .Y(_18602_));
 INVx3_ASAP7_75t_R _32614_ (.A(_18602_),
    .Y(_18604_));
 OR3x1_ASAP7_75t_R _32615_ (.A(_00152_),
    .B(_15104_),
    .C(_14650_),
    .Y(_15231_));
 OAI21x1_ASAP7_75t_R _32616_ (.A1(_14647_),
    .A2(_18604_),
    .B(_15231_),
    .Y(_18028_));
 INVx1_ASAP7_75t_R _32617_ (.A(_00160_),
    .Y(_15232_));
 AND3x4_ASAP7_75t_R _32618_ (.A(_13832_),
    .B(_14562_),
    .C(_14539_),
    .Y(_15233_));
 BUFx12f_ASAP7_75t_R _32619_ (.A(_15233_),
    .Y(_15234_));
 BUFx6f_ASAP7_75t_R _32620_ (.A(_15234_),
    .Y(_15235_));
 BUFx6f_ASAP7_75t_R _32621_ (.A(_15235_),
    .Y(_15236_));
 AND3x1_ASAP7_75t_R _32622_ (.A(_15232_),
    .B(_15236_),
    .C(_14907_),
    .Y(_15237_));
 AO21x1_ASAP7_75t_R _32623_ (.A1(_18607_),
    .A2(_14648_),
    .B(_15237_),
    .Y(_18030_));
 OA21x2_ASAP7_75t_R _32624_ (.A1(net1950),
    .A2(_15165_),
    .B(_00778_),
    .Y(_15238_));
 OA21x2_ASAP7_75t_R _32625_ (.A1(net1942),
    .A2(_15238_),
    .B(_00780_),
    .Y(_15239_));
 XNOR2x1_ASAP7_75t_R _32626_ (.B(_15239_),
    .Y(_15240_),
    .A(net1944));
 INVx3_ASAP7_75t_R _32627_ (.A(_15240_),
    .Y(\alu_adder_result_ex[11] ));
 BUFx12f_ASAP7_75t_R _32628_ (.A(net1953),
    .Y(_15241_));
 OA21x2_ASAP7_75t_R _32629_ (.A1(net1950),
    .A2(_15164_),
    .B(_00778_),
    .Y(_15242_));
 AND3x1_ASAP7_75t_R _32630_ (.A(_14626_),
    .B(_15043_),
    .C(_15242_),
    .Y(_15243_));
 AND2x2_ASAP7_75t_R _32631_ (.A(_00770_),
    .B(_15047_),
    .Y(_15244_));
 OR3x1_ASAP7_75t_R _32632_ (.A(net1949),
    .B(net1950),
    .C(_15167_),
    .Y(_15245_));
 OA21x2_ASAP7_75t_R _32633_ (.A1(_15244_),
    .A2(_15245_),
    .B(_15242_),
    .Y(_15246_));
 AO21x2_ASAP7_75t_R _32634_ (.A1(_15241_),
    .A2(_15243_),
    .B(_15246_),
    .Y(_15247_));
 XNOR2x1_ASAP7_75t_R _32635_ (.B(_15247_),
    .Y(_15248_),
    .A(net1943));
 INVx2_ASAP7_75t_R _32636_ (.A(_15248_),
    .Y(\alu_adder_result_ex[10] ));
 OR3x1_ASAP7_75t_R _32637_ (.A(_00168_),
    .B(_15104_),
    .C(_14650_),
    .Y(_15249_));
 OAI21x1_ASAP7_75t_R _32638_ (.A1(_18613_),
    .A2(_14647_),
    .B(_15249_),
    .Y(_18032_));
 BUFx12f_ASAP7_75t_R _32639_ (.A(_13969_),
    .Y(_15250_));
 BUFx6f_ASAP7_75t_R _32640_ (.A(_13764_),
    .Y(_15251_));
 BUFx12f_ASAP7_75t_R _32641_ (.A(_13669_),
    .Y(_15252_));
 BUFx6f_ASAP7_75t_R _32642_ (.A(_15252_),
    .Y(_15253_));
 BUFx12f_ASAP7_75t_R _32643_ (.A(_13688_),
    .Y(_15254_));
 BUFx6f_ASAP7_75t_R _32644_ (.A(_15254_),
    .Y(_15255_));
 BUFx12f_ASAP7_75t_R _32645_ (.A(_13813_),
    .Y(_15256_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 BUFx12f_ASAP7_75t_R _32647_ (.A(_15256_),
    .Y(_15258_));
 BUFx12f_ASAP7_75t_R _32648_ (.A(_15258_),
    .Y(_15259_));
 BUFx6f_ASAP7_75t_R _32649_ (.A(_15259_),
    .Y(_15260_));
 BUFx12f_ASAP7_75t_R _32650_ (.A(_15258_),
    .Y(_15261_));
 BUFx12f_ASAP7_75t_R _32651_ (.A(_15261_),
    .Y(_15262_));
 NAND2x1_ASAP7_75t_R _32652_ (.A(_00348_),
    .B(_15262_),
    .Y(_15263_));
 BUFx6f_ASAP7_75t_R _32653_ (.A(_13434_),
    .Y(_15264_));
 BUFx12f_ASAP7_75t_R _32654_ (.A(_15264_),
    .Y(_15265_));
 BUFx12f_ASAP7_75t_R _32655_ (.A(_15265_),
    .Y(_15266_));
 BUFx6f_ASAP7_75t_R _32656_ (.A(_15266_),
    .Y(_15267_));
 OA211x2_ASAP7_75t_R _32657_ (.A1(_13134_),
    .A2(_15260_),
    .B(_15263_),
    .C(_15267_),
    .Y(_15268_));
 BUFx6f_ASAP7_75t_R _32658_ (.A(_15259_),
    .Y(_15269_));
 BUFx12f_ASAP7_75t_R _32659_ (.A(_15261_),
    .Y(_15270_));
 NAND2x1_ASAP7_75t_R _32660_ (.A(_00347_),
    .B(_15270_),
    .Y(_15271_));
 BUFx6f_ASAP7_75t_R _32661_ (.A(_14191_),
    .Y(_15272_));
 BUFx12f_ASAP7_75t_R _32662_ (.A(_15272_),
    .Y(_15273_));
 BUFx12f_ASAP7_75t_R _32663_ (.A(_15273_),
    .Y(_15274_));
 BUFx6f_ASAP7_75t_R _32664_ (.A(_15274_),
    .Y(_15275_));
 OA211x2_ASAP7_75t_R _32665_ (.A1(_13144_),
    .A2(_15269_),
    .B(_15271_),
    .C(_15275_),
    .Y(_15276_));
 OR3x1_ASAP7_75t_R _32666_ (.A(_15255_),
    .B(_15268_),
    .C(_15276_),
    .Y(_15277_));
 BUFx12f_ASAP7_75t_R _32667_ (.A(_13724_),
    .Y(_15278_));
 BUFx6f_ASAP7_75t_R _32668_ (.A(_15278_),
    .Y(_15279_));
 NAND2x1_ASAP7_75t_R _32669_ (.A(_00356_),
    .B(_15262_),
    .Y(_15280_));
 OA211x2_ASAP7_75t_R _32670_ (.A1(_13154_),
    .A2(_15260_),
    .B(_15280_),
    .C(_15267_),
    .Y(_15281_));
 NAND2x1_ASAP7_75t_R _32671_ (.A(_00355_),
    .B(_15270_),
    .Y(_15282_));
 BUFx6f_ASAP7_75t_R _32672_ (.A(_15274_),
    .Y(_15283_));
 OA211x2_ASAP7_75t_R _32673_ (.A1(_13157_),
    .A2(_15269_),
    .B(_15282_),
    .C(_15283_),
    .Y(_15284_));
 OR3x1_ASAP7_75t_R _32674_ (.A(_15279_),
    .B(_15281_),
    .C(_15284_),
    .Y(_15285_));
 AND3x4_ASAP7_75t_R _32675_ (.A(_15253_),
    .B(_15277_),
    .C(_15285_),
    .Y(_15286_));
 BUFx6f_ASAP7_75t_R _32676_ (.A(_15254_),
    .Y(_15287_));
 BUFx6f_ASAP7_75t_R _32677_ (.A(_15287_),
    .Y(_15288_));
 BUFx12f_ASAP7_75t_R _32678_ (.A(_13670_),
    .Y(_15289_));
 BUFx6f_ASAP7_75t_R _32679_ (.A(_13328_),
    .Y(_15290_));
 BUFx12f_ASAP7_75t_R _32680_ (.A(net1968),
    .Y(_15291_));
 AND2x2_ASAP7_75t_R _32681_ (.A(_15291_),
    .B(_01784_),
    .Y(_15292_));
 AO21x1_ASAP7_75t_R _32682_ (.A1(_00346_),
    .A2(_15290_),
    .B(_15292_),
    .Y(_15293_));
 BUFx6f_ASAP7_75t_R _32683_ (.A(_15273_),
    .Y(_15294_));
 BUFx6f_ASAP7_75t_R _32684_ (.A(_15294_),
    .Y(_15295_));
 BUFx12f_ASAP7_75t_R _32685_ (.A(_15295_),
    .Y(_15296_));
 OAI22x1_ASAP7_75t_R _32686_ (.A1(_00345_),
    .A2(_15289_),
    .B1(_15293_),
    .B2(_15296_),
    .Y(_15297_));
 BUFx12f_ASAP7_75t_R _32687_ (.A(_15278_),
    .Y(_15298_));
 BUFx12f_ASAP7_75t_R _32688_ (.A(_15258_),
    .Y(_15299_));
 BUFx12f_ASAP7_75t_R _32689_ (.A(_15299_),
    .Y(_15300_));
 BUFx12f_ASAP7_75t_R _32690_ (.A(_15258_),
    .Y(_15301_));
 BUFx6f_ASAP7_75t_R _32691_ (.A(_15301_),
    .Y(_15302_));
 NAND2x1_ASAP7_75t_R _32692_ (.A(_00352_),
    .B(_15302_),
    .Y(_15303_));
 BUFx6f_ASAP7_75t_R _32693_ (.A(_15265_),
    .Y(_15304_));
 OA211x2_ASAP7_75t_R _32694_ (.A1(_13108_),
    .A2(_15300_),
    .B(_15303_),
    .C(_15304_),
    .Y(_15305_));
 BUFx12f_ASAP7_75t_R _32695_ (.A(_15258_),
    .Y(_15306_));
 BUFx6f_ASAP7_75t_R _32696_ (.A(_15306_),
    .Y(_15307_));
 NAND2x1_ASAP7_75t_R _32697_ (.A(_00351_),
    .B(_15302_),
    .Y(_15308_));
 BUFx6f_ASAP7_75t_R _32698_ (.A(_15273_),
    .Y(_15309_));
 OA211x2_ASAP7_75t_R _32699_ (.A1(_13117_),
    .A2(_15307_),
    .B(_15308_),
    .C(_15309_),
    .Y(_15310_));
 OR3x1_ASAP7_75t_R _32700_ (.A(_15298_),
    .B(_15305_),
    .C(_15310_),
    .Y(_15311_));
 BUFx12f_ASAP7_75t_R _32701_ (.A(_13814_),
    .Y(_15312_));
 BUFx6f_ASAP7_75t_R _32702_ (.A(_15312_),
    .Y(_15313_));
 OA211x2_ASAP7_75t_R _32703_ (.A1(_15288_),
    .A2(_15297_),
    .B(_15311_),
    .C(_15313_),
    .Y(_15314_));
 OR3x2_ASAP7_75t_R _32704_ (.A(_15251_),
    .B(_15286_),
    .C(_15314_),
    .Y(_15315_));
 BUFx6f_ASAP7_75t_R _32705_ (.A(_13306_),
    .Y(_15316_));
 BUFx6f_ASAP7_75t_R _32706_ (.A(_15252_),
    .Y(_15317_));
 BUFx6f_ASAP7_75t_R _32707_ (.A(_15254_),
    .Y(_15318_));
 BUFx12f_ASAP7_75t_R _32708_ (.A(_15258_),
    .Y(_15319_));
 BUFx6f_ASAP7_75t_R _32709_ (.A(_15319_),
    .Y(_15320_));
 BUFx12f_ASAP7_75t_R _32710_ (.A(_15299_),
    .Y(_15321_));
 NAND2x1_ASAP7_75t_R _32711_ (.A(_00364_),
    .B(_15321_),
    .Y(_15322_));
 BUFx6f_ASAP7_75t_R _32712_ (.A(_15266_),
    .Y(_15323_));
 OA211x2_ASAP7_75t_R _32713_ (.A1(_13167_),
    .A2(_15320_),
    .B(_15322_),
    .C(_15323_),
    .Y(_15324_));
 BUFx6f_ASAP7_75t_R _32714_ (.A(_15259_),
    .Y(_15325_));
 BUFx12f_ASAP7_75t_R _32715_ (.A(_15299_),
    .Y(_15326_));
 NAND2x1_ASAP7_75t_R _32716_ (.A(_00363_),
    .B(_15326_),
    .Y(_15327_));
 OA211x2_ASAP7_75t_R _32717_ (.A1(_13171_),
    .A2(_15325_),
    .B(_15327_),
    .C(_15275_),
    .Y(_15328_));
 OR3x1_ASAP7_75t_R _32718_ (.A(_15318_),
    .B(_15324_),
    .C(_15328_),
    .Y(_15329_));
 NAND2x1_ASAP7_75t_R _32719_ (.A(_00372_),
    .B(_15321_),
    .Y(_15330_));
 OA211x2_ASAP7_75t_R _32720_ (.A1(_13177_),
    .A2(_15325_),
    .B(_15330_),
    .C(_15323_),
    .Y(_15331_));
 NAND2x1_ASAP7_75t_R _32721_ (.A(_00371_),
    .B(_15326_),
    .Y(_15332_));
 OA211x2_ASAP7_75t_R _32722_ (.A1(_13180_),
    .A2(_15325_),
    .B(_15332_),
    .C(_15275_),
    .Y(_15333_));
 OR3x1_ASAP7_75t_R _32723_ (.A(_15279_),
    .B(_15331_),
    .C(_15333_),
    .Y(_15334_));
 AND3x1_ASAP7_75t_R _32724_ (.A(_15317_),
    .B(_15329_),
    .C(_15334_),
    .Y(_15335_));
 BUFx6f_ASAP7_75t_R _32725_ (.A(_15278_),
    .Y(_15336_));
 BUFx6f_ASAP7_75t_R _32726_ (.A(_15336_),
    .Y(_15337_));
 BUFx6f_ASAP7_75t_R _32727_ (.A(_15274_),
    .Y(_15338_));
 BUFx6f_ASAP7_75t_R _32728_ (.A(_15338_),
    .Y(_15339_));
 BUFx12f_ASAP7_75t_R _32729_ (.A(_15301_),
    .Y(_15340_));
 BUFx6f_ASAP7_75t_R _32730_ (.A(_15340_),
    .Y(_15341_));
 BUFx12f_ASAP7_75t_R _32731_ (.A(_15258_),
    .Y(_15342_));
 BUFx6f_ASAP7_75t_R _32732_ (.A(_15342_),
    .Y(_15343_));
 NOR2x1_ASAP7_75t_R _32733_ (.A(_00369_),
    .B(_15343_),
    .Y(_15344_));
 AO21x1_ASAP7_75t_R _32734_ (.A1(_13191_),
    .A2(_15341_),
    .B(_15344_),
    .Y(_15345_));
 BUFx6f_ASAP7_75t_R _32735_ (.A(_15319_),
    .Y(_15346_));
 BUFx12f_ASAP7_75t_R _32736_ (.A(net1957),
    .Y(_15347_));
 NAND2x1_ASAP7_75t_R _32737_ (.A(_00368_),
    .B(_15347_),
    .Y(_15348_));
 BUFx6f_ASAP7_75t_R _32738_ (.A(_15266_),
    .Y(_15349_));
 OA211x2_ASAP7_75t_R _32739_ (.A1(_13198_),
    .A2(_15346_),
    .B(_15348_),
    .C(_15349_),
    .Y(_15350_));
 AO21x1_ASAP7_75t_R _32740_ (.A1(_15339_),
    .A2(_15345_),
    .B(_15350_),
    .Y(_15351_));
 BUFx6f_ASAP7_75t_R _32741_ (.A(_15254_),
    .Y(_15352_));
 BUFx6f_ASAP7_75t_R _32742_ (.A(_15306_),
    .Y(_15353_));
 BUFx12f_ASAP7_75t_R _32743_ (.A(_15301_),
    .Y(_15354_));
 NAND2x1_ASAP7_75t_R _32744_ (.A(_00360_),
    .B(_15354_),
    .Y(_15355_));
 OA211x2_ASAP7_75t_R _32745_ (.A1(_13207_),
    .A2(_15353_),
    .B(_15355_),
    .C(_15304_),
    .Y(_15356_));
 NAND2x1_ASAP7_75t_R _32746_ (.A(_00359_),
    .B(_15354_),
    .Y(_15357_));
 OA211x2_ASAP7_75t_R _32747_ (.A1(_13210_),
    .A2(_15353_),
    .B(_15357_),
    .C(_15309_),
    .Y(_15358_));
 OR3x1_ASAP7_75t_R _32748_ (.A(_15352_),
    .B(_15356_),
    .C(_15358_),
    .Y(_15359_));
 BUFx6f_ASAP7_75t_R _32749_ (.A(_15312_),
    .Y(_15360_));
 OA211x2_ASAP7_75t_R _32750_ (.A1(_15337_),
    .A2(_15351_),
    .B(_15359_),
    .C(_15360_),
    .Y(_15361_));
 OR3x2_ASAP7_75t_R _32751_ (.A(_15316_),
    .B(_15335_),
    .C(_15361_),
    .Y(_15362_));
 NAND2x2_ASAP7_75t_R _32752_ (.A(_15315_),
    .B(_15362_),
    .Y(_15363_));
 NAND2x2_ASAP7_75t_R _32753_ (.A(_14262_),
    .B(_14263_),
    .Y(_15364_));
 OR3x2_ASAP7_75t_R _32754_ (.A(_14262_),
    .B(_13444_),
    .C(_14263_),
    .Y(_15365_));
 AND2x6_ASAP7_75t_R _32755_ (.A(_15364_),
    .B(_15365_),
    .Y(_15366_));
 INVx2_ASAP7_75t_R _32756_ (.A(_14099_),
    .Y(_15367_));
 AO32x2_ASAP7_75t_R _32757_ (.A1(_13296_),
    .A2(_13260_),
    .A3(_13437_),
    .B1(_13439_),
    .B2(_13444_),
    .Y(_15368_));
 NAND2x2_ASAP7_75t_R _32758_ (.A(_15367_),
    .B(_15368_),
    .Y(_15369_));
 BUFx6f_ASAP7_75t_R _32759_ (.A(_13763_),
    .Y(_15370_));
 OA211x2_ASAP7_75t_R _32760_ (.A1(_14272_),
    .A2(_15366_),
    .B(_15369_),
    .C(_15370_),
    .Y(_15371_));
 AOI21x1_ASAP7_75t_R _32761_ (.A1(_15250_),
    .A2(_15363_),
    .B(_15371_),
    .Y(_18614_));
 INVx1_ASAP7_75t_R _32762_ (.A(_18614_),
    .Y(_18612_));
 AND2x2_ASAP7_75t_R _32763_ (.A(_13107_),
    .B(_01783_),
    .Y(_15372_));
 AO21x1_ASAP7_75t_R _32764_ (.A1(_14286_),
    .A2(_00784_),
    .B(_15372_),
    .Y(_15373_));
 OAI22x1_ASAP7_75t_R _32765_ (.A1(_00783_),
    .A2(_14284_),
    .B1(_15373_),
    .B2(_14289_),
    .Y(_15374_));
 INVx2_ASAP7_75t_R _32766_ (.A(_00792_),
    .Y(_15375_));
 NAND2x1_ASAP7_75t_R _32767_ (.A(_14450_),
    .B(_00790_),
    .Y(_15376_));
 OA211x2_ASAP7_75t_R _32768_ (.A1(_14985_),
    .A2(_15375_),
    .B(_15376_),
    .C(_14369_),
    .Y(_15377_));
 INVx1_ASAP7_75t_R _32769_ (.A(_00791_),
    .Y(_15378_));
 NAND2x1_ASAP7_75t_R _32770_ (.A(_14752_),
    .B(_00789_),
    .Y(_15379_));
 OA211x2_ASAP7_75t_R _32771_ (.A1(_14921_),
    .A2(_15378_),
    .B(_15379_),
    .C(_14372_),
    .Y(_15380_));
 OR3x1_ASAP7_75t_R _32772_ (.A(_14291_),
    .B(_15377_),
    .C(_15380_),
    .Y(_15381_));
 OA211x2_ASAP7_75t_R _32773_ (.A1(_14283_),
    .A2(_15374_),
    .B(_15381_),
    .C(_14305_),
    .Y(_15382_));
 INVx2_ASAP7_75t_R _32774_ (.A(_00788_),
    .Y(_15383_));
 NAND2x1_ASAP7_75t_R _32775_ (.A(_14756_),
    .B(_00786_),
    .Y(_15384_));
 OA211x2_ASAP7_75t_R _32776_ (.A1(_14886_),
    .A2(_15383_),
    .B(_15384_),
    .C(_14652_),
    .Y(_15385_));
 INVx2_ASAP7_75t_R _32777_ (.A(_00787_),
    .Y(_15386_));
 NAND2x1_ASAP7_75t_R _32778_ (.A(_14782_),
    .B(_00785_),
    .Y(_15387_));
 OA211x2_ASAP7_75t_R _32779_ (.A1(_14886_),
    .A2(_15386_),
    .B(_15387_),
    .C(_15122_),
    .Y(_15388_));
 OR3x1_ASAP7_75t_R _32780_ (.A(_15117_),
    .B(_15385_),
    .C(_15388_),
    .Y(_15389_));
 INVx1_ASAP7_75t_R _32781_ (.A(_00796_),
    .Y(_15390_));
 NAND2x1_ASAP7_75t_R _32782_ (.A(_14888_),
    .B(_00794_),
    .Y(_15391_));
 OA211x2_ASAP7_75t_R _32783_ (.A1(_14886_),
    .A2(_15390_),
    .B(_15391_),
    .C(_14652_),
    .Y(_15392_));
 INVx1_ASAP7_75t_R _32784_ (.A(_00795_),
    .Y(_15393_));
 NAND2x1_ASAP7_75t_R _32785_ (.A(_14782_),
    .B(_00793_),
    .Y(_15394_));
 OA211x2_ASAP7_75t_R _32786_ (.A1(_14711_),
    .A2(_15393_),
    .B(_15394_),
    .C(_15122_),
    .Y(_15395_));
 OR3x1_ASAP7_75t_R _32787_ (.A(_14877_),
    .B(_15392_),
    .C(_15395_),
    .Y(_15396_));
 AND3x4_ASAP7_75t_R _32788_ (.A(_14340_),
    .B(_15389_),
    .C(_15396_),
    .Y(_15397_));
 OR3x2_ASAP7_75t_R _32789_ (.A(_14281_),
    .B(_15382_),
    .C(_15397_),
    .Y(_15398_));
 INVx2_ASAP7_75t_R _32790_ (.A(_00804_),
    .Y(_15399_));
 NAND2x1_ASAP7_75t_R _32791_ (.A(_14756_),
    .B(_00802_),
    .Y(_15400_));
 OA211x2_ASAP7_75t_R _32792_ (.A1(_14331_),
    .A2(_15399_),
    .B(_15400_),
    .C(_14329_),
    .Y(_15401_));
 INVx2_ASAP7_75t_R _32793_ (.A(_00803_),
    .Y(_15402_));
 NAND2x1_ASAP7_75t_R _32794_ (.A(_14888_),
    .B(_00801_),
    .Y(_15403_));
 OA211x2_ASAP7_75t_R _32795_ (.A1(_14886_),
    .A2(_15402_),
    .B(_15403_),
    .C(_14323_),
    .Y(_15404_));
 OR3x1_ASAP7_75t_R _32796_ (.A(_15117_),
    .B(_15401_),
    .C(_15404_),
    .Y(_15405_));
 INVx1_ASAP7_75t_R _32797_ (.A(_00812_),
    .Y(_15406_));
 NAND2x1_ASAP7_75t_R _32798_ (.A(_14756_),
    .B(_00810_),
    .Y(_15407_));
 OA211x2_ASAP7_75t_R _32799_ (.A1(_14331_),
    .A2(_15406_),
    .B(_15407_),
    .C(_14329_),
    .Y(_15408_));
 INVx2_ASAP7_75t_R _32800_ (.A(_00811_),
    .Y(_15409_));
 NAND2x1_ASAP7_75t_R _32801_ (.A(_14888_),
    .B(_00809_),
    .Y(_15410_));
 OA211x2_ASAP7_75t_R _32802_ (.A1(_14886_),
    .A2(_15409_),
    .B(_15410_),
    .C(_14323_),
    .Y(_15411_));
 OR3x1_ASAP7_75t_R _32803_ (.A(_14327_),
    .B(_15408_),
    .C(_15411_),
    .Y(_15412_));
 AND3x1_ASAP7_75t_R _32804_ (.A(_14340_),
    .B(_15405_),
    .C(_15412_),
    .Y(_15413_));
 INVx2_ASAP7_75t_R _32805_ (.A(_00805_),
    .Y(_15414_));
 NOR2x1_ASAP7_75t_R _32806_ (.A(_14299_),
    .B(_00807_),
    .Y(_15415_));
 AO21x1_ASAP7_75t_R _32807_ (.A1(_14278_),
    .A2(_15414_),
    .B(_15415_),
    .Y(_15416_));
 INVx2_ASAP7_75t_R _32808_ (.A(_00808_),
    .Y(_15417_));
 NAND2x1_ASAP7_75t_R _32809_ (.A(_14312_),
    .B(_00806_),
    .Y(_15418_));
 OA211x2_ASAP7_75t_R _32810_ (.A1(_14311_),
    .A2(_15417_),
    .B(_15418_),
    .C(_14329_),
    .Y(_15419_));
 AO21x1_ASAP7_75t_R _32811_ (.A1(_14975_),
    .A2(_15416_),
    .B(_15419_),
    .Y(_15420_));
 INVx2_ASAP7_75t_R _32812_ (.A(_00800_),
    .Y(_15421_));
 NAND2x1_ASAP7_75t_R _32813_ (.A(_14808_),
    .B(_00798_),
    .Y(_15422_));
 OA211x2_ASAP7_75t_R _32814_ (.A1(_14943_),
    .A2(_15421_),
    .B(_15422_),
    .C(_14494_),
    .Y(_15423_));
 INVx2_ASAP7_75t_R _32815_ (.A(_00799_),
    .Y(_15424_));
 NAND2x1_ASAP7_75t_R _32816_ (.A(_14502_),
    .B(_00797_),
    .Y(_15425_));
 OA211x2_ASAP7_75t_R _32817_ (.A1(_14501_),
    .A2(_15424_),
    .B(_15425_),
    .C(_14498_),
    .Y(_15426_));
 OR3x1_ASAP7_75t_R _32818_ (.A(_14489_),
    .B(_15423_),
    .C(_15426_),
    .Y(_15427_));
 OA211x2_ASAP7_75t_R _32819_ (.A1(_14354_),
    .A2(_15420_),
    .B(_15427_),
    .C(_14852_),
    .Y(_15428_));
 OR3x2_ASAP7_75t_R _32820_ (.A(_14339_),
    .B(_15413_),
    .C(_15428_),
    .Y(_15429_));
 AO21x2_ASAP7_75t_R _32821_ (.A1(_15398_),
    .A2(_15429_),
    .B(_13268_),
    .Y(_15430_));
 AND2x2_ASAP7_75t_R _32822_ (.A(_01473_),
    .B(_15100_),
    .Y(_15431_));
 OAI22x1_ASAP7_75t_R _32823_ (.A1(_01502_),
    .A2(_14382_),
    .B1(_14385_),
    .B2(_15431_),
    .Y(_15432_));
 NAND2x2_ASAP7_75t_R _32824_ (.A(_15430_),
    .B(_15432_),
    .Y(_18618_));
 INVx1_ASAP7_75t_R _32825_ (.A(_18618_),
    .Y(_18620_));
 OR3x1_ASAP7_75t_R _32826_ (.A(_00175_),
    .B(_15104_),
    .C(_14650_),
    .Y(_15433_));
 OAI21x1_ASAP7_75t_R _32827_ (.A1(_14647_),
    .A2(_18618_),
    .B(_15433_),
    .Y(_18034_));
 BUFx6f_ASAP7_75t_R _32828_ (.A(_15251_),
    .Y(_15434_));
 BUFx12f_ASAP7_75t_R _32829_ (.A(_15289_),
    .Y(_15435_));
 BUFx6f_ASAP7_75t_R _32830_ (.A(_15290_),
    .Y(_15436_));
 BUFx6f_ASAP7_75t_R _32831_ (.A(_15299_),
    .Y(_15437_));
 AND2x2_ASAP7_75t_R _32832_ (.A(_15437_),
    .B(_01783_),
    .Y(_15438_));
 AO21x1_ASAP7_75t_R _32833_ (.A1(_15436_),
    .A2(_00784_),
    .B(_15438_),
    .Y(_15439_));
 OAI22x1_ASAP7_75t_R _32834_ (.A1(_00783_),
    .A2(_15435_),
    .B1(_15439_),
    .B2(_15296_),
    .Y(_15440_));
 BUFx6f_ASAP7_75t_R _32835_ (.A(_15342_),
    .Y(_15441_));
 NAND2x1_ASAP7_75t_R _32836_ (.A(_15302_),
    .B(_00790_),
    .Y(_15442_));
 BUFx6f_ASAP7_75t_R _32837_ (.A(_15265_),
    .Y(_15443_));
 OA211x2_ASAP7_75t_R _32838_ (.A1(_15441_),
    .A2(_15375_),
    .B(_15442_),
    .C(_15443_),
    .Y(_15444_));
 BUFx6f_ASAP7_75t_R _32839_ (.A(_15306_),
    .Y(_15445_));
 NAND2x1_ASAP7_75t_R _32840_ (.A(_15302_),
    .B(_00789_),
    .Y(_15446_));
 OA211x2_ASAP7_75t_R _32841_ (.A1(_15445_),
    .A2(_15378_),
    .B(_15446_),
    .C(_15309_),
    .Y(_15447_));
 OR3x1_ASAP7_75t_R _32842_ (.A(_15298_),
    .B(_15444_),
    .C(_15447_),
    .Y(_15448_));
 OA211x2_ASAP7_75t_R _32843_ (.A1(_15288_),
    .A2(_15440_),
    .B(_15448_),
    .C(_15360_),
    .Y(_15449_));
 BUFx6f_ASAP7_75t_R _32844_ (.A(_15319_),
    .Y(_15450_));
 BUFx12f_ASAP7_75t_R _32845_ (.A(_15301_),
    .Y(_15451_));
 NAND2x1_ASAP7_75t_R _32846_ (.A(_15451_),
    .B(_00786_),
    .Y(_15452_));
 OA211x2_ASAP7_75t_R _32847_ (.A1(_15450_),
    .A2(_15383_),
    .B(_15452_),
    .C(_15323_),
    .Y(_15453_));
 BUFx12f_ASAP7_75t_R _32848_ (.A(_15261_),
    .Y(_15454_));
 NAND2x1_ASAP7_75t_R _32849_ (.A(_15454_),
    .B(_00785_),
    .Y(_15455_));
 BUFx6f_ASAP7_75t_R _32850_ (.A(_15274_),
    .Y(_15456_));
 OA211x2_ASAP7_75t_R _32851_ (.A1(_15320_),
    .A2(_15386_),
    .B(_15455_),
    .C(_15456_),
    .Y(_15457_));
 OR3x1_ASAP7_75t_R _32852_ (.A(_15318_),
    .B(_15453_),
    .C(_15457_),
    .Y(_15458_));
 NAND2x1_ASAP7_75t_R _32853_ (.A(_15454_),
    .B(_00794_),
    .Y(_15459_));
 OA211x2_ASAP7_75t_R _32854_ (.A1(_15450_),
    .A2(_15390_),
    .B(_15459_),
    .C(_15323_),
    .Y(_15460_));
 NAND2x1_ASAP7_75t_R _32855_ (.A(_15454_),
    .B(_00793_),
    .Y(_15461_));
 OA211x2_ASAP7_75t_R _32856_ (.A1(_15320_),
    .A2(_15393_),
    .B(_15461_),
    .C(_15275_),
    .Y(_15462_));
 OR3x1_ASAP7_75t_R _32857_ (.A(_15279_),
    .B(_15460_),
    .C(_15462_),
    .Y(_15463_));
 AND3x4_ASAP7_75t_R _32858_ (.A(_15317_),
    .B(_15458_),
    .C(_15463_),
    .Y(_15464_));
 OR3x2_ASAP7_75t_R _32859_ (.A(_15434_),
    .B(_15449_),
    .C(_15464_),
    .Y(_15465_));
 BUFx12f_ASAP7_75t_R _32860_ (.A(_15316_),
    .Y(_15466_));
 BUFx12f_ASAP7_75t_R _32861_ (.A(_15319_),
    .Y(_15467_));
 NAND2x1_ASAP7_75t_R _32862_ (.A(_15326_),
    .B(_00802_),
    .Y(_15468_));
 BUFx6f_ASAP7_75t_R _32863_ (.A(_15266_),
    .Y(_15469_));
 OA211x2_ASAP7_75t_R _32864_ (.A1(_15467_),
    .A2(_15399_),
    .B(_15468_),
    .C(_15469_),
    .Y(_15470_));
 BUFx6f_ASAP7_75t_R _32865_ (.A(_15319_),
    .Y(_15471_));
 NAND2x1_ASAP7_75t_R _32866_ (.A(_15326_),
    .B(_00801_),
    .Y(_15472_));
 OA211x2_ASAP7_75t_R _32867_ (.A1(_15471_),
    .A2(_15402_),
    .B(_15472_),
    .C(_15338_),
    .Y(_15473_));
 OR3x1_ASAP7_75t_R _32868_ (.A(_15318_),
    .B(_15470_),
    .C(_15473_),
    .Y(_15474_));
 BUFx6f_ASAP7_75t_R _32869_ (.A(_15278_),
    .Y(_15475_));
 NAND2x1_ASAP7_75t_R _32870_ (.A(_15326_),
    .B(_00810_),
    .Y(_15476_));
 OA211x2_ASAP7_75t_R _32871_ (.A1(_15467_),
    .A2(_15406_),
    .B(_15476_),
    .C(_15349_),
    .Y(_15477_));
 NAND2x1_ASAP7_75t_R _32872_ (.A(_15262_),
    .B(_00809_),
    .Y(_15478_));
 OA211x2_ASAP7_75t_R _32873_ (.A1(_15471_),
    .A2(_15409_),
    .B(_15478_),
    .C(_15338_),
    .Y(_15479_));
 OR3x1_ASAP7_75t_R _32874_ (.A(_15475_),
    .B(_15477_),
    .C(_15479_),
    .Y(_15480_));
 AND3x1_ASAP7_75t_R _32875_ (.A(_15317_),
    .B(_15474_),
    .C(_15480_),
    .Y(_15481_));
 BUFx12f_ASAP7_75t_R _32876_ (.A(_15298_),
    .Y(_15482_));
 BUFx12f_ASAP7_75t_R _32877_ (.A(_15301_),
    .Y(_15483_));
 BUFx6f_ASAP7_75t_R _32878_ (.A(_15483_),
    .Y(_15484_));
 BUFx12f_ASAP7_75t_R _32879_ (.A(_15258_),
    .Y(_15485_));
 BUFx12f_ASAP7_75t_R _32880_ (.A(_15485_),
    .Y(_15486_));
 NOR2x1_ASAP7_75t_R _32881_ (.A(_15486_),
    .B(_00807_),
    .Y(_15487_));
 AO21x1_ASAP7_75t_R _32882_ (.A1(_15484_),
    .A2(_15414_),
    .B(_15487_),
    .Y(_15488_));
 BUFx12f_ASAP7_75t_R _32883_ (.A(_15301_),
    .Y(_15489_));
 BUFx6f_ASAP7_75t_R _32884_ (.A(_15489_),
    .Y(_15490_));
 NAND2x1_ASAP7_75t_R _32885_ (.A(_15347_),
    .B(_00806_),
    .Y(_15491_));
 OA211x2_ASAP7_75t_R _32886_ (.A1(_15490_),
    .A2(_15417_),
    .B(_15491_),
    .C(_15469_),
    .Y(_15492_));
 AO21x1_ASAP7_75t_R _32887_ (.A1(_15339_),
    .A2(_15488_),
    .B(_15492_),
    .Y(_15493_));
 NAND2x1_ASAP7_75t_R _32888_ (.A(_15354_),
    .B(_00798_),
    .Y(_15494_));
 OA211x2_ASAP7_75t_R _32889_ (.A1(_15441_),
    .A2(_15421_),
    .B(_15494_),
    .C(_15443_),
    .Y(_15495_));
 NAND2x1_ASAP7_75t_R _32890_ (.A(_15354_),
    .B(_00797_),
    .Y(_15496_));
 BUFx6f_ASAP7_75t_R _32891_ (.A(_15273_),
    .Y(_15497_));
 OA211x2_ASAP7_75t_R _32892_ (.A1(_15441_),
    .A2(_15424_),
    .B(_15496_),
    .C(_15497_),
    .Y(_15498_));
 OR3x1_ASAP7_75t_R _32893_ (.A(_15352_),
    .B(_15495_),
    .C(_15498_),
    .Y(_15499_));
 OA211x2_ASAP7_75t_R _32894_ (.A1(_15482_),
    .A2(_15493_),
    .B(_15499_),
    .C(_15360_),
    .Y(_15500_));
 OR3x2_ASAP7_75t_R _32895_ (.A(_15466_),
    .B(_15481_),
    .C(_15500_),
    .Y(_15501_));
 NAND2x2_ASAP7_75t_R _32896_ (.A(_15501_),
    .B(_15465_),
    .Y(_15502_));
 BUFx3_ASAP7_75t_R _32897_ (.A(_15370_),
    .Y(_15503_));
 OA211x2_ASAP7_75t_R _32898_ (.A1(_14112_),
    .A2(_15366_),
    .B(_15369_),
    .C(_15503_),
    .Y(_15504_));
 AOI21x1_ASAP7_75t_R _32899_ (.A1(_14090_),
    .A2(net1970),
    .B(_15504_),
    .Y(_18619_));
 INVx1_ASAP7_75t_R _32900_ (.A(_18619_),
    .Y(_18617_));
 OR4x1_ASAP7_75t_R _32901_ (.A(net1950),
    .B(net1942),
    .C(net1945),
    .D(net1938),
    .Y(_15505_));
 OA21x2_ASAP7_75t_R _32902_ (.A1(_00774_),
    .A2(net1948),
    .B(_00776_),
    .Y(_15506_));
 OAI21x1_ASAP7_75t_R _32903_ (.A1(_15505_),
    .A2(_15506_),
    .B(net1955),
    .Y(_15507_));
 OR2x6_ASAP7_75t_R _32904_ (.A(net1942),
    .B(net1944),
    .Y(_15508_));
 OR3x1_ASAP7_75t_R _32905_ (.A(net1948),
    .B(net1950),
    .C(_15508_),
    .Y(_15509_));
 BUFx6f_ASAP7_75t_R _32906_ (.A(_15509_),
    .Y(_15510_));
 OR4x1_ASAP7_75t_R _32907_ (.A(_15031_),
    .B(_15037_),
    .C(_15167_),
    .D(_15510_),
    .Y(_15511_));
 OA21x2_ASAP7_75t_R _32908_ (.A1(_00778_),
    .A2(net1942),
    .B(_00780_),
    .Y(_15512_));
 OA21x2_ASAP7_75t_R _32909_ (.A1(net1945),
    .A2(_15512_),
    .B(_00782_),
    .Y(_15513_));
 OR3x1_ASAP7_75t_R _32910_ (.A(_00772_),
    .B(_00771_),
    .C(_15510_),
    .Y(_15514_));
 AND2x2_ASAP7_75t_R _32911_ (.A(_15513_),
    .B(_15514_),
    .Y(_15515_));
 AOI21x1_ASAP7_75t_R _32912_ (.A1(_15511_),
    .A2(_15515_),
    .B(net1939),
    .Y(_15516_));
 NOR2x1_ASAP7_75t_R _32913_ (.A(_15507_),
    .B(_15516_),
    .Y(_15517_));
 XNOR2x1_ASAP7_75t_R _32914_ (.B(_15517_),
    .Y(_15518_),
    .A(net1937));
 INVx5_ASAP7_75t_R _32915_ (.A(_15518_),
    .Y(\alu_adder_result_ex[13] ));
 OR2x2_ASAP7_75t_R _32916_ (.A(_15169_),
    .B(_15510_),
    .Y(_15519_));
 OA21x2_ASAP7_75t_R _32917_ (.A1(_00776_),
    .A2(net1950),
    .B(_00778_),
    .Y(_15520_));
 OA21x2_ASAP7_75t_R _32918_ (.A1(_00780_),
    .A2(net1945),
    .B(_00782_),
    .Y(_15521_));
 OA21x2_ASAP7_75t_R _32919_ (.A1(_15508_),
    .A2(_15520_),
    .B(_15521_),
    .Y(_15522_));
 OA21x2_ASAP7_75t_R _32920_ (.A1(_15176_),
    .A2(_15519_),
    .B(_15522_),
    .Y(_15523_));
 XNOR2x1_ASAP7_75t_R _32921_ (.B(_15523_),
    .Y(_15524_),
    .A(net1938));
 INVx4_ASAP7_75t_R _32922_ (.A(_15524_),
    .Y(\alu_adder_result_ex[12] ));
 AND2x2_ASAP7_75t_R _32923_ (.A(_14888_),
    .B(_01782_),
    .Y(_15525_));
 AO21x1_ASAP7_75t_R _32924_ (.A1(_13092_),
    .A2(_00816_),
    .B(_15525_),
    .Y(_15526_));
 OAI22x1_ASAP7_75t_R _32925_ (.A1(_00815_),
    .A2(_13102_),
    .B1(_15526_),
    .B2(_14975_),
    .Y(_15527_));
 INVx1_ASAP7_75t_R _32926_ (.A(_00824_),
    .Y(_15528_));
 NAND2x1_ASAP7_75t_R _32927_ (.A(_14697_),
    .B(_00822_),
    .Y(_15529_));
 OA211x2_ASAP7_75t_R _32928_ (.A1(_14360_),
    .A2(_15528_),
    .B(_15529_),
    .C(_14914_),
    .Y(_15530_));
 INVx2_ASAP7_75t_R _32929_ (.A(_00823_),
    .Y(_15531_));
 NAND2x1_ASAP7_75t_R _32930_ (.A(_14697_),
    .B(_00821_),
    .Y(_15532_));
 OA211x2_ASAP7_75t_R _32931_ (.A1(_14360_),
    .A2(_15531_),
    .B(_15532_),
    .C(_14463_),
    .Y(_15533_));
 OR3x1_ASAP7_75t_R _32932_ (.A(_13105_),
    .B(_15530_),
    .C(_15533_),
    .Y(_15534_));
 OA211x2_ASAP7_75t_R _32933_ (.A1(_14448_),
    .A2(_15527_),
    .B(_15534_),
    .C(_14466_),
    .Y(_15535_));
 INVx1_ASAP7_75t_R _32934_ (.A(_00820_),
    .Y(_15536_));
 NAND2x1_ASAP7_75t_R _32935_ (.A(_14502_),
    .B(_00818_),
    .Y(_15537_));
 OA211x2_ASAP7_75t_R _32936_ (.A1(_14496_),
    .A2(_15536_),
    .B(_15537_),
    .C(_14504_),
    .Y(_15538_));
 INVx1_ASAP7_75t_R _32937_ (.A(_00819_),
    .Y(_15539_));
 NAND2x1_ASAP7_75t_R _32938_ (.A(_14507_),
    .B(_00817_),
    .Y(_15540_));
 OA211x2_ASAP7_75t_R _32939_ (.A1(_14506_),
    .A2(_15539_),
    .B(_15540_),
    .C(_14509_),
    .Y(_15541_));
 OR3x1_ASAP7_75t_R _32940_ (.A(_14469_),
    .B(_15538_),
    .C(_15541_),
    .Y(_15542_));
 INVx1_ASAP7_75t_R _32941_ (.A(_00828_),
    .Y(_15543_));
 NAND2x1_ASAP7_75t_R _32942_ (.A(_13189_),
    .B(_00826_),
    .Y(_15544_));
 OA211x2_ASAP7_75t_R _32943_ (.A1(_14496_),
    .A2(_15543_),
    .B(_15544_),
    .C(_14504_),
    .Y(_15545_));
 INVx2_ASAP7_75t_R _32944_ (.A(_00827_),
    .Y(_15546_));
 NAND2x1_ASAP7_75t_R _32945_ (.A(_14517_),
    .B(_00825_),
    .Y(_15547_));
 OA211x2_ASAP7_75t_R _32946_ (.A1(_14516_),
    .A2(_15546_),
    .B(_15547_),
    .C(_14509_),
    .Y(_15548_));
 OR3x1_ASAP7_75t_R _32947_ (.A(_14353_),
    .B(_15545_),
    .C(_15548_),
    .Y(_15549_));
 AND3x1_ASAP7_75t_R _32948_ (.A(_14468_),
    .B(_15542_),
    .C(_15549_),
    .Y(_15550_));
 OR3x2_ASAP7_75t_R _32949_ (.A(_14447_),
    .B(_15535_),
    .C(_15550_),
    .Y(_15551_));
 INVx2_ASAP7_75t_R _32950_ (.A(_00836_),
    .Y(_15552_));
 NAND2x1_ASAP7_75t_R _32951_ (.A(_14450_),
    .B(_00834_),
    .Y(_15553_));
 OA211x2_ASAP7_75t_R _32952_ (.A1(_14366_),
    .A2(_15552_),
    .B(_15553_),
    .C(_14369_),
    .Y(_15554_));
 INVx2_ASAP7_75t_R _32953_ (.A(_00835_),
    .Y(_15555_));
 NAND2x1_ASAP7_75t_R _32954_ (.A(_14450_),
    .B(_00833_),
    .Y(_15556_));
 OA211x2_ASAP7_75t_R _32955_ (.A1(_14985_),
    .A2(_15555_),
    .B(_15556_),
    .C(_14372_),
    .Y(_15557_));
 OR3x1_ASAP7_75t_R _32956_ (.A(_14282_),
    .B(_15554_),
    .C(_15557_),
    .Y(_15558_));
 INVx1_ASAP7_75t_R _32957_ (.A(_00844_),
    .Y(_15559_));
 NAND2x1_ASAP7_75t_R _32958_ (.A(_14450_),
    .B(_00842_),
    .Y(_15560_));
 OA211x2_ASAP7_75t_R _32959_ (.A1(_14985_),
    .A2(_15559_),
    .B(_15560_),
    .C(_14369_),
    .Y(_15561_));
 INVx2_ASAP7_75t_R _32960_ (.A(_00843_),
    .Y(_15562_));
 NAND2x1_ASAP7_75t_R _32961_ (.A(_14752_),
    .B(_00841_),
    .Y(_15563_));
 OA211x2_ASAP7_75t_R _32962_ (.A1(_14985_),
    .A2(_15562_),
    .B(_15563_),
    .C(_14372_),
    .Y(_15564_));
 OR3x1_ASAP7_75t_R _32963_ (.A(_14291_),
    .B(_15561_),
    .C(_15564_),
    .Y(_15565_));
 AND3x1_ASAP7_75t_R _32964_ (.A(_14488_),
    .B(_15558_),
    .C(_15565_),
    .Y(_15566_));
 INVx2_ASAP7_75t_R _32965_ (.A(_00837_),
    .Y(_15567_));
 NOR2x1_ASAP7_75t_R _32966_ (.A(_13206_),
    .B(_00839_),
    .Y(_15568_));
 AO21x1_ASAP7_75t_R _32967_ (.A1(_14358_),
    .A2(_15567_),
    .B(_15568_),
    .Y(_15569_));
 INVx2_ASAP7_75t_R _32968_ (.A(_00840_),
    .Y(_15570_));
 NAND2x1_ASAP7_75t_R _32969_ (.A(_14277_),
    .B(_00838_),
    .Y(_15571_));
 OA211x2_ASAP7_75t_R _32970_ (.A1(_14293_),
    .A2(_15570_),
    .B(_15571_),
    .C(_14296_),
    .Y(_15572_));
 AO21x1_ASAP7_75t_R _32971_ (.A1(_13187_),
    .A2(_15569_),
    .B(_15572_),
    .Y(_15573_));
 INVx2_ASAP7_75t_R _32972_ (.A(_00832_),
    .Y(_15574_));
 NAND2x1_ASAP7_75t_R _32973_ (.A(_13165_),
    .B(_00830_),
    .Y(_15575_));
 OA211x2_ASAP7_75t_R _32974_ (.A1(_13097_),
    .A2(_15574_),
    .B(_15575_),
    .C(_14914_),
    .Y(_15576_));
 INVx1_ASAP7_75t_R _32975_ (.A(_00831_),
    .Y(_15577_));
 NAND2x1_ASAP7_75t_R _32976_ (.A(_14697_),
    .B(_00829_),
    .Y(_15578_));
 OA211x2_ASAP7_75t_R _32977_ (.A1(_14360_),
    .A2(_15577_),
    .B(_15578_),
    .C(_14463_),
    .Y(_15579_));
 OR3x1_ASAP7_75t_R _32978_ (.A(_13085_),
    .B(_15576_),
    .C(_15579_),
    .Y(_15580_));
 OA211x2_ASAP7_75t_R _32979_ (.A1(_13186_),
    .A2(_15573_),
    .B(_15580_),
    .C(_14466_),
    .Y(_15581_));
 OR3x2_ASAP7_75t_R _32980_ (.A(_13164_),
    .B(_15566_),
    .C(_15581_),
    .Y(_15582_));
 NAND2x2_ASAP7_75t_R _32981_ (.A(_15551_),
    .B(_15582_),
    .Y(_15583_));
 AO21x2_ASAP7_75t_R _32982_ (.A1(_01501_),
    .A2(_14968_),
    .B(_14967_),
    .Y(_15584_));
 OR2x6_ASAP7_75t_R _32983_ (.A(_01472_),
    .B(_14384_),
    .Y(_15585_));
 AOI22x1_ASAP7_75t_R _32984_ (.A1(_14446_),
    .A2(_15583_),
    .B1(_15584_),
    .B2(_15585_),
    .Y(_18625_));
 INVx3_ASAP7_75t_R _32985_ (.A(_18625_),
    .Y(_18623_));
 OR3x1_ASAP7_75t_R _32986_ (.A(_00180_),
    .B(_15104_),
    .C(_14650_),
    .Y(_15586_));
 OAI21x1_ASAP7_75t_R _32987_ (.A1(_14647_),
    .A2(_18623_),
    .B(_15586_),
    .Y(_18036_));
 BUFx12f_ASAP7_75t_R _32988_ (.A(_15312_),
    .Y(_15587_));
 BUFx6f_ASAP7_75t_R _32989_ (.A(_15352_),
    .Y(_15588_));
 BUFx12f_ASAP7_75t_R _32990_ (.A(_15485_),
    .Y(_15589_));
 AND2x2_ASAP7_75t_R _32991_ (.A(_15589_),
    .B(_01782_),
    .Y(_15590_));
 AO21x1_ASAP7_75t_R _32992_ (.A1(_15436_),
    .A2(_00816_),
    .B(_15590_),
    .Y(_15591_));
 BUFx6f_ASAP7_75t_R _32993_ (.A(_15273_),
    .Y(_15592_));
 BUFx12f_ASAP7_75t_R _32994_ (.A(_15592_),
    .Y(_15593_));
 BUFx12f_ASAP7_75t_R _32995_ (.A(_15593_),
    .Y(_15594_));
 OAI22x1_ASAP7_75t_R _32996_ (.A1(_00815_),
    .A2(_15435_),
    .B1(_15591_),
    .B2(_15594_),
    .Y(_15595_));
 BUFx6f_ASAP7_75t_R _32997_ (.A(_15278_),
    .Y(_15596_));
 BUFx6f_ASAP7_75t_R _32998_ (.A(_15258_),
    .Y(_15597_));
 BUFx6f_ASAP7_75t_R _32999_ (.A(_15597_),
    .Y(_15598_));
 NAND2x1_ASAP7_75t_R _33000_ (.A(_15291_),
    .B(_00822_),
    .Y(_15599_));
 BUFx6f_ASAP7_75t_R _33001_ (.A(_15266_),
    .Y(_15600_));
 OA211x2_ASAP7_75t_R _33002_ (.A1(_15598_),
    .A2(_15528_),
    .B(_15599_),
    .C(_15600_),
    .Y(_15601_));
 NAND2x1_ASAP7_75t_R _33003_ (.A(_15347_),
    .B(_00821_),
    .Y(_15602_));
 OA211x2_ASAP7_75t_R _33004_ (.A1(_15598_),
    .A2(_15531_),
    .B(_15602_),
    .C(_15338_),
    .Y(_15603_));
 OR3x1_ASAP7_75t_R _33005_ (.A(_15596_),
    .B(_15601_),
    .C(_15603_),
    .Y(_15604_));
 OA21x2_ASAP7_75t_R _33006_ (.A1(_15588_),
    .A2(_15595_),
    .B(_15604_),
    .Y(_15605_));
 NAND2x1_ASAP7_75t_R _33007_ (.A(_15326_),
    .B(_00818_),
    .Y(_15606_));
 OA211x2_ASAP7_75t_R _33008_ (.A1(_15471_),
    .A2(_15536_),
    .B(_15606_),
    .C(_15349_),
    .Y(_15607_));
 NAND2x1_ASAP7_75t_R _33009_ (.A(_15262_),
    .B(_00817_),
    .Y(_15608_));
 OA211x2_ASAP7_75t_R _33010_ (.A1(_15471_),
    .A2(_15539_),
    .B(_15608_),
    .C(_15456_),
    .Y(_15609_));
 OR3x1_ASAP7_75t_R _33011_ (.A(_15318_),
    .B(_15607_),
    .C(_15609_),
    .Y(_15610_));
 NAND2x1_ASAP7_75t_R _33012_ (.A(_15326_),
    .B(_00826_),
    .Y(_15611_));
 OA211x2_ASAP7_75t_R _33013_ (.A1(_15471_),
    .A2(_15543_),
    .B(_15611_),
    .C(_15349_),
    .Y(_15612_));
 NAND2x1_ASAP7_75t_R _33014_ (.A(_15262_),
    .B(_00825_),
    .Y(_15613_));
 OA211x2_ASAP7_75t_R _33015_ (.A1(_15346_),
    .A2(_15546_),
    .B(_15613_),
    .C(_15456_),
    .Y(_15614_));
 OR3x1_ASAP7_75t_R _33016_ (.A(_15475_),
    .B(_15612_),
    .C(_15614_),
    .Y(_15615_));
 AND3x1_ASAP7_75t_R _33017_ (.A(_15317_),
    .B(_15610_),
    .C(_15615_),
    .Y(_15616_));
 AO21x1_ASAP7_75t_R _33018_ (.A1(_15587_),
    .A2(_15605_),
    .B(_15616_),
    .Y(_15617_));
 BUFx12f_ASAP7_75t_R _33019_ (.A(_15261_),
    .Y(_15618_));
 NAND2x1_ASAP7_75t_R _33020_ (.A(_15618_),
    .B(_00834_),
    .Y(_15619_));
 BUFx6f_ASAP7_75t_R _33021_ (.A(_15266_),
    .Y(_15620_));
 OA211x2_ASAP7_75t_R _33022_ (.A1(_15269_),
    .A2(_15552_),
    .B(_15619_),
    .C(_15620_),
    .Y(_15621_));
 BUFx6f_ASAP7_75t_R _33023_ (.A(_15259_),
    .Y(_15622_));
 NAND2x1_ASAP7_75t_R _33024_ (.A(_15618_),
    .B(_00833_),
    .Y(_15623_));
 OA211x2_ASAP7_75t_R _33025_ (.A1(_15622_),
    .A2(_15555_),
    .B(_15623_),
    .C(_15283_),
    .Y(_15624_));
 OR3x1_ASAP7_75t_R _33026_ (.A(_15255_),
    .B(_15621_),
    .C(_15624_),
    .Y(_15625_));
 NAND2x1_ASAP7_75t_R _33027_ (.A(_15618_),
    .B(_00842_),
    .Y(_15626_));
 OA211x2_ASAP7_75t_R _33028_ (.A1(_15269_),
    .A2(_15559_),
    .B(_15626_),
    .C(_15620_),
    .Y(_15627_));
 NAND2x1_ASAP7_75t_R _33029_ (.A(_15340_),
    .B(_00841_),
    .Y(_15628_));
 OA211x2_ASAP7_75t_R _33030_ (.A1(_15622_),
    .A2(_15562_),
    .B(_15628_),
    .C(_15283_),
    .Y(_15629_));
 OR3x1_ASAP7_75t_R _33031_ (.A(_15279_),
    .B(_15627_),
    .C(_15629_),
    .Y(_15630_));
 AND3x1_ASAP7_75t_R _33032_ (.A(_15253_),
    .B(_15625_),
    .C(_15630_),
    .Y(_15631_));
 BUFx6f_ASAP7_75t_R _33033_ (.A(_15301_),
    .Y(_15632_));
 BUFx6f_ASAP7_75t_R _33034_ (.A(_15632_),
    .Y(_15633_));
 NOR2x1_ASAP7_75t_R _33035_ (.A(_15445_),
    .B(_00839_),
    .Y(_15634_));
 AO21x1_ASAP7_75t_R _33036_ (.A1(_15633_),
    .A2(_15567_),
    .B(_15634_),
    .Y(_15635_));
 NAND2x1_ASAP7_75t_R _33037_ (.A(_15454_),
    .B(_00838_),
    .Y(_15636_));
 OA211x2_ASAP7_75t_R _33038_ (.A1(_15320_),
    .A2(_15570_),
    .B(_15636_),
    .C(_15267_),
    .Y(_15637_));
 AO21x1_ASAP7_75t_R _33039_ (.A1(_15339_),
    .A2(_15635_),
    .B(_15637_),
    .Y(_15638_));
 NAND2x1_ASAP7_75t_R _33040_ (.A(_15489_),
    .B(_00830_),
    .Y(_15639_));
 OA211x2_ASAP7_75t_R _33041_ (.A1(_15307_),
    .A2(_15574_),
    .B(_15639_),
    .C(_15304_),
    .Y(_15640_));
 NAND2x1_ASAP7_75t_R _33042_ (.A(_15597_),
    .B(_00829_),
    .Y(_15641_));
 OA211x2_ASAP7_75t_R _33043_ (.A1(_15307_),
    .A2(_15577_),
    .B(_15641_),
    .C(_15309_),
    .Y(_15642_));
 OR3x1_ASAP7_75t_R _33044_ (.A(_15352_),
    .B(_15640_),
    .C(_15642_),
    .Y(_15643_));
 OA211x2_ASAP7_75t_R _33045_ (.A1(_15337_),
    .A2(_15638_),
    .B(_15643_),
    .C(_15313_),
    .Y(_15644_));
 OR3x2_ASAP7_75t_R _33046_ (.A(_15316_),
    .B(_15631_),
    .C(_15644_),
    .Y(_15645_));
 OAI21x1_ASAP7_75t_R _33047_ (.A1(_15434_),
    .A2(_15617_),
    .B(_15645_),
    .Y(_15646_));
 OA211x2_ASAP7_75t_R _33048_ (.A1(_14534_),
    .A2(_15366_),
    .B(_15369_),
    .C(_15370_),
    .Y(_15647_));
 AOI21x1_ASAP7_75t_R _33049_ (.A1(_15250_),
    .A2(net1947),
    .B(_15647_),
    .Y(_18624_));
 INVx1_ASAP7_75t_R _33050_ (.A(_18624_),
    .Y(_18622_));
 AND2x2_ASAP7_75t_R _33051_ (.A(_13192_),
    .B(_01781_),
    .Y(_15648_));
 AO21x1_ASAP7_75t_R _33052_ (.A1(_14285_),
    .A2(_00848_),
    .B(_15648_),
    .Y(_15649_));
 OAI22x1_ASAP7_75t_R _33053_ (.A1(_00847_),
    .A2(_13101_),
    .B1(_15649_),
    .B2(_13089_),
    .Y(_15650_));
 INVx2_ASAP7_75t_R _33054_ (.A(_00856_),
    .Y(_15651_));
 NAND2x1_ASAP7_75t_R _33055_ (.A(_13199_),
    .B(_00854_),
    .Y(_15652_));
 OA211x2_ASAP7_75t_R _33056_ (.A1(_14298_),
    .A2(_15651_),
    .B(_15652_),
    .C(_13139_),
    .Y(_15653_));
 INVx2_ASAP7_75t_R _33057_ (.A(_00855_),
    .Y(_15654_));
 NAND2x1_ASAP7_75t_R _33058_ (.A(_14300_),
    .B(_00853_),
    .Y(_15655_));
 OA211x2_ASAP7_75t_R _33059_ (.A1(_14403_),
    .A2(_15654_),
    .B(_15655_),
    .C(_13148_),
    .Y(_15656_));
 OR3x1_ASAP7_75t_R _33060_ (.A(_13152_),
    .B(_15653_),
    .C(_15656_),
    .Y(_15657_));
 OA211x2_ASAP7_75t_R _33061_ (.A1(_14282_),
    .A2(_15650_),
    .B(_15657_),
    .C(_13124_),
    .Y(_15658_));
 INVx2_ASAP7_75t_R _33062_ (.A(_00852_),
    .Y(_15659_));
 NAND2x1_ASAP7_75t_R _33063_ (.A(_14319_),
    .B(_00850_),
    .Y(_15660_));
 OA211x2_ASAP7_75t_R _33064_ (.A1(_13211_),
    .A2(_15659_),
    .B(_15660_),
    .C(_14362_),
    .Y(_15661_));
 INVx2_ASAP7_75t_R _33065_ (.A(_00851_),
    .Y(_15662_));
 NAND2x1_ASAP7_75t_R _33066_ (.A(_14319_),
    .B(_00849_),
    .Y(_15663_));
 OA211x2_ASAP7_75t_R _33067_ (.A1(_13211_),
    .A2(_15662_),
    .B(_15663_),
    .C(_14322_),
    .Y(_15664_));
 OR3x1_ASAP7_75t_R _33068_ (.A(_14308_),
    .B(_15661_),
    .C(_15664_),
    .Y(_15665_));
 INVx2_ASAP7_75t_R _33069_ (.A(_00860_),
    .Y(_15666_));
 NAND2x1_ASAP7_75t_R _33070_ (.A(_14319_),
    .B(_00858_),
    .Y(_15667_));
 OA211x2_ASAP7_75t_R _33071_ (.A1(_13211_),
    .A2(_15666_),
    .B(_15667_),
    .C(_14362_),
    .Y(_15668_));
 INVx2_ASAP7_75t_R _33072_ (.A(_00859_),
    .Y(_15669_));
 NAND2x1_ASAP7_75t_R _33073_ (.A(_14319_),
    .B(_00857_),
    .Y(_15670_));
 OA211x2_ASAP7_75t_R _33074_ (.A1(_13211_),
    .A2(_15669_),
    .B(_15670_),
    .C(_14322_),
    .Y(_15671_));
 OR3x1_ASAP7_75t_R _33075_ (.A(_14326_),
    .B(_15668_),
    .C(_15671_),
    .Y(_15672_));
 AND3x1_ASAP7_75t_R _33076_ (.A(_14807_),
    .B(_15665_),
    .C(_15672_),
    .Y(_15673_));
 OR3x2_ASAP7_75t_R _33077_ (.A(_13081_),
    .B(_15658_),
    .C(_15673_),
    .Y(_15674_));
 BUFx6f_ASAP7_75t_R _33078_ (.A(_13188_),
    .Y(_15675_));
 INVx2_ASAP7_75t_R _33079_ (.A(_00868_),
    .Y(_15676_));
 NAND2x1_ASAP7_75t_R _33080_ (.A(_14460_),
    .B(_00866_),
    .Y(_15677_));
 OA211x2_ASAP7_75t_R _33081_ (.A1(_15675_),
    .A2(_15676_),
    .B(_15677_),
    .C(_14362_),
    .Y(_15678_));
 INVx2_ASAP7_75t_R _33082_ (.A(_00867_),
    .Y(_15679_));
 NAND2x1_ASAP7_75t_R _33083_ (.A(_14319_),
    .B(_00865_),
    .Y(_15680_));
 OA211x2_ASAP7_75t_R _33084_ (.A1(_13118_),
    .A2(_15679_),
    .B(_15680_),
    .C(_13088_),
    .Y(_15681_));
 OR3x1_ASAP7_75t_R _33085_ (.A(_14308_),
    .B(_15678_),
    .C(_15681_),
    .Y(_15682_));
 INVx1_ASAP7_75t_R _33086_ (.A(_00876_),
    .Y(_15683_));
 NAND2x1_ASAP7_75t_R _33087_ (.A(_14460_),
    .B(_00874_),
    .Y(_15684_));
 OA211x2_ASAP7_75t_R _33088_ (.A1(_13118_),
    .A2(_15683_),
    .B(_15684_),
    .C(_14362_),
    .Y(_15685_));
 INVx2_ASAP7_75t_R _33089_ (.A(_00875_),
    .Y(_15686_));
 NAND2x1_ASAP7_75t_R _33090_ (.A(_14319_),
    .B(_00873_),
    .Y(_15687_));
 OA211x2_ASAP7_75t_R _33091_ (.A1(_13211_),
    .A2(_15686_),
    .B(_15687_),
    .C(_13088_),
    .Y(_15688_));
 OR3x1_ASAP7_75t_R _33092_ (.A(_14326_),
    .B(_15685_),
    .C(_15688_),
    .Y(_15689_));
 AND3x1_ASAP7_75t_R _33093_ (.A(_14807_),
    .B(_15682_),
    .C(_15689_),
    .Y(_15690_));
 INVx2_ASAP7_75t_R _33094_ (.A(_00869_),
    .Y(_15691_));
 NOR2x1_ASAP7_75t_R _33095_ (.A(_13142_),
    .B(_00871_),
    .Y(_15692_));
 AO21x1_ASAP7_75t_R _33096_ (.A1(_14888_),
    .A2(_15691_),
    .B(_15692_),
    .Y(_15693_));
 INVx2_ASAP7_75t_R _33097_ (.A(_00872_),
    .Y(_15694_));
 NAND2x1_ASAP7_75t_R _33098_ (.A(_13096_),
    .B(_00870_),
    .Y(_15695_));
 OA211x2_ASAP7_75t_R _33099_ (.A1(_14470_),
    .A2(_15694_),
    .B(_15695_),
    .C(_14762_),
    .Y(_15696_));
 AO21x1_ASAP7_75t_R _33100_ (.A1(_13089_),
    .A2(_15693_),
    .B(_15696_),
    .Y(_15697_));
 INVx1_ASAP7_75t_R _33101_ (.A(_00864_),
    .Y(_15698_));
 NAND2x1_ASAP7_75t_R _33102_ (.A(_14300_),
    .B(_00862_),
    .Y(_15699_));
 OA211x2_ASAP7_75t_R _33103_ (.A1(_14403_),
    .A2(_15698_),
    .B(_15699_),
    .C(_14295_),
    .Y(_15700_));
 INVx1_ASAP7_75t_R _33104_ (.A(_00863_),
    .Y(_15701_));
 NAND2x1_ASAP7_75t_R _33105_ (.A(_13145_),
    .B(_00861_),
    .Y(_15702_));
 OA211x2_ASAP7_75t_R _33106_ (.A1(_14437_),
    .A2(_15701_),
    .B(_15702_),
    .C(_13148_),
    .Y(_15703_));
 OR3x1_ASAP7_75t_R _33107_ (.A(_13084_),
    .B(_15700_),
    .C(_15703_),
    .Y(_15704_));
 OA211x2_ASAP7_75t_R _33108_ (.A1(_14291_),
    .A2(_15697_),
    .B(_15704_),
    .C(_13124_),
    .Y(_15705_));
 OR3x2_ASAP7_75t_R _33109_ (.A(_13163_),
    .B(_15690_),
    .C(_15705_),
    .Y(_15706_));
 AND2x6_ASAP7_75t_R _33110_ (.A(_15674_),
    .B(_15706_),
    .Y(_15707_));
 BUFx6f_ASAP7_75t_R _33111_ (.A(_01500_),
    .Y(_15708_));
 AND2x2_ASAP7_75t_R _33112_ (.A(_01471_),
    .B(_14380_),
    .Y(_15709_));
 OAI22x1_ASAP7_75t_R _33113_ (.A1(_15708_),
    .A2(_15100_),
    .B1(_14384_),
    .B2(_15709_),
    .Y(_15710_));
 OA21x2_ASAP7_75t_R _33114_ (.A1(_14709_),
    .A2(_15707_),
    .B(_15710_),
    .Y(_15711_));
 BUFx3_ASAP7_75t_R _33115_ (.A(_15711_),
    .Y(_18630_));
 INVx3_ASAP7_75t_R _33116_ (.A(_18630_),
    .Y(_18628_));
 OR3x1_ASAP7_75t_R _33117_ (.A(_00187_),
    .B(_15104_),
    .C(_14649_),
    .Y(_15712_));
 OAI21x1_ASAP7_75t_R _33118_ (.A1(_14646_),
    .A2(_18628_),
    .B(_15712_),
    .Y(_18038_));
 AND2x2_ASAP7_75t_R _33119_ (.A(_15441_),
    .B(_01781_),
    .Y(_15713_));
 AO21x1_ASAP7_75t_R _33120_ (.A1(_15436_),
    .A2(_00848_),
    .B(_15713_),
    .Y(_15714_));
 OAI22x1_ASAP7_75t_R _33121_ (.A1(_00847_),
    .A2(_15435_),
    .B1(_15714_),
    .B2(_15296_),
    .Y(_15715_));
 NAND2x1_ASAP7_75t_R _33122_ (.A(_15347_),
    .B(_00854_),
    .Y(_15716_));
 OA211x2_ASAP7_75t_R _33123_ (.A1(_15490_),
    .A2(_15651_),
    .B(_15716_),
    .C(_15469_),
    .Y(_15717_));
 NAND2x1_ASAP7_75t_R _33124_ (.A(_15347_),
    .B(_00853_),
    .Y(_15718_));
 OA211x2_ASAP7_75t_R _33125_ (.A1(_15490_),
    .A2(_15654_),
    .B(_15718_),
    .C(_15338_),
    .Y(_15719_));
 OR3x1_ASAP7_75t_R _33126_ (.A(_15475_),
    .B(_15717_),
    .C(_15719_),
    .Y(_15720_));
 OA21x2_ASAP7_75t_R _33127_ (.A1(_15588_),
    .A2(_15715_),
    .B(_15720_),
    .Y(_15721_));
 NAND2x1_ASAP7_75t_R _33128_ (.A(_15451_),
    .B(_00850_),
    .Y(_15722_));
 OA211x2_ASAP7_75t_R _33129_ (.A1(_15346_),
    .A2(_15659_),
    .B(_15722_),
    .C(_15323_),
    .Y(_15723_));
 NAND2x1_ASAP7_75t_R _33130_ (.A(_15454_),
    .B(_00849_),
    .Y(_15724_));
 OA211x2_ASAP7_75t_R _33131_ (.A1(_15450_),
    .A2(_15662_),
    .B(_15724_),
    .C(_15456_),
    .Y(_15725_));
 OR3x1_ASAP7_75t_R _33132_ (.A(_15318_),
    .B(_15723_),
    .C(_15725_),
    .Y(_15726_));
 NAND2x1_ASAP7_75t_R _33133_ (.A(_15451_),
    .B(_00858_),
    .Y(_15727_));
 OA211x2_ASAP7_75t_R _33134_ (.A1(_15450_),
    .A2(_15666_),
    .B(_15727_),
    .C(_15323_),
    .Y(_15728_));
 NAND2x1_ASAP7_75t_R _33135_ (.A(_15454_),
    .B(_00857_),
    .Y(_15729_));
 OA211x2_ASAP7_75t_R _33136_ (.A1(_15320_),
    .A2(_15669_),
    .B(_15729_),
    .C(_15275_),
    .Y(_15730_));
 OR3x1_ASAP7_75t_R _33137_ (.A(_15475_),
    .B(_15728_),
    .C(_15730_),
    .Y(_15731_));
 AND3x1_ASAP7_75t_R _33138_ (.A(_15317_),
    .B(_15726_),
    .C(_15731_),
    .Y(_15732_));
 AO21x1_ASAP7_75t_R _33139_ (.A1(_15587_),
    .A2(_15721_),
    .B(_15732_),
    .Y(_15733_));
 BUFx6f_ASAP7_75t_R _33140_ (.A(_15301_),
    .Y(_15734_));
 NAND2x1_ASAP7_75t_R _33141_ (.A(_15734_),
    .B(_00866_),
    .Y(_15735_));
 OA211x2_ASAP7_75t_R _33142_ (.A1(_15486_),
    .A2(_15676_),
    .B(_15735_),
    .C(_15620_),
    .Y(_15736_));
 NAND2x1_ASAP7_75t_R _33143_ (.A(_15483_),
    .B(_00865_),
    .Y(_15737_));
 OA211x2_ASAP7_75t_R _33144_ (.A1(_15486_),
    .A2(_15679_),
    .B(_15737_),
    .C(_15497_),
    .Y(_15738_));
 OR3x1_ASAP7_75t_R _33145_ (.A(_15255_),
    .B(_15736_),
    .C(_15738_),
    .Y(_15739_));
 NAND2x1_ASAP7_75t_R _33146_ (.A(_15483_),
    .B(_00874_),
    .Y(_15740_));
 OA211x2_ASAP7_75t_R _33147_ (.A1(_15486_),
    .A2(_15683_),
    .B(_15740_),
    .C(_15443_),
    .Y(_15741_));
 NAND2x1_ASAP7_75t_R _33148_ (.A(_15483_),
    .B(_00873_),
    .Y(_15742_));
 OA211x2_ASAP7_75t_R _33149_ (.A1(_15589_),
    .A2(_15686_),
    .B(_15742_),
    .C(_15497_),
    .Y(_15743_));
 OR3x1_ASAP7_75t_R _33150_ (.A(_15298_),
    .B(_15741_),
    .C(_15743_),
    .Y(_15744_));
 AND3x1_ASAP7_75t_R _33151_ (.A(_15253_),
    .B(_15739_),
    .C(_15744_),
    .Y(_15745_));
 NOR2x1_ASAP7_75t_R _33152_ (.A(_15307_),
    .B(_00871_),
    .Y(_15746_));
 AO21x1_ASAP7_75t_R _33153_ (.A1(_15598_),
    .A2(_15691_),
    .B(_15746_),
    .Y(_15747_));
 NAND2x1_ASAP7_75t_R _33154_ (.A(_15618_),
    .B(_00870_),
    .Y(_15748_));
 OA211x2_ASAP7_75t_R _33155_ (.A1(_15622_),
    .A2(_15694_),
    .B(_15748_),
    .C(_15620_),
    .Y(_15749_));
 AO21x1_ASAP7_75t_R _33156_ (.A1(_15593_),
    .A2(_15747_),
    .B(_15749_),
    .Y(_15750_));
 NAND2x1_ASAP7_75t_R _33157_ (.A(_15319_),
    .B(_00862_),
    .Y(_15751_));
 BUFx6f_ASAP7_75t_R _33158_ (.A(_15265_),
    .Y(_15752_));
 OA211x2_ASAP7_75t_R _33159_ (.A1(_15437_),
    .A2(_15698_),
    .B(_15751_),
    .C(_15752_),
    .Y(_15753_));
 NAND2x1_ASAP7_75t_R _33160_ (.A(_15319_),
    .B(_00861_),
    .Y(_15754_));
 OA211x2_ASAP7_75t_R _33161_ (.A1(_15291_),
    .A2(_15701_),
    .B(_15754_),
    .C(_15592_),
    .Y(_15755_));
 OR3x1_ASAP7_75t_R _33162_ (.A(_15287_),
    .B(_15753_),
    .C(_15755_),
    .Y(_15756_));
 OA211x2_ASAP7_75t_R _33163_ (.A1(_15337_),
    .A2(_15750_),
    .B(_15756_),
    .C(_15313_),
    .Y(_15757_));
 OR3x1_ASAP7_75t_R _33164_ (.A(_15316_),
    .B(_15745_),
    .C(_15757_),
    .Y(_15758_));
 OAI21x1_ASAP7_75t_R _33165_ (.A1(_15434_),
    .A2(_15733_),
    .B(_15758_),
    .Y(_15759_));
 OA211x2_ASAP7_75t_R _33166_ (.A1(_14289_),
    .A2(_15366_),
    .B(_15369_),
    .C(_15370_),
    .Y(_15760_));
 AOI21x1_ASAP7_75t_R _33167_ (.A1(_15250_),
    .A2(_15759_),
    .B(_15760_),
    .Y(_18629_));
 INVx1_ASAP7_75t_R _33168_ (.A(_18629_),
    .Y(_18627_));
 OR2x2_ASAP7_75t_R _33169_ (.A(net1937),
    .B(_00845_),
    .Y(_15761_));
 OA21x2_ASAP7_75t_R _33170_ (.A1(_00846_),
    .A2(net1935),
    .B(_00878_),
    .Y(_15762_));
 OA21x2_ASAP7_75t_R _33171_ (.A1(_15517_),
    .A2(_15761_),
    .B(_15762_),
    .Y(_15763_));
 XNOR2x1_ASAP7_75t_R _33172_ (.B(_15763_),
    .Y(_15764_),
    .A(net1941));
 INVx5_ASAP7_75t_R _33173_ (.A(_15764_),
    .Y(\alu_adder_result_ex[15] ));
 OA21x2_ASAP7_75t_R _33174_ (.A1(net1938),
    .A2(_15521_),
    .B(net1955),
    .Y(_15765_));
 OA21x2_ASAP7_75t_R _33175_ (.A1(net1937),
    .A2(_15765_),
    .B(_00846_),
    .Y(_15766_));
 INVx1_ASAP7_75t_R _33176_ (.A(_15766_),
    .Y(_15767_));
 OR3x2_ASAP7_75t_R _33177_ (.A(net1939),
    .B(net1937),
    .C(_15508_),
    .Y(_15768_));
 AOI211x1_ASAP7_75t_R _33178_ (.A1(_15241_),
    .A2(_15243_),
    .B(_15768_),
    .C(_15246_),
    .Y(_15769_));
 OA21x2_ASAP7_75t_R _33179_ (.A1(_15767_),
    .A2(_15769_),
    .B(net1936),
    .Y(_15770_));
 NOR3x1_ASAP7_75t_R _33180_ (.A(net1936),
    .B(_15767_),
    .C(_15769_),
    .Y(_15771_));
 NOR2x2_ASAP7_75t_R _33181_ (.A(_15770_),
    .B(_15771_),
    .Y(_15772_));
 INVx4_ASAP7_75t_R _33182_ (.A(_15772_),
    .Y(\alu_adder_result_ex[14] ));
 INVx2_ASAP7_75t_R _33183_ (.A(_00901_),
    .Y(_15773_));
 NOR2x1_ASAP7_75t_R _33184_ (.A(_14858_),
    .B(_00903_),
    .Y(_15774_));
 AO21x1_ASAP7_75t_R _33185_ (.A1(_14293_),
    .A2(_15773_),
    .B(_15774_),
    .Y(_15775_));
 INVx2_ASAP7_75t_R _33186_ (.A(_00904_),
    .Y(_15776_));
 NAND2x1_ASAP7_75t_R _33187_ (.A(_14678_),
    .B(_00902_),
    .Y(_15777_));
 OA211x2_ASAP7_75t_R _33188_ (.A1(_14717_),
    .A2(_15776_),
    .B(_15777_),
    .C(_14914_),
    .Y(_15778_));
 AO21x1_ASAP7_75t_R _33189_ (.A1(_14710_),
    .A2(_15775_),
    .B(_15778_),
    .Y(_15779_));
 INVx2_ASAP7_75t_R _33190_ (.A(_00896_),
    .Y(_15780_));
 NAND2x1_ASAP7_75t_R _33191_ (.A(_14292_),
    .B(_00894_),
    .Y(_15781_));
 OA211x2_ASAP7_75t_R _33192_ (.A1(_14320_),
    .A2(_15780_),
    .B(_15781_),
    .C(_14458_),
    .Y(_15782_));
 INVx1_ASAP7_75t_R _33193_ (.A(_00895_),
    .Y(_15783_));
 NAND2x1_ASAP7_75t_R _33194_ (.A(_14298_),
    .B(_00893_),
    .Y(_15784_));
 OA211x2_ASAP7_75t_R _33195_ (.A1(_14333_),
    .A2(_15783_),
    .B(_15784_),
    .C(_14743_),
    .Y(_15785_));
 OA21x2_ASAP7_75t_R _33196_ (.A1(_15782_),
    .A2(_15785_),
    .B(_13105_),
    .Y(_15786_));
 AO21x1_ASAP7_75t_R _33197_ (.A1(_14448_),
    .A2(_15779_),
    .B(_15786_),
    .Y(_15787_));
 INVx2_ASAP7_75t_R _33198_ (.A(_00900_),
    .Y(_15788_));
 NAND2x1_ASAP7_75t_R _33199_ (.A(_13205_),
    .B(_00898_),
    .Y(_15789_));
 OA211x2_ASAP7_75t_R _33200_ (.A1(_14367_),
    .A2(_15788_),
    .B(_15789_),
    .C(_14729_),
    .Y(_15790_));
 INVx2_ASAP7_75t_R _33201_ (.A(_00899_),
    .Y(_15791_));
 NAND2x1_ASAP7_75t_R _33202_ (.A(_13205_),
    .B(_00897_),
    .Y(_15792_));
 OA211x2_ASAP7_75t_R _33203_ (.A1(_14367_),
    .A2(_15791_),
    .B(_15792_),
    .C(_14765_),
    .Y(_15793_));
 OR3x1_ASAP7_75t_R _33204_ (.A(_14737_),
    .B(_15790_),
    .C(_15793_),
    .Y(_15794_));
 INVx1_ASAP7_75t_R _33205_ (.A(_00908_),
    .Y(_15795_));
 NAND2x1_ASAP7_75t_R _33206_ (.A(_13205_),
    .B(_00906_),
    .Y(_15796_));
 OA211x2_ASAP7_75t_R _33207_ (.A1(_14367_),
    .A2(_15795_),
    .B(_15796_),
    .C(_14729_),
    .Y(_15797_));
 INVx2_ASAP7_75t_R _33208_ (.A(_00907_),
    .Y(_15798_));
 NAND2x1_ASAP7_75t_R _33209_ (.A(_13205_),
    .B(_00905_),
    .Y(_15799_));
 OA211x2_ASAP7_75t_R _33210_ (.A1(_14450_),
    .A2(_15798_),
    .B(_15799_),
    .C(_14765_),
    .Y(_15800_));
 OR3x1_ASAP7_75t_R _33211_ (.A(_13185_),
    .B(_15797_),
    .C(_15800_),
    .Y(_15801_));
 AND3x1_ASAP7_75t_R _33212_ (.A(_14807_),
    .B(_15794_),
    .C(_15801_),
    .Y(_15802_));
 AO21x1_ASAP7_75t_R _33213_ (.A1(_14778_),
    .A2(_15787_),
    .B(_15802_),
    .Y(_15803_));
 AND2x2_ASAP7_75t_R _33214_ (.A(_13192_),
    .B(_01780_),
    .Y(_15804_));
 AO21x1_ASAP7_75t_R _33215_ (.A1(_14285_),
    .A2(_00880_),
    .B(_15804_),
    .Y(_15805_));
 OAI22x1_ASAP7_75t_R _33216_ (.A1(_00879_),
    .A2(_13101_),
    .B1(_15805_),
    .B2(_14710_),
    .Y(_15806_));
 INVx1_ASAP7_75t_R _33217_ (.A(_00888_),
    .Y(_15807_));
 NAND2x1_ASAP7_75t_R _33218_ (.A(_14755_),
    .B(_00886_),
    .Y(_15808_));
 OA211x2_ASAP7_75t_R _33219_ (.A1(_14292_),
    .A2(_15807_),
    .B(_15808_),
    .C(_13139_),
    .Y(_15809_));
 INVx1_ASAP7_75t_R _33220_ (.A(_00887_),
    .Y(_15810_));
 NAND2x1_ASAP7_75t_R _33221_ (.A(_14755_),
    .B(_00885_),
    .Y(_15811_));
 OA211x2_ASAP7_75t_R _33222_ (.A1(_14298_),
    .A2(_15810_),
    .B(_15811_),
    .C(_13173_),
    .Y(_15812_));
 OR3x1_ASAP7_75t_R _33223_ (.A(_13152_),
    .B(_15809_),
    .C(_15812_),
    .Y(_15813_));
 OA211x2_ASAP7_75t_R _33224_ (.A1(_13131_),
    .A2(_15806_),
    .B(_15813_),
    .C(_14428_),
    .Y(_15814_));
 INVx1_ASAP7_75t_R _33225_ (.A(_00884_),
    .Y(_15815_));
 NAND2x1_ASAP7_75t_R _33226_ (.A(_14760_),
    .B(_00882_),
    .Y(_15816_));
 OA211x2_ASAP7_75t_R _33227_ (.A1(_14317_),
    .A2(_15815_),
    .B(_15816_),
    .C(_14762_),
    .Y(_15817_));
 INVx1_ASAP7_75t_R _33228_ (.A(_00883_),
    .Y(_15818_));
 NAND2x1_ASAP7_75t_R _33229_ (.A(_14391_),
    .B(_00881_),
    .Y(_15819_));
 OA211x2_ASAP7_75t_R _33230_ (.A1(_13110_),
    .A2(_15818_),
    .B(_15819_),
    .C(_14765_),
    .Y(_15820_));
 OR3x1_ASAP7_75t_R _33231_ (.A(_14308_),
    .B(_15817_),
    .C(_15820_),
    .Y(_15821_));
 INVx1_ASAP7_75t_R _33232_ (.A(_00892_),
    .Y(_15822_));
 NAND2x1_ASAP7_75t_R _33233_ (.A(_14760_),
    .B(_00890_),
    .Y(_15823_));
 OA211x2_ASAP7_75t_R _33234_ (.A1(_13110_),
    .A2(_15822_),
    .B(_15823_),
    .C(_14762_),
    .Y(_15824_));
 INVx1_ASAP7_75t_R _33235_ (.A(_00891_),
    .Y(_15825_));
 NAND2x1_ASAP7_75t_R _33236_ (.A(_14391_),
    .B(_00889_),
    .Y(_15826_));
 OA211x2_ASAP7_75t_R _33237_ (.A1(_15675_),
    .A2(_15825_),
    .B(_15826_),
    .C(_13088_),
    .Y(_15827_));
 OR3x1_ASAP7_75t_R _33238_ (.A(_13185_),
    .B(_15824_),
    .C(_15827_),
    .Y(_15828_));
 AND3x1_ASAP7_75t_R _33239_ (.A(_14807_),
    .B(_15821_),
    .C(_15828_),
    .Y(_15829_));
 OR3x1_ASAP7_75t_R _33240_ (.A(_14447_),
    .B(_15814_),
    .C(_15829_),
    .Y(_15830_));
 OA21x2_ASAP7_75t_R _33241_ (.A1(_13164_),
    .A2(_15803_),
    .B(_15830_),
    .Y(_15831_));
 BUFx6f_ASAP7_75t_R _33242_ (.A(_01499_),
    .Y(_15832_));
 AND2x2_ASAP7_75t_R _33243_ (.A(_01470_),
    .B(_14380_),
    .Y(_15833_));
 OAI22x1_ASAP7_75t_R _33244_ (.A1(_15832_),
    .A2(_15100_),
    .B1(_14384_),
    .B2(_15833_),
    .Y(_15834_));
 OA21x2_ASAP7_75t_R _33245_ (.A1(_14377_),
    .A2(_15831_),
    .B(_15834_),
    .Y(_15835_));
 BUFx6f_ASAP7_75t_R _33246_ (.A(_15835_),
    .Y(_18635_));
 INVx3_ASAP7_75t_R _33247_ (.A(_18635_),
    .Y(_18633_));
 BUFx6f_ASAP7_75t_R _33248_ (.A(_00063_),
    .Y(_15836_));
 OR3x1_ASAP7_75t_R _33249_ (.A(_15836_),
    .B(_15104_),
    .C(_14649_),
    .Y(_15837_));
 OAI21x1_ASAP7_75t_R _33250_ (.A1(_14646_),
    .A2(_18633_),
    .B(_15837_),
    .Y(_18040_));
 AND2x2_ASAP7_75t_R _33251_ (.A(net1973),
    .B(_01780_),
    .Y(_15838_));
 AO21x1_ASAP7_75t_R _33252_ (.A1(_13328_),
    .A2(_00880_),
    .B(_15838_),
    .Y(_15839_));
 OAI22x1_ASAP7_75t_R _33253_ (.A1(_00879_),
    .A2(_15289_),
    .B1(_15839_),
    .B2(_15272_),
    .Y(_15840_));
 BUFx12f_ASAP7_75t_R _33254_ (.A(_13813_),
    .Y(_15841_));
 NAND2x1_ASAP7_75t_R _33255_ (.A(_15841_),
    .B(_00886_),
    .Y(_15842_));
 OA211x2_ASAP7_75t_R _33256_ (.A1(net1973),
    .A2(_15807_),
    .B(_15842_),
    .C(_15264_),
    .Y(_15843_));
 NAND2x1_ASAP7_75t_R _33257_ (.A(_13813_),
    .B(_00885_),
    .Y(_15844_));
 OA211x2_ASAP7_75t_R _33258_ (.A1(net1973),
    .A2(_15810_),
    .B(_15844_),
    .C(_14191_),
    .Y(_15845_));
 OR3x1_ASAP7_75t_R _33259_ (.A(_13724_),
    .B(_15843_),
    .C(_15845_),
    .Y(_15846_));
 OA211x2_ASAP7_75t_R _33260_ (.A1(_13688_),
    .A2(_15840_),
    .B(_15846_),
    .C(_13814_),
    .Y(_15847_));
 BUFx6f_ASAP7_75t_R _33261_ (.A(_13813_),
    .Y(_15848_));
 NAND2x1_ASAP7_75t_R _33262_ (.A(_15841_),
    .B(_00882_),
    .Y(_15849_));
 OA211x2_ASAP7_75t_R _33263_ (.A1(_15848_),
    .A2(_15815_),
    .B(_15849_),
    .C(_15264_),
    .Y(_15850_));
 NAND2x1_ASAP7_75t_R _33264_ (.A(_15841_),
    .B(_00881_),
    .Y(_15851_));
 OA211x2_ASAP7_75t_R _33265_ (.A1(_15848_),
    .A2(_15818_),
    .B(_15851_),
    .C(_15272_),
    .Y(_15852_));
 OR3x1_ASAP7_75t_R _33266_ (.A(_13688_),
    .B(_15850_),
    .C(_15852_),
    .Y(_15853_));
 NAND2x1_ASAP7_75t_R _33267_ (.A(_15841_),
    .B(_00890_),
    .Y(_15854_));
 OA211x2_ASAP7_75t_R _33268_ (.A1(_15848_),
    .A2(_15822_),
    .B(_15854_),
    .C(_15264_),
    .Y(_15855_));
 NAND2x1_ASAP7_75t_R _33269_ (.A(_15841_),
    .B(_00889_),
    .Y(_15856_));
 OA211x2_ASAP7_75t_R _33270_ (.A1(_15848_),
    .A2(_15825_),
    .B(_15856_),
    .C(_15272_),
    .Y(_15857_));
 OR3x1_ASAP7_75t_R _33271_ (.A(_13724_),
    .B(_15855_),
    .C(_15857_),
    .Y(_15858_));
 AND3x1_ASAP7_75t_R _33272_ (.A(_13669_),
    .B(_15853_),
    .C(_15858_),
    .Y(_15859_));
 OR3x1_ASAP7_75t_R _33273_ (.A(_13764_),
    .B(_15847_),
    .C(_15859_),
    .Y(_15860_));
 NAND2x1_ASAP7_75t_R _33274_ (.A(net1972),
    .B(_00898_),
    .Y(_15861_));
 OA211x2_ASAP7_75t_R _33275_ (.A1(_15848_),
    .A2(_15788_),
    .B(_15861_),
    .C(_15264_),
    .Y(_15862_));
 NAND2x1_ASAP7_75t_R _33276_ (.A(_15841_),
    .B(_00897_),
    .Y(_15863_));
 OA211x2_ASAP7_75t_R _33277_ (.A1(_15848_),
    .A2(_15791_),
    .B(_15863_),
    .C(_15272_),
    .Y(_15864_));
 OR3x1_ASAP7_75t_R _33278_ (.A(_13688_),
    .B(_15862_),
    .C(_15864_),
    .Y(_15865_));
 NAND2x1_ASAP7_75t_R _33279_ (.A(_15841_),
    .B(_00906_),
    .Y(_15866_));
 OA211x2_ASAP7_75t_R _33280_ (.A1(_15848_),
    .A2(_15795_),
    .B(_15866_),
    .C(_15264_),
    .Y(_15867_));
 NAND2x1_ASAP7_75t_R _33281_ (.A(_15841_),
    .B(_00905_),
    .Y(_15868_));
 OA211x2_ASAP7_75t_R _33282_ (.A1(_15848_),
    .A2(_15798_),
    .B(_15868_),
    .C(_15272_),
    .Y(_15869_));
 OR3x1_ASAP7_75t_R _33283_ (.A(_13724_),
    .B(_15867_),
    .C(_15869_),
    .Y(_15870_));
 AND3x1_ASAP7_75t_R _33284_ (.A(_13669_),
    .B(_15865_),
    .C(_15870_),
    .Y(_15871_));
 NOR2x1_ASAP7_75t_R _33285_ (.A(net1972),
    .B(_00903_),
    .Y(_15872_));
 AO21x1_ASAP7_75t_R _33286_ (.A1(_15848_),
    .A2(_15773_),
    .B(_15872_),
    .Y(_15873_));
 NAND2x1_ASAP7_75t_R _33287_ (.A(net1972),
    .B(_00902_),
    .Y(_15874_));
 OA211x2_ASAP7_75t_R _33288_ (.A1(_15848_),
    .A2(_15776_),
    .B(_15874_),
    .C(_15264_),
    .Y(_15875_));
 AO21x1_ASAP7_75t_R _33289_ (.A1(_15272_),
    .A2(_15873_),
    .B(_15875_),
    .Y(_15876_));
 NAND2x1_ASAP7_75t_R _33290_ (.A(_15841_),
    .B(_00894_),
    .Y(_15877_));
 OA211x2_ASAP7_75t_R _33291_ (.A1(_15256_),
    .A2(_15780_),
    .B(_15877_),
    .C(_15264_),
    .Y(_15878_));
 NAND2x1_ASAP7_75t_R _33292_ (.A(_15841_),
    .B(_00893_),
    .Y(_15879_));
 OA211x2_ASAP7_75t_R _33293_ (.A1(_15256_),
    .A2(_15783_),
    .B(_15879_),
    .C(_14191_),
    .Y(_15880_));
 OR3x1_ASAP7_75t_R _33294_ (.A(_13688_),
    .B(_15878_),
    .C(_15880_),
    .Y(_15881_));
 OA211x2_ASAP7_75t_R _33295_ (.A1(_13724_),
    .A2(_15876_),
    .B(_15881_),
    .C(_13814_),
    .Y(_15882_));
 OR3x2_ASAP7_75t_R _33296_ (.A(_13306_),
    .B(_15871_),
    .C(_15882_),
    .Y(_15883_));
 NAND2x2_ASAP7_75t_R _33297_ (.A(_15860_),
    .B(_15883_),
    .Y(_15884_));
 OA211x2_ASAP7_75t_R _33298_ (.A1(_14278_),
    .A2(_15366_),
    .B(_15369_),
    .C(_15503_),
    .Y(_15885_));
 AOI21x1_ASAP7_75t_R _33299_ (.A1(_14090_),
    .A2(_15884_),
    .B(_15885_),
    .Y(_18634_));
 INVx1_ASAP7_75t_R _33300_ (.A(_18634_),
    .Y(_18632_));
 AND2x2_ASAP7_75t_R _33301_ (.A(_14496_),
    .B(_01779_),
    .Y(_15886_));
 AO21x1_ASAP7_75t_R _33302_ (.A1(_14286_),
    .A2(_00912_),
    .B(_15886_),
    .Y(_15887_));
 OAI22x1_ASAP7_75t_R _33303_ (.A1(_00911_),
    .A2(_14284_),
    .B1(_15887_),
    .B2(_14289_),
    .Y(_15888_));
 INVx1_ASAP7_75t_R _33304_ (.A(_00920_),
    .Y(_15889_));
 NAND2x1_ASAP7_75t_R _33305_ (.A(_13146_),
    .B(_00918_),
    .Y(_15890_));
 OA211x2_ASAP7_75t_R _33306_ (.A1(_14293_),
    .A2(_15889_),
    .B(_15890_),
    .C(_14296_),
    .Y(_15891_));
 INVx1_ASAP7_75t_R _33307_ (.A(_00919_),
    .Y(_15892_));
 NAND2x1_ASAP7_75t_R _33308_ (.A(_14794_),
    .B(_00917_),
    .Y(_15893_));
 OA211x2_ASAP7_75t_R _33309_ (.A1(_14293_),
    .A2(_15892_),
    .B(_15893_),
    .C(_13149_),
    .Y(_15894_));
 OR3x1_ASAP7_75t_R _33310_ (.A(_13153_),
    .B(_15891_),
    .C(_15894_),
    .Y(_15895_));
 OA211x2_ASAP7_75t_R _33311_ (.A1(_14283_),
    .A2(_15888_),
    .B(_15895_),
    .C(_14778_),
    .Y(_15896_));
 INVx1_ASAP7_75t_R _33312_ (.A(_00916_),
    .Y(_15897_));
 NAND2x1_ASAP7_75t_R _33313_ (.A(_14455_),
    .B(_00914_),
    .Y(_15898_));
 OA211x2_ASAP7_75t_R _33314_ (.A1(_14358_),
    .A2(_15897_),
    .B(_15898_),
    .C(_14363_),
    .Y(_15899_));
 INVx1_ASAP7_75t_R _33315_ (.A(_00915_),
    .Y(_15900_));
 NAND2x1_ASAP7_75t_R _33316_ (.A(_14461_),
    .B(_00913_),
    .Y(_15901_));
 OA211x2_ASAP7_75t_R _33317_ (.A1(_15191_),
    .A2(_15900_),
    .B(_15901_),
    .C(_13089_),
    .Y(_15902_));
 OR3x1_ASAP7_75t_R _33318_ (.A(_14309_),
    .B(_15899_),
    .C(_15902_),
    .Y(_15903_));
 INVx1_ASAP7_75t_R _33319_ (.A(_00924_),
    .Y(_15904_));
 NAND2x1_ASAP7_75t_R _33320_ (.A(_14455_),
    .B(_00922_),
    .Y(_15905_));
 OA211x2_ASAP7_75t_R _33321_ (.A1(_14358_),
    .A2(_15904_),
    .B(_15905_),
    .C(_14363_),
    .Y(_15906_));
 INVx1_ASAP7_75t_R _33322_ (.A(_00923_),
    .Y(_15907_));
 NAND2x1_ASAP7_75t_R _33323_ (.A(_15052_),
    .B(_00921_),
    .Y(_15908_));
 OA211x2_ASAP7_75t_R _33324_ (.A1(_15191_),
    .A2(_15907_),
    .B(_15908_),
    .C(_15195_),
    .Y(_15909_));
 OR3x1_ASAP7_75t_R _33325_ (.A(_14327_),
    .B(_15906_),
    .C(_15909_),
    .Y(_15910_));
 AND3x1_ASAP7_75t_R _33326_ (.A(_14307_),
    .B(_15903_),
    .C(_15910_),
    .Y(_15911_));
 OR3x1_ASAP7_75t_R _33327_ (.A(_14281_),
    .B(_15896_),
    .C(_15911_),
    .Y(_15912_));
 INVx2_ASAP7_75t_R _33328_ (.A(_00932_),
    .Y(_15913_));
 NAND2x1_ASAP7_75t_R _33329_ (.A(_14455_),
    .B(_00930_),
    .Y(_15914_));
 OA211x2_ASAP7_75t_R _33330_ (.A1(_14358_),
    .A2(_15913_),
    .B(_15914_),
    .C(_14363_),
    .Y(_15915_));
 INVx2_ASAP7_75t_R _33331_ (.A(_00931_),
    .Y(_15916_));
 NAND2x1_ASAP7_75t_R _33332_ (.A(_14461_),
    .B(_00929_),
    .Y(_15917_));
 OA211x2_ASAP7_75t_R _33333_ (.A1(_15191_),
    .A2(_15916_),
    .B(_15917_),
    .C(_15195_),
    .Y(_15918_));
 OR3x1_ASAP7_75t_R _33334_ (.A(_14309_),
    .B(_15915_),
    .C(_15918_),
    .Y(_15919_));
 INVx1_ASAP7_75t_R _33335_ (.A(_00940_),
    .Y(_15920_));
 NAND2x1_ASAP7_75t_R _33336_ (.A(_14461_),
    .B(_00938_),
    .Y(_15921_));
 OA211x2_ASAP7_75t_R _33337_ (.A1(_15191_),
    .A2(_15920_),
    .B(_15921_),
    .C(_14315_),
    .Y(_15922_));
 INVx2_ASAP7_75t_R _33338_ (.A(_00939_),
    .Y(_15923_));
 NAND2x1_ASAP7_75t_R _33339_ (.A(_15052_),
    .B(_00937_),
    .Y(_15924_));
 OA211x2_ASAP7_75t_R _33340_ (.A1(_14311_),
    .A2(_15923_),
    .B(_15924_),
    .C(_15195_),
    .Y(_15925_));
 OR3x1_ASAP7_75t_R _33341_ (.A(_14327_),
    .B(_15922_),
    .C(_15925_),
    .Y(_15926_));
 AND3x1_ASAP7_75t_R _33342_ (.A(_14307_),
    .B(_15919_),
    .C(_15926_),
    .Y(_15927_));
 INVx2_ASAP7_75t_R _33343_ (.A(_00933_),
    .Y(_15928_));
 NOR2x1_ASAP7_75t_R _33344_ (.A(_13133_),
    .B(_00935_),
    .Y(_15929_));
 AO21x1_ASAP7_75t_R _33345_ (.A1(_14278_),
    .A2(_15928_),
    .B(_15929_),
    .Y(_15930_));
 INVx2_ASAP7_75t_R _33346_ (.A(_00936_),
    .Y(_15931_));
 NAND2x1_ASAP7_75t_R _33347_ (.A(_13097_),
    .B(_00934_),
    .Y(_15932_));
 OA211x2_ASAP7_75t_R _33348_ (.A1(_13190_),
    .A2(_15931_),
    .B(_15932_),
    .C(_14363_),
    .Y(_15933_));
 AO21x1_ASAP7_75t_R _33349_ (.A1(_13090_),
    .A2(_15930_),
    .B(_15933_),
    .Y(_15934_));
 INVx2_ASAP7_75t_R _33350_ (.A(_00928_),
    .Y(_15935_));
 NAND2x1_ASAP7_75t_R _33351_ (.A(_14277_),
    .B(_00926_),
    .Y(_15936_));
 OA211x2_ASAP7_75t_R _33352_ (.A1(_14299_),
    .A2(_15935_),
    .B(_15936_),
    .C(_14296_),
    .Y(_15937_));
 INVx1_ASAP7_75t_R _33353_ (.A(_00927_),
    .Y(_15938_));
 NAND2x1_ASAP7_75t_R _33354_ (.A(_14301_),
    .B(_00925_),
    .Y(_15939_));
 OA211x2_ASAP7_75t_R _33355_ (.A1(_14299_),
    .A2(_15938_),
    .B(_15939_),
    .C(_14372_),
    .Y(_15940_));
 OR3x1_ASAP7_75t_R _33356_ (.A(_14282_),
    .B(_15937_),
    .C(_15940_),
    .Y(_15941_));
 OA211x2_ASAP7_75t_R _33357_ (.A1(_14354_),
    .A2(_15934_),
    .B(_15941_),
    .C(_14305_),
    .Y(_15942_));
 OR3x2_ASAP7_75t_R _33358_ (.A(_14339_),
    .B(_15927_),
    .C(_15942_),
    .Y(_15943_));
 AO21x2_ASAP7_75t_R _33359_ (.A1(_15912_),
    .A2(_15943_),
    .B(_13268_),
    .Y(_15944_));
 AND2x2_ASAP7_75t_R _33360_ (.A(_01469_),
    .B(_15100_),
    .Y(_15945_));
 OAI22x1_ASAP7_75t_R _33361_ (.A1(_01498_),
    .A2(_14382_),
    .B1(_14385_),
    .B2(_15945_),
    .Y(_15946_));
 NAND2x2_ASAP7_75t_R _33362_ (.A(_15944_),
    .B(_15946_),
    .Y(_18638_));
 INVx1_ASAP7_75t_R _33363_ (.A(_18638_),
    .Y(_18640_));
 BUFx6f_ASAP7_75t_R _33364_ (.A(_00098_),
    .Y(_15947_));
 OR3x1_ASAP7_75t_R _33365_ (.A(_15947_),
    .B(_15104_),
    .C(_14649_),
    .Y(_15948_));
 OAI21x1_ASAP7_75t_R _33366_ (.A1(_14646_),
    .A2(_18638_),
    .B(_15948_),
    .Y(_18042_));
 BUFx6f_ASAP7_75t_R _33367_ (.A(net1972),
    .Y(_15949_));
 AND2x2_ASAP7_75t_R _33368_ (.A(_15949_),
    .B(_01779_),
    .Y(_15950_));
 AO21x1_ASAP7_75t_R _33369_ (.A1(_15290_),
    .A2(_00912_),
    .B(_15950_),
    .Y(_15951_));
 OAI22x1_ASAP7_75t_R _33370_ (.A1(_00911_),
    .A2(_15289_),
    .B1(_15951_),
    .B2(_15273_),
    .Y(_15952_));
 BUFx6f_ASAP7_75t_R _33371_ (.A(net1972),
    .Y(_15953_));
 NAND2x1_ASAP7_75t_R _33372_ (.A(_15949_),
    .B(_00918_),
    .Y(_15954_));
 OA211x2_ASAP7_75t_R _33373_ (.A1(_15953_),
    .A2(_15889_),
    .B(_15954_),
    .C(_15265_),
    .Y(_15955_));
 NAND2x1_ASAP7_75t_R _33374_ (.A(_15949_),
    .B(_00917_),
    .Y(_15956_));
 OA211x2_ASAP7_75t_R _33375_ (.A1(_15953_),
    .A2(_15892_),
    .B(_15956_),
    .C(_15273_),
    .Y(_15957_));
 OR3x1_ASAP7_75t_R _33376_ (.A(_15278_),
    .B(_15955_),
    .C(_15957_),
    .Y(_15958_));
 OA21x2_ASAP7_75t_R _33377_ (.A1(_15254_),
    .A2(_15952_),
    .B(_15958_),
    .Y(_15959_));
 NAND2x1_ASAP7_75t_R _33378_ (.A(_15949_),
    .B(_00914_),
    .Y(_15960_));
 OA211x2_ASAP7_75t_R _33379_ (.A1(_15953_),
    .A2(_15897_),
    .B(_15960_),
    .C(_15265_),
    .Y(_15961_));
 NAND2x1_ASAP7_75t_R _33380_ (.A(_15949_),
    .B(_00913_),
    .Y(_15962_));
 OA211x2_ASAP7_75t_R _33381_ (.A1(_15953_),
    .A2(_15900_),
    .B(_15962_),
    .C(_15273_),
    .Y(_15963_));
 OR3x1_ASAP7_75t_R _33382_ (.A(_15254_),
    .B(_15961_),
    .C(_15963_),
    .Y(_15964_));
 NAND2x1_ASAP7_75t_R _33383_ (.A(_15949_),
    .B(_00922_),
    .Y(_15965_));
 OA211x2_ASAP7_75t_R _33384_ (.A1(_15953_),
    .A2(_15904_),
    .B(_15965_),
    .C(_15265_),
    .Y(_15966_));
 NAND2x1_ASAP7_75t_R _33385_ (.A(net1973),
    .B(_00921_),
    .Y(_15967_));
 OA211x2_ASAP7_75t_R _33386_ (.A1(_15953_),
    .A2(_15907_),
    .B(_15967_),
    .C(_15273_),
    .Y(_15968_));
 OR3x1_ASAP7_75t_R _33387_ (.A(_15278_),
    .B(_15966_),
    .C(_15968_),
    .Y(_15969_));
 AND3x1_ASAP7_75t_R _33388_ (.A(_15252_),
    .B(_15964_),
    .C(_15969_),
    .Y(_15970_));
 AO21x1_ASAP7_75t_R _33389_ (.A1(_15312_),
    .A2(_15959_),
    .B(_15970_),
    .Y(_15971_));
 NAND2x1_ASAP7_75t_R _33390_ (.A(net1972),
    .B(_00930_),
    .Y(_15972_));
 OA211x2_ASAP7_75t_R _33391_ (.A1(_15953_),
    .A2(_15913_),
    .B(_15972_),
    .C(_15265_),
    .Y(_15973_));
 NAND2x1_ASAP7_75t_R _33392_ (.A(net1972),
    .B(_00929_),
    .Y(_15974_));
 OA211x2_ASAP7_75t_R _33393_ (.A1(_15953_),
    .A2(_15916_),
    .B(_15974_),
    .C(_15272_),
    .Y(_15975_));
 OR3x1_ASAP7_75t_R _33394_ (.A(_15254_),
    .B(_15973_),
    .C(_15975_),
    .Y(_15976_));
 NAND2x1_ASAP7_75t_R _33395_ (.A(net1972),
    .B(_00938_),
    .Y(_15977_));
 OA211x2_ASAP7_75t_R _33396_ (.A1(_15953_),
    .A2(_15920_),
    .B(_15977_),
    .C(_15264_),
    .Y(_15978_));
 NAND2x1_ASAP7_75t_R _33397_ (.A(net1972),
    .B(_00937_),
    .Y(_15979_));
 OA211x2_ASAP7_75t_R _33398_ (.A1(_15949_),
    .A2(_15923_),
    .B(_15979_),
    .C(_15272_),
    .Y(_15980_));
 OR3x1_ASAP7_75t_R _33399_ (.A(_13724_),
    .B(_15978_),
    .C(_15980_),
    .Y(_15981_));
 AND3x1_ASAP7_75t_R _33400_ (.A(_15252_),
    .B(_15976_),
    .C(_15981_),
    .Y(_15982_));
 NOR2x1_ASAP7_75t_R _33401_ (.A(_15949_),
    .B(_00935_),
    .Y(_15983_));
 AO21x1_ASAP7_75t_R _33402_ (.A1(_15258_),
    .A2(_15928_),
    .B(_15983_),
    .Y(_15984_));
 NAND2x1_ASAP7_75t_R _33403_ (.A(net1972),
    .B(_00934_),
    .Y(_15985_));
 OA211x2_ASAP7_75t_R _33404_ (.A1(_15953_),
    .A2(_15931_),
    .B(_15985_),
    .C(_15265_),
    .Y(_15986_));
 AO21x1_ASAP7_75t_R _33405_ (.A1(_15273_),
    .A2(_15984_),
    .B(_15986_),
    .Y(_15987_));
 NAND2x1_ASAP7_75t_R _33406_ (.A(net1972),
    .B(_00926_),
    .Y(_15988_));
 OA211x2_ASAP7_75t_R _33407_ (.A1(_15949_),
    .A2(_15935_),
    .B(_15988_),
    .C(_15264_),
    .Y(_15989_));
 NAND2x1_ASAP7_75t_R _33408_ (.A(net1972),
    .B(_00925_),
    .Y(_15990_));
 OA211x2_ASAP7_75t_R _33409_ (.A1(_15949_),
    .A2(_15938_),
    .B(_15990_),
    .C(_15272_),
    .Y(_15991_));
 OR3x1_ASAP7_75t_R _33410_ (.A(_15254_),
    .B(_15989_),
    .C(_15991_),
    .Y(_15992_));
 OA211x2_ASAP7_75t_R _33411_ (.A1(_15278_),
    .A2(_15987_),
    .B(_15992_),
    .C(_13814_),
    .Y(_15993_));
 OR3x1_ASAP7_75t_R _33412_ (.A(_13306_),
    .B(_15982_),
    .C(_15993_),
    .Y(_15994_));
 OAI21x1_ASAP7_75t_R _33413_ (.A1(_15251_),
    .A2(_15971_),
    .B(_15994_),
    .Y(_15995_));
 OA211x2_ASAP7_75t_R _33414_ (.A1(_14778_),
    .A2(_15366_),
    .B(_15369_),
    .C(_15503_),
    .Y(_15996_));
 AOI21x1_ASAP7_75t_R _33415_ (.A1(_14090_),
    .A2(_15995_),
    .B(_15996_),
    .Y(_18639_));
 INVx1_ASAP7_75t_R _33416_ (.A(_18639_),
    .Y(_18637_));
 BUFx6f_ASAP7_75t_R _33417_ (.A(_00909_),
    .Y(_15997_));
 OA21x2_ASAP7_75t_R _33418_ (.A1(net1941),
    .A2(_15762_),
    .B(_00910_),
    .Y(_15998_));
 OAI21x1_ASAP7_75t_R _33419_ (.A1(_15997_),
    .A2(_15998_),
    .B(_00942_),
    .Y(_15999_));
 OR4x1_ASAP7_75t_R _33420_ (.A(net1937),
    .B(net1935),
    .C(net1941),
    .D(_15997_),
    .Y(_16000_));
 INVx1_ASAP7_75t_R _33421_ (.A(_16000_),
    .Y(_16001_));
 OA21x2_ASAP7_75t_R _33422_ (.A1(_15507_),
    .A2(_15516_),
    .B(_16001_),
    .Y(_16002_));
 NOR2x1_ASAP7_75t_R _33423_ (.A(_15999_),
    .B(_16002_),
    .Y(_16003_));
 XNOR2x1_ASAP7_75t_R _33424_ (.B(_16003_),
    .Y(_16004_),
    .A(net1940));
 INVx4_ASAP7_75t_R _33425_ (.A(_16004_),
    .Y(\alu_adder_result_ex[17] ));
 INVx1_ASAP7_75t_R _33426_ (.A(_15997_),
    .Y(_16005_));
 OR4x1_ASAP7_75t_R _33427_ (.A(net1935),
    .B(net1937),
    .C(net1938),
    .D(net1941),
    .Y(_16006_));
 OR5x2_ASAP7_75t_R _33428_ (.A(_16005_),
    .B(_15169_),
    .C(_15176_),
    .D(_15510_),
    .E(net1956),
    .Y(_16007_));
 OR2x2_ASAP7_75t_R _33429_ (.A(net1935),
    .B(net1941),
    .Y(_16008_));
 OA21x2_ASAP7_75t_R _33430_ (.A1(_00814_),
    .A2(net1937),
    .B(_00846_),
    .Y(_16009_));
 OA21x2_ASAP7_75t_R _33431_ (.A1(_00878_),
    .A2(net1941),
    .B(_00910_),
    .Y(_16010_));
 OA21x2_ASAP7_75t_R _33432_ (.A1(_16008_),
    .A2(_16009_),
    .B(_16010_),
    .Y(_16011_));
 NAND3x1_ASAP7_75t_R _33433_ (.A(_16005_),
    .B(_15522_),
    .C(_16011_),
    .Y(_16012_));
 INVx1_ASAP7_75t_R _33434_ (.A(_16012_),
    .Y(_16013_));
 OAI21x1_ASAP7_75t_R _33435_ (.A1(_15169_),
    .A2(_15176_),
    .B(_16013_),
    .Y(_16014_));
 AO21x1_ASAP7_75t_R _33436_ (.A1(_15510_),
    .A2(_15522_),
    .B(net1956),
    .Y(_16015_));
 NAND2x1_ASAP7_75t_R _33437_ (.A(_16011_),
    .B(_16015_),
    .Y(_16016_));
 OA211x2_ASAP7_75t_R _33438_ (.A1(_15522_),
    .A2(net1956),
    .B(_16011_),
    .C(_15997_),
    .Y(_16017_));
 AO21x1_ASAP7_75t_R _33439_ (.A1(_16005_),
    .A2(_16016_),
    .B(_16017_),
    .Y(_16018_));
 AND3x4_ASAP7_75t_R _33440_ (.A(_16007_),
    .B(_16014_),
    .C(_16018_),
    .Y(_16019_));
 INVx3_ASAP7_75t_R _33441_ (.A(_16019_),
    .Y(\alu_adder_result_ex[16] ));
 INVx2_ASAP7_75t_R _33442_ (.A(_00965_),
    .Y(_16020_));
 NOR2x1_ASAP7_75t_R _33443_ (.A(_14360_),
    .B(_00967_),
    .Y(_16021_));
 AO21x1_ASAP7_75t_R _33444_ (.A1(_14331_),
    .A2(_16020_),
    .B(_16021_),
    .Y(_16022_));
 INVx2_ASAP7_75t_R _33445_ (.A(_00968_),
    .Y(_16023_));
 NAND2x1_ASAP7_75t_R _33446_ (.A(_14808_),
    .B(_00966_),
    .Y(_16024_));
 OA211x2_ASAP7_75t_R _33447_ (.A1(_14943_),
    .A2(_16023_),
    .B(_16024_),
    .C(_14494_),
    .Y(_16025_));
 AO21x1_ASAP7_75t_R _33448_ (.A1(_14710_),
    .A2(_16022_),
    .B(_16025_),
    .Y(_16026_));
 INVx2_ASAP7_75t_R _33449_ (.A(_00960_),
    .Y(_16027_));
 NAND2x1_ASAP7_75t_R _33450_ (.A(_13118_),
    .B(_00958_),
    .Y(_16028_));
 OA211x2_ASAP7_75t_R _33451_ (.A1(_13206_),
    .A2(_16027_),
    .B(_16028_),
    .C(_13115_),
    .Y(_16029_));
 INVx2_ASAP7_75t_R _33452_ (.A(_00959_),
    .Y(_16030_));
 NAND2x1_ASAP7_75t_R _33453_ (.A(_13211_),
    .B(_00957_),
    .Y(_16031_));
 OA211x2_ASAP7_75t_R _33454_ (.A1(_13206_),
    .A2(_16030_),
    .B(_16031_),
    .C(_13120_),
    .Y(_16032_));
 OA21x2_ASAP7_75t_R _33455_ (.A1(_16029_),
    .A2(_16032_),
    .B(_14353_),
    .Y(_16033_));
 AO21x1_ASAP7_75t_R _33456_ (.A1(_14448_),
    .A2(_16026_),
    .B(_16033_),
    .Y(_16034_));
 INVx2_ASAP7_75t_R _33457_ (.A(_00964_),
    .Y(_16035_));
 NAND2x1_ASAP7_75t_R _33458_ (.A(_14403_),
    .B(_00962_),
    .Y(_16036_));
 OA211x2_ASAP7_75t_R _33459_ (.A1(_14756_),
    .A2(_16035_),
    .B(_16036_),
    .C(_14458_),
    .Y(_16037_));
 INVx2_ASAP7_75t_R _33460_ (.A(_00963_),
    .Y(_16038_));
 NAND2x1_ASAP7_75t_R _33461_ (.A(_13132_),
    .B(_00961_),
    .Y(_16039_));
 OA211x2_ASAP7_75t_R _33462_ (.A1(_14756_),
    .A2(_16038_),
    .B(_16039_),
    .C(_14743_),
    .Y(_16040_));
 OR3x1_ASAP7_75t_R _33463_ (.A(_14737_),
    .B(_16037_),
    .C(_16040_),
    .Y(_16041_));
 INVx1_ASAP7_75t_R _33464_ (.A(_00972_),
    .Y(_16042_));
 NAND2x1_ASAP7_75t_R _33465_ (.A(_13132_),
    .B(_00970_),
    .Y(_16043_));
 OA211x2_ASAP7_75t_R _33466_ (.A1(_14756_),
    .A2(_16042_),
    .B(_16043_),
    .C(_14458_),
    .Y(_16044_));
 INVx2_ASAP7_75t_R _33467_ (.A(_00971_),
    .Y(_16045_));
 NAND2x1_ASAP7_75t_R _33468_ (.A(_14437_),
    .B(_00969_),
    .Y(_16046_));
 OA211x2_ASAP7_75t_R _33469_ (.A1(_14888_),
    .A2(_16045_),
    .B(_16046_),
    .C(_14743_),
    .Y(_16047_));
 OR3x1_ASAP7_75t_R _33470_ (.A(_14454_),
    .B(_16044_),
    .C(_16047_),
    .Y(_16048_));
 AND3x1_ASAP7_75t_R _33471_ (.A(_14468_),
    .B(_16041_),
    .C(_16048_),
    .Y(_16049_));
 AO21x1_ASAP7_75t_R _33472_ (.A1(_14778_),
    .A2(_16034_),
    .B(_16049_),
    .Y(_16050_));
 AND2x2_ASAP7_75t_R _33473_ (.A(_13165_),
    .B(_01778_),
    .Y(_16051_));
 AO21x1_ASAP7_75t_R _33474_ (.A1(_14285_),
    .A2(_00944_),
    .B(_16051_),
    .Y(_16052_));
 OAI22x1_ASAP7_75t_R _33475_ (.A1(_00943_),
    .A2(_13101_),
    .B1(_16052_),
    .B2(_14710_),
    .Y(_16053_));
 INVx2_ASAP7_75t_R _33476_ (.A(_00952_),
    .Y(_16054_));
 NAND2x1_ASAP7_75t_R _33477_ (.A(_14391_),
    .B(_00950_),
    .Y(_16055_));
 OA211x2_ASAP7_75t_R _33478_ (.A1(_15675_),
    .A2(_16054_),
    .B(_16055_),
    .C(_14362_),
    .Y(_16056_));
 INVx2_ASAP7_75t_R _33479_ (.A(_00951_),
    .Y(_16057_));
 NAND2x1_ASAP7_75t_R _33480_ (.A(_14460_),
    .B(_00949_),
    .Y(_16058_));
 OA211x2_ASAP7_75t_R _33481_ (.A1(_13118_),
    .A2(_16057_),
    .B(_16058_),
    .C(_13088_),
    .Y(_16059_));
 OR3x1_ASAP7_75t_R _33482_ (.A(_14326_),
    .B(_16056_),
    .C(_16059_),
    .Y(_16060_));
 OA211x2_ASAP7_75t_R _33483_ (.A1(_14309_),
    .A2(_16053_),
    .B(_16060_),
    .C(_14428_),
    .Y(_16061_));
 INVx2_ASAP7_75t_R _33484_ (.A(_00948_),
    .Y(_16062_));
 NAND2x1_ASAP7_75t_R _33485_ (.A(_13106_),
    .B(_00946_),
    .Y(_16063_));
 OA211x2_ASAP7_75t_R _33486_ (.A1(_13137_),
    .A2(_16062_),
    .B(_16063_),
    .C(_14740_),
    .Y(_16064_));
 INVx2_ASAP7_75t_R _33487_ (.A(_00947_),
    .Y(_16065_));
 NAND2x1_ASAP7_75t_R _33488_ (.A(_13106_),
    .B(_00945_),
    .Y(_16066_));
 OA211x2_ASAP7_75t_R _33489_ (.A1(_13146_),
    .A2(_16065_),
    .B(_16066_),
    .C(_14732_),
    .Y(_16067_));
 OR3x1_ASAP7_75t_R _33490_ (.A(_14737_),
    .B(_16064_),
    .C(_16067_),
    .Y(_16068_));
 INVx2_ASAP7_75t_R _33491_ (.A(_00956_),
    .Y(_16069_));
 NAND2x1_ASAP7_75t_R _33492_ (.A(_13106_),
    .B(_00954_),
    .Y(_16070_));
 OA211x2_ASAP7_75t_R _33493_ (.A1(_13146_),
    .A2(_16069_),
    .B(_16070_),
    .C(_14740_),
    .Y(_16071_));
 INVx2_ASAP7_75t_R _33494_ (.A(_00955_),
    .Y(_16072_));
 NAND2x1_ASAP7_75t_R _33495_ (.A(_13106_),
    .B(_00953_),
    .Y(_16073_));
 OA211x2_ASAP7_75t_R _33496_ (.A1(_14794_),
    .A2(_16072_),
    .B(_16073_),
    .C(_14732_),
    .Y(_16074_));
 OR3x1_ASAP7_75t_R _33497_ (.A(_14454_),
    .B(_16071_),
    .C(_16074_),
    .Y(_16075_));
 AND3x1_ASAP7_75t_R _33498_ (.A(_14468_),
    .B(_16068_),
    .C(_16075_),
    .Y(_16076_));
 OR3x1_ASAP7_75t_R _33499_ (.A(_14447_),
    .B(_16061_),
    .C(_16076_),
    .Y(_16077_));
 OA21x2_ASAP7_75t_R _33500_ (.A1(_14339_),
    .A2(_16050_),
    .B(_16077_),
    .Y(_16078_));
 BUFx6f_ASAP7_75t_R _33501_ (.A(_00020_),
    .Y(_16079_));
 AND2x2_ASAP7_75t_R _33502_ (.A(_01468_),
    .B(_14772_),
    .Y(_16080_));
 OAI22x1_ASAP7_75t_R _33503_ (.A1(_16079_),
    .A2(_14967_),
    .B1(_14968_),
    .B2(_16080_),
    .Y(_16081_));
 OA21x2_ASAP7_75t_R _33504_ (.A1(_13268_),
    .A2(_16078_),
    .B(_16081_),
    .Y(_16082_));
 BUFx6f_ASAP7_75t_R _33505_ (.A(_16082_),
    .Y(_18645_));
 INVx3_ASAP7_75t_R _33506_ (.A(_18645_),
    .Y(_18643_));
 BUFx6f_ASAP7_75t_R _33507_ (.A(_00101_),
    .Y(_16083_));
 OR3x1_ASAP7_75t_R _33508_ (.A(_16083_),
    .B(_15104_),
    .C(_14649_),
    .Y(_16084_));
 OAI21x1_ASAP7_75t_R _33509_ (.A1(_14646_),
    .A2(_18643_),
    .B(_16084_),
    .Y(_18044_));
 AND2x2_ASAP7_75t_R _33510_ (.A(_15291_),
    .B(_01778_),
    .Y(_16085_));
 AO21x1_ASAP7_75t_R _33511_ (.A1(_15290_),
    .A2(_00944_),
    .B(_16085_),
    .Y(_16086_));
 OAI22x1_ASAP7_75t_R _33512_ (.A1(_00943_),
    .A2(_15289_),
    .B1(_16086_),
    .B2(_15296_),
    .Y(_16087_));
 NAND2x1_ASAP7_75t_R _33513_ (.A(_15489_),
    .B(_00950_),
    .Y(_16088_));
 OA211x2_ASAP7_75t_R _33514_ (.A1(_15300_),
    .A2(_16054_),
    .B(_16088_),
    .C(_15304_),
    .Y(_16089_));
 NAND2x1_ASAP7_75t_R _33515_ (.A(_15489_),
    .B(_00949_),
    .Y(_16090_));
 OA211x2_ASAP7_75t_R _33516_ (.A1(_15307_),
    .A2(_16057_),
    .B(_16090_),
    .C(_15309_),
    .Y(_16091_));
 OR3x1_ASAP7_75t_R _33517_ (.A(_15298_),
    .B(_16089_),
    .C(_16091_),
    .Y(_16092_));
 OA211x2_ASAP7_75t_R _33518_ (.A1(_15288_),
    .A2(_16087_),
    .B(_16092_),
    .C(_15313_),
    .Y(_16093_));
 NAND2x1_ASAP7_75t_R _33519_ (.A(_15618_),
    .B(_00946_),
    .Y(_16094_));
 OA211x2_ASAP7_75t_R _33520_ (.A1(_15269_),
    .A2(_16062_),
    .B(_16094_),
    .C(_15620_),
    .Y(_16095_));
 NAND2x1_ASAP7_75t_R _33521_ (.A(_15340_),
    .B(_00945_),
    .Y(_16096_));
 OA211x2_ASAP7_75t_R _33522_ (.A1(_15622_),
    .A2(_16065_),
    .B(_16096_),
    .C(_15283_),
    .Y(_16097_));
 OR3x1_ASAP7_75t_R _33523_ (.A(_15255_),
    .B(_16095_),
    .C(_16097_),
    .Y(_16098_));
 NAND2x1_ASAP7_75t_R _33524_ (.A(_15618_),
    .B(_00954_),
    .Y(_16099_));
 OA211x2_ASAP7_75t_R _33525_ (.A1(_15622_),
    .A2(_16069_),
    .B(_16099_),
    .C(_15620_),
    .Y(_16100_));
 NAND2x1_ASAP7_75t_R _33526_ (.A(_15340_),
    .B(_00953_),
    .Y(_16101_));
 OA211x2_ASAP7_75t_R _33527_ (.A1(_15343_),
    .A2(_16072_),
    .B(_16101_),
    .C(_15283_),
    .Y(_16102_));
 OR3x1_ASAP7_75t_R _33528_ (.A(_15279_),
    .B(_16100_),
    .C(_16102_),
    .Y(_16103_));
 AND3x1_ASAP7_75t_R _33529_ (.A(_15253_),
    .B(_16098_),
    .C(_16103_),
    .Y(_16104_));
 OR3x2_ASAP7_75t_R _33530_ (.A(_15251_),
    .B(_16093_),
    .C(_16104_),
    .Y(_16105_));
 BUFx12f_ASAP7_75t_R _33531_ (.A(_15301_),
    .Y(_16106_));
 NAND2x1_ASAP7_75t_R _33532_ (.A(_16106_),
    .B(_00962_),
    .Y(_16107_));
 OA211x2_ASAP7_75t_R _33533_ (.A1(_15325_),
    .A2(_16035_),
    .B(_16107_),
    .C(_15267_),
    .Y(_16108_));
 BUFx12f_ASAP7_75t_R _33534_ (.A(_15301_),
    .Y(_16109_));
 NAND2x1_ASAP7_75t_R _33535_ (.A(_16109_),
    .B(_00961_),
    .Y(_16110_));
 OA211x2_ASAP7_75t_R _33536_ (.A1(_15260_),
    .A2(_16038_),
    .B(_16110_),
    .C(_15275_),
    .Y(_16111_));
 OR3x1_ASAP7_75t_R _33537_ (.A(_15255_),
    .B(_16108_),
    .C(_16111_),
    .Y(_16112_));
 NAND2x1_ASAP7_75t_R _33538_ (.A(_16106_),
    .B(_00970_),
    .Y(_16113_));
 OA211x2_ASAP7_75t_R _33539_ (.A1(_15325_),
    .A2(_16042_),
    .B(_16113_),
    .C(_15267_),
    .Y(_16114_));
 NAND2x1_ASAP7_75t_R _33540_ (.A(_16109_),
    .B(_00969_),
    .Y(_16115_));
 OA211x2_ASAP7_75t_R _33541_ (.A1(_15260_),
    .A2(_16045_),
    .B(_16115_),
    .C(_15275_),
    .Y(_16116_));
 OR3x1_ASAP7_75t_R _33542_ (.A(_15279_),
    .B(_16114_),
    .C(_16116_),
    .Y(_16117_));
 AND3x1_ASAP7_75t_R _33543_ (.A(_15317_),
    .B(_16112_),
    .C(_16117_),
    .Y(_16118_));
 NOR2x1_ASAP7_75t_R _33544_ (.A(_15445_),
    .B(_00967_),
    .Y(_16119_));
 AO21x1_ASAP7_75t_R _33545_ (.A1(_15341_),
    .A2(_16020_),
    .B(_16119_),
    .Y(_16120_));
 NAND2x1_ASAP7_75t_R _33546_ (.A(_15270_),
    .B(_00966_),
    .Y(_16121_));
 OA211x2_ASAP7_75t_R _33547_ (.A1(_15346_),
    .A2(_16023_),
    .B(_16121_),
    .C(_15349_),
    .Y(_16122_));
 AO21x1_ASAP7_75t_R _33548_ (.A1(_15339_),
    .A2(_16120_),
    .B(_16122_),
    .Y(_16123_));
 NAND2x1_ASAP7_75t_R _33549_ (.A(_15632_),
    .B(_00958_),
    .Y(_16124_));
 OA211x2_ASAP7_75t_R _33550_ (.A1(_15353_),
    .A2(_16027_),
    .B(_16124_),
    .C(_15304_),
    .Y(_16125_));
 NAND2x1_ASAP7_75t_R _33551_ (.A(_15489_),
    .B(_00957_),
    .Y(_16126_));
 OA211x2_ASAP7_75t_R _33552_ (.A1(_15300_),
    .A2(_16030_),
    .B(_16126_),
    .C(_15309_),
    .Y(_16127_));
 OR3x1_ASAP7_75t_R _33553_ (.A(_15352_),
    .B(_16125_),
    .C(_16127_),
    .Y(_16128_));
 OA211x2_ASAP7_75t_R _33554_ (.A1(_15337_),
    .A2(_16123_),
    .B(_16128_),
    .C(_15313_),
    .Y(_16129_));
 OR3x2_ASAP7_75t_R _33555_ (.A(_15316_),
    .B(_16118_),
    .C(_16129_),
    .Y(_16130_));
 NAND2x2_ASAP7_75t_R _33556_ (.A(_16130_),
    .B(_16105_),
    .Y(_16131_));
 OA211x2_ASAP7_75t_R _33557_ (.A1(_14354_),
    .A2(_15366_),
    .B(_15369_),
    .C(_15503_),
    .Y(_16132_));
 AOI21x1_ASAP7_75t_R _33558_ (.A1(_14090_),
    .A2(net1966),
    .B(_16132_),
    .Y(_18644_));
 INVx1_ASAP7_75t_R _33559_ (.A(_18644_),
    .Y(_18642_));
 AND2x2_ASAP7_75t_R _33560_ (.A(_14717_),
    .B(_01777_),
    .Y(_16133_));
 AO21x1_ASAP7_75t_R _33561_ (.A1(_13092_),
    .A2(_00976_),
    .B(_16133_),
    .Y(_16134_));
 OAI22x1_ASAP7_75t_R _33562_ (.A1(_00975_),
    .A2(_13102_),
    .B1(_16134_),
    .B2(_13090_),
    .Y(_16135_));
 INVx2_ASAP7_75t_R _33563_ (.A(_00984_),
    .Y(_16136_));
 NAND2x1_ASAP7_75t_R _33564_ (.A(_14317_),
    .B(_00982_),
    .Y(_16137_));
 OA211x2_ASAP7_75t_R _33565_ (.A1(_13107_),
    .A2(_16136_),
    .B(_16137_),
    .C(_13115_),
    .Y(_16138_));
 INVx2_ASAP7_75t_R _33566_ (.A(_00983_),
    .Y(_16139_));
 NAND2x1_ASAP7_75t_R _33567_ (.A(_13110_),
    .B(_00981_),
    .Y(_16140_));
 OA211x2_ASAP7_75t_R _33568_ (.A1(_13107_),
    .A2(_16139_),
    .B(_16140_),
    .C(_13120_),
    .Y(_16141_));
 OR3x1_ASAP7_75t_R _33569_ (.A(_13105_),
    .B(_16138_),
    .C(_16141_),
    .Y(_16142_));
 OA211x2_ASAP7_75t_R _33570_ (.A1(_13086_),
    .A2(_16135_),
    .B(_16142_),
    .C(_13125_),
    .Y(_16143_));
 INVx2_ASAP7_75t_R _33571_ (.A(_00980_),
    .Y(_16144_));
 NAND2x1_ASAP7_75t_R _33572_ (.A(_13168_),
    .B(_00978_),
    .Y(_16145_));
 OA211x2_ASAP7_75t_R _33573_ (.A1(_13166_),
    .A2(_16144_),
    .B(_16145_),
    .C(_13140_),
    .Y(_16146_));
 INVx2_ASAP7_75t_R _33574_ (.A(_00979_),
    .Y(_16147_));
 NAND2x1_ASAP7_75t_R _33575_ (.A(_13137_),
    .B(_00977_),
    .Y(_16148_));
 OA211x2_ASAP7_75t_R _33576_ (.A1(_13143_),
    .A2(_16147_),
    .B(_16148_),
    .C(_13174_),
    .Y(_16149_));
 OR3x1_ASAP7_75t_R _33577_ (.A(_13131_),
    .B(_16146_),
    .C(_16149_),
    .Y(_16150_));
 INVx2_ASAP7_75t_R _33578_ (.A(_00988_),
    .Y(_16151_));
 NAND2x1_ASAP7_75t_R _33579_ (.A(_13168_),
    .B(_00986_),
    .Y(_16152_));
 OA211x2_ASAP7_75t_R _33580_ (.A1(_13133_),
    .A2(_16151_),
    .B(_16152_),
    .C(_13140_),
    .Y(_16153_));
 INVx2_ASAP7_75t_R _33581_ (.A(_00987_),
    .Y(_16154_));
 NAND2x1_ASAP7_75t_R _33582_ (.A(_13146_),
    .B(_00985_),
    .Y(_16155_));
 OA211x2_ASAP7_75t_R _33583_ (.A1(_13143_),
    .A2(_16154_),
    .B(_16155_),
    .C(_13149_),
    .Y(_16156_));
 OR3x1_ASAP7_75t_R _33584_ (.A(_13153_),
    .B(_16153_),
    .C(_16156_),
    .Y(_16157_));
 AND3x4_ASAP7_75t_R _33585_ (.A(_13129_),
    .B(_16150_),
    .C(_16157_),
    .Y(_16158_));
 OR3x2_ASAP7_75t_R _33586_ (.A(_13082_),
    .B(_16143_),
    .C(_16158_),
    .Y(_16159_));
 INVx2_ASAP7_75t_R _33587_ (.A(_00996_),
    .Y(_16160_));
 NAND2x1_ASAP7_75t_R _33588_ (.A(_13168_),
    .B(_00994_),
    .Y(_16161_));
 OA211x2_ASAP7_75t_R _33589_ (.A1(_13166_),
    .A2(_16160_),
    .B(_16161_),
    .C(_13140_),
    .Y(_16162_));
 INVx1_ASAP7_75t_R _33590_ (.A(_00995_),
    .Y(_16163_));
 NAND2x1_ASAP7_75t_R _33591_ (.A(_13137_),
    .B(_00993_),
    .Y(_16164_));
 OA211x2_ASAP7_75t_R _33592_ (.A1(_13133_),
    .A2(_16163_),
    .B(_16164_),
    .C(_13174_),
    .Y(_16165_));
 OR3x1_ASAP7_75t_R _33593_ (.A(_13131_),
    .B(_16162_),
    .C(_16165_),
    .Y(_16166_));
 INVx1_ASAP7_75t_R _33594_ (.A(_01004_),
    .Y(_16167_));
 NAND2x1_ASAP7_75t_R _33595_ (.A(_13168_),
    .B(_01002_),
    .Y(_16168_));
 OA211x2_ASAP7_75t_R _33596_ (.A1(_13133_),
    .A2(_16167_),
    .B(_16168_),
    .C(_13140_),
    .Y(_16169_));
 INVx2_ASAP7_75t_R _33597_ (.A(_01003_),
    .Y(_16170_));
 NAND2x1_ASAP7_75t_R _33598_ (.A(_13137_),
    .B(_01001_),
    .Y(_16171_));
 OA211x2_ASAP7_75t_R _33599_ (.A1(_13143_),
    .A2(_16170_),
    .B(_16171_),
    .C(_13174_),
    .Y(_16172_));
 OR3x1_ASAP7_75t_R _33600_ (.A(_13153_),
    .B(_16169_),
    .C(_16172_),
    .Y(_16173_));
 AND3x1_ASAP7_75t_R _33601_ (.A(_13129_),
    .B(_16166_),
    .C(_16173_),
    .Y(_16174_));
 INVx2_ASAP7_75t_R _33602_ (.A(_00997_),
    .Y(_16175_));
 NOR2x1_ASAP7_75t_R _33603_ (.A(_14516_),
    .B(_00999_),
    .Y(_16176_));
 AO21x1_ASAP7_75t_R _33604_ (.A1(_13190_),
    .A2(_16175_),
    .B(_16176_),
    .Y(_16177_));
 INVx2_ASAP7_75t_R _33605_ (.A(_01000_),
    .Y(_16178_));
 NAND2x1_ASAP7_75t_R _33606_ (.A(_13200_),
    .B(_00998_),
    .Y(_16179_));
 OA211x2_ASAP7_75t_R _33607_ (.A1(_13197_),
    .A2(_16178_),
    .B(_16179_),
    .C(_13202_),
    .Y(_16180_));
 AO21x1_ASAP7_75t_R _33608_ (.A1(_13187_),
    .A2(_16177_),
    .B(_16180_),
    .Y(_16181_));
 INVx2_ASAP7_75t_R _33609_ (.A(_00992_),
    .Y(_16182_));
 NAND2x1_ASAP7_75t_R _33610_ (.A(_13118_),
    .B(_00990_),
    .Y(_16183_));
 OA211x2_ASAP7_75t_R _33611_ (.A1(_13107_),
    .A2(_16182_),
    .B(_16183_),
    .C(_13115_),
    .Y(_16184_));
 INVx2_ASAP7_75t_R _33612_ (.A(_00991_),
    .Y(_16185_));
 NAND2x1_ASAP7_75t_R _33613_ (.A(_13211_),
    .B(_00989_),
    .Y(_16186_));
 OA211x2_ASAP7_75t_R _33614_ (.A1(_13206_),
    .A2(_16185_),
    .B(_16186_),
    .C(_13120_),
    .Y(_16187_));
 OR3x1_ASAP7_75t_R _33615_ (.A(_13085_),
    .B(_16184_),
    .C(_16187_),
    .Y(_16188_));
 OA211x2_ASAP7_75t_R _33616_ (.A1(_13186_),
    .A2(_16181_),
    .B(_16188_),
    .C(_13125_),
    .Y(_16189_));
 OR3x2_ASAP7_75t_R _33617_ (.A(_13164_),
    .B(_16174_),
    .C(_16189_),
    .Y(_16190_));
 AO21x2_ASAP7_75t_R _33618_ (.A1(_16159_),
    .A2(_16190_),
    .B(_13268_),
    .Y(_16191_));
 BUFx6f_ASAP7_75t_R _33619_ (.A(_01497_),
    .Y(_16192_));
 AND2x2_ASAP7_75t_R _33620_ (.A(_01467_),
    .B(_15100_),
    .Y(_16193_));
 OAI22x1_ASAP7_75t_R _33621_ (.A1(_16192_),
    .A2(_14382_),
    .B1(_14385_),
    .B2(_16193_),
    .Y(_16194_));
 NAND2x2_ASAP7_75t_R _33622_ (.A(_16191_),
    .B(_16194_),
    .Y(_18648_));
 INVx1_ASAP7_75t_R _33623_ (.A(_18648_),
    .Y(_18650_));
 BUFx6f_ASAP7_75t_R _33624_ (.A(_00105_),
    .Y(_16195_));
 OR3x1_ASAP7_75t_R _33625_ (.A(_16195_),
    .B(_14627_),
    .C(_14649_),
    .Y(_16196_));
 OAI21x1_ASAP7_75t_R _33626_ (.A1(_14646_),
    .A2(_18648_),
    .B(_16196_),
    .Y(_18046_));
 AND2x2_ASAP7_75t_R _33627_ (.A(_15307_),
    .B(_01777_),
    .Y(_16197_));
 AO21x1_ASAP7_75t_R _33628_ (.A1(_15436_),
    .A2(_00976_),
    .B(_16197_),
    .Y(_16198_));
 OAI22x1_ASAP7_75t_R _33629_ (.A1(_00975_),
    .A2(_15435_),
    .B1(_16198_),
    .B2(_15296_),
    .Y(_16199_));
 NAND2x1_ASAP7_75t_R _33630_ (.A(_15354_),
    .B(_00982_),
    .Y(_16200_));
 OA211x2_ASAP7_75t_R _33631_ (.A1(_15441_),
    .A2(_16136_),
    .B(_16200_),
    .C(_15443_),
    .Y(_16201_));
 NAND2x1_ASAP7_75t_R _33632_ (.A(_15302_),
    .B(_00981_),
    .Y(_16202_));
 OA211x2_ASAP7_75t_R _33633_ (.A1(_15441_),
    .A2(_16139_),
    .B(_16202_),
    .C(_15497_),
    .Y(_16203_));
 OR3x1_ASAP7_75t_R _33634_ (.A(_15298_),
    .B(_16201_),
    .C(_16203_),
    .Y(_16204_));
 OA211x2_ASAP7_75t_R _33635_ (.A1(_15588_),
    .A2(_16199_),
    .B(_16204_),
    .C(_15360_),
    .Y(_16205_));
 NAND2x1_ASAP7_75t_R _33636_ (.A(_15270_),
    .B(_00978_),
    .Y(_16206_));
 OA211x2_ASAP7_75t_R _33637_ (.A1(_15346_),
    .A2(_16144_),
    .B(_16206_),
    .C(_15349_),
    .Y(_16207_));
 NAND2x1_ASAP7_75t_R _33638_ (.A(_15451_),
    .B(_00977_),
    .Y(_16208_));
 OA211x2_ASAP7_75t_R _33639_ (.A1(_15346_),
    .A2(_16147_),
    .B(_16208_),
    .C(_15456_),
    .Y(_16209_));
 OR3x1_ASAP7_75t_R _33640_ (.A(_15318_),
    .B(_16207_),
    .C(_16209_),
    .Y(_16210_));
 NAND2x1_ASAP7_75t_R _33641_ (.A(_15270_),
    .B(_00986_),
    .Y(_16211_));
 OA211x2_ASAP7_75t_R _33642_ (.A1(_15346_),
    .A2(_16151_),
    .B(_16211_),
    .C(_15349_),
    .Y(_16212_));
 NAND2x1_ASAP7_75t_R _33643_ (.A(_15451_),
    .B(_00985_),
    .Y(_16213_));
 OA211x2_ASAP7_75t_R _33644_ (.A1(_15450_),
    .A2(_16154_),
    .B(_16213_),
    .C(_15456_),
    .Y(_16214_));
 OR3x1_ASAP7_75t_R _33645_ (.A(_15475_),
    .B(_16212_),
    .C(_16214_),
    .Y(_16215_));
 AND3x4_ASAP7_75t_R _33646_ (.A(_15317_),
    .B(_16210_),
    .C(_16215_),
    .Y(_16216_));
 OR3x2_ASAP7_75t_R _33647_ (.A(_15434_),
    .B(_16205_),
    .C(_16216_),
    .Y(_16217_));
 BUFx6f_ASAP7_75t_R _33648_ (.A(_15252_),
    .Y(_16218_));
 NAND2x1_ASAP7_75t_R _33649_ (.A(_15321_),
    .B(_00994_),
    .Y(_16219_));
 OA211x2_ASAP7_75t_R _33650_ (.A1(_15490_),
    .A2(_16160_),
    .B(_16219_),
    .C(_15469_),
    .Y(_16220_));
 NAND2x1_ASAP7_75t_R _33651_ (.A(_15321_),
    .B(_00993_),
    .Y(_16221_));
 OA211x2_ASAP7_75t_R _33652_ (.A1(_15467_),
    .A2(_16163_),
    .B(_16221_),
    .C(_15338_),
    .Y(_16222_));
 OR3x1_ASAP7_75t_R _33653_ (.A(_15318_),
    .B(_16220_),
    .C(_16222_),
    .Y(_16223_));
 NAND2x1_ASAP7_75t_R _33654_ (.A(_15321_),
    .B(_01002_),
    .Y(_16224_));
 OA211x2_ASAP7_75t_R _33655_ (.A1(_15490_),
    .A2(_16167_),
    .B(_16224_),
    .C(_15469_),
    .Y(_16225_));
 NAND2x1_ASAP7_75t_R _33656_ (.A(_15326_),
    .B(_01001_),
    .Y(_16226_));
 OA211x2_ASAP7_75t_R _33657_ (.A1(_15467_),
    .A2(_16170_),
    .B(_16226_),
    .C(_15338_),
    .Y(_16227_));
 OR3x1_ASAP7_75t_R _33658_ (.A(_15475_),
    .B(_16225_),
    .C(_16227_),
    .Y(_16228_));
 AND3x1_ASAP7_75t_R _33659_ (.A(_16218_),
    .B(_16223_),
    .C(_16228_),
    .Y(_16229_));
 NOR2x1_ASAP7_75t_R _33660_ (.A(_15343_),
    .B(_00999_),
    .Y(_16230_));
 AO21x1_ASAP7_75t_R _33661_ (.A1(_15484_),
    .A2(_16175_),
    .B(_16230_),
    .Y(_16231_));
 NAND2x1_ASAP7_75t_R _33662_ (.A(_15347_),
    .B(_00998_),
    .Y(_16232_));
 OA211x2_ASAP7_75t_R _33663_ (.A1(_15598_),
    .A2(_16178_),
    .B(_16232_),
    .C(_15469_),
    .Y(_16233_));
 AO21x1_ASAP7_75t_R _33664_ (.A1(_15339_),
    .A2(_16231_),
    .B(_16233_),
    .Y(_16234_));
 NAND2x1_ASAP7_75t_R _33665_ (.A(_15483_),
    .B(_00990_),
    .Y(_16235_));
 OA211x2_ASAP7_75t_R _33666_ (.A1(_15441_),
    .A2(_16182_),
    .B(_16235_),
    .C(_15443_),
    .Y(_16236_));
 NAND2x1_ASAP7_75t_R _33667_ (.A(_15354_),
    .B(_00989_),
    .Y(_16237_));
 OA211x2_ASAP7_75t_R _33668_ (.A1(_15441_),
    .A2(_16185_),
    .B(_16237_),
    .C(_15497_),
    .Y(_16238_));
 OR3x1_ASAP7_75t_R _33669_ (.A(_15352_),
    .B(_16236_),
    .C(_16238_),
    .Y(_16239_));
 OA211x2_ASAP7_75t_R _33670_ (.A1(_15482_),
    .A2(_16234_),
    .B(_16239_),
    .C(_15360_),
    .Y(_16240_));
 OR3x2_ASAP7_75t_R _33671_ (.A(_15466_),
    .B(_16229_),
    .C(_16240_),
    .Y(_16241_));
 NAND2x2_ASAP7_75t_R _33672_ (.A(_16217_),
    .B(_16241_),
    .Y(_16242_));
 OA211x2_ASAP7_75t_R _33673_ (.A1(_14339_),
    .A2(_15366_),
    .B(_15369_),
    .C(_15503_),
    .Y(_16243_));
 AOI21x1_ASAP7_75t_R _33674_ (.A1(_14090_),
    .A2(_16242_),
    .B(_16243_),
    .Y(_18649_));
 INVx1_ASAP7_75t_R _33675_ (.A(_18649_),
    .Y(_18647_));
 INVx2_ASAP7_75t_R _33676_ (.A(net1951),
    .Y(_16244_));
 AND3x1_ASAP7_75t_R _33677_ (.A(_00974_),
    .B(_01006_),
    .C(_16244_),
    .Y(_16245_));
 BUFx6f_ASAP7_75t_R _33678_ (.A(_00973_),
    .Y(_16246_));
 OAI21x1_ASAP7_75t_R _33679_ (.A1(_00974_),
    .A2(_16246_),
    .B(_01006_),
    .Y(_16247_));
 AO21x1_ASAP7_75t_R _33680_ (.A1(net1940),
    .A2(_00974_),
    .B(_16246_),
    .Y(_16248_));
 AND3x1_ASAP7_75t_R _33681_ (.A(_01006_),
    .B(_16244_),
    .C(_16248_),
    .Y(_16249_));
 AO21x1_ASAP7_75t_R _33682_ (.A1(net1951),
    .A2(_16247_),
    .B(_16249_),
    .Y(_16250_));
 NOR2x1_ASAP7_75t_R _33683_ (.A(net1940),
    .B(_16246_),
    .Y(_16251_));
 OA211x2_ASAP7_75t_R _33684_ (.A1(_15999_),
    .A2(_16002_),
    .B(_16251_),
    .C(net1951),
    .Y(_16252_));
 AOI211x1_ASAP7_75t_R _33685_ (.A1(_16003_),
    .A2(_16245_),
    .B(_16250_),
    .C(_16252_),
    .Y(_16253_));
 INVx3_ASAP7_75t_R _33686_ (.A(_16253_),
    .Y(\alu_adder_result_ex[19] ));
 INVx2_ASAP7_75t_R _33687_ (.A(_16246_),
    .Y(_16254_));
 OA21x2_ASAP7_75t_R _33688_ (.A1(_15997_),
    .A2(_16010_),
    .B(_00942_),
    .Y(_16255_));
 OA21x2_ASAP7_75t_R _33689_ (.A1(net1940),
    .A2(_16255_),
    .B(_00974_),
    .Y(_16256_));
 AND4x1_ASAP7_75t_R _33690_ (.A(_16254_),
    .B(_15247_),
    .C(_15766_),
    .D(_16256_),
    .Y(_16257_));
 OR3x1_ASAP7_75t_R _33691_ (.A(_15997_),
    .B(net1940),
    .C(_16008_),
    .Y(_16258_));
 OR3x1_ASAP7_75t_R _33692_ (.A(_16254_),
    .B(_15768_),
    .C(_16258_),
    .Y(_16259_));
 NOR2x1_ASAP7_75t_R _33693_ (.A(_15247_),
    .B(_16259_),
    .Y(_16260_));
 INVx1_ASAP7_75t_R _33694_ (.A(_16256_),
    .Y(_16261_));
 AND3x1_ASAP7_75t_R _33695_ (.A(_16254_),
    .B(_16256_),
    .C(_16258_),
    .Y(_16262_));
 AND4x1_ASAP7_75t_R _33696_ (.A(_16254_),
    .B(_15766_),
    .C(_15768_),
    .D(_16256_),
    .Y(_16263_));
 AOI211x1_ASAP7_75t_R _33697_ (.A1(_16246_),
    .A2(_16261_),
    .B(_16262_),
    .C(_16263_),
    .Y(_16264_));
 OR3x1_ASAP7_75t_R _33698_ (.A(_16254_),
    .B(_15766_),
    .C(_16258_),
    .Y(_16265_));
 NAND2x1_ASAP7_75t_R _33699_ (.A(_16264_),
    .B(_16265_),
    .Y(_16266_));
 NOR3x2_ASAP7_75t_R _33700_ (.B(_16260_),
    .C(_16266_),
    .Y(_16267_),
    .A(_16257_));
 INVx4_ASAP7_75t_R _33701_ (.A(_16267_),
    .Y(\alu_adder_result_ex[18] ));
 AND2x2_ASAP7_75t_R _33702_ (.A(_13206_),
    .B(_01776_),
    .Y(_16268_));
 AO21x1_ASAP7_75t_R _33703_ (.A1(_14286_),
    .A2(_01008_),
    .B(_16268_),
    .Y(_16269_));
 OAI22x1_ASAP7_75t_R _33704_ (.A1(_01007_),
    .A2(_14284_),
    .B1(_16269_),
    .B2(_13090_),
    .Y(_16270_));
 INVx2_ASAP7_75t_R _33705_ (.A(_01016_),
    .Y(_16271_));
 NAND2x1_ASAP7_75t_R _33706_ (.A(_14492_),
    .B(_01014_),
    .Y(_16272_));
 OA211x2_ASAP7_75t_R _33707_ (.A1(_14501_),
    .A2(_16271_),
    .B(_16272_),
    .C(_14504_),
    .Y(_16273_));
 INVx2_ASAP7_75t_R _33708_ (.A(_01015_),
    .Y(_16274_));
 NAND2x1_ASAP7_75t_R _33709_ (.A(_14507_),
    .B(_01013_),
    .Y(_16275_));
 OA211x2_ASAP7_75t_R _33710_ (.A1(_14506_),
    .A2(_16274_),
    .B(_16275_),
    .C(_14509_),
    .Y(_16276_));
 OR3x1_ASAP7_75t_R _33711_ (.A(_14353_),
    .B(_16273_),
    .C(_16276_),
    .Y(_16277_));
 OA211x2_ASAP7_75t_R _33712_ (.A1(_13086_),
    .A2(_16270_),
    .B(_16277_),
    .C(_14852_),
    .Y(_16278_));
 INVx2_ASAP7_75t_R _33713_ (.A(_01012_),
    .Y(_16279_));
 NAND2x1_ASAP7_75t_R _33714_ (.A(_15061_),
    .B(_01010_),
    .Y(_16280_));
 OA211x2_ASAP7_75t_R _33715_ (.A1(_15120_),
    .A2(_16279_),
    .B(_16280_),
    .C(_13202_),
    .Y(_16281_));
 INVx2_ASAP7_75t_R _33716_ (.A(_01011_),
    .Y(_16282_));
 NAND2x1_ASAP7_75t_R _33717_ (.A(_14738_),
    .B(_01009_),
    .Y(_16283_));
 OA211x2_ASAP7_75t_R _33718_ (.A1(_13197_),
    .A2(_16282_),
    .B(_16283_),
    .C(_14874_),
    .Y(_16284_));
 OR3x1_ASAP7_75t_R _33719_ (.A(_15117_),
    .B(_16281_),
    .C(_16284_),
    .Y(_16285_));
 INVx2_ASAP7_75t_R _33720_ (.A(_01020_),
    .Y(_16286_));
 NAND2x1_ASAP7_75t_R _33721_ (.A(_15061_),
    .B(_01018_),
    .Y(_16287_));
 OA211x2_ASAP7_75t_R _33722_ (.A1(_15120_),
    .A2(_16286_),
    .B(_16287_),
    .C(_13202_),
    .Y(_16288_));
 INVx2_ASAP7_75t_R _33723_ (.A(_01019_),
    .Y(_16289_));
 NAND2x1_ASAP7_75t_R _33724_ (.A(_13200_),
    .B(_01017_),
    .Y(_16290_));
 OA211x2_ASAP7_75t_R _33725_ (.A1(_13197_),
    .A2(_16289_),
    .B(_16290_),
    .C(_14874_),
    .Y(_16291_));
 OR3x1_ASAP7_75t_R _33726_ (.A(_14877_),
    .B(_16288_),
    .C(_16291_),
    .Y(_16292_));
 AND3x4_ASAP7_75t_R _33727_ (.A(_14340_),
    .B(_16285_),
    .C(_16292_),
    .Y(_16293_));
 OR3x2_ASAP7_75t_R _33728_ (.A(_13082_),
    .B(_16278_),
    .C(_16293_),
    .Y(_16294_));
 INVx2_ASAP7_75t_R _33729_ (.A(_01028_),
    .Y(_16295_));
 NAND2x1_ASAP7_75t_R _33730_ (.A(_14782_),
    .B(_01026_),
    .Y(_16296_));
 OA211x2_ASAP7_75t_R _33731_ (.A1(_14711_),
    .A2(_16295_),
    .B(_16296_),
    .C(_13202_),
    .Y(_16297_));
 INVx2_ASAP7_75t_R _33732_ (.A(_01027_),
    .Y(_16298_));
 NAND2x1_ASAP7_75t_R _33733_ (.A(_14738_),
    .B(_01025_),
    .Y(_16299_));
 OA211x2_ASAP7_75t_R _33734_ (.A1(_15120_),
    .A2(_16298_),
    .B(_16299_),
    .C(_15122_),
    .Y(_16300_));
 OR3x1_ASAP7_75t_R _33735_ (.A(_15117_),
    .B(_16297_),
    .C(_16300_),
    .Y(_16301_));
 INVx2_ASAP7_75t_R _33736_ (.A(_01036_),
    .Y(_16302_));
 NAND2x1_ASAP7_75t_R _33737_ (.A(_15061_),
    .B(_01034_),
    .Y(_16303_));
 OA211x2_ASAP7_75t_R _33738_ (.A1(_14711_),
    .A2(_16302_),
    .B(_16303_),
    .C(_13202_),
    .Y(_16304_));
 INVx2_ASAP7_75t_R _33739_ (.A(_01035_),
    .Y(_16305_));
 NAND2x1_ASAP7_75t_R _33740_ (.A(_14738_),
    .B(_01033_),
    .Y(_16306_));
 OA211x2_ASAP7_75t_R _33741_ (.A1(_15120_),
    .A2(_16305_),
    .B(_16306_),
    .C(_14874_),
    .Y(_16307_));
 OR3x1_ASAP7_75t_R _33742_ (.A(_14877_),
    .B(_16304_),
    .C(_16307_),
    .Y(_16308_));
 AND3x1_ASAP7_75t_R _33743_ (.A(_14340_),
    .B(_16301_),
    .C(_16308_),
    .Y(_16309_));
 INVx2_ASAP7_75t_R _33744_ (.A(_01029_),
    .Y(_16310_));
 NOR2x1_ASAP7_75t_R _33745_ (.A(_14366_),
    .B(_01031_),
    .Y(_16311_));
 AO21x1_ASAP7_75t_R _33746_ (.A1(_13190_),
    .A2(_16310_),
    .B(_16311_),
    .Y(_16312_));
 INVx2_ASAP7_75t_R _33747_ (.A(_01032_),
    .Y(_16313_));
 NAND2x1_ASAP7_75t_R _33748_ (.A(_14333_),
    .B(_01030_),
    .Y(_16314_));
 OA211x2_ASAP7_75t_R _33749_ (.A1(_14331_),
    .A2(_16313_),
    .B(_16314_),
    .C(_14329_),
    .Y(_16315_));
 AO21x1_ASAP7_75t_R _33750_ (.A1(_14975_),
    .A2(_16312_),
    .B(_16315_),
    .Y(_16316_));
 INVx2_ASAP7_75t_R _33751_ (.A(_01024_),
    .Y(_16317_));
 NAND2x1_ASAP7_75t_R _33752_ (.A(_14507_),
    .B(_01022_),
    .Y(_16318_));
 OA211x2_ASAP7_75t_R _33753_ (.A1(_14506_),
    .A2(_16317_),
    .B(_16318_),
    .C(_14472_),
    .Y(_16319_));
 INVx2_ASAP7_75t_R _33754_ (.A(_01023_),
    .Y(_16320_));
 NAND2x1_ASAP7_75t_R _33755_ (.A(_14517_),
    .B(_01021_),
    .Y(_16321_));
 OA211x2_ASAP7_75t_R _33756_ (.A1(_13193_),
    .A2(_16320_),
    .B(_16321_),
    .C(_14509_),
    .Y(_16322_));
 OR3x1_ASAP7_75t_R _33757_ (.A(_14469_),
    .B(_16319_),
    .C(_16322_),
    .Y(_16323_));
 OA211x2_ASAP7_75t_R _33758_ (.A1(_14354_),
    .A2(_16316_),
    .B(_16323_),
    .C(_14852_),
    .Y(_16324_));
 OR3x2_ASAP7_75t_R _33759_ (.A(_13164_),
    .B(_16309_),
    .C(_16324_),
    .Y(_16325_));
 AO21x2_ASAP7_75t_R _33760_ (.A1(_16294_),
    .A2(_16325_),
    .B(_14377_),
    .Y(_16326_));
 AND2x2_ASAP7_75t_R _33761_ (.A(_01465_),
    .B(_15100_),
    .Y(_16327_));
 OAI22x1_ASAP7_75t_R _33762_ (.A1(_01495_),
    .A2(_14382_),
    .B1(_14385_),
    .B2(_16327_),
    .Y(_16328_));
 AND2x4_ASAP7_75t_R _33763_ (.A(_16326_),
    .B(_16328_),
    .Y(_18655_));
 INVx2_ASAP7_75t_R _33764_ (.A(_18655_),
    .Y(_18653_));
 BUFx6f_ASAP7_75t_R _33765_ (.A(_00110_),
    .Y(_16329_));
 INVx1_ASAP7_75t_R _33766_ (.A(_16329_),
    .Y(_16330_));
 AND3x1_ASAP7_75t_R _33767_ (.A(_16330_),
    .B(_15236_),
    .C(_14907_),
    .Y(_16331_));
 AO21x1_ASAP7_75t_R _33768_ (.A1(_14903_),
    .A2(_18655_),
    .B(_16331_),
    .Y(_18048_));
 BUFx12f_ASAP7_75t_R _33769_ (.A(_15486_),
    .Y(_16332_));
 BUFx6f_ASAP7_75t_R _33770_ (.A(_15291_),
    .Y(_16333_));
 NOR2x1_ASAP7_75t_R _33771_ (.A(_16333_),
    .B(_01031_),
    .Y(_16334_));
 AO21x1_ASAP7_75t_R _33772_ (.A1(_16332_),
    .A2(_16310_),
    .B(_16334_),
    .Y(_16335_));
 NAND2x1_ASAP7_75t_R _33773_ (.A(_15484_),
    .B(_01030_),
    .Y(_16336_));
 BUFx12f_ASAP7_75t_R _33774_ (.A(_15752_),
    .Y(_16337_));
 OA211x2_ASAP7_75t_R _33775_ (.A1(_16332_),
    .A2(_16313_),
    .B(_16336_),
    .C(_16337_),
    .Y(_16338_));
 AO21x1_ASAP7_75t_R _33776_ (.A1(_15594_),
    .A2(_16335_),
    .B(_16338_),
    .Y(_16339_));
 NAND2x1_ASAP7_75t_R _33777_ (.A(_15341_),
    .B(_01022_),
    .Y(_16340_));
 OA211x2_ASAP7_75t_R _33778_ (.A1(_16332_),
    .A2(_16317_),
    .B(_16340_),
    .C(_16337_),
    .Y(_16341_));
 NAND2x1_ASAP7_75t_R _33779_ (.A(_15633_),
    .B(_01021_),
    .Y(_16342_));
 OA211x2_ASAP7_75t_R _33780_ (.A1(_16332_),
    .A2(_16320_),
    .B(_16342_),
    .C(_15593_),
    .Y(_16343_));
 OA21x2_ASAP7_75t_R _33781_ (.A1(_16341_),
    .A2(_16343_),
    .B(_15482_),
    .Y(_16344_));
 AO21x1_ASAP7_75t_R _33782_ (.A1(_15588_),
    .A2(_16339_),
    .B(_16344_),
    .Y(_16345_));
 NAND2x1_ASAP7_75t_R _33783_ (.A(_15467_),
    .B(_01026_),
    .Y(_16346_));
 OA211x2_ASAP7_75t_R _33784_ (.A1(_16333_),
    .A2(_16295_),
    .B(_16346_),
    .C(_16337_),
    .Y(_16347_));
 NAND2x1_ASAP7_75t_R _33785_ (.A(_15467_),
    .B(_01025_),
    .Y(_16348_));
 OA211x2_ASAP7_75t_R _33786_ (.A1(_16333_),
    .A2(_16298_),
    .B(_16348_),
    .C(_15593_),
    .Y(_16349_));
 OR3x1_ASAP7_75t_R _33787_ (.A(_15288_),
    .B(_16347_),
    .C(_16349_),
    .Y(_16350_));
 NAND2x1_ASAP7_75t_R _33788_ (.A(_15467_),
    .B(_01034_),
    .Y(_16351_));
 OA211x2_ASAP7_75t_R _33789_ (.A1(_16333_),
    .A2(_16302_),
    .B(_16351_),
    .C(_16337_),
    .Y(_16352_));
 NAND2x1_ASAP7_75t_R _33790_ (.A(_15471_),
    .B(_01033_),
    .Y(_16353_));
 BUFx6f_ASAP7_75t_R _33791_ (.A(_15592_),
    .Y(_16354_));
 OA211x2_ASAP7_75t_R _33792_ (.A1(_16333_),
    .A2(_16305_),
    .B(_16353_),
    .C(_16354_),
    .Y(_16355_));
 OR3x1_ASAP7_75t_R _33793_ (.A(_15337_),
    .B(_16352_),
    .C(_16355_),
    .Y(_16356_));
 AND3x1_ASAP7_75t_R _33794_ (.A(_16218_),
    .B(_16350_),
    .C(_16356_),
    .Y(_16357_));
 AO21x1_ASAP7_75t_R _33795_ (.A1(_15587_),
    .A2(_16345_),
    .B(_16357_),
    .Y(_16358_));
 AND2x2_ASAP7_75t_R _33796_ (.A(_15598_),
    .B(_01776_),
    .Y(_16359_));
 AO21x1_ASAP7_75t_R _33797_ (.A1(_15436_),
    .A2(_01008_),
    .B(_16359_),
    .Y(_16360_));
 OAI22x1_ASAP7_75t_R _33798_ (.A1(_01007_),
    .A2(_15435_),
    .B1(_16360_),
    .B2(_15594_),
    .Y(_16361_));
 NAND2x1_ASAP7_75t_R _33799_ (.A(_15300_),
    .B(_01014_),
    .Y(_16362_));
 OA211x2_ASAP7_75t_R _33800_ (.A1(_15341_),
    .A2(_16271_),
    .B(_16362_),
    .C(_15600_),
    .Y(_16363_));
 NAND2x1_ASAP7_75t_R _33801_ (.A(_15300_),
    .B(_01013_),
    .Y(_16364_));
 OA211x2_ASAP7_75t_R _33802_ (.A1(_15633_),
    .A2(_16274_),
    .B(_16364_),
    .C(_15295_),
    .Y(_16365_));
 OR3x1_ASAP7_75t_R _33803_ (.A(_15596_),
    .B(_16363_),
    .C(_16365_),
    .Y(_16366_));
 OA211x2_ASAP7_75t_R _33804_ (.A1(_15588_),
    .A2(_16361_),
    .B(_16366_),
    .C(_15587_),
    .Y(_16367_));
 BUFx6f_ASAP7_75t_R _33805_ (.A(_15254_),
    .Y(_16368_));
 BUFx6f_ASAP7_75t_R _33806_ (.A(_15291_),
    .Y(_16369_));
 NAND2x1_ASAP7_75t_R _33807_ (.A(_15269_),
    .B(_01010_),
    .Y(_16370_));
 BUFx6f_ASAP7_75t_R _33808_ (.A(_15752_),
    .Y(_16371_));
 OA211x2_ASAP7_75t_R _33809_ (.A1(_16369_),
    .A2(_16279_),
    .B(_16370_),
    .C(_16371_),
    .Y(_16372_));
 BUFx6f_ASAP7_75t_R _33810_ (.A(_15321_),
    .Y(_16373_));
 NAND2x1_ASAP7_75t_R _33811_ (.A(_15622_),
    .B(_01009_),
    .Y(_16374_));
 OA211x2_ASAP7_75t_R _33812_ (.A1(_16373_),
    .A2(_16282_),
    .B(_16374_),
    .C(_16354_),
    .Y(_16375_));
 OR3x1_ASAP7_75t_R _33813_ (.A(_16368_),
    .B(_16372_),
    .C(_16375_),
    .Y(_16376_));
 NAND2x1_ASAP7_75t_R _33814_ (.A(_15269_),
    .B(_01018_),
    .Y(_16377_));
 OA211x2_ASAP7_75t_R _33815_ (.A1(_16369_),
    .A2(_16286_),
    .B(_16377_),
    .C(_16371_),
    .Y(_16378_));
 NAND2x1_ASAP7_75t_R _33816_ (.A(_15622_),
    .B(_01017_),
    .Y(_16379_));
 OA211x2_ASAP7_75t_R _33817_ (.A1(_16373_),
    .A2(_16289_),
    .B(_16379_),
    .C(_16354_),
    .Y(_16380_));
 OR3x1_ASAP7_75t_R _33818_ (.A(_15596_),
    .B(_16378_),
    .C(_16380_),
    .Y(_16381_));
 AND3x1_ASAP7_75t_R _33819_ (.A(_16218_),
    .B(_16376_),
    .C(_16381_),
    .Y(_16382_));
 OR3x1_ASAP7_75t_R _33820_ (.A(_15434_),
    .B(_16367_),
    .C(_16382_),
    .Y(_16383_));
 OA21x2_ASAP7_75t_R _33821_ (.A1(_15466_),
    .A2(_16358_),
    .B(_16383_),
    .Y(_16384_));
 INVx2_ASAP7_75t_R _33822_ (.A(_16384_),
    .Y(_16385_));
 BUFx6f_ASAP7_75t_R _33823_ (.A(_15364_),
    .Y(_16386_));
 OR3x2_ASAP7_75t_R _33824_ (.A(_13272_),
    .B(_14267_),
    .C(_13535_),
    .Y(_16387_));
 OR2x2_ASAP7_75t_R _33825_ (.A(_14099_),
    .B(_16387_),
    .Y(_16388_));
 BUFx3_ASAP7_75t_R _33826_ (.A(_16388_),
    .Y(_16389_));
 OA211x2_ASAP7_75t_R _33827_ (.A1(_15594_),
    .A2(_16386_),
    .B(_16389_),
    .C(_15503_),
    .Y(_16390_));
 AOI21x1_ASAP7_75t_R _33828_ (.A1(_14090_),
    .A2(_16385_),
    .B(_16390_),
    .Y(_18654_));
 INVx1_ASAP7_75t_R _33829_ (.A(_18654_),
    .Y(_18652_));
 AND2x2_ASAP7_75t_R _33830_ (.A(_14506_),
    .B(_01775_),
    .Y(_16391_));
 AO21x1_ASAP7_75t_R _33831_ (.A1(_14286_),
    .A2(_01040_),
    .B(_16391_),
    .Y(_16392_));
 OAI22x1_ASAP7_75t_R _33832_ (.A1(_01039_),
    .A2(_14284_),
    .B1(_16392_),
    .B2(_14289_),
    .Y(_16393_));
 INVx2_ASAP7_75t_R _33833_ (.A(_01048_),
    .Y(_16394_));
 NAND2x1_ASAP7_75t_R _33834_ (.A(_14794_),
    .B(_01046_),
    .Y(_16395_));
 OA211x2_ASAP7_75t_R _33835_ (.A1(_14293_),
    .A2(_16394_),
    .B(_16395_),
    .C(_14296_),
    .Y(_16396_));
 INVx2_ASAP7_75t_R _33836_ (.A(_01047_),
    .Y(_16397_));
 NAND2x1_ASAP7_75t_R _33837_ (.A(_14794_),
    .B(_01045_),
    .Y(_16398_));
 OA211x2_ASAP7_75t_R _33838_ (.A1(_14293_),
    .A2(_16397_),
    .B(_16398_),
    .C(_13149_),
    .Y(_16399_));
 OR3x1_ASAP7_75t_R _33839_ (.A(_13153_),
    .B(_16396_),
    .C(_16399_),
    .Y(_16400_));
 OA211x2_ASAP7_75t_R _33840_ (.A1(_14283_),
    .A2(_16393_),
    .B(_16400_),
    .C(_14305_),
    .Y(_16401_));
 INVx2_ASAP7_75t_R _33841_ (.A(_01044_),
    .Y(_16402_));
 NAND2x1_ASAP7_75t_R _33842_ (.A(_14455_),
    .B(_01042_),
    .Y(_16403_));
 OA211x2_ASAP7_75t_R _33843_ (.A1(_14358_),
    .A2(_16402_),
    .B(_16403_),
    .C(_14363_),
    .Y(_16404_));
 INVx2_ASAP7_75t_R _33844_ (.A(_01043_),
    .Y(_16405_));
 NAND2x1_ASAP7_75t_R _33845_ (.A(_15052_),
    .B(_01041_),
    .Y(_16406_));
 OA211x2_ASAP7_75t_R _33846_ (.A1(_15191_),
    .A2(_16405_),
    .B(_16406_),
    .C(_15195_),
    .Y(_16407_));
 OR3x1_ASAP7_75t_R _33847_ (.A(_14309_),
    .B(_16404_),
    .C(_16407_),
    .Y(_16408_));
 INVx2_ASAP7_75t_R _33848_ (.A(_01052_),
    .Y(_16409_));
 NAND2x1_ASAP7_75t_R _33849_ (.A(_14461_),
    .B(_01050_),
    .Y(_16410_));
 OA211x2_ASAP7_75t_R _33850_ (.A1(_15191_),
    .A2(_16409_),
    .B(_16410_),
    .C(_14315_),
    .Y(_16411_));
 INVx2_ASAP7_75t_R _33851_ (.A(_01051_),
    .Y(_16412_));
 NAND2x1_ASAP7_75t_R _33852_ (.A(_14312_),
    .B(_01049_),
    .Y(_16413_));
 OA211x2_ASAP7_75t_R _33853_ (.A1(_14311_),
    .A2(_16412_),
    .B(_16413_),
    .C(_15195_),
    .Y(_16414_));
 OR3x1_ASAP7_75t_R _33854_ (.A(_14327_),
    .B(_16411_),
    .C(_16414_),
    .Y(_16415_));
 AND3x4_ASAP7_75t_R _33855_ (.A(_14307_),
    .B(_16408_),
    .C(_16415_),
    .Y(_16416_));
 OR3x1_ASAP7_75t_R _33856_ (.A(_14281_),
    .B(_16401_),
    .C(_16416_),
    .Y(_16417_));
 INVx2_ASAP7_75t_R _33857_ (.A(_01060_),
    .Y(_16418_));
 NAND2x1_ASAP7_75t_R _33858_ (.A(_14461_),
    .B(_01058_),
    .Y(_16419_));
 OA211x2_ASAP7_75t_R _33859_ (.A1(_14358_),
    .A2(_16418_),
    .B(_16419_),
    .C(_14363_),
    .Y(_16420_));
 INVx2_ASAP7_75t_R _33860_ (.A(_01059_),
    .Y(_16421_));
 NAND2x1_ASAP7_75t_R _33861_ (.A(_15052_),
    .B(_01057_),
    .Y(_16422_));
 OA211x2_ASAP7_75t_R _33862_ (.A1(_14311_),
    .A2(_16421_),
    .B(_16422_),
    .C(_15195_),
    .Y(_16423_));
 OR3x1_ASAP7_75t_R _33863_ (.A(_14309_),
    .B(_16420_),
    .C(_16423_),
    .Y(_16424_));
 INVx2_ASAP7_75t_R _33864_ (.A(_01068_),
    .Y(_16425_));
 NAND2x1_ASAP7_75t_R _33865_ (.A(_14461_),
    .B(_01066_),
    .Y(_16426_));
 OA211x2_ASAP7_75t_R _33866_ (.A1(_15191_),
    .A2(_16425_),
    .B(_16426_),
    .C(_14315_),
    .Y(_16427_));
 INVx2_ASAP7_75t_R _33867_ (.A(_01067_),
    .Y(_16428_));
 NAND2x1_ASAP7_75t_R _33868_ (.A(_14312_),
    .B(_01065_),
    .Y(_16429_));
 OA211x2_ASAP7_75t_R _33869_ (.A1(_14311_),
    .A2(_16428_),
    .B(_16429_),
    .C(_15195_),
    .Y(_16430_));
 OR3x1_ASAP7_75t_R _33870_ (.A(_14327_),
    .B(_16427_),
    .C(_16430_),
    .Y(_16431_));
 AND3x1_ASAP7_75t_R _33871_ (.A(_14307_),
    .B(_16424_),
    .C(_16431_),
    .Y(_16432_));
 INVx2_ASAP7_75t_R _33872_ (.A(_01061_),
    .Y(_16433_));
 NOR2x1_ASAP7_75t_R _33873_ (.A(_13133_),
    .B(_01063_),
    .Y(_16434_));
 AO21x1_ASAP7_75t_R _33874_ (.A1(_14278_),
    .A2(_16433_),
    .B(_16434_),
    .Y(_16435_));
 INVx2_ASAP7_75t_R _33875_ (.A(_01064_),
    .Y(_16436_));
 NAND2x1_ASAP7_75t_R _33876_ (.A(_14360_),
    .B(_01062_),
    .Y(_16437_));
 OA211x2_ASAP7_75t_R _33877_ (.A1(_13190_),
    .A2(_16436_),
    .B(_16437_),
    .C(_14363_),
    .Y(_16438_));
 AO21x1_ASAP7_75t_R _33878_ (.A1(_13090_),
    .A2(_16435_),
    .B(_16438_),
    .Y(_16439_));
 INVx2_ASAP7_75t_R _33879_ (.A(_01056_),
    .Y(_16440_));
 NAND2x1_ASAP7_75t_R _33880_ (.A(_14301_),
    .B(_01054_),
    .Y(_16441_));
 OA211x2_ASAP7_75t_R _33881_ (.A1(_14299_),
    .A2(_16440_),
    .B(_16441_),
    .C(_14296_),
    .Y(_16442_));
 INVx2_ASAP7_75t_R _33882_ (.A(_01055_),
    .Y(_16443_));
 NAND2x1_ASAP7_75t_R _33883_ (.A(_14367_),
    .B(_01053_),
    .Y(_16444_));
 OA211x2_ASAP7_75t_R _33884_ (.A1(_14366_),
    .A2(_16443_),
    .B(_16444_),
    .C(_14372_),
    .Y(_16445_));
 OR3x1_ASAP7_75t_R _33885_ (.A(_14282_),
    .B(_16442_),
    .C(_16445_),
    .Y(_16446_));
 OA211x2_ASAP7_75t_R _33886_ (.A1(_14354_),
    .A2(_16439_),
    .B(_16446_),
    .C(_14305_),
    .Y(_16447_));
 OR3x2_ASAP7_75t_R _33887_ (.A(_14339_),
    .B(_16432_),
    .C(_16447_),
    .Y(_16448_));
 AO21x2_ASAP7_75t_R _33888_ (.A1(_16417_),
    .A2(_16448_),
    .B(_13268_),
    .Y(_16449_));
 AND2x2_ASAP7_75t_R _33889_ (.A(_01464_),
    .B(_15100_),
    .Y(_16450_));
 OAI22x1_ASAP7_75t_R _33890_ (.A1(_01494_),
    .A2(_14382_),
    .B1(_14385_),
    .B2(_16450_),
    .Y(_16451_));
 AND2x4_ASAP7_75t_R _33891_ (.A(_16449_),
    .B(_16451_),
    .Y(_18660_));
 INVx2_ASAP7_75t_R _33892_ (.A(_18660_),
    .Y(_18658_));
 INVx2_ASAP7_75t_R _33893_ (.A(_00115_),
    .Y(_16452_));
 AND3x1_ASAP7_75t_R _33894_ (.A(_16452_),
    .B(_15236_),
    .C(_14907_),
    .Y(_16453_));
 AO21x1_ASAP7_75t_R _33895_ (.A1(_14903_),
    .A2(_18660_),
    .B(_16453_),
    .Y(_18050_));
 AND2x2_ASAP7_75t_R _33896_ (.A(_15484_),
    .B(_01775_),
    .Y(_16454_));
 AO21x1_ASAP7_75t_R _33897_ (.A1(_15436_),
    .A2(_01040_),
    .B(_16454_),
    .Y(_16455_));
 OAI22x1_ASAP7_75t_R _33898_ (.A1(_01039_),
    .A2(_15435_),
    .B1(_16455_),
    .B2(_15594_),
    .Y(_16456_));
 NAND2x1_ASAP7_75t_R _33899_ (.A(_15467_),
    .B(_01046_),
    .Y(_16457_));
 OA211x2_ASAP7_75t_R _33900_ (.A1(_16333_),
    .A2(_16394_),
    .B(_16457_),
    .C(_16337_),
    .Y(_16458_));
 NAND2x1_ASAP7_75t_R _33901_ (.A(_15471_),
    .B(_01045_),
    .Y(_16459_));
 OA211x2_ASAP7_75t_R _33902_ (.A1(_16333_),
    .A2(_16397_),
    .B(_16459_),
    .C(_15593_),
    .Y(_16460_));
 OR3x1_ASAP7_75t_R _33903_ (.A(_15337_),
    .B(_16458_),
    .C(_16460_),
    .Y(_16461_));
 OA21x2_ASAP7_75t_R _33904_ (.A1(_15588_),
    .A2(_16456_),
    .B(_16461_),
    .Y(_16462_));
 NAND2x1_ASAP7_75t_R _33905_ (.A(_15325_),
    .B(_01042_),
    .Y(_16463_));
 OA211x2_ASAP7_75t_R _33906_ (.A1(_16369_),
    .A2(_16402_),
    .B(_16463_),
    .C(_16371_),
    .Y(_16464_));
 NAND2x1_ASAP7_75t_R _33907_ (.A(_15260_),
    .B(_01041_),
    .Y(_16465_));
 OA211x2_ASAP7_75t_R _33908_ (.A1(_16369_),
    .A2(_16405_),
    .B(_16465_),
    .C(_16354_),
    .Y(_16466_));
 OR3x1_ASAP7_75t_R _33909_ (.A(_15288_),
    .B(_16464_),
    .C(_16466_),
    .Y(_16467_));
 NAND2x1_ASAP7_75t_R _33910_ (.A(_15325_),
    .B(_01050_),
    .Y(_16468_));
 OA211x2_ASAP7_75t_R _33911_ (.A1(_16369_),
    .A2(_16409_),
    .B(_16468_),
    .C(_16371_),
    .Y(_16469_));
 NAND2x1_ASAP7_75t_R _33912_ (.A(_15260_),
    .B(_01049_),
    .Y(_16470_));
 OA211x2_ASAP7_75t_R _33913_ (.A1(_16369_),
    .A2(_16412_),
    .B(_16470_),
    .C(_16354_),
    .Y(_16471_));
 OR3x1_ASAP7_75t_R _33914_ (.A(_15337_),
    .B(_16469_),
    .C(_16471_),
    .Y(_16472_));
 AND3x1_ASAP7_75t_R _33915_ (.A(_16218_),
    .B(_16467_),
    .C(_16472_),
    .Y(_16473_));
 AO21x1_ASAP7_75t_R _33916_ (.A1(_15587_),
    .A2(_16462_),
    .B(_16473_),
    .Y(_16474_));
 NAND2x1_ASAP7_75t_R _33917_ (.A(_15589_),
    .B(_01058_),
    .Y(_16475_));
 OA211x2_ASAP7_75t_R _33918_ (.A1(_16373_),
    .A2(_16418_),
    .B(_16475_),
    .C(_16371_),
    .Y(_16476_));
 NAND2x1_ASAP7_75t_R _33919_ (.A(_15589_),
    .B(_01057_),
    .Y(_16477_));
 OA211x2_ASAP7_75t_R _33920_ (.A1(_16373_),
    .A2(_16421_),
    .B(_16477_),
    .C(_15295_),
    .Y(_16478_));
 OR3x1_ASAP7_75t_R _33921_ (.A(_16368_),
    .B(_16476_),
    .C(_16478_),
    .Y(_16479_));
 NAND2x1_ASAP7_75t_R _33922_ (.A(_15589_),
    .B(_01066_),
    .Y(_16480_));
 OA211x2_ASAP7_75t_R _33923_ (.A1(_16373_),
    .A2(_16425_),
    .B(_16480_),
    .C(_15600_),
    .Y(_16481_));
 NAND2x1_ASAP7_75t_R _33924_ (.A(_15589_),
    .B(_01065_),
    .Y(_16482_));
 OA211x2_ASAP7_75t_R _33925_ (.A1(_15484_),
    .A2(_16428_),
    .B(_16482_),
    .C(_15295_),
    .Y(_16483_));
 OR3x1_ASAP7_75t_R _33926_ (.A(_15596_),
    .B(_16481_),
    .C(_16483_),
    .Y(_16484_));
 AND3x1_ASAP7_75t_R _33927_ (.A(_16218_),
    .B(_16479_),
    .C(_16484_),
    .Y(_16485_));
 NOR2x1_ASAP7_75t_R _33928_ (.A(_15633_),
    .B(_01063_),
    .Y(_16486_));
 AO21x1_ASAP7_75t_R _33929_ (.A1(_16333_),
    .A2(_16433_),
    .B(_16486_),
    .Y(_16487_));
 NAND2x1_ASAP7_75t_R _33930_ (.A(_15343_),
    .B(_01062_),
    .Y(_16488_));
 OA211x2_ASAP7_75t_R _33931_ (.A1(_16373_),
    .A2(_16436_),
    .B(_16488_),
    .C(_16371_),
    .Y(_16489_));
 AO21x1_ASAP7_75t_R _33932_ (.A1(_15296_),
    .A2(_16487_),
    .B(_16489_),
    .Y(_16490_));
 NAND2x1_ASAP7_75t_R _33933_ (.A(_15291_),
    .B(_01054_),
    .Y(_16491_));
 OA211x2_ASAP7_75t_R _33934_ (.A1(_15598_),
    .A2(_16440_),
    .B(_16491_),
    .C(_15600_),
    .Y(_16492_));
 NAND2x1_ASAP7_75t_R _33935_ (.A(_15291_),
    .B(_01053_),
    .Y(_16493_));
 OA211x2_ASAP7_75t_R _33936_ (.A1(_15598_),
    .A2(_16443_),
    .B(_16493_),
    .C(_15338_),
    .Y(_16494_));
 OR3x1_ASAP7_75t_R _33937_ (.A(_16368_),
    .B(_16492_),
    .C(_16494_),
    .Y(_16495_));
 OA211x2_ASAP7_75t_R _33938_ (.A1(_15482_),
    .A2(_16490_),
    .B(_16495_),
    .C(_15587_),
    .Y(_16496_));
 OR3x1_ASAP7_75t_R _33939_ (.A(_15466_),
    .B(_16485_),
    .C(_16496_),
    .Y(_16497_));
 OA21x2_ASAP7_75t_R _33940_ (.A1(_15434_),
    .A2(_16474_),
    .B(_16497_),
    .Y(_16498_));
 INVx2_ASAP7_75t_R _33941_ (.A(_16498_),
    .Y(_16499_));
 OA211x2_ASAP7_75t_R _33942_ (.A1(_16332_),
    .A2(_16386_),
    .B(_16389_),
    .C(_15503_),
    .Y(_16500_));
 AOI21x1_ASAP7_75t_R _33943_ (.A1(_14090_),
    .A2(_16499_),
    .B(_16500_),
    .Y(_18659_));
 INVx1_ASAP7_75t_R _33944_ (.A(_18659_),
    .Y(_18657_));
 OR3x1_ASAP7_75t_R _33945_ (.A(net1940),
    .B(_16246_),
    .C(net1951),
    .Y(_16501_));
 OR3x2_ASAP7_75t_R _33946_ (.A(_16006_),
    .B(_15997_),
    .C(_16501_),
    .Y(_16502_));
 OR3x1_ASAP7_75t_R _33947_ (.A(_15167_),
    .B(_15510_),
    .C(_16502_),
    .Y(_16503_));
 OR3x1_ASAP7_75t_R _33948_ (.A(_15031_),
    .B(_15037_),
    .C(_16503_),
    .Y(_16504_));
 AO21x1_ASAP7_75t_R _33949_ (.A1(_15513_),
    .A2(_15514_),
    .B(_16502_),
    .Y(_16505_));
 NAND3x1_ASAP7_75t_R _33950_ (.A(_16244_),
    .B(_15999_),
    .C(_16251_),
    .Y(_16506_));
 AND3x1_ASAP7_75t_R _33951_ (.A(_16504_),
    .B(_16505_),
    .C(_16506_),
    .Y(_16507_));
 INVx3_ASAP7_75t_R _33952_ (.A(_01037_),
    .Y(_16508_));
 NOR2x1_ASAP7_75t_R _33953_ (.A(_16000_),
    .B(_16501_),
    .Y(_16509_));
 INVx1_ASAP7_75t_R _33954_ (.A(_01038_),
    .Y(_16510_));
 AO221x1_ASAP7_75t_R _33955_ (.A1(_16244_),
    .A2(_16247_),
    .B1(_16509_),
    .B2(_15507_),
    .C(_16510_),
    .Y(_16511_));
 INVx1_ASAP7_75t_R _33956_ (.A(_01070_),
    .Y(_16512_));
 AOI21x1_ASAP7_75t_R _33957_ (.A1(_16508_),
    .A2(_16511_),
    .B(_16512_),
    .Y(_16513_));
 OA21x2_ASAP7_75t_R _33958_ (.A1(_01037_),
    .A2(_16507_),
    .B(_16513_),
    .Y(_16514_));
 XNOR2x1_ASAP7_75t_R _33959_ (.B(_16514_),
    .Y(_16515_),
    .A(_01069_));
 INVx4_ASAP7_75t_R _33960_ (.A(_16515_),
    .Y(\alu_adder_result_ex[21] ));
 OA21x2_ASAP7_75t_R _33961_ (.A1(_15997_),
    .A2(_16011_),
    .B(_00942_),
    .Y(_16516_));
 OA21x2_ASAP7_75t_R _33962_ (.A1(net1940),
    .A2(_16516_),
    .B(_00974_),
    .Y(_16517_));
 OA21x2_ASAP7_75t_R _33963_ (.A1(_16246_),
    .A2(_16517_),
    .B(_01006_),
    .Y(_16518_));
 OA21x2_ASAP7_75t_R _33964_ (.A1(net1951),
    .A2(_16518_),
    .B(_01038_),
    .Y(_16519_));
 AND3x1_ASAP7_75t_R _33965_ (.A(_16508_),
    .B(_15522_),
    .C(_16519_),
    .Y(_16520_));
 OA21x2_ASAP7_75t_R _33966_ (.A1(_15169_),
    .A2(_15176_),
    .B(_16520_),
    .Y(_16521_));
 OA21x2_ASAP7_75t_R _33967_ (.A1(_15522_),
    .A2(net1954),
    .B(_16519_),
    .Y(_16522_));
 AO21x1_ASAP7_75t_R _33968_ (.A1(_15510_),
    .A2(_15522_),
    .B(net1954),
    .Y(_16523_));
 NAND3x1_ASAP7_75t_R _33969_ (.A(_16508_),
    .B(_16519_),
    .C(_16523_),
    .Y(_16524_));
 OAI21x1_ASAP7_75t_R _33970_ (.A1(_16508_),
    .A2(_16522_),
    .B(_16524_),
    .Y(_16525_));
 OR3x1_ASAP7_75t_R _33971_ (.A(_16508_),
    .B(_15510_),
    .C(net1954),
    .Y(_16526_));
 NOR3x1_ASAP7_75t_R _33972_ (.A(_15169_),
    .B(_15176_),
    .C(_16526_),
    .Y(_16527_));
 NOR3x2_ASAP7_75t_R _33973_ (.B(_16525_),
    .C(_16527_),
    .Y(_16528_),
    .A(_16521_));
 INVx6_ASAP7_75t_R _33974_ (.A(_16528_),
    .Y(\alu_adder_result_ex[20] ));
 AND2x2_ASAP7_75t_R _33975_ (.A(_13192_),
    .B(_01774_),
    .Y(_16529_));
 AO21x1_ASAP7_75t_R _33976_ (.A1(_14285_),
    .A2(_01072_),
    .B(_16529_),
    .Y(_16530_));
 OAI22x1_ASAP7_75t_R _33977_ (.A1(_01071_),
    .A2(_13101_),
    .B1(_16530_),
    .B2(_14710_),
    .Y(_16531_));
 INVx2_ASAP7_75t_R _33978_ (.A(_01080_),
    .Y(_16532_));
 NAND2x1_ASAP7_75t_R _33979_ (.A(_14755_),
    .B(_01078_),
    .Y(_16533_));
 OA211x2_ASAP7_75t_R _33980_ (.A1(_14292_),
    .A2(_16532_),
    .B(_16533_),
    .C(_13139_),
    .Y(_16534_));
 INVx2_ASAP7_75t_R _33981_ (.A(_01079_),
    .Y(_16535_));
 NAND2x1_ASAP7_75t_R _33982_ (.A(_14755_),
    .B(_01077_),
    .Y(_16536_));
 OA211x2_ASAP7_75t_R _33983_ (.A1(_14298_),
    .A2(_16535_),
    .B(_16536_),
    .C(_13173_),
    .Y(_16537_));
 OR3x1_ASAP7_75t_R _33984_ (.A(_13152_),
    .B(_16534_),
    .C(_16537_),
    .Y(_16538_));
 OA211x2_ASAP7_75t_R _33985_ (.A1(_13131_),
    .A2(_16531_),
    .B(_16538_),
    .C(_14428_),
    .Y(_16539_));
 INVx2_ASAP7_75t_R _33986_ (.A(_01076_),
    .Y(_16540_));
 NAND2x1_ASAP7_75t_R _33987_ (.A(_14760_),
    .B(_01074_),
    .Y(_16541_));
 OA211x2_ASAP7_75t_R _33988_ (.A1(_13110_),
    .A2(_16540_),
    .B(_16541_),
    .C(_14762_),
    .Y(_16542_));
 INVx1_ASAP7_75t_R _33989_ (.A(_01075_),
    .Y(_16543_));
 NAND2x1_ASAP7_75t_R _33990_ (.A(_14391_),
    .B(_01073_),
    .Y(_16544_));
 OA211x2_ASAP7_75t_R _33991_ (.A1(_15675_),
    .A2(_16543_),
    .B(_16544_),
    .C(_13088_),
    .Y(_16545_));
 OR3x1_ASAP7_75t_R _33992_ (.A(_14308_),
    .B(_16542_),
    .C(_16545_),
    .Y(_16546_));
 INVx2_ASAP7_75t_R _33993_ (.A(_01084_),
    .Y(_16547_));
 NAND2x1_ASAP7_75t_R _33994_ (.A(_14391_),
    .B(_01082_),
    .Y(_16548_));
 OA211x2_ASAP7_75t_R _33995_ (.A1(_13110_),
    .A2(_16547_),
    .B(_16548_),
    .C(_14362_),
    .Y(_16549_));
 INVx2_ASAP7_75t_R _33996_ (.A(_01083_),
    .Y(_16550_));
 NAND2x1_ASAP7_75t_R _33997_ (.A(_14460_),
    .B(_01081_),
    .Y(_16551_));
 OA211x2_ASAP7_75t_R _33998_ (.A1(_15675_),
    .A2(_16550_),
    .B(_16551_),
    .C(_13088_),
    .Y(_16552_));
 OR3x1_ASAP7_75t_R _33999_ (.A(_14326_),
    .B(_16549_),
    .C(_16552_),
    .Y(_16553_));
 AND3x1_ASAP7_75t_R _34000_ (.A(_14807_),
    .B(_16546_),
    .C(_16553_),
    .Y(_16554_));
 OR3x2_ASAP7_75t_R _34001_ (.A(_14447_),
    .B(_16539_),
    .C(_16554_),
    .Y(_16555_));
 INVx2_ASAP7_75t_R _34002_ (.A(_01092_),
    .Y(_16556_));
 NAND2x1_ASAP7_75t_R _34003_ (.A(_14760_),
    .B(_01090_),
    .Y(_16557_));
 OA211x2_ASAP7_75t_R _34004_ (.A1(_14310_),
    .A2(_16556_),
    .B(_16557_),
    .C(_14762_),
    .Y(_16558_));
 INVx2_ASAP7_75t_R _34005_ (.A(_01091_),
    .Y(_16559_));
 NAND2x1_ASAP7_75t_R _34006_ (.A(_14760_),
    .B(_01089_),
    .Y(_16560_));
 OA211x2_ASAP7_75t_R _34007_ (.A1(_13110_),
    .A2(_16559_),
    .B(_16560_),
    .C(_14765_),
    .Y(_16561_));
 OR3x1_ASAP7_75t_R _34008_ (.A(_14308_),
    .B(_16558_),
    .C(_16561_),
    .Y(_16562_));
 INVx2_ASAP7_75t_R _34009_ (.A(_01100_),
    .Y(_16563_));
 NAND2x1_ASAP7_75t_R _34010_ (.A(_14760_),
    .B(_01098_),
    .Y(_16564_));
 OA211x2_ASAP7_75t_R _34011_ (.A1(_14317_),
    .A2(_16563_),
    .B(_16564_),
    .C(_14762_),
    .Y(_16565_));
 INVx2_ASAP7_75t_R _34012_ (.A(_01099_),
    .Y(_16566_));
 NAND2x1_ASAP7_75t_R _34013_ (.A(_14391_),
    .B(_01097_),
    .Y(_16567_));
 OA211x2_ASAP7_75t_R _34014_ (.A1(_13110_),
    .A2(_16566_),
    .B(_16567_),
    .C(_14765_),
    .Y(_16568_));
 OR3x1_ASAP7_75t_R _34015_ (.A(_13185_),
    .B(_16565_),
    .C(_16568_),
    .Y(_16569_));
 AND3x1_ASAP7_75t_R _34016_ (.A(_14807_),
    .B(_16562_),
    .C(_16569_),
    .Y(_16570_));
 INVx2_ASAP7_75t_R _34017_ (.A(_01093_),
    .Y(_16571_));
 NOR2x1_ASAP7_75t_R _34018_ (.A(_13142_),
    .B(_01095_),
    .Y(_16572_));
 AO21x1_ASAP7_75t_R _34019_ (.A1(_14333_),
    .A2(_16571_),
    .B(_16572_),
    .Y(_16573_));
 INVx2_ASAP7_75t_R _34020_ (.A(_01096_),
    .Y(_16574_));
 NAND2x1_ASAP7_75t_R _34021_ (.A(_13096_),
    .B(_01094_),
    .Y(_16575_));
 OA211x2_ASAP7_75t_R _34022_ (.A1(_13189_),
    .A2(_16574_),
    .B(_16575_),
    .C(_14729_),
    .Y(_16576_));
 AO21x1_ASAP7_75t_R _34023_ (.A1(_13089_),
    .A2(_16573_),
    .B(_16576_),
    .Y(_16577_));
 INVx2_ASAP7_75t_R _34024_ (.A(_01088_),
    .Y(_16578_));
 NAND2x1_ASAP7_75t_R _34025_ (.A(_14755_),
    .B(_01086_),
    .Y(_16579_));
 OA211x2_ASAP7_75t_R _34026_ (.A1(_14298_),
    .A2(_16578_),
    .B(_16579_),
    .C(_13139_),
    .Y(_16580_));
 INVx2_ASAP7_75t_R _34027_ (.A(_01087_),
    .Y(_16581_));
 NAND2x1_ASAP7_75t_R _34028_ (.A(_13199_),
    .B(_01085_),
    .Y(_16582_));
 OA211x2_ASAP7_75t_R _34029_ (.A1(_14298_),
    .A2(_16581_),
    .B(_16582_),
    .C(_13173_),
    .Y(_16583_));
 OR3x1_ASAP7_75t_R _34030_ (.A(_13130_),
    .B(_16580_),
    .C(_16583_),
    .Y(_16584_));
 OA211x2_ASAP7_75t_R _34031_ (.A1(_14291_),
    .A2(_16577_),
    .B(_16584_),
    .C(_14428_),
    .Y(_16585_));
 OR3x2_ASAP7_75t_R _34032_ (.A(_14487_),
    .B(_16570_),
    .C(_16585_),
    .Y(_16586_));
 AND2x6_ASAP7_75t_R _34033_ (.A(_16555_),
    .B(_16586_),
    .Y(_16587_));
 AND2x2_ASAP7_75t_R _34034_ (.A(_01463_),
    .B(_14772_),
    .Y(_16588_));
 OAI22x1_ASAP7_75t_R _34035_ (.A1(_01493_),
    .A2(_15100_),
    .B1(_14384_),
    .B2(_16588_),
    .Y(_16589_));
 OA21x2_ASAP7_75t_R _34036_ (.A1(_13268_),
    .A2(_16587_),
    .B(_16589_),
    .Y(_16590_));
 BUFx6f_ASAP7_75t_R _34037_ (.A(_16590_),
    .Y(_18665_));
 INVx3_ASAP7_75t_R _34038_ (.A(_18665_),
    .Y(_18663_));
 BUFx6f_ASAP7_75t_R _34039_ (.A(_00122_),
    .Y(_16591_));
 OR3x1_ASAP7_75t_R _34040_ (.A(_16591_),
    .B(_14627_),
    .C(_14649_),
    .Y(_16592_));
 OAI21x1_ASAP7_75t_R _34041_ (.A1(_14646_),
    .A2(_18663_),
    .B(_16592_),
    .Y(_18052_));
 AND2x2_ASAP7_75t_R _34042_ (.A(_15291_),
    .B(_01774_),
    .Y(_16593_));
 AO21x1_ASAP7_75t_R _34043_ (.A1(_15290_),
    .A2(_01072_),
    .B(_16593_),
    .Y(_16594_));
 OAI22x1_ASAP7_75t_R _34044_ (.A1(_01071_),
    .A2(_15289_),
    .B1(_16594_),
    .B2(_15296_),
    .Y(_16595_));
 NAND2x1_ASAP7_75t_R _34045_ (.A(_15489_),
    .B(_01078_),
    .Y(_16596_));
 OA211x2_ASAP7_75t_R _34046_ (.A1(_15307_),
    .A2(_16532_),
    .B(_16596_),
    .C(_15304_),
    .Y(_16597_));
 NAND2x1_ASAP7_75t_R _34047_ (.A(_15597_),
    .B(_01077_),
    .Y(_16598_));
 OA211x2_ASAP7_75t_R _34048_ (.A1(_15437_),
    .A2(_16535_),
    .B(_16598_),
    .C(_15592_),
    .Y(_16599_));
 OR3x1_ASAP7_75t_R _34049_ (.A(_15336_),
    .B(_16597_),
    .C(_16599_),
    .Y(_16600_));
 OA211x2_ASAP7_75t_R _34050_ (.A1(_15288_),
    .A2(_16595_),
    .B(_16600_),
    .C(_15313_),
    .Y(_16601_));
 NAND2x1_ASAP7_75t_R _34051_ (.A(_15340_),
    .B(_01074_),
    .Y(_16602_));
 OA211x2_ASAP7_75t_R _34052_ (.A1(_15343_),
    .A2(_16540_),
    .B(_16602_),
    .C(_15620_),
    .Y(_16603_));
 NAND2x1_ASAP7_75t_R _34053_ (.A(_15734_),
    .B(_01073_),
    .Y(_16604_));
 OA211x2_ASAP7_75t_R _34054_ (.A1(_15343_),
    .A2(_16543_),
    .B(_16604_),
    .C(_15497_),
    .Y(_16605_));
 OR3x1_ASAP7_75t_R _34055_ (.A(_15255_),
    .B(_16603_),
    .C(_16605_),
    .Y(_16606_));
 NAND2x1_ASAP7_75t_R _34056_ (.A(_15340_),
    .B(_01082_),
    .Y(_16607_));
 OA211x2_ASAP7_75t_R _34057_ (.A1(_15343_),
    .A2(_16547_),
    .B(_16607_),
    .C(_15620_),
    .Y(_16608_));
 NAND2x1_ASAP7_75t_R _34058_ (.A(_15734_),
    .B(_01081_),
    .Y(_16609_));
 OA211x2_ASAP7_75t_R _34059_ (.A1(_15343_),
    .A2(_16550_),
    .B(_16609_),
    .C(_15497_),
    .Y(_16610_));
 OR3x1_ASAP7_75t_R _34060_ (.A(_15298_),
    .B(_16608_),
    .C(_16610_),
    .Y(_16611_));
 AND3x1_ASAP7_75t_R _34061_ (.A(_15253_),
    .B(_16606_),
    .C(_16611_),
    .Y(_16612_));
 OR3x2_ASAP7_75t_R _34062_ (.A(_15251_),
    .B(_16601_),
    .C(_16612_),
    .Y(_16613_));
 NAND2x1_ASAP7_75t_R _34063_ (.A(_16109_),
    .B(_01090_),
    .Y(_16614_));
 OA211x2_ASAP7_75t_R _34064_ (.A1(_15260_),
    .A2(_16556_),
    .B(_16614_),
    .C(_15267_),
    .Y(_16615_));
 NAND2x1_ASAP7_75t_R _34065_ (.A(_15618_),
    .B(_01089_),
    .Y(_16616_));
 OA211x2_ASAP7_75t_R _34066_ (.A1(_15269_),
    .A2(_16559_),
    .B(_16616_),
    .C(_15283_),
    .Y(_16617_));
 OR3x1_ASAP7_75t_R _34067_ (.A(_15255_),
    .B(_16615_),
    .C(_16617_),
    .Y(_16618_));
 NAND2x1_ASAP7_75t_R _34068_ (.A(_16109_),
    .B(_01098_),
    .Y(_16619_));
 OA211x2_ASAP7_75t_R _34069_ (.A1(_15269_),
    .A2(_16563_),
    .B(_16619_),
    .C(_15267_),
    .Y(_16620_));
 NAND2x1_ASAP7_75t_R _34070_ (.A(_15618_),
    .B(_01097_),
    .Y(_16621_));
 OA211x2_ASAP7_75t_R _34071_ (.A1(_15269_),
    .A2(_16566_),
    .B(_16621_),
    .C(_15283_),
    .Y(_16622_));
 OR3x1_ASAP7_75t_R _34072_ (.A(_15279_),
    .B(_16620_),
    .C(_16622_),
    .Y(_16623_));
 AND3x1_ASAP7_75t_R _34073_ (.A(_15253_),
    .B(_16618_),
    .C(_16623_),
    .Y(_16624_));
 NOR2x1_ASAP7_75t_R _34074_ (.A(_15445_),
    .B(_01095_),
    .Y(_16625_));
 AO21x1_ASAP7_75t_R _34075_ (.A1(_15633_),
    .A2(_16571_),
    .B(_16625_),
    .Y(_16626_));
 NAND2x1_ASAP7_75t_R _34076_ (.A(_15454_),
    .B(_01094_),
    .Y(_16627_));
 OA211x2_ASAP7_75t_R _34077_ (.A1(_15320_),
    .A2(_16574_),
    .B(_16627_),
    .C(_15323_),
    .Y(_16628_));
 AO21x1_ASAP7_75t_R _34078_ (.A1(_15339_),
    .A2(_16626_),
    .B(_16628_),
    .Y(_16629_));
 NAND2x1_ASAP7_75t_R _34079_ (.A(_15489_),
    .B(_01086_),
    .Y(_16630_));
 OA211x2_ASAP7_75t_R _34080_ (.A1(_15300_),
    .A2(_16578_),
    .B(_16630_),
    .C(_15304_),
    .Y(_16631_));
 NAND2x1_ASAP7_75t_R _34081_ (.A(_15489_),
    .B(_01085_),
    .Y(_16632_));
 OA211x2_ASAP7_75t_R _34082_ (.A1(_15307_),
    .A2(_16581_),
    .B(_16632_),
    .C(_15309_),
    .Y(_16633_));
 OR3x1_ASAP7_75t_R _34083_ (.A(_15352_),
    .B(_16631_),
    .C(_16633_),
    .Y(_16634_));
 OA211x2_ASAP7_75t_R _34084_ (.A1(_15337_),
    .A2(_16629_),
    .B(_16634_),
    .C(_15313_),
    .Y(_16635_));
 OR3x2_ASAP7_75t_R _34085_ (.A(_15316_),
    .B(_16624_),
    .C(_16635_),
    .Y(_16636_));
 NAND2x2_ASAP7_75t_R _34086_ (.A(_16613_),
    .B(_16636_),
    .Y(_16637_));
 OA211x2_ASAP7_75t_R _34087_ (.A1(_15587_),
    .A2(_16386_),
    .B(_16389_),
    .C(_15503_),
    .Y(_16638_));
 AOI21x1_ASAP7_75t_R _34088_ (.A1(_15250_),
    .A2(_16637_),
    .B(_16638_),
    .Y(_18664_));
 INVx1_ASAP7_75t_R _34089_ (.A(_18664_),
    .Y(_18662_));
 AND2x2_ASAP7_75t_R _34090_ (.A(_13206_),
    .B(_01773_),
    .Y(_16639_));
 AO21x1_ASAP7_75t_R _34091_ (.A1(_14286_),
    .A2(_01104_),
    .B(_16639_),
    .Y(_16640_));
 OAI22x1_ASAP7_75t_R _34092_ (.A1(_01103_),
    .A2(_14284_),
    .B1(_16640_),
    .B2(_14289_),
    .Y(_16641_));
 INVx2_ASAP7_75t_R _34093_ (.A(_01112_),
    .Y(_16642_));
 NAND2x1_ASAP7_75t_R _34094_ (.A(_14450_),
    .B(_01110_),
    .Y(_16643_));
 OA211x2_ASAP7_75t_R _34095_ (.A1(_14985_),
    .A2(_16642_),
    .B(_16643_),
    .C(_14923_),
    .Y(_16644_));
 INVx2_ASAP7_75t_R _34096_ (.A(_01111_),
    .Y(_16645_));
 NAND2x1_ASAP7_75t_R _34097_ (.A(_14815_),
    .B(_01109_),
    .Y(_16646_));
 OA211x2_ASAP7_75t_R _34098_ (.A1(_14943_),
    .A2(_16645_),
    .B(_16646_),
    .C(_14372_),
    .Y(_16647_));
 OR3x1_ASAP7_75t_R _34099_ (.A(_14929_),
    .B(_16644_),
    .C(_16647_),
    .Y(_16648_));
 OA211x2_ASAP7_75t_R _34100_ (.A1(_14283_),
    .A2(_16641_),
    .B(_16648_),
    .C(_14852_),
    .Y(_16649_));
 INVx2_ASAP7_75t_R _34101_ (.A(_01108_),
    .Y(_16650_));
 NAND2x1_ASAP7_75t_R _34102_ (.A(_14888_),
    .B(_01106_),
    .Y(_16651_));
 OA211x2_ASAP7_75t_R _34103_ (.A1(_14886_),
    .A2(_16650_),
    .B(_16651_),
    .C(_14652_),
    .Y(_16652_));
 INVx2_ASAP7_75t_R _34104_ (.A(_01107_),
    .Y(_16653_));
 NAND2x1_ASAP7_75t_R _34105_ (.A(_14782_),
    .B(_01105_),
    .Y(_16654_));
 OA211x2_ASAP7_75t_R _34106_ (.A1(_14711_),
    .A2(_16653_),
    .B(_16654_),
    .C(_15122_),
    .Y(_16655_));
 OR3x1_ASAP7_75t_R _34107_ (.A(_15117_),
    .B(_16652_),
    .C(_16655_),
    .Y(_16656_));
 INVx2_ASAP7_75t_R _34108_ (.A(_01116_),
    .Y(_16657_));
 NAND2x1_ASAP7_75t_R _34109_ (.A(_14782_),
    .B(_01114_),
    .Y(_16658_));
 OA211x2_ASAP7_75t_R _34110_ (.A1(_14886_),
    .A2(_16657_),
    .B(_16658_),
    .C(_14652_),
    .Y(_16659_));
 INVx2_ASAP7_75t_R _34111_ (.A(_01115_),
    .Y(_16660_));
 NAND2x1_ASAP7_75t_R _34112_ (.A(_15061_),
    .B(_01113_),
    .Y(_16661_));
 OA211x2_ASAP7_75t_R _34113_ (.A1(_15120_),
    .A2(_16660_),
    .B(_16661_),
    .C(_15122_),
    .Y(_16662_));
 OR3x1_ASAP7_75t_R _34114_ (.A(_14877_),
    .B(_16659_),
    .C(_16662_),
    .Y(_16663_));
 AND3x4_ASAP7_75t_R _34115_ (.A(_14340_),
    .B(_16656_),
    .C(_16663_),
    .Y(_16664_));
 OR3x1_ASAP7_75t_R _34116_ (.A(_14281_),
    .B(_16649_),
    .C(_16664_),
    .Y(_16665_));
 INVx2_ASAP7_75t_R _34117_ (.A(_01124_),
    .Y(_16666_));
 NAND2x1_ASAP7_75t_R _34118_ (.A(_14888_),
    .B(_01122_),
    .Y(_16667_));
 OA211x2_ASAP7_75t_R _34119_ (.A1(_14886_),
    .A2(_16666_),
    .B(_16667_),
    .C(_14652_),
    .Y(_16668_));
 INVx2_ASAP7_75t_R _34120_ (.A(_01123_),
    .Y(_16669_));
 NAND2x1_ASAP7_75t_R _34121_ (.A(_14782_),
    .B(_01121_),
    .Y(_16670_));
 OA211x2_ASAP7_75t_R _34122_ (.A1(_14711_),
    .A2(_16669_),
    .B(_16670_),
    .C(_15122_),
    .Y(_16671_));
 OR3x1_ASAP7_75t_R _34123_ (.A(_15117_),
    .B(_16668_),
    .C(_16671_),
    .Y(_16672_));
 INVx2_ASAP7_75t_R _34124_ (.A(_01132_),
    .Y(_16673_));
 NAND2x1_ASAP7_75t_R _34125_ (.A(_14782_),
    .B(_01130_),
    .Y(_16674_));
 OA211x2_ASAP7_75t_R _34126_ (.A1(_14711_),
    .A2(_16673_),
    .B(_16674_),
    .C(_14652_),
    .Y(_16675_));
 INVx2_ASAP7_75t_R _34127_ (.A(_01131_),
    .Y(_16676_));
 NAND2x1_ASAP7_75t_R _34128_ (.A(_15061_),
    .B(_01129_),
    .Y(_16677_));
 OA211x2_ASAP7_75t_R _34129_ (.A1(_15120_),
    .A2(_16676_),
    .B(_16677_),
    .C(_15122_),
    .Y(_16678_));
 OR3x1_ASAP7_75t_R _34130_ (.A(_14877_),
    .B(_16675_),
    .C(_16678_),
    .Y(_16679_));
 AND3x1_ASAP7_75t_R _34131_ (.A(_14340_),
    .B(_16672_),
    .C(_16679_),
    .Y(_16680_));
 INVx2_ASAP7_75t_R _34132_ (.A(_01125_),
    .Y(_16681_));
 NOR2x1_ASAP7_75t_R _34133_ (.A(_14366_),
    .B(_01127_),
    .Y(_16682_));
 AO21x1_ASAP7_75t_R _34134_ (.A1(_14278_),
    .A2(_16681_),
    .B(_16682_),
    .Y(_16683_));
 INVx2_ASAP7_75t_R _34135_ (.A(_01128_),
    .Y(_16684_));
 NAND2x1_ASAP7_75t_R _34136_ (.A(_14333_),
    .B(_01126_),
    .Y(_16685_));
 OA211x2_ASAP7_75t_R _34137_ (.A1(_14331_),
    .A2(_16684_),
    .B(_16685_),
    .C(_14329_),
    .Y(_16686_));
 AO21x1_ASAP7_75t_R _34138_ (.A1(_14975_),
    .A2(_16683_),
    .B(_16686_),
    .Y(_16687_));
 INVx2_ASAP7_75t_R _34139_ (.A(_01120_),
    .Y(_16688_));
 NAND2x1_ASAP7_75t_R _34140_ (.A(_13189_),
    .B(_01118_),
    .Y(_16689_));
 OA211x2_ASAP7_75t_R _34141_ (.A1(_14496_),
    .A2(_16688_),
    .B(_16689_),
    .C(_14504_),
    .Y(_16690_));
 INVx2_ASAP7_75t_R _34142_ (.A(_01119_),
    .Y(_16691_));
 NAND2x1_ASAP7_75t_R _34143_ (.A(_14517_),
    .B(_01117_),
    .Y(_16692_));
 OA211x2_ASAP7_75t_R _34144_ (.A1(_14516_),
    .A2(_16691_),
    .B(_16692_),
    .C(_14509_),
    .Y(_16693_));
 OR3x1_ASAP7_75t_R _34145_ (.A(_14469_),
    .B(_16690_),
    .C(_16693_),
    .Y(_16694_));
 OA211x2_ASAP7_75t_R _34146_ (.A1(_14354_),
    .A2(_16687_),
    .B(_16694_),
    .C(_14852_),
    .Y(_16695_));
 OR3x2_ASAP7_75t_R _34147_ (.A(_13164_),
    .B(_16680_),
    .C(_16695_),
    .Y(_16696_));
 AO21x2_ASAP7_75t_R _34148_ (.A1(_16665_),
    .A2(_16696_),
    .B(_14377_),
    .Y(_16697_));
 BUFx6f_ASAP7_75t_R _34149_ (.A(_01492_),
    .Y(_16698_));
 AND2x2_ASAP7_75t_R _34150_ (.A(_01462_),
    .B(_14381_),
    .Y(_16699_));
 OAI22x1_ASAP7_75t_R _34151_ (.A1(_16698_),
    .A2(_14382_),
    .B1(_14385_),
    .B2(_16699_),
    .Y(_16700_));
 NAND2x2_ASAP7_75t_R _34152_ (.A(_16697_),
    .B(_16700_),
    .Y(_18668_));
 INVx1_ASAP7_75t_R _34153_ (.A(_18668_),
    .Y(_18670_));
 BUFx6f_ASAP7_75t_R _34154_ (.A(_00129_),
    .Y(_16701_));
 OR3x1_ASAP7_75t_R _34155_ (.A(_16701_),
    .B(_14627_),
    .C(_14649_),
    .Y(_16702_));
 OAI21x1_ASAP7_75t_R _34156_ (.A1(_14646_),
    .A2(_18668_),
    .B(_16702_),
    .Y(_18054_));
 AND2x2_ASAP7_75t_R _34157_ (.A(_15291_),
    .B(_01773_),
    .Y(_16703_));
 AO21x1_ASAP7_75t_R _34158_ (.A1(_15290_),
    .A2(_01104_),
    .B(_16703_),
    .Y(_16704_));
 OAI22x1_ASAP7_75t_R _34159_ (.A1(_01103_),
    .A2(_15435_),
    .B1(_16704_),
    .B2(_15296_),
    .Y(_16705_));
 NAND2x1_ASAP7_75t_R _34160_ (.A(_15632_),
    .B(_01110_),
    .Y(_16706_));
 OA211x2_ASAP7_75t_R _34161_ (.A1(_15353_),
    .A2(_16642_),
    .B(_16706_),
    .C(_15304_),
    .Y(_16707_));
 NAND2x1_ASAP7_75t_R _34162_ (.A(_15632_),
    .B(_01109_),
    .Y(_16708_));
 OA211x2_ASAP7_75t_R _34163_ (.A1(_15353_),
    .A2(_16645_),
    .B(_16708_),
    .C(_15309_),
    .Y(_16709_));
 OR3x1_ASAP7_75t_R _34164_ (.A(_15298_),
    .B(_16707_),
    .C(_16709_),
    .Y(_16710_));
 OA211x2_ASAP7_75t_R _34165_ (.A1(_15288_),
    .A2(_16705_),
    .B(_16710_),
    .C(_15313_),
    .Y(_16711_));
 NAND2x1_ASAP7_75t_R _34166_ (.A(_16106_),
    .B(_01106_),
    .Y(_16712_));
 OA211x2_ASAP7_75t_R _34167_ (.A1(_15325_),
    .A2(_16650_),
    .B(_16712_),
    .C(_15267_),
    .Y(_16713_));
 NAND2x1_ASAP7_75t_R _34168_ (.A(_16109_),
    .B(_01105_),
    .Y(_16714_));
 OA211x2_ASAP7_75t_R _34169_ (.A1(_15260_),
    .A2(_16653_),
    .B(_16714_),
    .C(_15275_),
    .Y(_16715_));
 OR3x1_ASAP7_75t_R _34170_ (.A(_15255_),
    .B(_16713_),
    .C(_16715_),
    .Y(_16716_));
 NAND2x1_ASAP7_75t_R _34171_ (.A(_16106_),
    .B(_01114_),
    .Y(_16717_));
 OA211x2_ASAP7_75t_R _34172_ (.A1(_15260_),
    .A2(_16657_),
    .B(_16717_),
    .C(_15267_),
    .Y(_16718_));
 NAND2x1_ASAP7_75t_R _34173_ (.A(_16109_),
    .B(_01113_),
    .Y(_16719_));
 OA211x2_ASAP7_75t_R _34174_ (.A1(_15260_),
    .A2(_16660_),
    .B(_16719_),
    .C(_15283_),
    .Y(_16720_));
 OR3x1_ASAP7_75t_R _34175_ (.A(_15279_),
    .B(_16718_),
    .C(_16720_),
    .Y(_16721_));
 AND3x4_ASAP7_75t_R _34176_ (.A(_15253_),
    .B(_16716_),
    .C(_16721_),
    .Y(_16722_));
 OR3x2_ASAP7_75t_R _34177_ (.A(_15251_),
    .B(_16711_),
    .C(_16722_),
    .Y(_16723_));
 NAND2x1_ASAP7_75t_R _34178_ (.A(_15270_),
    .B(_01122_),
    .Y(_16724_));
 OA211x2_ASAP7_75t_R _34179_ (.A1(_15346_),
    .A2(_16666_),
    .B(_16724_),
    .C(_15349_),
    .Y(_16725_));
 NAND2x1_ASAP7_75t_R _34180_ (.A(_15451_),
    .B(_01121_),
    .Y(_16726_));
 OA211x2_ASAP7_75t_R _34181_ (.A1(_15450_),
    .A2(_16669_),
    .B(_16726_),
    .C(_15456_),
    .Y(_16727_));
 OR3x1_ASAP7_75t_R _34182_ (.A(_15318_),
    .B(_16725_),
    .C(_16727_),
    .Y(_16728_));
 NAND2x1_ASAP7_75t_R _34183_ (.A(_15451_),
    .B(_01130_),
    .Y(_16729_));
 OA211x2_ASAP7_75t_R _34184_ (.A1(_15346_),
    .A2(_16673_),
    .B(_16729_),
    .C(_15323_),
    .Y(_16730_));
 NAND2x1_ASAP7_75t_R _34185_ (.A(_15454_),
    .B(_01129_),
    .Y(_16731_));
 OA211x2_ASAP7_75t_R _34186_ (.A1(_15450_),
    .A2(_16676_),
    .B(_16731_),
    .C(_15456_),
    .Y(_16732_));
 OR3x1_ASAP7_75t_R _34187_ (.A(_15475_),
    .B(_16730_),
    .C(_16732_),
    .Y(_16733_));
 AND3x1_ASAP7_75t_R _34188_ (.A(_15317_),
    .B(_16728_),
    .C(_16733_),
    .Y(_16734_));
 NOR2x1_ASAP7_75t_R _34189_ (.A(_15589_),
    .B(_01127_),
    .Y(_16735_));
 AO21x1_ASAP7_75t_R _34190_ (.A1(_15484_),
    .A2(_16681_),
    .B(_16735_),
    .Y(_16736_));
 NAND2x1_ASAP7_75t_R _34191_ (.A(_15321_),
    .B(_01126_),
    .Y(_16737_));
 OA211x2_ASAP7_75t_R _34192_ (.A1(_15467_),
    .A2(_16684_),
    .B(_16737_),
    .C(_15469_),
    .Y(_16738_));
 AO21x1_ASAP7_75t_R _34193_ (.A1(_15339_),
    .A2(_16736_),
    .B(_16738_),
    .Y(_16739_));
 NAND2x1_ASAP7_75t_R _34194_ (.A(_15632_),
    .B(_01118_),
    .Y(_16740_));
 OA211x2_ASAP7_75t_R _34195_ (.A1(_15445_),
    .A2(_16688_),
    .B(_16740_),
    .C(_15443_),
    .Y(_16741_));
 NAND2x1_ASAP7_75t_R _34196_ (.A(_15632_),
    .B(_01117_),
    .Y(_16742_));
 OA211x2_ASAP7_75t_R _34197_ (.A1(_15445_),
    .A2(_16691_),
    .B(_16742_),
    .C(_15309_),
    .Y(_16743_));
 OR3x1_ASAP7_75t_R _34198_ (.A(_15352_),
    .B(_16741_),
    .C(_16743_),
    .Y(_16744_));
 OA211x2_ASAP7_75t_R _34199_ (.A1(_15482_),
    .A2(_16739_),
    .B(_16744_),
    .C(_15360_),
    .Y(_16745_));
 OR3x2_ASAP7_75t_R _34200_ (.A(_15466_),
    .B(_16734_),
    .C(_16745_),
    .Y(_16746_));
 NAND2x2_ASAP7_75t_R _34201_ (.A(_16723_),
    .B(_16746_),
    .Y(_16747_));
 OA211x2_ASAP7_75t_R _34202_ (.A1(_15482_),
    .A2(_16386_),
    .B(_16389_),
    .C(_15370_),
    .Y(_16748_));
 AOI21x1_ASAP7_75t_R _34203_ (.A1(_15250_),
    .A2(_16747_),
    .B(_16748_),
    .Y(_18669_));
 INVx1_ASAP7_75t_R _34204_ (.A(_18669_),
    .Y(_18667_));
 AO21x1_ASAP7_75t_R _34205_ (.A1(_01037_),
    .A2(_01070_),
    .B(_01069_),
    .Y(_16749_));
 AND2x2_ASAP7_75t_R _34206_ (.A(_01102_),
    .B(_16513_),
    .Y(_16750_));
 AO221x1_ASAP7_75t_R _34207_ (.A1(_01102_),
    .A2(_16749_),
    .B1(_16750_),
    .B2(_16507_),
    .C(_01101_),
    .Y(_16751_));
 AND2x2_ASAP7_75t_R _34208_ (.A(_01134_),
    .B(_16751_),
    .Y(_16752_));
 XNOR2x1_ASAP7_75t_R _34209_ (.B(_16752_),
    .Y(_16753_),
    .A(_01133_));
 INVx4_ASAP7_75t_R _34210_ (.A(_16753_),
    .Y(\alu_adder_result_ex[23] ));
 NOR2x1_ASAP7_75t_R _34211_ (.A(_15510_),
    .B(net1954),
    .Y(_16754_));
 INVx1_ASAP7_75t_R _34212_ (.A(_16754_),
    .Y(_16755_));
 OA31x2_ASAP7_75t_R _34213_ (.A1(_15169_),
    .A2(_15176_),
    .A3(_16755_),
    .B1(_16522_),
    .Y(_16756_));
 OR2x2_ASAP7_75t_R _34214_ (.A(_01037_),
    .B(_01069_),
    .Y(_16757_));
 BUFx6f_ASAP7_75t_R _34215_ (.A(_16757_),
    .Y(_16758_));
 OA21x2_ASAP7_75t_R _34216_ (.A1(_01070_),
    .A2(_01069_),
    .B(_01102_),
    .Y(_16759_));
 OA21x2_ASAP7_75t_R _34217_ (.A1(_16756_),
    .A2(_16758_),
    .B(_16759_),
    .Y(_16760_));
 XNOR2x1_ASAP7_75t_R _34218_ (.B(_16760_),
    .Y(_16761_),
    .A(_01101_));
 INVx4_ASAP7_75t_R _34219_ (.A(_16761_),
    .Y(\alu_adder_result_ex[22] ));
 AND2x2_ASAP7_75t_R _34220_ (.A(_14756_),
    .B(_01772_),
    .Y(_16762_));
 AO21x1_ASAP7_75t_R _34221_ (.A1(_13092_),
    .A2(_01136_),
    .B(_16762_),
    .Y(_16763_));
 OAI22x1_ASAP7_75t_R _34222_ (.A1(_01135_),
    .A2(_13102_),
    .B1(_16763_),
    .B2(_14975_),
    .Y(_16764_));
 INVx2_ASAP7_75t_R _34223_ (.A(_01144_),
    .Y(_16765_));
 NAND2x1_ASAP7_75t_R _34224_ (.A(_13196_),
    .B(_01142_),
    .Y(_16766_));
 OA211x2_ASAP7_75t_R _34225_ (.A1(_13097_),
    .A2(_16765_),
    .B(_16766_),
    .C(_14914_),
    .Y(_16767_));
 INVx2_ASAP7_75t_R _34226_ (.A(_01143_),
    .Y(_16768_));
 NAND2x1_ASAP7_75t_R _34227_ (.A(_13165_),
    .B(_01141_),
    .Y(_16769_));
 OA211x2_ASAP7_75t_R _34228_ (.A1(_14360_),
    .A2(_16768_),
    .B(_16769_),
    .C(_14463_),
    .Y(_16770_));
 OR3x1_ASAP7_75t_R _34229_ (.A(_13105_),
    .B(_16767_),
    .C(_16770_),
    .Y(_16771_));
 OA211x2_ASAP7_75t_R _34230_ (.A1(_13086_),
    .A2(_16764_),
    .B(_16771_),
    .C(_13125_),
    .Y(_16772_));
 INVx2_ASAP7_75t_R _34231_ (.A(_01140_),
    .Y(_16773_));
 NAND2x1_ASAP7_75t_R _34232_ (.A(_14808_),
    .B(_01138_),
    .Y(_16774_));
 OA211x2_ASAP7_75t_R _34233_ (.A1(_14921_),
    .A2(_16773_),
    .B(_16774_),
    .C(_14494_),
    .Y(_16775_));
 INVx2_ASAP7_75t_R _34234_ (.A(_01139_),
    .Y(_16776_));
 NAND2x1_ASAP7_75t_R _34235_ (.A(_14502_),
    .B(_01137_),
    .Y(_16777_));
 OA211x2_ASAP7_75t_R _34236_ (.A1(_14501_),
    .A2(_16776_),
    .B(_16777_),
    .C(_14926_),
    .Y(_16778_));
 OR3x1_ASAP7_75t_R _34237_ (.A(_14489_),
    .B(_16775_),
    .C(_16778_),
    .Y(_16779_));
 INVx2_ASAP7_75t_R _34238_ (.A(_01148_),
    .Y(_16780_));
 NAND2x1_ASAP7_75t_R _34239_ (.A(_14815_),
    .B(_01146_),
    .Y(_16781_));
 OA211x2_ASAP7_75t_R _34240_ (.A1(_14943_),
    .A2(_16780_),
    .B(_16781_),
    .C(_14494_),
    .Y(_16782_));
 INVx2_ASAP7_75t_R _34241_ (.A(_01147_),
    .Y(_16783_));
 NAND2x1_ASAP7_75t_R _34242_ (.A(_14502_),
    .B(_01145_),
    .Y(_16784_));
 OA211x2_ASAP7_75t_R _34243_ (.A1(_14496_),
    .A2(_16783_),
    .B(_16784_),
    .C(_14498_),
    .Y(_16785_));
 OR3x1_ASAP7_75t_R _34244_ (.A(_14929_),
    .B(_16782_),
    .C(_16785_),
    .Y(_16786_));
 AND3x1_ASAP7_75t_R _34245_ (.A(_14488_),
    .B(_16779_),
    .C(_16786_),
    .Y(_16787_));
 OR3x2_ASAP7_75t_R _34246_ (.A(_13082_),
    .B(_16772_),
    .C(_16787_),
    .Y(_16788_));
 INVx2_ASAP7_75t_R _34247_ (.A(_01156_),
    .Y(_16789_));
 NAND2x1_ASAP7_75t_R _34248_ (.A(_14752_),
    .B(_01154_),
    .Y(_16790_));
 OA211x2_ASAP7_75t_R _34249_ (.A1(_14985_),
    .A2(_16789_),
    .B(_16790_),
    .C(_14923_),
    .Y(_16791_));
 INVx2_ASAP7_75t_R _34250_ (.A(_01155_),
    .Y(_16792_));
 NAND2x1_ASAP7_75t_R _34251_ (.A(_14815_),
    .B(_01153_),
    .Y(_16793_));
 OA211x2_ASAP7_75t_R _34252_ (.A1(_14491_),
    .A2(_16792_),
    .B(_16793_),
    .C(_14926_),
    .Y(_16794_));
 OR3x1_ASAP7_75t_R _34253_ (.A(_14489_),
    .B(_16791_),
    .C(_16794_),
    .Y(_16795_));
 INVx2_ASAP7_75t_R _34254_ (.A(_01164_),
    .Y(_16796_));
 NAND2x1_ASAP7_75t_R _34255_ (.A(_14808_),
    .B(_01162_),
    .Y(_16797_));
 OA211x2_ASAP7_75t_R _34256_ (.A1(_14921_),
    .A2(_16796_),
    .B(_16797_),
    .C(_14923_),
    .Y(_16798_));
 INVx2_ASAP7_75t_R _34257_ (.A(_01163_),
    .Y(_16799_));
 NAND2x1_ASAP7_75t_R _34258_ (.A(_14492_),
    .B(_01161_),
    .Y(_16800_));
 OA211x2_ASAP7_75t_R _34259_ (.A1(_14501_),
    .A2(_16799_),
    .B(_16800_),
    .C(_14926_),
    .Y(_16801_));
 OR3x1_ASAP7_75t_R _34260_ (.A(_14929_),
    .B(_16798_),
    .C(_16801_),
    .Y(_16802_));
 AND3x1_ASAP7_75t_R _34261_ (.A(_14488_),
    .B(_16795_),
    .C(_16802_),
    .Y(_16803_));
 INVx2_ASAP7_75t_R _34262_ (.A(_01157_),
    .Y(_16804_));
 NOR2x1_ASAP7_75t_R _34263_ (.A(_14717_),
    .B(_01159_),
    .Y(_16805_));
 AO21x1_ASAP7_75t_R _34264_ (.A1(_14358_),
    .A2(_16804_),
    .B(_16805_),
    .Y(_16806_));
 INVx2_ASAP7_75t_R _34265_ (.A(_01160_),
    .Y(_16807_));
 NAND2x1_ASAP7_75t_R _34266_ (.A(_14367_),
    .B(_01158_),
    .Y(_16808_));
 OA211x2_ASAP7_75t_R _34267_ (.A1(_14366_),
    .A2(_16807_),
    .B(_16808_),
    .C(_14369_),
    .Y(_16809_));
 AO21x1_ASAP7_75t_R _34268_ (.A1(_13187_),
    .A2(_16806_),
    .B(_16809_),
    .Y(_16810_));
 INVx2_ASAP7_75t_R _34269_ (.A(_01152_),
    .Y(_16811_));
 NAND2x1_ASAP7_75t_R _34270_ (.A(_14697_),
    .B(_01150_),
    .Y(_16812_));
 OA211x2_ASAP7_75t_R _34271_ (.A1(_14360_),
    .A2(_16811_),
    .B(_16812_),
    .C(_14914_),
    .Y(_16813_));
 INVx2_ASAP7_75t_R _34272_ (.A(_01151_),
    .Y(_16814_));
 NAND2x1_ASAP7_75t_R _34273_ (.A(_14697_),
    .B(_01149_),
    .Y(_16815_));
 OA211x2_ASAP7_75t_R _34274_ (.A1(_14455_),
    .A2(_16814_),
    .B(_16815_),
    .C(_14463_),
    .Y(_16816_));
 OR3x1_ASAP7_75t_R _34275_ (.A(_13085_),
    .B(_16813_),
    .C(_16816_),
    .Y(_16817_));
 OA211x2_ASAP7_75t_R _34276_ (.A1(_13186_),
    .A2(_16810_),
    .B(_16817_),
    .C(_14466_),
    .Y(_16818_));
 OR3x2_ASAP7_75t_R _34277_ (.A(_14487_),
    .B(_16803_),
    .C(_16818_),
    .Y(_16819_));
 AO21x2_ASAP7_75t_R _34278_ (.A1(_16788_),
    .A2(_16819_),
    .B(_13267_),
    .Y(_16820_));
 AND2x2_ASAP7_75t_R _34279_ (.A(_01461_),
    .B(_14772_),
    .Y(_16821_));
 OAI22x1_ASAP7_75t_R _34280_ (.A1(_01491_),
    .A2(_14967_),
    .B1(_14968_),
    .B2(_16821_),
    .Y(_16822_));
 NAND2x2_ASAP7_75t_R _34281_ (.A(_16820_),
    .B(_16822_),
    .Y(_18673_));
 INVx1_ASAP7_75t_R _34282_ (.A(_18673_),
    .Y(_18675_));
 BUFx6f_ASAP7_75t_R _34283_ (.A(_00136_),
    .Y(_16823_));
 INVx1_ASAP7_75t_R _34284_ (.A(_16823_),
    .Y(_16824_));
 AND3x1_ASAP7_75t_R _34285_ (.A(_16824_),
    .B(_15236_),
    .C(_14907_),
    .Y(_16825_));
 AO21x1_ASAP7_75t_R _34286_ (.A1(_14903_),
    .A2(_18675_),
    .B(_16825_),
    .Y(_18056_));
 NOR2x1_ASAP7_75t_R _34287_ (.A(_16333_),
    .B(_01159_),
    .Y(_16826_));
 AO21x1_ASAP7_75t_R _34288_ (.A1(_16332_),
    .A2(_16804_),
    .B(_16826_),
    .Y(_16827_));
 NAND2x1_ASAP7_75t_R _34289_ (.A(_15484_),
    .B(_01158_),
    .Y(_16828_));
 OA211x2_ASAP7_75t_R _34290_ (.A1(_16332_),
    .A2(_16807_),
    .B(_16828_),
    .C(_16337_),
    .Y(_16829_));
 AO21x1_ASAP7_75t_R _34291_ (.A1(_15594_),
    .A2(_16827_),
    .B(_16829_),
    .Y(_16830_));
 NAND2x1_ASAP7_75t_R _34292_ (.A(_15633_),
    .B(_01150_),
    .Y(_16831_));
 OA211x2_ASAP7_75t_R _34293_ (.A1(_16332_),
    .A2(_16811_),
    .B(_16831_),
    .C(_16337_),
    .Y(_16832_));
 NAND2x1_ASAP7_75t_R _34294_ (.A(_15598_),
    .B(_01149_),
    .Y(_16833_));
 OA211x2_ASAP7_75t_R _34295_ (.A1(_16332_),
    .A2(_16814_),
    .B(_16833_),
    .C(_15593_),
    .Y(_16834_));
 OA21x2_ASAP7_75t_R _34296_ (.A1(_16832_),
    .A2(_16834_),
    .B(_15482_),
    .Y(_16835_));
 AO21x1_ASAP7_75t_R _34297_ (.A1(_15588_),
    .A2(_16830_),
    .B(_16835_),
    .Y(_16836_));
 NAND2x1_ASAP7_75t_R _34298_ (.A(_15346_),
    .B(_01154_),
    .Y(_16837_));
 OA211x2_ASAP7_75t_R _34299_ (.A1(_16369_),
    .A2(_16789_),
    .B(_16837_),
    .C(_16371_),
    .Y(_16838_));
 NAND2x1_ASAP7_75t_R _34300_ (.A(_15320_),
    .B(_01153_),
    .Y(_16839_));
 OA211x2_ASAP7_75t_R _34301_ (.A1(_16369_),
    .A2(_16792_),
    .B(_16839_),
    .C(_16354_),
    .Y(_16840_));
 OR3x1_ASAP7_75t_R _34302_ (.A(_15288_),
    .B(_16838_),
    .C(_16840_),
    .Y(_16841_));
 NAND2x1_ASAP7_75t_R _34303_ (.A(_15450_),
    .B(_01162_),
    .Y(_16842_));
 OA211x2_ASAP7_75t_R _34304_ (.A1(_16369_),
    .A2(_16796_),
    .B(_16842_),
    .C(_16371_),
    .Y(_16843_));
 NAND2x1_ASAP7_75t_R _34305_ (.A(_15320_),
    .B(_01161_),
    .Y(_16844_));
 OA211x2_ASAP7_75t_R _34306_ (.A1(_16369_),
    .A2(_16799_),
    .B(_16844_),
    .C(_16354_),
    .Y(_16845_));
 OR3x1_ASAP7_75t_R _34307_ (.A(_15337_),
    .B(_16843_),
    .C(_16845_),
    .Y(_16846_));
 AND3x1_ASAP7_75t_R _34308_ (.A(_16218_),
    .B(_16841_),
    .C(_16846_),
    .Y(_16847_));
 AO21x1_ASAP7_75t_R _34309_ (.A1(_15587_),
    .A2(_16836_),
    .B(_16847_),
    .Y(_16848_));
 AND2x2_ASAP7_75t_R _34310_ (.A(_15598_),
    .B(_01772_),
    .Y(_16849_));
 AO21x1_ASAP7_75t_R _34311_ (.A1(_15436_),
    .A2(_01136_),
    .B(_16849_),
    .Y(_16850_));
 OAI22x1_ASAP7_75t_R _34312_ (.A1(_01135_),
    .A2(_15435_),
    .B1(_16850_),
    .B2(_15594_),
    .Y(_16851_));
 NAND2x1_ASAP7_75t_R _34313_ (.A(_15437_),
    .B(_01142_),
    .Y(_16852_));
 OA211x2_ASAP7_75t_R _34314_ (.A1(_15633_),
    .A2(_16765_),
    .B(_16852_),
    .C(_15600_),
    .Y(_16853_));
 NAND2x1_ASAP7_75t_R _34315_ (.A(_15437_),
    .B(_01141_),
    .Y(_16854_));
 OA211x2_ASAP7_75t_R _34316_ (.A1(_15633_),
    .A2(_16768_),
    .B(_16854_),
    .C(_15295_),
    .Y(_16855_));
 OR3x1_ASAP7_75t_R _34317_ (.A(_15596_),
    .B(_16853_),
    .C(_16855_),
    .Y(_16856_));
 OA211x2_ASAP7_75t_R _34318_ (.A1(_15588_),
    .A2(_16851_),
    .B(_16856_),
    .C(_15587_),
    .Y(_16857_));
 NAND2x1_ASAP7_75t_R _34319_ (.A(_15343_),
    .B(_01138_),
    .Y(_16858_));
 OA211x2_ASAP7_75t_R _34320_ (.A1(_16373_),
    .A2(_16773_),
    .B(_16858_),
    .C(_16371_),
    .Y(_16859_));
 NAND2x1_ASAP7_75t_R _34321_ (.A(_15486_),
    .B(_01137_),
    .Y(_16860_));
 OA211x2_ASAP7_75t_R _34322_ (.A1(_16373_),
    .A2(_16776_),
    .B(_16860_),
    .C(_16354_),
    .Y(_16861_));
 OR3x1_ASAP7_75t_R _34323_ (.A(_16368_),
    .B(_16859_),
    .C(_16861_),
    .Y(_16862_));
 NAND2x1_ASAP7_75t_R _34324_ (.A(_15486_),
    .B(_01146_),
    .Y(_16863_));
 OA211x2_ASAP7_75t_R _34325_ (.A1(_16373_),
    .A2(_16780_),
    .B(_16863_),
    .C(_16371_),
    .Y(_16864_));
 NAND2x1_ASAP7_75t_R _34326_ (.A(_15589_),
    .B(_01145_),
    .Y(_16865_));
 OA211x2_ASAP7_75t_R _34327_ (.A1(_16373_),
    .A2(_16783_),
    .B(_16865_),
    .C(_15295_),
    .Y(_16866_));
 OR3x1_ASAP7_75t_R _34328_ (.A(_15596_),
    .B(_16864_),
    .C(_16866_),
    .Y(_16867_));
 AND3x1_ASAP7_75t_R _34329_ (.A(_16218_),
    .B(_16862_),
    .C(_16867_),
    .Y(_16868_));
 OR3x1_ASAP7_75t_R _34330_ (.A(_15434_),
    .B(_16857_),
    .C(_16868_),
    .Y(_16869_));
 OA21x2_ASAP7_75t_R _34331_ (.A1(_15466_),
    .A2(_16848_),
    .B(_16869_),
    .Y(_16870_));
 INVx2_ASAP7_75t_R _34332_ (.A(_16870_),
    .Y(_16871_));
 OA211x2_ASAP7_75t_R _34333_ (.A1(_15466_),
    .A2(_16386_),
    .B(_16389_),
    .C(_15503_),
    .Y(_16872_));
 AOI21x1_ASAP7_75t_R _34334_ (.A1(_14090_),
    .A2(_16871_),
    .B(_16872_),
    .Y(_18674_));
 INVx1_ASAP7_75t_R _34335_ (.A(_18674_),
    .Y(_18672_));
 INVx2_ASAP7_75t_R _34336_ (.A(_01189_),
    .Y(_16873_));
 NOR2x1_ASAP7_75t_R _34337_ (.A(_13197_),
    .B(_01191_),
    .Y(_16874_));
 AO21x1_ASAP7_75t_R _34338_ (.A1(_14278_),
    .A2(_16873_),
    .B(_16874_),
    .Y(_16875_));
 INVx2_ASAP7_75t_R _34339_ (.A(_01192_),
    .Y(_16876_));
 NAND2x1_ASAP7_75t_R _34340_ (.A(_14717_),
    .B(_01190_),
    .Y(_16877_));
 OA211x2_ASAP7_75t_R _34341_ (.A1(_13190_),
    .A2(_16876_),
    .B(_16877_),
    .C(_14363_),
    .Y(_16878_));
 AO21x1_ASAP7_75t_R _34342_ (.A1(_13090_),
    .A2(_16875_),
    .B(_16878_),
    .Y(_16879_));
 INVx2_ASAP7_75t_R _34343_ (.A(_01184_),
    .Y(_16880_));
 NAND2x1_ASAP7_75t_R _34344_ (.A(_14461_),
    .B(_01182_),
    .Y(_16881_));
 OA211x2_ASAP7_75t_R _34345_ (.A1(_15191_),
    .A2(_16880_),
    .B(_16881_),
    .C(_14315_),
    .Y(_16882_));
 INVx2_ASAP7_75t_R _34346_ (.A(_01183_),
    .Y(_16883_));
 NAND2x1_ASAP7_75t_R _34347_ (.A(_15052_),
    .B(_01181_),
    .Y(_16884_));
 OA211x2_ASAP7_75t_R _34348_ (.A1(_15191_),
    .A2(_16883_),
    .B(_16884_),
    .C(_15195_),
    .Y(_16885_));
 OA21x2_ASAP7_75t_R _34349_ (.A1(_16882_),
    .A2(_16885_),
    .B(_13186_),
    .Y(_16886_));
 AO21x1_ASAP7_75t_R _34350_ (.A1(_14283_),
    .A2(_16879_),
    .B(_16886_),
    .Y(_16887_));
 INVx2_ASAP7_75t_R _34351_ (.A(_01188_),
    .Y(_16888_));
 NAND2x1_ASAP7_75t_R _34352_ (.A(_14277_),
    .B(_01186_),
    .Y(_16889_));
 OA211x2_ASAP7_75t_R _34353_ (.A1(_14293_),
    .A2(_16888_),
    .B(_16889_),
    .C(_14296_),
    .Y(_16890_));
 INVx2_ASAP7_75t_R _34354_ (.A(_01187_),
    .Y(_16891_));
 NAND2x1_ASAP7_75t_R _34355_ (.A(_14301_),
    .B(_01185_),
    .Y(_16892_));
 OA211x2_ASAP7_75t_R _34356_ (.A1(_14299_),
    .A2(_16891_),
    .B(_16892_),
    .C(_13149_),
    .Y(_16893_));
 OR3x1_ASAP7_75t_R _34357_ (.A(_14282_),
    .B(_16890_),
    .C(_16893_),
    .Y(_16894_));
 INVx2_ASAP7_75t_R _34358_ (.A(_01196_),
    .Y(_16895_));
 NAND2x1_ASAP7_75t_R _34359_ (.A(_14277_),
    .B(_01194_),
    .Y(_16896_));
 OA211x2_ASAP7_75t_R _34360_ (.A1(_14299_),
    .A2(_16895_),
    .B(_16896_),
    .C(_14296_),
    .Y(_16897_));
 INVx2_ASAP7_75t_R _34361_ (.A(_01195_),
    .Y(_16898_));
 NAND2x1_ASAP7_75t_R _34362_ (.A(_14301_),
    .B(_01193_),
    .Y(_16899_));
 OA211x2_ASAP7_75t_R _34363_ (.A1(_14299_),
    .A2(_16898_),
    .B(_16899_),
    .C(_14372_),
    .Y(_16900_));
 OR3x1_ASAP7_75t_R _34364_ (.A(_14291_),
    .B(_16897_),
    .C(_16900_),
    .Y(_16901_));
 AND3x1_ASAP7_75t_R _34365_ (.A(_13129_),
    .B(_16894_),
    .C(_16901_),
    .Y(_16902_));
 AO21x1_ASAP7_75t_R _34366_ (.A1(_14778_),
    .A2(_16887_),
    .B(_16902_),
    .Y(_16903_));
 AND2x2_ASAP7_75t_R _34367_ (.A(_15061_),
    .B(_01771_),
    .Y(_16904_));
 AO21x1_ASAP7_75t_R _34368_ (.A1(_13092_),
    .A2(_01168_),
    .B(_16904_),
    .Y(_16905_));
 OAI22x1_ASAP7_75t_R _34369_ (.A1(_01167_),
    .A2(_13102_),
    .B1(_16905_),
    .B2(_14975_),
    .Y(_16906_));
 INVx2_ASAP7_75t_R _34370_ (.A(_01176_),
    .Y(_16907_));
 NAND2x1_ASAP7_75t_R _34371_ (.A(_13142_),
    .B(_01174_),
    .Y(_16908_));
 OA211x2_ASAP7_75t_R _34372_ (.A1(_14455_),
    .A2(_16907_),
    .B(_16908_),
    .C(_14914_),
    .Y(_16909_));
 INVx2_ASAP7_75t_R _34373_ (.A(_01175_),
    .Y(_16910_));
 NAND2x1_ASAP7_75t_R _34374_ (.A(_13142_),
    .B(_01173_),
    .Y(_16911_));
 OA211x2_ASAP7_75t_R _34375_ (.A1(_14461_),
    .A2(_16910_),
    .B(_16911_),
    .C(_14463_),
    .Y(_16912_));
 OR3x1_ASAP7_75t_R _34376_ (.A(_14454_),
    .B(_16909_),
    .C(_16912_),
    .Y(_16913_));
 OA211x2_ASAP7_75t_R _34377_ (.A1(_14448_),
    .A2(_16906_),
    .B(_16913_),
    .C(_14466_),
    .Y(_16914_));
 INVx2_ASAP7_75t_R _34378_ (.A(_01172_),
    .Y(_16915_));
 NAND2x1_ASAP7_75t_R _34379_ (.A(_14470_),
    .B(_01170_),
    .Y(_16916_));
 OA211x2_ASAP7_75t_R _34380_ (.A1(_13193_),
    .A2(_16915_),
    .B(_16916_),
    .C(_14472_),
    .Y(_16917_));
 INVx2_ASAP7_75t_R _34381_ (.A(_01171_),
    .Y(_16918_));
 NAND2x1_ASAP7_75t_R _34382_ (.A(_14310_),
    .B(_01169_),
    .Y(_16919_));
 OA211x2_ASAP7_75t_R _34383_ (.A1(_14474_),
    .A2(_16918_),
    .B(_16919_),
    .C(_14476_),
    .Y(_16920_));
 OR3x1_ASAP7_75t_R _34384_ (.A(_14469_),
    .B(_16917_),
    .C(_16920_),
    .Y(_16921_));
 INVx2_ASAP7_75t_R _34385_ (.A(_01180_),
    .Y(_16922_));
 NAND2x1_ASAP7_75t_R _34386_ (.A(_14470_),
    .B(_01178_),
    .Y(_16923_));
 OA211x2_ASAP7_75t_R _34387_ (.A1(_13193_),
    .A2(_16922_),
    .B(_16923_),
    .C(_14472_),
    .Y(_16924_));
 INVx2_ASAP7_75t_R _34388_ (.A(_01179_),
    .Y(_16925_));
 NAND2x1_ASAP7_75t_R _34389_ (.A(_14310_),
    .B(_01177_),
    .Y(_16926_));
 OA211x2_ASAP7_75t_R _34390_ (.A1(_14474_),
    .A2(_16925_),
    .B(_16926_),
    .C(_14476_),
    .Y(_16927_));
 OR3x1_ASAP7_75t_R _34391_ (.A(_14353_),
    .B(_16924_),
    .C(_16927_),
    .Y(_16928_));
 AND3x1_ASAP7_75t_R _34392_ (.A(_14468_),
    .B(_16921_),
    .C(_16928_),
    .Y(_16929_));
 OR3x1_ASAP7_75t_R _34393_ (.A(_14447_),
    .B(_16914_),
    .C(_16929_),
    .Y(_16930_));
 OA21x2_ASAP7_75t_R _34394_ (.A1(_14339_),
    .A2(_16903_),
    .B(_16930_),
    .Y(_16931_));
 AND2x2_ASAP7_75t_R _34395_ (.A(_01460_),
    .B(_14772_),
    .Y(_16932_));
 OAI22x1_ASAP7_75t_R _34396_ (.A1(_01490_),
    .A2(_14967_),
    .B1(_14968_),
    .B2(_16932_),
    .Y(_16933_));
 OA21x2_ASAP7_75t_R _34397_ (.A1(_14709_),
    .A2(_16931_),
    .B(_16933_),
    .Y(_16934_));
 BUFx3_ASAP7_75t_R _34398_ (.A(_16934_),
    .Y(_18680_));
 INVx2_ASAP7_75t_R _34399_ (.A(_18680_),
    .Y(_18678_));
 BUFx6f_ASAP7_75t_R _34400_ (.A(_00145_),
    .Y(_16935_));
 INVx1_ASAP7_75t_R _34401_ (.A(_16935_),
    .Y(_16936_));
 AND3x1_ASAP7_75t_R _34402_ (.A(_16936_),
    .B(_15236_),
    .C(_14907_),
    .Y(_16937_));
 AO21x1_ASAP7_75t_R _34403_ (.A1(_14903_),
    .A2(_18680_),
    .B(_16937_),
    .Y(_18058_));
 AND2x2_ASAP7_75t_R _34404_ (.A(_15319_),
    .B(_01771_),
    .Y(_16938_));
 AO21x1_ASAP7_75t_R _34405_ (.A1(_15290_),
    .A2(_01168_),
    .B(_16938_),
    .Y(_16939_));
 OAI22x1_ASAP7_75t_R _34406_ (.A1(_01167_),
    .A2(_15289_),
    .B1(_16939_),
    .B2(_15593_),
    .Y(_16940_));
 NAND2x1_ASAP7_75t_R _34407_ (.A(net1971),
    .B(_01174_),
    .Y(_16941_));
 OA211x2_ASAP7_75t_R _34408_ (.A1(_15632_),
    .A2(_16907_),
    .B(_16941_),
    .C(_15266_),
    .Y(_16942_));
 NAND2x1_ASAP7_75t_R _34409_ (.A(net1971),
    .B(_01173_),
    .Y(_16943_));
 OA211x2_ASAP7_75t_R _34410_ (.A1(_15632_),
    .A2(_16910_),
    .B(_16943_),
    .C(_15274_),
    .Y(_16944_));
 OR3x1_ASAP7_75t_R _34411_ (.A(_15278_),
    .B(_16942_),
    .C(_16944_),
    .Y(_16945_));
 OA211x2_ASAP7_75t_R _34412_ (.A1(_16368_),
    .A2(_16940_),
    .B(_16945_),
    .C(_15312_),
    .Y(_16946_));
 NAND2x1_ASAP7_75t_R _34413_ (.A(_15342_),
    .B(_01170_),
    .Y(_16947_));
 BUFx6f_ASAP7_75t_R _34414_ (.A(_15265_),
    .Y(_16948_));
 OA211x2_ASAP7_75t_R _34415_ (.A1(_16106_),
    .A2(_16915_),
    .B(_16947_),
    .C(_16948_),
    .Y(_16949_));
 NAND2x1_ASAP7_75t_R _34416_ (.A(_15485_),
    .B(_01169_),
    .Y(_16950_));
 OA211x2_ASAP7_75t_R _34417_ (.A1(_16109_),
    .A2(_16918_),
    .B(_16950_),
    .C(_15294_),
    .Y(_16951_));
 OR3x1_ASAP7_75t_R _34418_ (.A(_15287_),
    .B(_16949_),
    .C(_16951_),
    .Y(_16952_));
 NAND2x1_ASAP7_75t_R _34419_ (.A(_15485_),
    .B(_01178_),
    .Y(_16953_));
 OA211x2_ASAP7_75t_R _34420_ (.A1(_16109_),
    .A2(_16922_),
    .B(_16953_),
    .C(_16948_),
    .Y(_16954_));
 NAND2x1_ASAP7_75t_R _34421_ (.A(_15485_),
    .B(_01177_),
    .Y(_16955_));
 OA211x2_ASAP7_75t_R _34422_ (.A1(_15618_),
    .A2(_16925_),
    .B(_16955_),
    .C(_15294_),
    .Y(_16956_));
 OR3x1_ASAP7_75t_R _34423_ (.A(_15336_),
    .B(_16954_),
    .C(_16956_),
    .Y(_16957_));
 AND3x1_ASAP7_75t_R _34424_ (.A(_15252_),
    .B(_16952_),
    .C(_16957_),
    .Y(_16958_));
 OR3x2_ASAP7_75t_R _34425_ (.A(_15251_),
    .B(_16946_),
    .C(_16958_),
    .Y(_16959_));
 NAND2x1_ASAP7_75t_R _34426_ (.A(_15342_),
    .B(_01186_),
    .Y(_16960_));
 OA211x2_ASAP7_75t_R _34427_ (.A1(_16106_),
    .A2(_16888_),
    .B(_16960_),
    .C(_15752_),
    .Y(_16961_));
 NAND2x1_ASAP7_75t_R _34428_ (.A(_15342_),
    .B(_01185_),
    .Y(_16962_));
 OA211x2_ASAP7_75t_R _34429_ (.A1(_16106_),
    .A2(_16891_),
    .B(_16962_),
    .C(_15294_),
    .Y(_16963_));
 OR3x1_ASAP7_75t_R _34430_ (.A(_15287_),
    .B(_16961_),
    .C(_16963_),
    .Y(_16964_));
 NAND2x1_ASAP7_75t_R _34431_ (.A(_15342_),
    .B(_01194_),
    .Y(_16965_));
 OA211x2_ASAP7_75t_R _34432_ (.A1(_16106_),
    .A2(_16895_),
    .B(_16965_),
    .C(_16948_),
    .Y(_16966_));
 NAND2x1_ASAP7_75t_R _34433_ (.A(_15485_),
    .B(_01193_),
    .Y(_16967_));
 OA211x2_ASAP7_75t_R _34434_ (.A1(_16109_),
    .A2(_16898_),
    .B(_16967_),
    .C(_15294_),
    .Y(_16968_));
 OR3x1_ASAP7_75t_R _34435_ (.A(_15336_),
    .B(_16966_),
    .C(_16968_),
    .Y(_16969_));
 AND3x1_ASAP7_75t_R _34436_ (.A(_15252_),
    .B(_16964_),
    .C(_16969_),
    .Y(_16970_));
 NOR2x1_ASAP7_75t_R _34437_ (.A(_15302_),
    .B(_01191_),
    .Y(_16971_));
 AO21x1_ASAP7_75t_R _34438_ (.A1(_15300_),
    .A2(_16873_),
    .B(_16971_),
    .Y(_16972_));
 NAND2x1_ASAP7_75t_R _34439_ (.A(_15259_),
    .B(_01190_),
    .Y(_16973_));
 OA211x2_ASAP7_75t_R _34440_ (.A1(_15270_),
    .A2(_16876_),
    .B(_16973_),
    .C(_15752_),
    .Y(_16974_));
 AO21x1_ASAP7_75t_R _34441_ (.A1(_16354_),
    .A2(_16972_),
    .B(_16974_),
    .Y(_16975_));
 NAND2x1_ASAP7_75t_R _34442_ (.A(net1969),
    .B(_01182_),
    .Y(_16976_));
 OA211x2_ASAP7_75t_R _34443_ (.A1(_15632_),
    .A2(_16880_),
    .B(_16976_),
    .C(_15266_),
    .Y(_16977_));
 NAND2x1_ASAP7_75t_R _34444_ (.A(net1969),
    .B(_01181_),
    .Y(_16978_));
 OA211x2_ASAP7_75t_R _34445_ (.A1(_15489_),
    .A2(_16883_),
    .B(_16978_),
    .C(_15274_),
    .Y(_16979_));
 OR3x1_ASAP7_75t_R _34446_ (.A(_15287_),
    .B(_16977_),
    .C(_16979_),
    .Y(_16980_));
 OA211x2_ASAP7_75t_R _34447_ (.A1(_15596_),
    .A2(_16975_),
    .B(_16980_),
    .C(_15312_),
    .Y(_16981_));
 OR3x2_ASAP7_75t_R _34448_ (.A(_15316_),
    .B(_16970_),
    .C(_16981_),
    .Y(_16982_));
 AND2x6_ASAP7_75t_R _34449_ (.A(_16959_),
    .B(_16982_),
    .Y(_16983_));
 INVx2_ASAP7_75t_R _34450_ (.A(_16983_),
    .Y(_16984_));
 OA211x2_ASAP7_75t_R _34451_ (.A1(_13831_),
    .A2(_16386_),
    .B(_16389_),
    .C(_15370_),
    .Y(_16985_));
 AOI21x1_ASAP7_75t_R _34452_ (.A1(_15250_),
    .A2(_16984_),
    .B(_16985_),
    .Y(_18679_));
 INVx1_ASAP7_75t_R _34453_ (.A(_18679_),
    .Y(_18677_));
 INVx1_ASAP7_75t_R _34454_ (.A(_01166_),
    .Y(_16986_));
 AOI21x1_ASAP7_75t_R _34455_ (.A1(_01134_),
    .A2(_16751_),
    .B(_01133_),
    .Y(_16987_));
 INVx1_ASAP7_75t_R _34456_ (.A(_01165_),
    .Y(_16988_));
 AND2x2_ASAP7_75t_R _34457_ (.A(_16988_),
    .B(_01197_),
    .Y(_16989_));
 OAI21x1_ASAP7_75t_R _34458_ (.A1(_16986_),
    .A2(_16987_),
    .B(_16989_),
    .Y(_16990_));
 INVx1_ASAP7_75t_R _34459_ (.A(_01198_),
    .Y(_16991_));
 OR4x1_ASAP7_75t_R _34460_ (.A(_16986_),
    .B(_16991_),
    .C(_01197_),
    .D(_16987_),
    .Y(_16992_));
 OR3x1_ASAP7_75t_R _34461_ (.A(_16988_),
    .B(_16991_),
    .C(_01197_),
    .Y(_16993_));
 NAND2x1_ASAP7_75t_R _34462_ (.A(_16991_),
    .B(_01197_),
    .Y(_16994_));
 AND4x1_ASAP7_75t_R _34463_ (.A(_16990_),
    .B(_16992_),
    .C(_16993_),
    .D(_16994_),
    .Y(_16995_));
 INVx4_ASAP7_75t_R _34464_ (.A(_16995_),
    .Y(\alu_adder_result_ex[25] ));
 OR2x2_ASAP7_75t_R _34465_ (.A(_01101_),
    .B(_01133_),
    .Y(_04242_));
 OA21x2_ASAP7_75t_R _34466_ (.A1(_01101_),
    .A2(_16759_),
    .B(_01134_),
    .Y(_04243_));
 OA21x2_ASAP7_75t_R _34467_ (.A1(_01133_),
    .A2(_04243_),
    .B(_01166_),
    .Y(_04244_));
 OA31x2_ASAP7_75t_R _34468_ (.A1(_16756_),
    .A2(_16758_),
    .A3(_04242_),
    .B1(_04244_),
    .Y(_04245_));
 XNOR2x1_ASAP7_75t_R _34469_ (.B(_04245_),
    .Y(_04246_),
    .A(_01165_));
 INVx6_ASAP7_75t_R _34470_ (.A(_04246_),
    .Y(\alu_adder_result_ex[24] ));
 AND2x2_ASAP7_75t_R _34471_ (.A(_13192_),
    .B(_01770_),
    .Y(_04247_));
 AO21x1_ASAP7_75t_R _34472_ (.A1(_14285_),
    .A2(_01200_),
    .B(_04247_),
    .Y(_04248_));
 OAI22x1_ASAP7_75t_R _34473_ (.A1(_01199_),
    .A2(_13101_),
    .B1(_04248_),
    .B2(_14710_),
    .Y(_04249_));
 INVx2_ASAP7_75t_R _34474_ (.A(_01208_),
    .Y(_04250_));
 NAND2x1_ASAP7_75t_R _34475_ (.A(_14755_),
    .B(_01206_),
    .Y(_04251_));
 OA211x2_ASAP7_75t_R _34476_ (.A1(_14292_),
    .A2(_04250_),
    .B(_04251_),
    .C(_13139_),
    .Y(_04252_));
 INVx2_ASAP7_75t_R _34477_ (.A(_01207_),
    .Y(_04253_));
 NAND2x1_ASAP7_75t_R _34478_ (.A(_14755_),
    .B(_01205_),
    .Y(_04254_));
 OA211x2_ASAP7_75t_R _34479_ (.A1(_14298_),
    .A2(_04253_),
    .B(_04254_),
    .C(_13173_),
    .Y(_04255_));
 OR3x1_ASAP7_75t_R _34480_ (.A(_13152_),
    .B(_04252_),
    .C(_04255_),
    .Y(_04256_));
 OA211x2_ASAP7_75t_R _34481_ (.A1(_14282_),
    .A2(_04249_),
    .B(_04256_),
    .C(_14428_),
    .Y(_04257_));
 INVx1_ASAP7_75t_R _34482_ (.A(_01204_),
    .Y(_04258_));
 NAND2x1_ASAP7_75t_R _34483_ (.A(_14391_),
    .B(_01202_),
    .Y(_04259_));
 OA211x2_ASAP7_75t_R _34484_ (.A1(_15675_),
    .A2(_04258_),
    .B(_04259_),
    .C(_14362_),
    .Y(_04260_));
 INVx1_ASAP7_75t_R _34485_ (.A(_01203_),
    .Y(_04261_));
 NAND2x1_ASAP7_75t_R _34486_ (.A(_14460_),
    .B(_01201_),
    .Y(_04262_));
 OA211x2_ASAP7_75t_R _34487_ (.A1(_13118_),
    .A2(_04261_),
    .B(_04262_),
    .C(_13088_),
    .Y(_04263_));
 OR3x1_ASAP7_75t_R _34488_ (.A(_14308_),
    .B(_04260_),
    .C(_04263_),
    .Y(_04264_));
 INVx1_ASAP7_75t_R _34489_ (.A(_01212_),
    .Y(_04265_));
 NAND2x1_ASAP7_75t_R _34490_ (.A(_14391_),
    .B(_01210_),
    .Y(_04266_));
 OA211x2_ASAP7_75t_R _34491_ (.A1(_15675_),
    .A2(_04265_),
    .B(_04266_),
    .C(_14362_),
    .Y(_04267_));
 INVx2_ASAP7_75t_R _34492_ (.A(_01211_),
    .Y(_04268_));
 NAND2x1_ASAP7_75t_R _34493_ (.A(_14319_),
    .B(_01209_),
    .Y(_04269_));
 OA211x2_ASAP7_75t_R _34494_ (.A1(_13118_),
    .A2(_04268_),
    .B(_04269_),
    .C(_13088_),
    .Y(_04270_));
 OR3x1_ASAP7_75t_R _34495_ (.A(_14326_),
    .B(_04267_),
    .C(_04270_),
    .Y(_04271_));
 AND3x1_ASAP7_75t_R _34496_ (.A(_14807_),
    .B(_04264_),
    .C(_04271_),
    .Y(_04272_));
 OR3x2_ASAP7_75t_R _34497_ (.A(_14447_),
    .B(_04257_),
    .C(_04272_),
    .Y(_04273_));
 INVx2_ASAP7_75t_R _34498_ (.A(_01220_),
    .Y(_04274_));
 NAND2x1_ASAP7_75t_R _34499_ (.A(_14760_),
    .B(_01218_),
    .Y(_04275_));
 OA211x2_ASAP7_75t_R _34500_ (.A1(_14317_),
    .A2(_04274_),
    .B(_04275_),
    .C(_14762_),
    .Y(_04276_));
 INVx2_ASAP7_75t_R _34501_ (.A(_01219_),
    .Y(_04277_));
 NAND2x1_ASAP7_75t_R _34502_ (.A(_14391_),
    .B(_01217_),
    .Y(_04278_));
 OA211x2_ASAP7_75t_R _34503_ (.A1(_15675_),
    .A2(_04277_),
    .B(_04278_),
    .C(_14765_),
    .Y(_04279_));
 OR3x1_ASAP7_75t_R _34504_ (.A(_14308_),
    .B(_04276_),
    .C(_04279_),
    .Y(_04280_));
 INVx2_ASAP7_75t_R _34505_ (.A(_01228_),
    .Y(_04281_));
 NAND2x1_ASAP7_75t_R _34506_ (.A(_14760_),
    .B(_01226_),
    .Y(_04282_));
 OA211x2_ASAP7_75t_R _34507_ (.A1(_13110_),
    .A2(_04281_),
    .B(_04282_),
    .C(_14362_),
    .Y(_04283_));
 INVx2_ASAP7_75t_R _34508_ (.A(_01227_),
    .Y(_04284_));
 NAND2x1_ASAP7_75t_R _34509_ (.A(_14460_),
    .B(_01225_),
    .Y(_04285_));
 OA211x2_ASAP7_75t_R _34510_ (.A1(_15675_),
    .A2(_04284_),
    .B(_04285_),
    .C(_13088_),
    .Y(_04286_));
 OR3x1_ASAP7_75t_R _34511_ (.A(_14326_),
    .B(_04283_),
    .C(_04286_),
    .Y(_04287_));
 AND3x1_ASAP7_75t_R _34512_ (.A(_14807_),
    .B(_04280_),
    .C(_04287_),
    .Y(_04288_));
 INVx2_ASAP7_75t_R _34513_ (.A(_01221_),
    .Y(_04289_));
 NOR2x1_ASAP7_75t_R _34514_ (.A(_13142_),
    .B(_01223_),
    .Y(_04290_));
 AO21x1_ASAP7_75t_R _34515_ (.A1(_14756_),
    .A2(_04289_),
    .B(_04290_),
    .Y(_04291_));
 INVx2_ASAP7_75t_R _34516_ (.A(_01224_),
    .Y(_04292_));
 NAND2x1_ASAP7_75t_R _34517_ (.A(_13096_),
    .B(_01222_),
    .Y(_04293_));
 OA211x2_ASAP7_75t_R _34518_ (.A1(_14507_),
    .A2(_04292_),
    .B(_04293_),
    .C(_14762_),
    .Y(_04294_));
 AO21x1_ASAP7_75t_R _34519_ (.A1(_13089_),
    .A2(_04291_),
    .B(_04294_),
    .Y(_04295_));
 INVx2_ASAP7_75t_R _34520_ (.A(_01216_),
    .Y(_04296_));
 NAND2x1_ASAP7_75t_R _34521_ (.A(_13199_),
    .B(_01214_),
    .Y(_04297_));
 OA211x2_ASAP7_75t_R _34522_ (.A1(_14298_),
    .A2(_04296_),
    .B(_04297_),
    .C(_13139_),
    .Y(_04298_));
 INVx2_ASAP7_75t_R _34523_ (.A(_01215_),
    .Y(_04299_));
 NAND2x1_ASAP7_75t_R _34524_ (.A(_14300_),
    .B(_01213_),
    .Y(_04300_));
 OA211x2_ASAP7_75t_R _34525_ (.A1(_14403_),
    .A2(_04299_),
    .B(_04300_),
    .C(_13173_),
    .Y(_04301_));
 OR3x1_ASAP7_75t_R _34526_ (.A(_13130_),
    .B(_04298_),
    .C(_04301_),
    .Y(_04302_));
 OA211x2_ASAP7_75t_R _34527_ (.A1(_14291_),
    .A2(_04295_),
    .B(_04302_),
    .C(_13124_),
    .Y(_04303_));
 OR3x2_ASAP7_75t_R _34528_ (.A(_14487_),
    .B(_04288_),
    .C(_04303_),
    .Y(_04304_));
 AND2x6_ASAP7_75t_R _34529_ (.A(_04273_),
    .B(_04304_),
    .Y(_04305_));
 BUFx6f_ASAP7_75t_R _34530_ (.A(_01489_),
    .Y(_04306_));
 AND2x2_ASAP7_75t_R _34531_ (.A(_01459_),
    .B(_14772_),
    .Y(_04307_));
 OAI22x1_ASAP7_75t_R _34532_ (.A1(_04306_),
    .A2(_15100_),
    .B1(_14384_),
    .B2(_04307_),
    .Y(_04308_));
 OA21x2_ASAP7_75t_R _34533_ (.A1(_13268_),
    .A2(_04305_),
    .B(_04308_),
    .Y(_04309_));
 BUFx12f_ASAP7_75t_R _34534_ (.A(_04309_),
    .Y(_18685_));
 INVx2_ASAP7_75t_R _34535_ (.A(_18685_),
    .Y(_18683_));
 BUFx6f_ASAP7_75t_R _34536_ (.A(_00153_),
    .Y(_04310_));
 INVx1_ASAP7_75t_R _34537_ (.A(_04310_),
    .Y(_04311_));
 AND3x1_ASAP7_75t_R _34538_ (.A(_04311_),
    .B(_15236_),
    .C(_14907_),
    .Y(_04312_));
 AO21x1_ASAP7_75t_R _34539_ (.A1(_14903_),
    .A2(_18685_),
    .B(_04312_),
    .Y(_18060_));
 AND2x2_ASAP7_75t_R _34540_ (.A(_15319_),
    .B(_01770_),
    .Y(_04313_));
 AO21x1_ASAP7_75t_R _34541_ (.A1(_15290_),
    .A2(_01200_),
    .B(_04313_),
    .Y(_04314_));
 OAI22x1_ASAP7_75t_R _34542_ (.A1(_01199_),
    .A2(_15289_),
    .B1(_04314_),
    .B2(_15593_),
    .Y(_04315_));
 NAND2x1_ASAP7_75t_R _34543_ (.A(net1958),
    .B(_01206_),
    .Y(_04316_));
 FAx1_ASAP7_75t_R _34544_ (.SN(\alu_adder_result_ex[0] ),
    .A(_16996_),
    .B(_16997_),
    .CI(_16998_),
    .CON(_00757_));
 FAx1_ASAP7_75t_R _34545_ (.SN(_18092_),
    .A(_17000_),
    .B(_17001_),
    .CI(_17002_),
    .CON(_17008_));
 FAx1_ASAP7_75t_R _34546_ (.SN(_17009_),
    .A(_17003_),
    .B(_17004_),
    .CI(_17005_),
    .CON(_18095_));
 FAx1_ASAP7_75t_R _34547_ (.SN(_00102_),
    .A(_17007_),
    .B(_17008_),
    .CI(_17009_),
    .CON(_00106_));
 FAx1_ASAP7_75t_R _34548_ (.SN(_18096_),
    .A(_17012_),
    .B(_17013_),
    .CI(_17014_),
    .CON(_18103_));
 FAx1_ASAP7_75t_R _34549_ (.SN(_18099_),
    .A(_17017_),
    .B(_17006_),
    .CI(_17016_),
    .CON(_17030_));
 FAx1_ASAP7_75t_R _34550_ (.SN(_18104_),
    .A(_17018_),
    .B(_17019_),
    .CI(_17020_),
    .CON(_18108_));
 FAx1_ASAP7_75t_R _34551_ (.SN(_17027_),
    .A(_17023_),
    .B(_17024_),
    .CI(_17025_),
    .CON(_00116_));
 FAx1_ASAP7_75t_R _34552_ (.SN(_17031_),
    .A(_17027_),
    .B(_17015_),
    .CI(_17022_),
    .CON(_18111_));
 FAx1_ASAP7_75t_R _34553_ (.SN(_00111_),
    .A(_17029_),
    .B(_17030_),
    .CI(_17031_),
    .CON(_00117_));
 FAx1_ASAP7_75t_R _34554_ (.SN(_18109_),
    .A(_17034_),
    .B(_17035_),
    .CI(_17036_),
    .CON(_18120_));
 FAx1_ASAP7_75t_R _34555_ (.SN(_18110_),
    .A(_17039_),
    .B(_17040_),
    .CI(_17041_),
    .CON(_18127_));
 FAx1_ASAP7_75t_R _34556_ (.SN(_18112_),
    .A(_17042_),
    .B(_17021_),
    .CI(_17038_),
    .CON(_18122_));
 FAx1_ASAP7_75t_R _34557_ (.SN(_18114_),
    .A(_17045_),
    .B(_17028_),
    .CI(_17044_),
    .CON(_17060_));
 FAx1_ASAP7_75t_R _34558_ (.SN(_18121_),
    .A(_17046_),
    .B(_17047_),
    .CI(_17048_),
    .CON(_18132_));
 FAx1_ASAP7_75t_R _34559_ (.SN(_17055_),
    .A(_17051_),
    .B(_17052_),
    .CI(_17053_),
    .CON(_00130_));
 FAx1_ASAP7_75t_R _34560_ (.SN(_18123_),
    .A(_17055_),
    .B(_17037_),
    .CI(_17050_),
    .CON(_18134_));
 FAx1_ASAP7_75t_R _34561_ (.SN(_17061_),
    .A(_17043_),
    .B(_17057_),
    .CI(_17058_),
    .CON(_17085_));
 FAx1_ASAP7_75t_R _34562_ (.SN(_00124_),
    .A(_17059_),
    .B(_17060_),
    .CI(_17061_),
    .CON(_00132_));
 FAx1_ASAP7_75t_R _34563_ (.SN(_18133_),
    .A(_17064_),
    .B(_17065_),
    .CI(_17066_),
    .CON(_18140_));
 FAx1_ASAP7_75t_R _34564_ (.SN(_17073_),
    .A(_17069_),
    .B(_17070_),
    .CI(_17071_),
    .CON(_00137_));
 FAx1_ASAP7_75t_R _34565_ (.SN(_18135_),
    .A(_17073_),
    .B(_17049_),
    .CI(_17068_),
    .CON(_18142_));
 FAx1_ASAP7_75t_R _34566_ (.SN(_17080_),
    .A(_17076_),
    .B(_17077_),
    .CI(_17078_),
    .CON(_17107_));
 FAx1_ASAP7_75t_R _34567_ (.SN(_17082_),
    .A(_17079_),
    .B(_17080_),
    .CI(_17054_),
    .CON(_00138_));
 FAx1_ASAP7_75t_R _34568_ (.SN(_17086_),
    .A(_17082_),
    .B(_17056_),
    .CI(_17075_),
    .CON(_18144_));
 FAx1_ASAP7_75t_R _34569_ (.SN(_00131_),
    .A(_17084_),
    .B(_17085_),
    .CI(_17086_),
    .CON(_00139_));
 FAx1_ASAP7_75t_R _34570_ (.SN(_02209_),
    .A(_17089_),
    .B(_17090_),
    .CI(_17091_),
    .CON(_00174_));
 FAx1_ASAP7_75t_R _34571_ (.SN(_18141_),
    .A(_17092_),
    .B(_17093_),
    .CI(_17094_),
    .CON(_18152_));
 FAx1_ASAP7_75t_R _34572_ (.SN(_17101_),
    .A(_17097_),
    .B(_17098_),
    .CI(_17099_),
    .CON(_00146_));
 FAx1_ASAP7_75t_R _34573_ (.SN(_18143_),
    .A(_17067_),
    .B(_17096_),
    .CI(_17101_),
    .CON(_18154_));
 FAx1_ASAP7_75t_R _34574_ (.SN(_17108_),
    .A(_17104_),
    .B(_17105_),
    .CI(_17106_),
    .CON(_17129_));
 FAx1_ASAP7_75t_R _34575_ (.SN(_17110_),
    .A(_17107_),
    .B(_17108_),
    .CI(_17072_),
    .CON(_02210_));
 FAx1_ASAP7_75t_R _34576_ (.SN(_18145_),
    .A(_17110_),
    .B(_17074_),
    .CI(_17103_),
    .CON(_18156_));
 FAx1_ASAP7_75t_R _34577_ (.SN(_18147_),
    .A(_17113_),
    .B(_17083_),
    .CI(_17112_),
    .CON(_17137_));
 FAx1_ASAP7_75t_R _34578_ (.SN(_18153_),
    .A(_17114_),
    .B(_17115_),
    .CI(_17116_),
    .CON(_18164_));
 FAx1_ASAP7_75t_R _34579_ (.SN(_17122_),
    .A(_17119_),
    .B(_17120_),
    .CI(_17121_),
    .CON(_17157_));
 FAx1_ASAP7_75t_R _34580_ (.SN(_18155_),
    .A(_17122_),
    .B(_17095_),
    .CI(_17118_),
    .CON(_18166_));
 FAx1_ASAP7_75t_R _34581_ (.SN(_17130_),
    .A(_17125_),
    .B(_17126_),
    .CI(_17127_),
    .CON(_18169_));
 FAx1_ASAP7_75t_R _34582_ (.SN(_17132_),
    .A(_17129_),
    .B(_17130_),
    .CI(_17100_),
    .CON(_02211_));
 FAx1_ASAP7_75t_R _34583_ (.SN(_18157_),
    .A(_17102_),
    .B(_17124_),
    .CI(_17132_),
    .CON(_18171_));
 FAx1_ASAP7_75t_R _34584_ (.SN(_17138_),
    .A(_17135_),
    .B(_17111_),
    .CI(_17134_),
    .CON(_17166_));
 FAx1_ASAP7_75t_R _34585_ (.SN(_00148_),
    .A(_17136_),
    .B(_17137_),
    .CI(_17138_),
    .CON(_00156_));
 FAx1_ASAP7_75t_R _34586_ (.SN(_18165_),
    .A(_17141_),
    .B(_17142_),
    .CI(_17143_),
    .CON(_18177_));
 FAx1_ASAP7_75t_R _34587_ (.SN(_17149_),
    .A(_17146_),
    .B(_17147_),
    .CI(_17148_),
    .CON(_17186_));
 FAx1_ASAP7_75t_R _34588_ (.SN(_18167_),
    .A(_17149_),
    .B(_17117_),
    .CI(_17145_),
    .CON(_18179_));
 FAx1_ASAP7_75t_R _34589_ (.SN(_18168_),
    .A(_17152_),
    .B(_17153_),
    .CI(_17154_),
    .CON(_18182_));
 FAx1_ASAP7_75t_R _34590_ (.SN(_18170_),
    .A(_17157_),
    .B(_17128_),
    .CI(_17156_),
    .CON(_17200_));
 FAx1_ASAP7_75t_R _34591_ (.SN(_18172_),
    .A(_17123_),
    .B(_17151_),
    .CI(_17158_),
    .CON(_18184_));
 FAx1_ASAP7_75t_R _34592_ (.SN(_18173_),
    .A(_17161_),
    .B(_17162_),
    .CI(_17163_),
    .CON(_17196_));
 FAx1_ASAP7_75t_R _34593_ (.SN(_17167_),
    .A(_17164_),
    .B(_17133_),
    .CI(_17160_),
    .CON(_17204_));
 FAx1_ASAP7_75t_R _34594_ (.SN(_00155_),
    .A(_17165_),
    .B(_17166_),
    .CI(_17167_),
    .CON(_00164_));
 FAx1_ASAP7_75t_R _34595_ (.SN(_18178_),
    .A(_17170_),
    .B(_17171_),
    .CI(_17172_),
    .CON(_18188_));
 FAx1_ASAP7_75t_R _34596_ (.SN(_17178_),
    .A(_17175_),
    .B(_17176_),
    .CI(_17177_),
    .CON(_17224_));
 FAx1_ASAP7_75t_R _34597_ (.SN(_18180_),
    .A(_17178_),
    .B(_17144_),
    .CI(_17174_),
    .CON(_18190_));
 FAx1_ASAP7_75t_R _34598_ (.SN(_18181_),
    .A(_17181_),
    .B(_17182_),
    .CI(_17183_),
    .CON(_18193_));
 FAx1_ASAP7_75t_R _34599_ (.SN(_18183_),
    .A(_17155_),
    .B(_17185_),
    .CI(_17186_),
    .CON(_18203_));
 FAx1_ASAP7_75t_R _34600_ (.SN(_18185_),
    .A(_17188_),
    .B(_17150_),
    .CI(_17180_),
    .CON(_18195_));
 FAx1_ASAP7_75t_R _34601_ (.SN(_17197_),
    .A(_17191_),
    .B(_17192_),
    .CI(_17193_),
    .CON(_18197_));
 FAx1_ASAP7_75t_R _34602_ (.SN(_00162_),
    .A(_17195_),
    .B(_17196_),
    .CI(_17197_),
    .CON(_17235_));
 FAx1_ASAP7_75t_R _34603_ (.SN(_17201_),
    .A(_17199_),
    .B(_17198_),
    .CI(_17200_),
    .CON(_17239_));
 FAx1_ASAP7_75t_R _34604_ (.SN(_17205_),
    .A(_17201_),
    .B(_17159_),
    .CI(_17190_),
    .CON(_18205_));
 FAx1_ASAP7_75t_R _34605_ (.SN(_00163_),
    .A(_17203_),
    .B(_17204_),
    .CI(_17205_),
    .CON(_00170_));
 FAx1_ASAP7_75t_R _34606_ (.SN(_18189_),
    .A(_17208_),
    .B(_17209_),
    .CI(_17210_),
    .CON(_18210_));
 FAx1_ASAP7_75t_R _34607_ (.SN(_17216_),
    .A(_17213_),
    .B(_17214_),
    .CI(_17215_),
    .CON(_17256_));
 FAx1_ASAP7_75t_R _34608_ (.SN(_18191_),
    .A(_17216_),
    .B(_17173_),
    .CI(_17212_),
    .CON(_18212_));
 FAx1_ASAP7_75t_R _34609_ (.SN(_18192_),
    .A(_17219_),
    .B(_17220_),
    .CI(_17221_),
    .CON(_18215_));
 FAx1_ASAP7_75t_R _34610_ (.SN(_18194_),
    .A(_17184_),
    .B(_17223_),
    .CI(_17224_),
    .CON(_17272_));
 FAx1_ASAP7_75t_R _34611_ (.SN(_18196_),
    .A(_17225_),
    .B(_17179_),
    .CI(_17218_),
    .CON(_18217_));
 FAx1_ASAP7_75t_R _34612_ (.SN(_18198_),
    .A(_17228_),
    .B(_17229_),
    .CI(_17230_),
    .CON(_18219_));
 FAx1_ASAP7_75t_R _34613_ (.SN(_18202_),
    .A(_17233_),
    .B(_17194_),
    .CI(_17232_),
    .CON(_17270_));
 FAx1_ASAP7_75t_R _34614_ (.SN(_18204_),
    .A(_17235_),
    .B(_17234_),
    .CI(_17187_),
    .CON(_18223_));
 FAx1_ASAP7_75t_R _34615_ (.SN(_18206_),
    .A(_17236_),
    .B(_17189_),
    .CI(_17227_),
    .CON(_18222_));
 FAx1_ASAP7_75t_R _34616_ (.SN(_18207_),
    .A(_17239_),
    .B(_17202_),
    .CI(_17238_),
    .CON(_18224_));
 FAx1_ASAP7_75t_R _34617_ (.SN(_18211_),
    .A(_17240_),
    .B(_17241_),
    .CI(_17242_),
    .CON(_18228_));
 FAx1_ASAP7_75t_R _34618_ (.SN(_17248_),
    .A(_17245_),
    .B(_17246_),
    .CI(_17247_),
    .CON(_17295_));
 FAx1_ASAP7_75t_R _34619_ (.SN(_18213_),
    .A(_17248_),
    .B(_17211_),
    .CI(_17244_),
    .CON(_18231_));
 FAx1_ASAP7_75t_R _34620_ (.SN(_18214_),
    .A(_17251_),
    .B(_17252_),
    .CI(_17253_),
    .CON(_18234_));
 FAx1_ASAP7_75t_R _34621_ (.SN(_18216_),
    .A(_17222_),
    .B(_17255_),
    .CI(_17256_),
    .CON(_17313_));
 FAx1_ASAP7_75t_R _34622_ (.SN(_18218_),
    .A(_17257_),
    .B(_17217_),
    .CI(_17250_),
    .CON(_18236_));
 FAx1_ASAP7_75t_R _34623_ (.SN(_18220_),
    .A(_17260_),
    .B(_17261_),
    .CI(_17262_),
    .CON(_18238_));
 FAx1_ASAP7_75t_R _34624_ (.SN(_17269_),
    .A(_17265_),
    .B(_17266_),
    .CI(_17267_),
    .CON(_00182_));
 FAx1_ASAP7_75t_R _34625_ (.SN(_17271_),
    .A(_17269_),
    .B(_17231_),
    .CI(_17264_),
    .CON(_17311_));
 FAx1_ASAP7_75t_R _34626_ (.SN(_17274_),
    .A(_17270_),
    .B(_17271_),
    .CI(_17272_),
    .CON(_02212_));
 FAx1_ASAP7_75t_R _34627_ (.SN(_18221_),
    .A(_17274_),
    .B(_17226_),
    .CI(_17259_),
    .CON(_18240_));
 FAx1_ASAP7_75t_R _34628_ (.SN(_18225_),
    .A(_17276_),
    .B(_17277_),
    .CI(_17237_),
    .CON(_17321_));
 FAx1_ASAP7_75t_R _34629_ (.SN(_18229_),
    .A(_17278_),
    .B(_17279_),
    .CI(_17280_),
    .CON(_18245_));
 FAx1_ASAP7_75t_R _34630_ (.SN(_18230_),
    .A(_17283_),
    .B(_17284_),
    .CI(_17285_),
    .CON(_18250_));
 FAx1_ASAP7_75t_R _34631_ (.SN(_18232_),
    .A(_17287_),
    .B(_17243_),
    .CI(_17282_),
    .CON(_18247_));
 FAx1_ASAP7_75t_R _34632_ (.SN(_18233_),
    .A(_17290_),
    .B(_17291_),
    .CI(_17292_),
    .CON(_18251_));
 FAx1_ASAP7_75t_R _34633_ (.SN(_18235_),
    .A(_17254_),
    .B(_17294_),
    .CI(_17295_),
    .CON(_18258_));
 FAx1_ASAP7_75t_R _34634_ (.SN(_18237_),
    .A(_17297_),
    .B(_17249_),
    .CI(_17289_),
    .CON(_18253_));
 FAx1_ASAP7_75t_R _34635_ (.SN(_18239_),
    .A(_17300_),
    .B(_17301_),
    .CI(_17302_),
    .CON(_18255_));
 FAx1_ASAP7_75t_R _34636_ (.SN(_17309_),
    .A(_17305_),
    .B(_17306_),
    .CI(_17307_),
    .CON(_00188_));
 FAx1_ASAP7_75t_R _34637_ (.SN(_17312_),
    .A(_17309_),
    .B(_17263_),
    .CI(_17304_),
    .CON(_18259_));
 FAx1_ASAP7_75t_R _34638_ (.SN(_17315_),
    .A(_17311_),
    .B(_17312_),
    .CI(_17313_),
    .CON(_02213_));
 FAx1_ASAP7_75t_R _34639_ (.SN(_18241_),
    .A(_17315_),
    .B(_17258_),
    .CI(_17299_),
    .CON(_18261_));
 FAx1_ASAP7_75t_R _34640_ (.SN(_17319_),
    .A(_17318_),
    .B(_17275_),
    .CI(_17317_),
    .CON(_17361_));
 FAx1_ASAP7_75t_R _34641_ (.SN(_00184_),
    .A(_17319_),
    .B(_17320_),
    .CI(_17321_),
    .CON(_00193_));
 FAx1_ASAP7_75t_R _34642_ (.SN(_18246_),
    .A(_17324_),
    .B(_17325_),
    .CI(_17326_),
    .CON(_18268_));
 FAx1_ASAP7_75t_R _34643_ (.SN(_17332_),
    .A(_17329_),
    .B(_17330_),
    .CI(_17331_),
    .CON(_17380_));
 FAx1_ASAP7_75t_R _34644_ (.SN(_18248_),
    .A(_17332_),
    .B(_17281_),
    .CI(_17328_),
    .CON(_18269_));
 FAx1_ASAP7_75t_R _34645_ (.SN(_18249_),
    .A(_17335_),
    .B(_17336_),
    .CI(_17337_),
    .CON(_18272_));
 FAx1_ASAP7_75t_R _34646_ (.SN(_18252_),
    .A(_17293_),
    .B(_17339_),
    .CI(_17286_),
    .CON(_18279_));
 FAx1_ASAP7_75t_R _34647_ (.SN(_18254_),
    .A(_17341_),
    .B(_17288_),
    .CI(_17334_),
    .CON(_18274_));
 FAx1_ASAP7_75t_R _34648_ (.SN(_18256_),
    .A(_17344_),
    .B(_17345_),
    .CI(_17346_),
    .CON(_18276_));
 FAx1_ASAP7_75t_R _34649_ (.SN(_17353_),
    .A(_17349_),
    .B(_17350_),
    .CI(_17351_),
    .CON(_00196_));
 FAx1_ASAP7_75t_R _34650_ (.SN(_18257_),
    .A(_17353_),
    .B(_17303_),
    .CI(_17348_),
    .CON(_18280_));
 FAx1_ASAP7_75t_R _34651_ (.SN(_18260_),
    .A(_17355_),
    .B(_17296_),
    .CI(_17310_),
    .CON(_17413_));
 FAx1_ASAP7_75t_R _34652_ (.SN(_18262_),
    .A(_17298_),
    .B(_17343_),
    .CI(_17356_),
    .CON(_18282_));
 FAx1_ASAP7_75t_R _34653_ (.SN(_17362_),
    .A(_17359_),
    .B(_17316_),
    .CI(_17358_),
    .CON(_17417_));
 FAx1_ASAP7_75t_R _34654_ (.SN(_00192_),
    .A(_17360_),
    .B(_17361_),
    .CI(_17362_),
    .CON(_00198_));
 FAx1_ASAP7_75t_R _34655_ (.SN(_17372_),
    .A(_17365_),
    .B(_17366_),
    .CI(_17367_),
    .CON(_17427_));
 FAx1_ASAP7_75t_R _34656_ (.SN(_17371_),
    .A(_17368_),
    .B(_17369_),
    .CI(_17370_),
    .CON(_17436_));
 FAx1_ASAP7_75t_R _34657_ (.SN(_18270_),
    .A(_17371_),
    .B(_17327_),
    .CI(_17372_),
    .CON(_18284_));
 FAx1_ASAP7_75t_R _34658_ (.SN(_18271_),
    .A(_17375_),
    .B(_17376_),
    .CI(_17377_),
    .CON(_18287_));
 FAx1_ASAP7_75t_R _34659_ (.SN(_18273_),
    .A(_17379_),
    .B(_17380_),
    .CI(_17338_),
    .CON(_18294_));
 FAx1_ASAP7_75t_R _34660_ (.SN(_18275_),
    .A(_17333_),
    .B(_17374_),
    .CI(_17382_),
    .CON(_18289_));
 FAx1_ASAP7_75t_R _34661_ (.SN(_18277_),
    .A(_17385_),
    .B(_17386_),
    .CI(_17387_),
    .CON(_18291_));
 FAx1_ASAP7_75t_R _34662_ (.SN(_17393_),
    .A(_17390_),
    .B(_17391_),
    .CI(_17392_),
    .CON(_17460_));
 FAx1_ASAP7_75t_R _34663_ (.SN(_18278_),
    .A(_17393_),
    .B(_17347_),
    .CI(_17389_),
    .CON(_18295_));
 FAx1_ASAP7_75t_R _34664_ (.SN(_18281_),
    .A(_17354_),
    .B(_17395_),
    .CI(_17340_),
    .CON(_18302_));
 FAx1_ASAP7_75t_R _34665_ (.SN(_18283_),
    .A(_17397_),
    .B(_17342_),
    .CI(_17384_),
    .CON(_18297_));
 FAx1_ASAP7_75t_R _34666_ (.SN(_17405_),
    .A(_17400_),
    .B(_17401_),
    .CI(_17402_),
    .CON(_18300_));
 FAx1_ASAP7_75t_R _34667_ (.SN(_17409_),
    .A(_17404_),
    .B(_17405_),
    .CI(_17352_),
    .CON(_00201_));
 FAx1_ASAP7_75t_R _34668_ (.SN(_17412_),
    .A(_17407_),
    .B(_17408_),
    .CI(_17409_),
    .CON(_18303_));
 FAx1_ASAP7_75t_R _34669_ (.SN(_17414_),
    .A(_17411_),
    .B(_17412_),
    .CI(_17413_),
    .CON(_17466_));
 FAx1_ASAP7_75t_R _34670_ (.SN(_17418_),
    .A(_17414_),
    .B(_17357_),
    .CI(_17399_),
    .CON(_18305_));
 FAx1_ASAP7_75t_R _34671_ (.SN(_00197_),
    .A(_17416_),
    .B(_17417_),
    .CI(_17418_),
    .CON(_00202_));
 FAx1_ASAP7_75t_R _34672_ (.SN(_17428_),
    .A(_17421_),
    .B(_17422_),
    .CI(_17365_),
    .CON(_17472_));
 FAx1_ASAP7_75t_R _34673_ (.SN(_17426_),
    .A(_17423_),
    .B(_17424_),
    .CI(_17425_),
    .CON(_17481_));
 FAx1_ASAP7_75t_R _34674_ (.SN(_18285_),
    .A(_17426_),
    .B(_17427_),
    .CI(_17428_),
    .CON(_18308_));
 FAx1_ASAP7_75t_R _34675_ (.SN(_18286_),
    .A(_17431_),
    .B(_17432_),
    .CI(_17433_),
    .CON(_18311_));
 FAx1_ASAP7_75t_R _34676_ (.SN(_18288_),
    .A(_17436_),
    .B(_17378_),
    .CI(_17435_),
    .CON(_18318_));
 FAx1_ASAP7_75t_R _34677_ (.SN(_18290_),
    .A(_17373_),
    .B(_17430_),
    .CI(_17438_),
    .CON(_18313_));
 FAx1_ASAP7_75t_R _34678_ (.SN(_18292_),
    .A(_17441_),
    .B(_17442_),
    .CI(_17443_),
    .CON(_18315_));
 FAx1_ASAP7_75t_R _34679_ (.SN(_17449_),
    .A(_17446_),
    .B(_17447_),
    .CI(_17448_),
    .CON(_17505_));
 FAx1_ASAP7_75t_R _34680_ (.SN(_18293_),
    .A(_17449_),
    .B(_17388_),
    .CI(_17445_),
    .CON(_18319_));
 FAx1_ASAP7_75t_R _34681_ (.SN(_18296_),
    .A(_17394_),
    .B(_17451_),
    .CI(_17381_),
    .CON(_17508_));
 FAx1_ASAP7_75t_R _34682_ (.SN(_18298_),
    .A(_17452_),
    .B(_17383_),
    .CI(_17440_),
    .CON(_18321_));
 FAx1_ASAP7_75t_R _34683_ (.SN(_18299_),
    .A(_17455_),
    .B(_17456_),
    .CI(_17457_),
    .CON(_18324_));
 FAx1_ASAP7_75t_R _34684_ (.SN(_18301_),
    .A(_17403_),
    .B(_17459_),
    .CI(_17460_),
    .CON(_18325_));
 FAx1_ASAP7_75t_R _34685_ (.SN(_18304_),
    .A(_17410_),
    .B(_17461_),
    .CI(_17396_),
    .CON(_18329_));
 FAx1_ASAP7_75t_R _34686_ (.SN(_18306_),
    .A(_17463_),
    .B(_17398_),
    .CI(_17454_),
    .CON(_18327_));
 FAx1_ASAP7_75t_R _34687_ (.SN(_18307_),
    .A(_17466_),
    .B(_17415_),
    .CI(_17465_),
    .CON(_18330_));
 FAx1_ASAP7_75t_R _34688_ (.SN(_17473_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17467_),
    .CON(_17517_));
 FAx1_ASAP7_75t_R _34689_ (.SN(_17471_),
    .A(_17468_),
    .B(_17469_),
    .CI(_17470_),
    .CON(_17526_));
 FAx1_ASAP7_75t_R _34690_ (.SN(_18309_),
    .A(_17471_),
    .B(_17472_),
    .CI(_17473_),
    .CON(_18332_));
 FAx1_ASAP7_75t_R _34691_ (.SN(_18310_),
    .A(_17476_),
    .B(_17477_),
    .CI(_17478_),
    .CON(_18335_));
 FAx1_ASAP7_75t_R _34692_ (.SN(_18312_),
    .A(_17480_),
    .B(_17481_),
    .CI(_17434_),
    .CON(_18342_));
 FAx1_ASAP7_75t_R _34693_ (.SN(_18314_),
    .A(_17429_),
    .B(_17475_),
    .CI(_17483_),
    .CON(_18337_));
 FAx1_ASAP7_75t_R _34694_ (.SN(_18316_),
    .A(_17486_),
    .B(_17487_),
    .CI(_17488_),
    .CON(_18339_));
 FAx1_ASAP7_75t_R _34695_ (.SN(_17494_),
    .A(_17491_),
    .B(_17492_),
    .CI(_17493_),
    .CON(_17550_));
 FAx1_ASAP7_75t_R _34696_ (.SN(_18317_),
    .A(_17494_),
    .B(_17444_),
    .CI(_17490_),
    .CON(_18343_));
 FAx1_ASAP7_75t_R _34697_ (.SN(_18320_),
    .A(_17450_),
    .B(_17496_),
    .CI(_17437_),
    .CON(_17553_));
 FAx1_ASAP7_75t_R _34698_ (.SN(_18322_),
    .A(_17497_),
    .B(_17439_),
    .CI(_17485_),
    .CON(_18345_));
 FAx1_ASAP7_75t_R _34699_ (.SN(_18323_),
    .A(_17500_),
    .B(_17501_),
    .CI(_17502_),
    .CON(_18348_));
 FAx1_ASAP7_75t_R _34700_ (.SN(_18326_),
    .A(_17458_),
    .B(_17504_),
    .CI(_17505_),
    .CON(_18349_));
 FAx1_ASAP7_75t_R _34701_ (.SN(_17509_),
    .A(_17506_),
    .B(_17507_),
    .CI(_17508_),
    .CON(_17557_));
 FAx1_ASAP7_75t_R _34702_ (.SN(_18328_),
    .A(_17509_),
    .B(_17453_),
    .CI(_17499_),
    .CON(_18351_));
 FAx1_ASAP7_75t_R _34703_ (.SN(_18331_),
    .A(_17462_),
    .B(_17464_),
    .CI(_17511_),
    .CON(_18353_));
 FAx1_ASAP7_75t_R _34704_ (.SN(_17518_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17512_),
    .CON(_17562_));
 FAx1_ASAP7_75t_R _34705_ (.SN(_17516_),
    .A(_17470_),
    .B(_17514_),
    .CI(_17515_),
    .CON(_17570_));
 FAx1_ASAP7_75t_R _34706_ (.SN(_18333_),
    .A(_17516_),
    .B(_17517_),
    .CI(_17518_),
    .CON(_18355_));
 FAx1_ASAP7_75t_R _34707_ (.SN(_18334_),
    .A(_17521_),
    .B(_17522_),
    .CI(_17523_),
    .CON(_18357_));
 FAx1_ASAP7_75t_R _34708_ (.SN(_18336_),
    .A(_17479_),
    .B(_17525_),
    .CI(_17526_),
    .CON(_18364_));
 FAx1_ASAP7_75t_R _34709_ (.SN(_18338_),
    .A(_17528_),
    .B(_17474_),
    .CI(_17520_),
    .CON(_18359_));
 FAx1_ASAP7_75t_R _34710_ (.SN(_18340_),
    .A(_17531_),
    .B(_17532_),
    .CI(_17533_),
    .CON(_18361_));
 FAx1_ASAP7_75t_R _34711_ (.SN(_17539_),
    .A(_17536_),
    .B(_17537_),
    .CI(_17538_),
    .CON(_17595_));
 FAx1_ASAP7_75t_R _34712_ (.SN(_18341_),
    .A(_17539_),
    .B(_17489_),
    .CI(_17535_),
    .CON(_18365_));
 FAx1_ASAP7_75t_R _34713_ (.SN(_18344_),
    .A(_17495_),
    .B(_17541_),
    .CI(_17482_),
    .CON(_17598_));
 FAx1_ASAP7_75t_R _34714_ (.SN(_18346_),
    .A(_17542_),
    .B(_17484_),
    .CI(_17530_),
    .CON(_18367_));
 FAx1_ASAP7_75t_R _34715_ (.SN(_18347_),
    .A(_17545_),
    .B(_17546_),
    .CI(_17547_),
    .CON(_18370_));
 FAx1_ASAP7_75t_R _34716_ (.SN(_18350_),
    .A(_17503_),
    .B(_17549_),
    .CI(_17550_),
    .CON(_18371_));
 FAx1_ASAP7_75t_R _34717_ (.SN(_17554_),
    .A(_17551_),
    .B(_17552_),
    .CI(_17553_),
    .CON(_17602_));
 FAx1_ASAP7_75t_R _34718_ (.SN(_18352_),
    .A(_17554_),
    .B(_17498_),
    .CI(_17544_),
    .CON(_18373_));
 FAx1_ASAP7_75t_R _34719_ (.SN(_18354_),
    .A(_17557_),
    .B(_17510_),
    .CI(_17556_),
    .CON(_18375_));
 FAx1_ASAP7_75t_R _34720_ (.SN(_17563_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17558_),
    .CON(_17604_));
 FAx1_ASAP7_75t_R _34721_ (.SN(_17564_),
    .A(_17560_),
    .B(_17470_),
    .CI(_17515_),
    .CON(_17612_));
 FAx1_ASAP7_75t_R _34722_ (.SN(_17573_),
    .A(_17561_),
    .B(_17559_),
    .CI(_17513_),
    .CON(_17615_));
 FAx1_ASAP7_75t_R _34723_ (.SN(_18356_),
    .A(_17565_),
    .B(_17566_),
    .CI(_17567_),
    .CON(_18378_));
 FAx1_ASAP7_75t_R _34724_ (.SN(_18358_),
    .A(_17524_),
    .B(_17569_),
    .CI(_17570_),
    .CON(_18385_));
 FAx1_ASAP7_75t_R _34725_ (.SN(_18360_),
    .A(_17572_),
    .B(_17519_),
    .CI(_17573_),
    .CON(_18380_));
 FAx1_ASAP7_75t_R _34726_ (.SN(_18362_),
    .A(_17576_),
    .B(_17577_),
    .CI(_17578_),
    .CON(_18382_));
 FAx1_ASAP7_75t_R _34727_ (.SN(_17584_),
    .A(_17581_),
    .B(_17582_),
    .CI(_17583_),
    .CON(_17637_));
 FAx1_ASAP7_75t_R _34728_ (.SN(_18363_),
    .A(_17584_),
    .B(_17534_),
    .CI(_17580_),
    .CON(_18386_));
 FAx1_ASAP7_75t_R _34729_ (.SN(_18366_),
    .A(_17540_),
    .B(_17586_),
    .CI(_17527_),
    .CON(_17640_));
 FAx1_ASAP7_75t_R _34730_ (.SN(_18368_),
    .A(_17587_),
    .B(_17529_),
    .CI(_17575_),
    .CON(_18388_));
 FAx1_ASAP7_75t_R _34731_ (.SN(_18369_),
    .A(_17590_),
    .B(_17591_),
    .CI(_17592_),
    .CON(_18391_));
 FAx1_ASAP7_75t_R _34732_ (.SN(_18372_),
    .A(_17548_),
    .B(_17594_),
    .CI(_17595_),
    .CON(_18392_));
 FAx1_ASAP7_75t_R _34733_ (.SN(_17599_),
    .A(_17596_),
    .B(_17597_),
    .CI(_17598_),
    .CON(_17644_));
 FAx1_ASAP7_75t_R _34734_ (.SN(_18374_),
    .A(_17599_),
    .B(_17543_),
    .CI(_17589_),
    .CON(_18395_));
 FAx1_ASAP7_75t_R _34735_ (.SN(_18376_),
    .A(_17602_),
    .B(_17555_),
    .CI(_17601_),
    .CON(_18396_));
 FAx1_ASAP7_75t_R _34736_ (.SN(_17605_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17603_),
    .CON(_17647_));
 FAx1_ASAP7_75t_R _34737_ (.SN(_18377_),
    .A(_17604_),
    .B(_17605_),
    .CI(_17564_),
    .CON(_18398_));
 FAx1_ASAP7_75t_R _34738_ (.SN(_17611_),
    .A(_17608_),
    .B(_17609_),
    .CI(_17610_),
    .CON(_17653_));
 FAx1_ASAP7_75t_R _34739_ (.SN(_18379_),
    .A(_17568_),
    .B(_17611_),
    .CI(_17612_),
    .CON(_18406_));
 FAx1_ASAP7_75t_R _34740_ (.SN(_18381_),
    .A(_17614_),
    .B(_17615_),
    .CI(_17607_),
    .CON(_18401_));
 FAx1_ASAP7_75t_R _34741_ (.SN(_18383_),
    .A(_17618_),
    .B(_17619_),
    .CI(_17620_),
    .CON(_18403_));
 FAx1_ASAP7_75t_R _34742_ (.SN(_17626_),
    .A(_17623_),
    .B(_17624_),
    .CI(_17625_),
    .CON(_17678_));
 FAx1_ASAP7_75t_R _34743_ (.SN(_18384_),
    .A(_17626_),
    .B(_17579_),
    .CI(_17622_),
    .CON(_18407_));
 FAx1_ASAP7_75t_R _34744_ (.SN(_18387_),
    .A(_17585_),
    .B(_17628_),
    .CI(_17571_),
    .CON(_17681_));
 FAx1_ASAP7_75t_R _34745_ (.SN(_18389_),
    .A(_17629_),
    .B(_17574_),
    .CI(_17617_),
    .CON(_18409_));
 FAx1_ASAP7_75t_R _34746_ (.SN(_18390_),
    .A(_17632_),
    .B(_17633_),
    .CI(_17634_),
    .CON(_18412_));
 FAx1_ASAP7_75t_R _34747_ (.SN(_18393_),
    .A(_17593_),
    .B(_17636_),
    .CI(_17637_),
    .CON(_18413_));
 FAx1_ASAP7_75t_R _34748_ (.SN(_17641_),
    .A(_17638_),
    .B(_17639_),
    .CI(_17640_),
    .CON(_17685_));
 FAx1_ASAP7_75t_R _34749_ (.SN(_18394_),
    .A(_17641_),
    .B(_17588_),
    .CI(_17631_),
    .CON(_18415_));
 FAx1_ASAP7_75t_R _34750_ (.SN(_18397_),
    .A(_17643_),
    .B(_17644_),
    .CI(_17600_),
    .CON(_18417_));
 FAx1_ASAP7_75t_R _34751_ (.SN(_17648_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17645_),
    .CON(_17690_));
 FAx1_ASAP7_75t_R _34752_ (.SN(_18399_),
    .A(_17647_),
    .B(_17648_),
    .CI(net32),
    .CON(_18419_));
 FAx1_ASAP7_75t_R _34753_ (.SN(_17654_),
    .A(_17610_),
    .B(_17651_),
    .CI(_17652_),
    .CON(_17693_));
 FAx1_ASAP7_75t_R _34754_ (.SN(_18400_),
    .A(_17612_),
    .B(_17653_),
    .CI(_17654_),
    .CON(_18426_));
 FAx1_ASAP7_75t_R _34755_ (.SN(_18402_),
    .A(_17656_),
    .B(_17606_),
    .CI(_17650_),
    .CON(_18421_));
 FAx1_ASAP7_75t_R _34756_ (.SN(_18404_),
    .A(_17659_),
    .B(_17660_),
    .CI(_17661_),
    .CON(_18423_));
 FAx1_ASAP7_75t_R _34757_ (.SN(_17667_),
    .A(_17664_),
    .B(_17665_),
    .CI(_17666_),
    .CON(_17719_));
 FAx1_ASAP7_75t_R _34758_ (.SN(_18405_),
    .A(_17667_),
    .B(_17621_),
    .CI(_17663_),
    .CON(_18427_));
 FAx1_ASAP7_75t_R _34759_ (.SN(_18408_),
    .A(_17627_),
    .B(_17669_),
    .CI(_17613_),
    .CON(_17722_));
 FAx1_ASAP7_75t_R _34760_ (.SN(_18410_),
    .A(_17670_),
    .B(_17616_),
    .CI(_17658_),
    .CON(_18429_));
 FAx1_ASAP7_75t_R _34761_ (.SN(_18411_),
    .A(_17673_),
    .B(_17674_),
    .CI(_17675_),
    .CON(_18432_));
 FAx1_ASAP7_75t_R _34762_ (.SN(_18414_),
    .A(_17635_),
    .B(_17677_),
    .CI(_17678_),
    .CON(_18433_));
 FAx1_ASAP7_75t_R _34763_ (.SN(_17682_),
    .A(_17679_),
    .B(_17680_),
    .CI(_17681_),
    .CON(_17726_));
 FAx1_ASAP7_75t_R _34764_ (.SN(_18416_),
    .A(_17682_),
    .B(_17630_),
    .CI(_17672_),
    .CON(_18435_));
 FAx1_ASAP7_75t_R _34765_ (.SN(_18418_),
    .A(_17685_),
    .B(_17642_),
    .CI(_17684_),
    .CON(_18437_));
 FAx1_ASAP7_75t_R _34766_ (.SN(_17691_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17686_),
    .CON(_17732_));
 FAx1_ASAP7_75t_R _34767_ (.SN(_17697_),
    .A(_17561_),
    .B(_17646_),
    .CI(_17688_),
    .CON(_17738_));
 FAx1_ASAP7_75t_R _34768_ (.SN(_17694_),
    .A(_17610_),
    .B(_17652_),
    .CI(_17692_),
    .CON(_17734_));
 FAx1_ASAP7_75t_R _34769_ (.SN(_18420_),
    .A(_17612_),
    .B(_17693_),
    .CI(_17694_),
    .CON(_18442_));
 FAx1_ASAP7_75t_R _34770_ (.SN(_18422_),
    .A(_17696_),
    .B(_17649_),
    .CI(_17697_),
    .CON(_18439_));
 FAx1_ASAP7_75t_R _34771_ (.SN(_18424_),
    .A(_17700_),
    .B(_17701_),
    .CI(_17702_),
    .CON(_18440_));
 FAx1_ASAP7_75t_R _34772_ (.SN(_17708_),
    .A(_17705_),
    .B(_17706_),
    .CI(_17707_),
    .CON(_17759_));
 FAx1_ASAP7_75t_R _34773_ (.SN(_18425_),
    .A(_17708_),
    .B(_17662_),
    .CI(_17704_),
    .CON(_18443_));
 FAx1_ASAP7_75t_R _34774_ (.SN(_18428_),
    .A(_17668_),
    .B(_17710_),
    .CI(_17655_),
    .CON(_17762_));
 FAx1_ASAP7_75t_R _34775_ (.SN(_18430_),
    .A(_17711_),
    .B(_17657_),
    .CI(_17699_),
    .CON(_18445_));
 FAx1_ASAP7_75t_R _34776_ (.SN(_18431_),
    .A(_17714_),
    .B(_17715_),
    .CI(_17716_),
    .CON(_18448_));
 FAx1_ASAP7_75t_R _34777_ (.SN(_18434_),
    .A(_17676_),
    .B(_17718_),
    .CI(_17719_),
    .CON(_18449_));
 FAx1_ASAP7_75t_R _34778_ (.SN(_17723_),
    .A(_17720_),
    .B(_17721_),
    .CI(_17722_),
    .CON(_17766_));
 FAx1_ASAP7_75t_R _34779_ (.SN(_18436_),
    .A(_17723_),
    .B(_17671_),
    .CI(_17713_),
    .CON(_18451_));
 FAx1_ASAP7_75t_R _34780_ (.SN(_18438_),
    .A(_17726_),
    .B(_17683_),
    .CI(_17725_),
    .CON(_18453_));
 FAx1_ASAP7_75t_R _34781_ (.SN(_17733_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17727_),
    .CON(_17771_));
 FAx1_ASAP7_75t_R _34782_ (.SN(_17739_),
    .A(_17561_),
    .B(_17687_),
    .CI(_17729_),
    .CON(_17773_));
 FAx1_ASAP7_75t_R _34783_ (.SN(_17737_),
    .A(_17734_),
    .B(_17612_),
    .CI(_17694_),
    .CON(_18456_));
 FAx1_ASAP7_75t_R _34784_ (.SN(_17751_),
    .A(net1962),
    .B(_17689_),
    .CI(_17731_),
    .CON(_17786_));
 FAx1_ASAP7_75t_R _34785_ (.SN(_17747_),
    .A(_17740_),
    .B(_17741_),
    .CI(_17742_),
    .CON(_17781_));
 FAx1_ASAP7_75t_R _34786_ (.SN(_17746_),
    .A(_17743_),
    .B(_17744_),
    .CI(_17745_),
    .CON(_17795_));
 FAx1_ASAP7_75t_R _34787_ (.SN(_18441_),
    .A(_17746_),
    .B(_17703_),
    .CI(_17747_),
    .CON(_18457_));
 FAx1_ASAP7_75t_R _34788_ (.SN(_18444_),
    .A(_17709_),
    .B(_17749_),
    .CI(_17695_),
    .CON(_17798_));
 FAx1_ASAP7_75t_R _34789_ (.SN(_18446_),
    .A(_17750_),
    .B(_17698_),
    .CI(_17751_),
    .CON(_18459_));
 FAx1_ASAP7_75t_R _34790_ (.SN(_18447_),
    .A(_17754_),
    .B(_17755_),
    .CI(_17756_),
    .CON(_18462_));
 FAx1_ASAP7_75t_R _34791_ (.SN(_18450_),
    .A(_17717_),
    .B(_17758_),
    .CI(_17759_),
    .CON(_18463_));
 FAx1_ASAP7_75t_R _34792_ (.SN(_17763_),
    .A(_17760_),
    .B(_17761_),
    .CI(_17762_),
    .CON(_17802_));
 FAx1_ASAP7_75t_R _34793_ (.SN(_18452_),
    .A(_17763_),
    .B(_17712_),
    .CI(_17753_),
    .CON(_18465_));
 FAx1_ASAP7_75t_R _34794_ (.SN(_18454_),
    .A(_17766_),
    .B(_17724_),
    .CI(_17765_),
    .CON(_18467_));
 FAx1_ASAP7_75t_R _34795_ (.SN(_17772_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17767_),
    .CON(_17806_));
 FAx1_ASAP7_75t_R _34796_ (.SN(_17774_),
    .A(_17561_),
    .B(_17728_),
    .CI(_17769_),
    .CON(_17808_));
 FAx1_ASAP7_75t_R _34797_ (.SN(_17787_),
    .A(net1962),
    .B(_17730_),
    .CI(_17770_),
    .CON(_17822_));
 FAx1_ASAP7_75t_R _34798_ (.SN(_17782_),
    .A(_17742_),
    .B(_17775_),
    .CI(_17776_),
    .CON(_17818_));
 FAx1_ASAP7_75t_R _34799_ (.SN(_17780_),
    .A(_17777_),
    .B(_17778_),
    .CI(_17779_),
    .CON(_17830_));
 FAx1_ASAP7_75t_R _34800_ (.SN(_18455_),
    .A(_17780_),
    .B(_17781_),
    .CI(_17782_),
    .CON(_18471_));
 FAx1_ASAP7_75t_R _34801_ (.SN(_18458_),
    .A(_17748_),
    .B(_17784_),
    .CI(_17735_),
    .CON(_17833_));
 FAx1_ASAP7_75t_R _34802_ (.SN(_18460_),
    .A(_17785_),
    .B(_17786_),
    .CI(_17787_),
    .CON(_18473_));
 FAx1_ASAP7_75t_R _34803_ (.SN(_18461_),
    .A(_17790_),
    .B(_17791_),
    .CI(_17792_),
    .CON(_18476_));
 FAx1_ASAP7_75t_R _34804_ (.SN(_18464_),
    .A(_17757_),
    .B(_17794_),
    .CI(_17795_),
    .CON(_18477_));
 FAx1_ASAP7_75t_R _34805_ (.SN(_17799_),
    .A(_17796_),
    .B(_17797_),
    .CI(_17798_),
    .CON(_17837_));
 FAx1_ASAP7_75t_R _34806_ (.SN(_18466_),
    .A(_17799_),
    .B(_17752_),
    .CI(_17789_),
    .CON(_18479_));
 FAx1_ASAP7_75t_R _34807_ (.SN(_18468_),
    .A(_17802_),
    .B(_17764_),
    .CI(_17801_),
    .CON(_18481_));
 FAx1_ASAP7_75t_R _34808_ (.SN(_17807_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17803_),
    .CON(_17841_));
 FAx1_ASAP7_75t_R _34809_ (.SN(_17809_),
    .A(_17805_),
    .B(_17768_),
    .CI(_17561_),
    .CON(_17843_));
 FAx1_ASAP7_75t_R _34810_ (.SN(_18469_),
    .A(_17809_),
    .B(_17808_),
    .CI(_17736_),
    .CON(_18483_));
 FAx1_ASAP7_75t_R _34811_ (.SN(_17816_),
    .A(_17812_),
    .B(_17742_),
    .CI(_17776_),
    .CON(_17850_));
 FAx1_ASAP7_75t_R _34812_ (.SN(_17817_),
    .A(_17813_),
    .B(_17814_),
    .CI(_17815_),
    .CON(_17862_));
 FAx1_ASAP7_75t_R _34813_ (.SN(_18470_),
    .A(_17816_),
    .B(_17817_),
    .CI(_17818_),
    .CON(_18486_));
 FAx1_ASAP7_75t_R _34814_ (.SN(_18472_),
    .A(_17783_),
    .B(_17820_),
    .CI(_17735_),
    .CON(_17865_));
 FAx1_ASAP7_75t_R _34815_ (.SN(_18474_),
    .A(_17822_),
    .B(_17811_),
    .CI(_17821_),
    .CON(_18488_));
 FAx1_ASAP7_75t_R _34816_ (.SN(_18475_),
    .A(_17825_),
    .B(_17826_),
    .CI(_17827_),
    .CON(_18491_));
 FAx1_ASAP7_75t_R _34817_ (.SN(_18478_),
    .A(_17793_),
    .B(_17829_),
    .CI(_17830_),
    .CON(_18492_));
 FAx1_ASAP7_75t_R _34818_ (.SN(_17834_),
    .A(_17831_),
    .B(_17832_),
    .CI(_17833_),
    .CON(_17869_));
 FAx1_ASAP7_75t_R _34819_ (.SN(_18480_),
    .A(_17834_),
    .B(_17788_),
    .CI(_17824_),
    .CON(_18494_));
 FAx1_ASAP7_75t_R _34820_ (.SN(_18482_),
    .A(_17837_),
    .B(_17836_),
    .CI(_17800_),
    .CON(_18496_));
 FAx1_ASAP7_75t_R _34821_ (.SN(_17842_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17838_),
    .CON(_17873_));
 FAx1_ASAP7_75t_R _34822_ (.SN(_17844_),
    .A(_17561_),
    .B(_17804_),
    .CI(_17840_),
    .CON(_17875_));
 FAx1_ASAP7_75t_R _34823_ (.SN(_18484_),
    .A(_17843_),
    .B(_17844_),
    .CI(_17736_),
    .CON(_18498_));
 FAx1_ASAP7_75t_R _34824_ (.SN(_17851_),
    .A(_17847_),
    .B(_17848_),
    .CI(_17849_),
    .CON(_17892_));
 FAx1_ASAP7_75t_R _34825_ (.SN(_18485_),
    .A(_17816_),
    .B(_17850_),
    .CI(_17851_),
    .CON(_18501_));
 FAx1_ASAP7_75t_R _34826_ (.SN(_18487_),
    .A(_17819_),
    .B(_17853_),
    .CI(_17735_),
    .CON(_17895_));
 FAx1_ASAP7_75t_R _34827_ (.SN(_18489_),
    .A(_17810_),
    .B(_17846_),
    .CI(_17854_),
    .CON(_18503_));
 FAx1_ASAP7_75t_R _34828_ (.SN(_18490_),
    .A(_17857_),
    .B(_17858_),
    .CI(_17859_),
    .CON(_18506_));
 FAx1_ASAP7_75t_R _34829_ (.SN(_18493_),
    .A(_17828_),
    .B(_17861_),
    .CI(_17862_),
    .CON(_18507_));
 FAx1_ASAP7_75t_R _34830_ (.SN(_17866_),
    .A(_17863_),
    .B(_17864_),
    .CI(_17865_),
    .CON(_17899_));
 FAx1_ASAP7_75t_R _34831_ (.SN(_18495_),
    .A(_17866_),
    .B(_17823_),
    .CI(_17856_),
    .CON(_18509_));
 FAx1_ASAP7_75t_R _34832_ (.SN(_18497_),
    .A(_17869_),
    .B(_17835_),
    .CI(_17868_),
    .CON(_18511_));
 FAx1_ASAP7_75t_R _34833_ (.SN(_17874_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17870_),
    .CON(_17902_));
 FAx1_ASAP7_75t_R _34834_ (.SN(_17876_),
    .A(_17561_),
    .B(_17839_),
    .CI(_17872_),
    .CON(_17904_));
 FAx1_ASAP7_75t_R _34835_ (.SN(_18499_),
    .A(_17875_),
    .B(_17876_),
    .CI(_17736_),
    .CON(_18513_));
 FAx1_ASAP7_75t_R _34836_ (.SN(_17881_),
    .A(_17879_),
    .B(_17880_),
    .CI(_17849_),
    .CON(_17920_));
 FAx1_ASAP7_75t_R _34837_ (.SN(_18500_),
    .A(_17816_),
    .B(_17850_),
    .CI(_17881_),
    .CON(_18516_));
 FAx1_ASAP7_75t_R _34838_ (.SN(_18502_),
    .A(_17883_),
    .B(_17735_),
    .CI(_17852_),
    .CON(_17923_));
 FAx1_ASAP7_75t_R _34839_ (.SN(_18504_),
    .A(_17845_),
    .B(_17878_),
    .CI(_17884_),
    .CON(_18518_));
 FAx1_ASAP7_75t_R _34840_ (.SN(_18505_),
    .A(_17887_),
    .B(_17888_),
    .CI(_17889_),
    .CON(_18521_));
 FAx1_ASAP7_75t_R _34841_ (.SN(_18508_),
    .A(_17860_),
    .B(_17891_),
    .CI(_17892_),
    .CON(_18522_));
 FAx1_ASAP7_75t_R _34842_ (.SN(_17896_),
    .A(_17893_),
    .B(_17894_),
    .CI(_17895_),
    .CON(_17927_));
 FAx1_ASAP7_75t_R _34843_ (.SN(_18510_),
    .A(_17896_),
    .B(_17855_),
    .CI(_17886_),
    .CON(_18524_));
 FAx1_ASAP7_75t_R _34844_ (.SN(_18512_),
    .A(_17899_),
    .B(_17867_),
    .CI(_17898_),
    .CON(_18526_));
 FAx1_ASAP7_75t_R _34845_ (.SN(_17903_),
    .A(_17421_),
    .B(_17365_),
    .CI(_17900_),
    .CON(_17929_));
 FAx1_ASAP7_75t_R _34846_ (.SN(_17905_),
    .A(_17561_),
    .B(_17871_),
    .CI(_17901_),
    .CON(_17933_));
 FAx1_ASAP7_75t_R _34847_ (.SN(_18514_),
    .A(_17904_),
    .B(_17905_),
    .CI(_17736_),
    .CON(_17938_));
 FAx1_ASAP7_75t_R _34848_ (.SN(_17909_),
    .A(_17880_),
    .B(_17907_),
    .CI(_17849_),
    .CON(_17944_));
 FAx1_ASAP7_75t_R _34849_ (.SN(_18515_),
    .A(_17816_),
    .B(_17850_),
    .CI(_17909_),
    .CON(_18528_));
 FAx1_ASAP7_75t_R _34850_ (.SN(_18517_),
    .A(_17882_),
    .B(_17911_),
    .CI(_17735_),
    .CON(_17947_));
 FAx1_ASAP7_75t_R _34851_ (.SN(_18519_),
    .A(_17912_),
    .B(_17877_),
    .CI(_17906_),
    .CON(_18529_));
 FAx1_ASAP7_75t_R _34852_ (.SN(_18520_),
    .A(_17915_),
    .B(_17916_),
    .CI(_17917_),
    .CON(_18530_));
 FAx1_ASAP7_75t_R _34853_ (.SN(_18523_),
    .A(_17890_),
    .B(_17919_),
    .CI(_17920_),
    .CON(_18531_));
 FAx1_ASAP7_75t_R _34854_ (.SN(_17924_),
    .A(_17921_),
    .B(_17922_),
    .CI(_17923_),
    .CON(_17952_));
 FAx1_ASAP7_75t_R _34855_ (.SN(_18525_),
    .A(_17924_),
    .B(_17885_),
    .CI(_17914_),
    .CON(_18533_));
 FAx1_ASAP7_75t_R _34856_ (.SN(_18527_),
    .A(_17927_),
    .B(_17897_),
    .CI(_17926_),
    .CON(_18535_));
 FAx1_ASAP7_75t_R _34857_ (.SN(_17930_),
    .A(_17928_),
    .B(_17421_),
    .CI(_17365_),
    .CON(_17954_));
 FAx1_ASAP7_75t_R _34858_ (.SN(_17935_),
    .A(_17929_),
    .B(_17930_),
    .CI(net32),
    .CON(_17960_));
 FAx1_ASAP7_75t_R _34859_ (.SN(_17939_),
    .A(_17933_),
    .B(_17932_),
    .CI(_17736_),
    .CON(_17964_));
 FAx1_ASAP7_75t_R _34860_ (.SN(_17937_),
    .A(_17910_),
    .B(_17911_),
    .CI(_17735_),
    .CON(_17973_));
 FAx1_ASAP7_75t_R _34861_ (.SN(_17949_),
    .A(_17937_),
    .B(_17938_),
    .CI(_17939_),
    .CON(_17975_));
 FAx1_ASAP7_75t_R _34862_ (.SN(_17943_),
    .A(_17940_),
    .B(_17941_),
    .CI(_17942_),
    .CON(_17969_));
 FAx1_ASAP7_75t_R _34863_ (.SN(_18532_),
    .A(_17918_),
    .B(_17943_),
    .CI(_17944_),
    .CON(_18538_));
 FAx1_ASAP7_75t_R _34864_ (.SN(_17948_),
    .A(_17945_),
    .B(_17946_),
    .CI(_17947_),
    .CON(_17978_));
 FAx1_ASAP7_75t_R _34865_ (.SN(_18534_),
    .A(_17948_),
    .B(_17913_),
    .CI(_17949_),
    .CON(_18540_));
 FAx1_ASAP7_75t_R _34866_ (.SN(_18536_),
    .A(_17952_),
    .B(_17925_),
    .CI(_17951_),
    .CON(_18542_));
 FAx1_ASAP7_75t_R _34867_ (.SN(_17955_),
    .A(_17953_),
    .B(_17421_),
    .CI(_17365_),
    .CON(_17980_));
 FAx1_ASAP7_75t_R _34868_ (.SN(_17961_),
    .A(_17954_),
    .B(_17955_),
    .CI(net32),
    .CON(_17984_));
 FAx1_ASAP7_75t_R _34869_ (.SN(_17965_),
    .A(_17931_),
    .B(_17957_),
    .CI(_17736_),
    .CON(_17987_));
 FAx1_ASAP7_75t_R _34870_ (.SN(_18537_),
    .A(_17934_),
    .B(_17959_),
    .CI(_17936_),
    .CON(_18544_));
 FAx1_ASAP7_75t_R _34871_ (.SN(_17970_),
    .A(_17966_),
    .B(_17967_),
    .CI(_17942_),
    .CON(_00250_));
 FAx1_ASAP7_75t_R _34872_ (.SN(_18539_),
    .A(_17969_),
    .B(_17970_),
    .CI(_17944_),
    .CON(_18546_));
 FAx1_ASAP7_75t_R _34873_ (.SN(_17974_),
    .A(_17971_),
    .B(_17972_),
    .CI(_17973_),
    .CON(_17996_));
 FAx1_ASAP7_75t_R _34874_ (.SN(_18541_),
    .A(_17974_),
    .B(_17975_),
    .CI(_17963_),
    .CON(_18547_));
 FAx1_ASAP7_75t_R _34875_ (.SN(_18543_),
    .A(_17978_),
    .B(_17950_),
    .CI(_17977_),
    .CON(_18549_));
 FAx1_ASAP7_75t_R _34876_ (.SN(_17981_),
    .A(_17979_),
    .B(_17421_),
    .CI(_17365_),
    .CON(_00254_));
 FAx1_ASAP7_75t_R _34877_ (.SN(_17985_),
    .A(_17980_),
    .B(_17981_),
    .CI(net32),
    .CON(_02214_));
 FAx1_ASAP7_75t_R _34878_ (.SN(_17988_),
    .A(_17956_),
    .B(_17982_),
    .CI(_17736_),
    .CON(_02215_));
 FAx1_ASAP7_75t_R _34879_ (.SN(_18545_),
    .A(_17958_),
    .B(_17983_),
    .CI(_17936_),
    .CON(_02216_));
 FAx1_ASAP7_75t_R _34880_ (.SN(_00248_),
    .A(_17989_),
    .B(_17967_),
    .CI(_17942_),
    .CON(_00255_));
 FAx1_ASAP7_75t_R _34881_ (.SN(_02217_),
    .A(_17968_),
    .B(_17990_),
    .CI(_17908_),
    .CON(_00257_));
 FAx1_ASAP7_75t_R _34882_ (.SN(_17994_),
    .A(_17992_),
    .B(_17993_),
    .CI(_17973_),
    .CON(_00258_));
 FAx1_ASAP7_75t_R _34883_ (.SN(_18548_),
    .A(_17994_),
    .B(_17962_),
    .CI(_17986_),
    .CON(_02218_));
 FAx1_ASAP7_75t_R _34884_ (.SN(_18550_),
    .A(_17996_),
    .B(_17976_),
    .CI(_17995_),
    .CON(_02219_));
 FAx1_ASAP7_75t_R _34885_ (.SN(_00265_),
    .A(_17997_),
    .B(_17998_),
    .CI(_17999_),
    .CON(_00267_));
 HAxp5_ASAP7_75t_R _34886_ (.A(_18000_),
    .B(_18001_),
    .CON(_01389_),
    .SN(_02220_));
 HAxp5_ASAP7_75t_R _34887_ (.A(_18000_),
    .B(_18002_),
    .CON(_02221_),
    .SN(_18003_));
 HAxp5_ASAP7_75t_R _34888_ (.A(_18004_),
    .B(_18001_),
    .CON(_02222_),
    .SN(_18005_));
 HAxp5_ASAP7_75t_R _34889_ (.A(_18002_),
    .B(_18004_),
    .CON(_00751_),
    .SN(_18006_));
 HAxp5_ASAP7_75t_R _34890_ (.A(_18007_),
    .B(_18008_),
    .CON(_00756_),
    .SN(_00754_));
 HAxp5_ASAP7_75t_R _34891_ (.A(_18009_),
    .B(_18010_),
    .CON(_00762_),
    .SN(_00755_));
 HAxp5_ASAP7_75t_R _34892_ (.A(_18011_),
    .B(_18012_),
    .CON(_00764_),
    .SN(_00761_));
 HAxp5_ASAP7_75t_R _34893_ (.A(_18013_),
    .B(_18014_),
    .CON(_00766_),
    .SN(_00763_));
 HAxp5_ASAP7_75t_R _34894_ (.A(_18015_),
    .B(_18016_),
    .CON(_00768_),
    .SN(_00765_));
 HAxp5_ASAP7_75t_R _34895_ (.A(_18017_),
    .B(_18018_),
    .CON(_00770_),
    .SN(_00767_));
 HAxp5_ASAP7_75t_R _34896_ (.A(_18019_),
    .B(_18020_),
    .CON(_00772_),
    .SN(_00769_));
 HAxp5_ASAP7_75t_R _34897_ (.A(_18021_),
    .B(_18022_),
    .CON(_00774_),
    .SN(_00771_));
 HAxp5_ASAP7_75t_R _34898_ (.A(_18024_),
    .B(_18023_),
    .CON(_00776_),
    .SN(_00773_));
 HAxp5_ASAP7_75t_R _34899_ (.A(_18026_),
    .B(_18025_),
    .CON(_00778_),
    .SN(_00775_));
 HAxp5_ASAP7_75t_R _34900_ (.A(_18028_),
    .B(_18027_),
    .CON(_00780_),
    .SN(_00777_));
 HAxp5_ASAP7_75t_R _34901_ (.A(_18030_),
    .B(_18029_),
    .CON(_00782_),
    .SN(_00779_));
 HAxp5_ASAP7_75t_R _34902_ (.A(_18032_),
    .B(_18031_),
    .CON(_00814_),
    .SN(_00781_));
 HAxp5_ASAP7_75t_R _34903_ (.A(_18034_),
    .B(_18033_),
    .CON(_00846_),
    .SN(_00813_));
 HAxp5_ASAP7_75t_R _34904_ (.A(_18036_),
    .B(_18035_),
    .CON(_00878_),
    .SN(_00845_));
 HAxp5_ASAP7_75t_R _34905_ (.A(_18038_),
    .B(_18037_),
    .CON(_00910_),
    .SN(_00877_));
 HAxp5_ASAP7_75t_R _34906_ (.A(_18039_),
    .B(_18040_),
    .CON(_00942_),
    .SN(_00909_));
 HAxp5_ASAP7_75t_R _34907_ (.A(_18042_),
    .B(_18041_),
    .CON(_00974_),
    .SN(_00941_));
 HAxp5_ASAP7_75t_R _34908_ (.A(_18043_),
    .B(_18044_),
    .CON(_01006_),
    .SN(_00973_));
 HAxp5_ASAP7_75t_R _34909_ (.A(_18046_),
    .B(_18045_),
    .CON(_01038_),
    .SN(_01005_));
 HAxp5_ASAP7_75t_R _34910_ (.A(_18047_),
    .B(_18048_),
    .CON(_01070_),
    .SN(_01037_));
 HAxp5_ASAP7_75t_R _34911_ (.A(_18049_),
    .B(_18050_),
    .CON(_01102_),
    .SN(_01069_));
 HAxp5_ASAP7_75t_R _34912_ (.A(_18051_),
    .B(_18052_),
    .CON(_01134_),
    .SN(_01101_));
 HAxp5_ASAP7_75t_R _34913_ (.A(_18053_),
    .B(_18054_),
    .CON(_01166_),
    .SN(_01133_));
 HAxp5_ASAP7_75t_R _34914_ (.A(_18055_),
    .B(_18056_),
    .CON(_01198_),
    .SN(_01165_));
 HAxp5_ASAP7_75t_R _34915_ (.A(_18057_),
    .B(_18058_),
    .CON(_01230_),
    .SN(_01197_));
 HAxp5_ASAP7_75t_R _34916_ (.A(_18059_),
    .B(_18060_),
    .CON(_01262_),
    .SN(_01229_));
 HAxp5_ASAP7_75t_R _34917_ (.A(_18061_),
    .B(_18062_),
    .CON(_01294_),
    .SN(_01261_));
 HAxp5_ASAP7_75t_R _34918_ (.A(_18063_),
    .B(_18064_),
    .CON(_01326_),
    .SN(_01293_));
 HAxp5_ASAP7_75t_R _34919_ (.A(_18065_),
    .B(_18066_),
    .CON(_01358_),
    .SN(_01325_));
 HAxp5_ASAP7_75t_R _34920_ (.A(_18067_),
    .B(_18068_),
    .CON(_02223_),
    .SN(_01357_));
 HAxp5_ASAP7_75t_R _34921_ (.A(_18069_),
    .B(_18070_),
    .CON(_02224_),
    .SN(_01390_));
 HAxp5_ASAP7_75t_R _34922_ (.A(_18071_),
    .B(_18072_),
    .CON(_00330_),
    .SN(_18073_));
 HAxp5_ASAP7_75t_R _34923_ (.A(_18074_),
    .B(_18075_),
    .CON(_02225_),
    .SN(_02226_));
 HAxp5_ASAP7_75t_R _34924_ (.A(_18074_),
    .B(_18076_),
    .CON(_02227_),
    .SN(_18077_));
 HAxp5_ASAP7_75t_R _34925_ (.A(_18078_),
    .B(_18075_),
    .CON(_02228_),
    .SN(_18079_));
 HAxp5_ASAP7_75t_R _34926_ (.A(_18080_),
    .B(_18081_),
    .CON(_02229_),
    .SN(_02230_));
 HAxp5_ASAP7_75t_R _34927_ (.A(\cs_registers_i.priv_mode_id_o[0] ),
    .B(_18082_),
    .CON(_02231_),
    .SN(_01392_));
 HAxp5_ASAP7_75t_R _34928_ (.A(\cs_registers_i.mhpmcounter[1856] ),
    .B(\cs_registers_i.mhpmcounter[1857] ),
    .CON(_02232_),
    .SN(_02233_));
 HAxp5_ASAP7_75t_R _34929_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .CON(_02234_),
    .SN(_02235_));
 HAxp5_ASAP7_75t_R _34930_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\cs_registers_i.pc_id_i[2] ),
    .CON(_02236_),
    .SN(_00017_));
 HAxp5_ASAP7_75t_R _34931_ (.A(_18083_),
    .B(_18084_),
    .CON(_00025_),
    .SN(_02237_));
 HAxp5_ASAP7_75t_R _34932_ (.A(_18083_),
    .B(_18084_),
    .CON(_02238_),
    .SN(_18085_));
 HAxp5_ASAP7_75t_R _34933_ (.A(_18083_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CON(_00032_),
    .SN(_18086_));
 HAxp5_ASAP7_75t_R _34934_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_18084_),
    .CON(_01395_),
    .SN(_18087_));
 HAxp5_ASAP7_75t_R _34935_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CON(_00024_),
    .SN(_18088_));
 HAxp5_ASAP7_75t_R _34936_ (.A(_18089_),
    .B(_18090_),
    .CON(_02239_),
    .SN(_00064_));
 HAxp5_ASAP7_75t_R _34937_ (.A(_18091_),
    .B(_18092_),
    .CON(_02240_),
    .SN(_00099_));
 HAxp5_ASAP7_75t_R _34938_ (.A(_18093_),
    .B(_17011_),
    .CON(_02241_),
    .SN(_00103_));
 HAxp5_ASAP7_75t_R _34939_ (.A(_18097_),
    .B(_18098_),
    .CON(_02242_),
    .SN(_17017_));
 HAxp5_ASAP7_75t_R _34940_ (.A(_17010_),
    .B(_18099_),
    .CON(_02243_),
    .SN(_00107_));
 HAxp5_ASAP7_75t_R _34941_ (.A(_18094_),
    .B(_18101_),
    .CON(_02244_),
    .SN(_00108_));
 HAxp5_ASAP7_75t_R _34942_ (.A(_18100_),
    .B(_17033_),
    .CON(_02245_),
    .SN(_00112_));
 HAxp5_ASAP7_75t_R _34943_ (.A(_18102_),
    .B(_18106_),
    .CON(_02246_),
    .SN(_00113_));
 HAxp5_ASAP7_75t_R _34944_ (.A(_18113_),
    .B(_17026_),
    .CON(_02247_),
    .SN(_17045_));
 HAxp5_ASAP7_75t_R _34945_ (.A(_17032_),
    .B(_18114_),
    .CON(_02248_),
    .SN(_00118_));
 HAxp5_ASAP7_75t_R _34946_ (.A(_18105_),
    .B(_18116_),
    .CON(_02249_),
    .SN(_00119_));
 HAxp5_ASAP7_75t_R _34947_ (.A(_18107_),
    .B(_18118_),
    .CON(_02250_),
    .SN(_00120_));
 HAxp5_ASAP7_75t_R _34948_ (.A(_18124_),
    .B(_18125_),
    .CON(_02251_),
    .SN(_00123_));
 HAxp5_ASAP7_75t_R _34949_ (.A(_18126_),
    .B(_18127_),
    .CON(_02252_),
    .SN(_17058_));
 HAxp5_ASAP7_75t_R _34950_ (.A(_18115_),
    .B(_17063_),
    .CON(_02253_),
    .SN(_00125_));
 HAxp5_ASAP7_75t_R _34951_ (.A(_18117_),
    .B(_18129_),
    .CON(_17090_),
    .SN(_00126_));
 HAxp5_ASAP7_75t_R _34952_ (.A(_18119_),
    .B(_18131_),
    .CON(_17089_),
    .SN(_00127_));
 HAxp5_ASAP7_75t_R _34953_ (.A(_17062_),
    .B(_17088_),
    .CON(_02254_),
    .SN(_00133_));
 HAxp5_ASAP7_75t_R _34954_ (.A(_18128_),
    .B(_18137_),
    .CON(_02255_),
    .SN(_17091_));
 HAxp5_ASAP7_75t_R _34955_ (.A(_18130_),
    .B(_18139_),
    .CON(_00143_),
    .SN(_00134_));
 HAxp5_ASAP7_75t_R _34956_ (.A(_18146_),
    .B(_17081_),
    .CON(_02256_),
    .SN(_17113_));
 HAxp5_ASAP7_75t_R _34957_ (.A(_17087_),
    .B(_18147_),
    .CON(_02257_),
    .SN(_00140_));
 HAxp5_ASAP7_75t_R _34958_ (.A(_18136_),
    .B(_18149_),
    .CON(_02258_),
    .SN(_00141_));
 HAxp5_ASAP7_75t_R _34959_ (.A(_18138_),
    .B(_18151_),
    .CON(_00151_),
    .SN(_00142_));
 HAxp5_ASAP7_75t_R _34960_ (.A(_18158_),
    .B(_18159_),
    .CON(_02259_),
    .SN(_00147_));
 HAxp5_ASAP7_75t_R _34961_ (.A(_18161_),
    .B(_17109_),
    .CON(_02260_),
    .SN(_17135_));
 HAxp5_ASAP7_75t_R _34962_ (.A(_18148_),
    .B(_17140_),
    .CON(_02261_),
    .SN(_00149_));
 HAxp5_ASAP7_75t_R _34963_ (.A(_18150_),
    .B(_18163_),
    .CON(_00159_),
    .SN(_00150_));
 HAxp5_ASAP7_75t_R _34964_ (.A(_18160_),
    .B(_18173_),
    .CON(_02262_),
    .SN(_00154_));
 HAxp5_ASAP7_75t_R _34965_ (.A(_18174_),
    .B(_17131_),
    .CON(_02263_),
    .SN(_17164_));
 HAxp5_ASAP7_75t_R _34966_ (.A(_17139_),
    .B(_17169_),
    .CON(_02264_),
    .SN(_00157_));
 HAxp5_ASAP7_75t_R _34967_ (.A(_18162_),
    .B(_18176_),
    .CON(_00167_),
    .SN(_00158_));
 HAxp5_ASAP7_75t_R _34968_ (.A(_17168_),
    .B(_17207_),
    .CON(_02265_),
    .SN(_00165_));
 HAxp5_ASAP7_75t_R _34969_ (.A(_18175_),
    .B(_18187_),
    .CON(_00173_),
    .SN(_00166_));
 HAxp5_ASAP7_75t_R _34970_ (.A(_18199_),
    .B(_18200_),
    .CON(_02266_),
    .SN(_17233_));
 HAxp5_ASAP7_75t_R _34971_ (.A(_17206_),
    .B(_18207_),
    .CON(_02267_),
    .SN(_00171_));
 HAxp5_ASAP7_75t_R _34972_ (.A(_18186_),
    .B(_18209_),
    .CON(_00179_),
    .SN(_00172_));
 HAxp5_ASAP7_75t_R _34973_ (.A(_18201_),
    .B(_18223_),
    .CON(_02268_),
    .SN(_17277_));
 HAxp5_ASAP7_75t_R _34974_ (.A(_18224_),
    .B(_18225_),
    .CON(_02269_),
    .SN(_00177_));
 HAxp5_ASAP7_75t_R _34975_ (.A(_18208_),
    .B(_18227_),
    .CON(_00186_),
    .SN(_00178_));
 HAxp5_ASAP7_75t_R _34976_ (.A(_18242_),
    .B(_17268_),
    .CON(_02270_),
    .SN(_00183_));
 HAxp5_ASAP7_75t_R _34977_ (.A(_18244_),
    .B(_17273_),
    .CON(_02271_),
    .SN(_17318_));
 HAxp5_ASAP7_75t_R _34978_ (.A(_17323_),
    .B(_18226_),
    .CON(_00195_),
    .SN(_00185_));
 HAxp5_ASAP7_75t_R _34979_ (.A(_18263_),
    .B(_18264_),
    .CON(_02272_),
    .SN(_00189_));
 HAxp5_ASAP7_75t_R _34980_ (.A(_18265_),
    .B(_17308_),
    .CON(_17408_),
    .SN(_00190_));
 HAxp5_ASAP7_75t_R _34981_ (.A(_18243_),
    .B(_18266_),
    .CON(_02273_),
    .SN(_00191_));
 HAxp5_ASAP7_75t_R _34982_ (.A(_18267_),
    .B(_17314_),
    .CON(_02274_),
    .SN(_17359_));
 HAxp5_ASAP7_75t_R _34983_ (.A(_17322_),
    .B(_17364_),
    .CON(_00200_),
    .SN(_00194_));
 HAxp5_ASAP7_75t_R _34984_ (.A(_17363_),
    .B(_17420_),
    .CON(_00204_),
    .SN(_00199_));
 HAxp5_ASAP7_75t_R _34985_ (.A(_17406_),
    .B(_18301_),
    .CON(_02275_),
    .SN(_17461_));
 HAxp5_ASAP7_75t_R _34986_ (.A(_17419_),
    .B(_18307_),
    .CON(_00208_),
    .SN(_00203_));
 HAxp5_ASAP7_75t_R _34987_ (.A(_18325_),
    .B(_18326_),
    .CON(_02276_),
    .SN(_00206_));
 HAxp5_ASAP7_75t_R _34988_ (.A(_18330_),
    .B(_18331_),
    .CON(_00211_),
    .SN(_00207_));
 HAxp5_ASAP7_75t_R _34989_ (.A(_18349_),
    .B(_18350_),
    .CON(_02277_),
    .SN(_00209_));
 HAxp5_ASAP7_75t_R _34990_ (.A(_18353_),
    .B(_18354_),
    .CON(_00214_),
    .SN(_00210_));
 HAxp5_ASAP7_75t_R _34991_ (.A(_18371_),
    .B(_18372_),
    .CON(_02278_),
    .SN(_00212_));
 HAxp5_ASAP7_75t_R _34992_ (.A(_18376_),
    .B(_18375_),
    .CON(_00217_),
    .SN(_00213_));
 HAxp5_ASAP7_75t_R _34993_ (.A(_18392_),
    .B(_18393_),
    .CON(_02279_),
    .SN(_00215_));
 HAxp5_ASAP7_75t_R _34994_ (.A(_18396_),
    .B(_18397_),
    .CON(_00220_),
    .SN(_00216_));
 HAxp5_ASAP7_75t_R _34995_ (.A(_18413_),
    .B(_18414_),
    .CON(_02280_),
    .SN(_00218_));
 HAxp5_ASAP7_75t_R _34996_ (.A(_18417_),
    .B(_18418_),
    .CON(_00223_),
    .SN(_00219_));
 HAxp5_ASAP7_75t_R _34997_ (.A(_18433_),
    .B(_18434_),
    .CON(_02281_),
    .SN(_00221_));
 HAxp5_ASAP7_75t_R _34998_ (.A(_18437_),
    .B(_18438_),
    .CON(_00226_),
    .SN(_00222_));
 HAxp5_ASAP7_75t_R _34999_ (.A(_18449_),
    .B(_18450_),
    .CON(_02282_),
    .SN(_00224_));
 HAxp5_ASAP7_75t_R _35000_ (.A(_18453_),
    .B(_18454_),
    .CON(_00229_),
    .SN(_00225_));
 HAxp5_ASAP7_75t_R _35001_ (.A(_18463_),
    .B(_18464_),
    .CON(_02283_),
    .SN(_00227_));
 HAxp5_ASAP7_75t_R _35002_ (.A(_18467_),
    .B(_18468_),
    .CON(_00232_),
    .SN(_00228_));
 HAxp5_ASAP7_75t_R _35003_ (.A(_18477_),
    .B(_18478_),
    .CON(_02284_),
    .SN(_00230_));
 HAxp5_ASAP7_75t_R _35004_ (.A(_18482_),
    .B(_18481_),
    .CON(_00235_),
    .SN(_00231_));
 HAxp5_ASAP7_75t_R _35005_ (.A(_18492_),
    .B(_18493_),
    .CON(_02285_),
    .SN(_00233_));
 HAxp5_ASAP7_75t_R _35006_ (.A(_18496_),
    .B(_18497_),
    .CON(_00238_),
    .SN(_00234_));
 HAxp5_ASAP7_75t_R _35007_ (.A(_18507_),
    .B(_18508_),
    .CON(_02286_),
    .SN(_00236_));
 HAxp5_ASAP7_75t_R _35008_ (.A(_18511_),
    .B(_18512_),
    .CON(_00241_),
    .SN(_00237_));
 HAxp5_ASAP7_75t_R _35009_ (.A(_18522_),
    .B(_18523_),
    .CON(_02287_),
    .SN(_00239_));
 HAxp5_ASAP7_75t_R _35010_ (.A(_18526_),
    .B(_18527_),
    .CON(_00244_),
    .SN(_00240_));
 HAxp5_ASAP7_75t_R _35011_ (.A(_18531_),
    .B(_18532_),
    .CON(_02288_),
    .SN(_00242_));
 HAxp5_ASAP7_75t_R _35012_ (.A(_18535_),
    .B(_18536_),
    .CON(_00247_),
    .SN(_00243_));
 HAxp5_ASAP7_75t_R _35013_ (.A(_18538_),
    .B(_18539_),
    .CON(_02289_),
    .SN(_00245_));
 HAxp5_ASAP7_75t_R _35014_ (.A(_18542_),
    .B(_18543_),
    .CON(_00253_),
    .SN(_00246_));
 HAxp5_ASAP7_75t_R _35015_ (.A(_17990_),
    .B(_17908_),
    .CON(_00256_),
    .SN(_00249_));
 HAxp5_ASAP7_75t_R _35016_ (.A(_18546_),
    .B(_17991_),
    .CON(_02290_),
    .SN(_00251_));
 HAxp5_ASAP7_75t_R _35017_ (.A(_18549_),
    .B(_18550_),
    .CON(_00259_),
    .SN(_00252_));
 HAxp5_ASAP7_75t_R _35018_ (.A(\cs_registers_i.pc_if_i[2] ),
    .B(_18551_),
    .CON(_00266_),
    .SN(_00264_));
 HAxp5_ASAP7_75t_R _35019_ (.A(_18552_),
    .B(_18553_),
    .CON(_02291_),
    .SN(_00268_));
 HAxp5_ASAP7_75t_R _35020_ (.A(_18554_),
    .B(_18555_),
    .CON(_00269_),
    .SN(_02292_));
 HAxp5_ASAP7_75t_R _35021_ (.A(_18556_),
    .B(_18553_),
    .CON(_02293_),
    .SN(_18557_));
 HAxp5_ASAP7_75t_R _35022_ (.A(_18558_),
    .B(_18559_),
    .CON(_00271_),
    .SN(_00270_));
 HAxp5_ASAP7_75t_R _35023_ (.A(_18560_),
    .B(_18552_),
    .CON(_02294_),
    .SN(_18561_));
 HAxp5_ASAP7_75t_R _35024_ (.A(_18562_),
    .B(_18563_),
    .CON(_00273_),
    .SN(_00272_));
 HAxp5_ASAP7_75t_R _35025_ (.A(_18564_),
    .B(_18565_),
    .CON(_02295_),
    .SN(_18566_));
 HAxp5_ASAP7_75t_R _35026_ (.A(_18567_),
    .B(_18568_),
    .CON(_00275_),
    .SN(_00274_));
 HAxp5_ASAP7_75t_R _35027_ (.A(_18569_),
    .B(_18570_),
    .CON(_02296_),
    .SN(_18571_));
 HAxp5_ASAP7_75t_R _35028_ (.A(_18572_),
    .B(_18573_),
    .CON(_00277_),
    .SN(_00276_));
 HAxp5_ASAP7_75t_R _35029_ (.A(_18574_),
    .B(_18575_),
    .CON(_02297_),
    .SN(_18576_));
 HAxp5_ASAP7_75t_R _35030_ (.A(_18577_),
    .B(_18578_),
    .CON(_00279_),
    .SN(_00278_));
 HAxp5_ASAP7_75t_R _35031_ (.A(_18579_),
    .B(_18580_),
    .CON(_02298_),
    .SN(_18581_));
 HAxp5_ASAP7_75t_R _35032_ (.A(_18582_),
    .B(_18583_),
    .CON(_00281_),
    .SN(_00280_));
 HAxp5_ASAP7_75t_R _35033_ (.A(_18584_),
    .B(_18585_),
    .CON(_02299_),
    .SN(_18586_));
 HAxp5_ASAP7_75t_R _35034_ (.A(_18587_),
    .B(_18588_),
    .CON(_00283_),
    .SN(_00282_));
 HAxp5_ASAP7_75t_R _35035_ (.A(_18589_),
    .B(_18590_),
    .CON(_02300_),
    .SN(_18591_));
 HAxp5_ASAP7_75t_R _35036_ (.A(_18592_),
    .B(_18593_),
    .CON(_00285_),
    .SN(_00284_));
 HAxp5_ASAP7_75t_R _35037_ (.A(_18594_),
    .B(_18595_),
    .CON(_02301_),
    .SN(_18596_));
 HAxp5_ASAP7_75t_R _35038_ (.A(_18597_),
    .B(_18598_),
    .CON(_00287_),
    .SN(_00286_));
 HAxp5_ASAP7_75t_R _35039_ (.A(_18599_),
    .B(_18600_),
    .CON(_02302_),
    .SN(_18601_));
 HAxp5_ASAP7_75t_R _35040_ (.A(_18602_),
    .B(_18603_),
    .CON(_00289_),
    .SN(_00288_));
 HAxp5_ASAP7_75t_R _35041_ (.A(_18604_),
    .B(_18605_),
    .CON(_02303_),
    .SN(_18606_));
 HAxp5_ASAP7_75t_R _35042_ (.A(_18607_),
    .B(_18608_),
    .CON(_00291_),
    .SN(_00290_));
 HAxp5_ASAP7_75t_R _35043_ (.A(_18609_),
    .B(_18610_),
    .CON(_02304_),
    .SN(_18611_));
 HAxp5_ASAP7_75t_R _35044_ (.A(_18612_),
    .B(_18613_),
    .CON(_02305_),
    .SN(_00292_));
 HAxp5_ASAP7_75t_R _35045_ (.A(_18614_),
    .B(_18615_),
    .CON(_00293_),
    .SN(_18616_));
 HAxp5_ASAP7_75t_R _35046_ (.A(_18617_),
    .B(_18618_),
    .CON(_02306_),
    .SN(_00294_));
 HAxp5_ASAP7_75t_R _35047_ (.A(_18619_),
    .B(_18620_),
    .CON(_00295_),
    .SN(_18621_));
 HAxp5_ASAP7_75t_R _35048_ (.A(_18622_),
    .B(_18623_),
    .CON(_02307_),
    .SN(_00296_));
 HAxp5_ASAP7_75t_R _35049_ (.A(_18624_),
    .B(_18625_),
    .CON(_00297_),
    .SN(_18626_));
 HAxp5_ASAP7_75t_R _35050_ (.A(_18627_),
    .B(_18628_),
    .CON(_02308_),
    .SN(_00298_));
 HAxp5_ASAP7_75t_R _35051_ (.A(_18629_),
    .B(_18630_),
    .CON(_00299_),
    .SN(_18631_));
 HAxp5_ASAP7_75t_R _35052_ (.A(_18632_),
    .B(_18633_),
    .CON(_02309_),
    .SN(_00300_));
 HAxp5_ASAP7_75t_R _35053_ (.A(_18634_),
    .B(_18635_),
    .CON(_00301_),
    .SN(_18636_));
 HAxp5_ASAP7_75t_R _35054_ (.A(_18637_),
    .B(_18638_),
    .CON(_02310_),
    .SN(_00302_));
 HAxp5_ASAP7_75t_R _35055_ (.A(_18639_),
    .B(_18640_),
    .CON(_00303_),
    .SN(_18641_));
 HAxp5_ASAP7_75t_R _35056_ (.A(_18642_),
    .B(_18643_),
    .CON(_02311_),
    .SN(_00304_));
 HAxp5_ASAP7_75t_R _35057_ (.A(_18644_),
    .B(_18645_),
    .CON(_00305_),
    .SN(_18646_));
 HAxp5_ASAP7_75t_R _35058_ (.A(_18647_),
    .B(_18648_),
    .CON(_02312_),
    .SN(_00306_));
 HAxp5_ASAP7_75t_R _35059_ (.A(_18649_),
    .B(_18650_),
    .CON(_00307_),
    .SN(_18651_));
 HAxp5_ASAP7_75t_R _35060_ (.A(_18652_),
    .B(_18653_),
    .CON(_02313_),
    .SN(_00308_));
 HAxp5_ASAP7_75t_R _35061_ (.A(_18654_),
    .B(_18655_),
    .CON(_00309_),
    .SN(_18656_));
 HAxp5_ASAP7_75t_R _35062_ (.A(_18657_),
    .B(_18658_),
    .CON(_02314_),
    .SN(_00310_));
 HAxp5_ASAP7_75t_R _35063_ (.A(_18659_),
    .B(_18660_),
    .CON(_00311_),
    .SN(_18661_));
 HAxp5_ASAP7_75t_R _35064_ (.A(_18662_),
    .B(_18663_),
    .CON(_02315_),
    .SN(_00312_));
 HAxp5_ASAP7_75t_R _35065_ (.A(_18664_),
    .B(_18665_),
    .CON(_00313_),
    .SN(_18666_));
 HAxp5_ASAP7_75t_R _35066_ (.A(_18667_),
    .B(_18668_),
    .CON(_02316_),
    .SN(_00314_));
 HAxp5_ASAP7_75t_R _35067_ (.A(_18669_),
    .B(_18670_),
    .CON(_00315_),
    .SN(_18671_));
 HAxp5_ASAP7_75t_R _35068_ (.A(_18672_),
    .B(_18673_),
    .CON(_02317_),
    .SN(_00316_));
 HAxp5_ASAP7_75t_R _35069_ (.A(_18674_),
    .B(_18675_),
    .CON(_00317_),
    .SN(_18676_));
 HAxp5_ASAP7_75t_R _35070_ (.A(_18677_),
    .B(_18678_),
    .CON(_02318_),
    .SN(_00318_));
 HAxp5_ASAP7_75t_R _35071_ (.A(_18679_),
    .B(_18680_),
    .CON(_00319_),
    .SN(_18681_));
 HAxp5_ASAP7_75t_R _35072_ (.A(_18682_),
    .B(_18683_),
    .CON(_02319_),
    .SN(_00320_));
 HAxp5_ASAP7_75t_R _35073_ (.A(_18684_),
    .B(_18685_),
    .CON(_00321_),
    .SN(_18686_));
 HAxp5_ASAP7_75t_R _35074_ (.A(_18687_),
    .B(_18688_),
    .CON(_02320_),
    .SN(_00322_));
 HAxp5_ASAP7_75t_R _35075_ (.A(_18689_),
    .B(_18690_),
    .CON(_00323_),
    .SN(_18691_));
 HAxp5_ASAP7_75t_R _35076_ (.A(_18692_),
    .B(_18693_),
    .CON(_02321_),
    .SN(_00324_));
 HAxp5_ASAP7_75t_R _35077_ (.A(_18694_),
    .B(_18695_),
    .CON(_00325_),
    .SN(_18696_));
 HAxp5_ASAP7_75t_R _35078_ (.A(_18697_),
    .B(_18698_),
    .CON(_02322_),
    .SN(_00326_));
 HAxp5_ASAP7_75t_R _35079_ (.A(_18699_),
    .B(_18700_),
    .CON(_00327_),
    .SN(_18701_));
 HAxp5_ASAP7_75t_R _35080_ (.A(_18702_),
    .B(_18703_),
    .CON(_02323_),
    .SN(_00328_));
 HAxp5_ASAP7_75t_R _35081_ (.A(_18704_),
    .B(_18705_),
    .CON(_00329_),
    .SN(_18706_));
 HAxp5_ASAP7_75t_R _35082_ (.A(_18707_),
    .B(_18708_),
    .CON(_02324_),
    .SN(_02325_));
 HAxp5_ASAP7_75t_R _35083_ (.A(\alu_adder_result_ex[1] ),
    .B(\alu_adder_result_ex[0] ),
    .CON(_00336_),
    .SN(_00338_));
 HAxp5_ASAP7_75t_R _35084_ (.A(\alu_adder_result_ex[1] ),
    .B(\alu_adder_result_ex[0] ),
    .CON(_02326_),
    .SN(_18709_));
 HAxp5_ASAP7_75t_R _35085_ (.A(\alu_adder_result_ex[1] ),
    .B(_16999_),
    .CON(_00337_),
    .SN(_18710_));
 HAxp5_ASAP7_75t_R _35086_ (.A(\alu_adder_result_ex[1] ),
    .B(_16999_),
    .CON(_02327_),
    .SN(_18711_));
 HAxp5_ASAP7_75t_R _35087_ (.A(_18712_),
    .B(\alu_adder_result_ex[0] ),
    .CON(_00335_),
    .SN(_18713_));
 HAxp5_ASAP7_75t_R _35088_ (.A(_18712_),
    .B(\alu_adder_result_ex[0] ),
    .CON(_02328_),
    .SN(_18714_));
 HAxp5_ASAP7_75t_R _35089_ (.A(_18712_),
    .B(_16999_),
    .CON(_18708_),
    .SN(_18715_));
 HAxp5_ASAP7_75t_R _35090_ (.A(_18716_),
    .B(_18717_),
    .CON(_02329_),
    .SN(_02330_));
 HAxp5_ASAP7_75t_R _35091_ (.A(_18719_),
    .B(_18718_),
    .CON(_02331_),
    .SN(_02332_));
 DFFASRHQNx1_ASAP7_75t_R _35092_ (.CLK(clknet_leaf_19_clk),
    .D(_02333_),
    .QN(_02195_),
    .RESETN(net277),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R _35093_ (.CLK(clknet_leaf_19_clk),
    .D(_02334_),
    .QN(_02194_),
    .RESETN(net278),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R _35094_ (.CLK(clknet_leaf_17_clk),
    .D(_02335_),
    .QN(_00753_),
    .RESETN(net279),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R _35095_ (.CLK(clknet_leaf_17_clk),
    .D(_02336_),
    .QN(_02193_),
    .RESETN(net280),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R _35096_ (.CLK(clknet_leaf_17_clk),
    .D(_02337_),
    .QN(_02192_),
    .RESETN(net52),
    .SETN(net281));
 DFFASRHQNx1_ASAP7_75t_R _35097_ (.CLK(clknet_leaf_0_clk),
    .D(_02338_),
    .QN(_02191_),
    .RESETN(net282),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R _35098_ (.CLK(clknet_leaf_0_clk),
    .D(_02339_),
    .QN(_02196_),
    .RESETN(net283),
    .SETN(net36));
 BUFx16f_ASAP7_75t_R clkbuf_regs_0_core_clock (.A(clk_i),
    .Y(delaynet_0_core_clock));
 TIEHIx1_ASAP7_75t_R _35092__256 (.H(net277));
 BUFx2_ASAP7_75t_R _35101_ (.A(net271),
    .Y(alert_major_o));
 BUFx2_ASAP7_75t_R _35102_ (.A(net272),
    .Y(alert_minor_o));
 BUFx2_ASAP7_75t_R _35103_ (.A(net273),
    .Y(data_addr_o[0]));
 BUFx2_ASAP7_75t_R _35104_ (.A(net274),
    .Y(data_addr_o[1]));
 BUFx3_ASAP7_75t_R _35105_ (.A(\alu_adder_result_ex[2] ),
    .Y(net192));
 BUFx3_ASAP7_75t_R _35106_ (.A(\alu_adder_result_ex[3] ),
    .Y(net195));
 BUFx3_ASAP7_75t_R _35107_ (.A(\alu_adder_result_ex[4] ),
    .Y(net196));
 BUFx3_ASAP7_75t_R _35108_ (.A(\alu_adder_result_ex[5] ),
    .Y(net197));
 BUFx3_ASAP7_75t_R _35109_ (.A(\alu_adder_result_ex[6] ),
    .Y(net198));
 BUFx3_ASAP7_75t_R _35110_ (.A(\alu_adder_result_ex[7] ),
    .Y(net199));
 BUFx3_ASAP7_75t_R _35111_ (.A(\alu_adder_result_ex[8] ),
    .Y(net200));
 BUFx3_ASAP7_75t_R _35112_ (.A(\alu_adder_result_ex[9] ),
    .Y(net201));
 BUFx3_ASAP7_75t_R _35113_ (.A(\alu_adder_result_ex[10] ),
    .Y(net172));
 BUFx3_ASAP7_75t_R _35114_ (.A(\alu_adder_result_ex[11] ),
    .Y(net173));
 BUFx3_ASAP7_75t_R _35115_ (.A(\alu_adder_result_ex[12] ),
    .Y(net174));
 BUFx3_ASAP7_75t_R _35116_ (.A(\alu_adder_result_ex[13] ),
    .Y(net175));
 BUFx3_ASAP7_75t_R _35117_ (.A(\alu_adder_result_ex[14] ),
    .Y(net176));
 BUFx3_ASAP7_75t_R _35118_ (.A(\alu_adder_result_ex[15] ),
    .Y(net177));
 BUFx3_ASAP7_75t_R _35119_ (.A(\alu_adder_result_ex[16] ),
    .Y(net178));
 BUFx3_ASAP7_75t_R _35120_ (.A(\alu_adder_result_ex[17] ),
    .Y(net179));
 BUFx3_ASAP7_75t_R _35121_ (.A(\alu_adder_result_ex[18] ),
    .Y(net180));
 BUFx3_ASAP7_75t_R _35122_ (.A(\alu_adder_result_ex[19] ),
    .Y(net181));
 BUFx3_ASAP7_75t_R _35123_ (.A(\alu_adder_result_ex[20] ),
    .Y(net182));
 BUFx3_ASAP7_75t_R _35124_ (.A(\alu_adder_result_ex[21] ),
    .Y(net183));
 BUFx3_ASAP7_75t_R _35125_ (.A(\alu_adder_result_ex[22] ),
    .Y(net184));
 BUFx3_ASAP7_75t_R _35126_ (.A(\alu_adder_result_ex[23] ),
    .Y(net185));
 BUFx3_ASAP7_75t_R _35127_ (.A(\alu_adder_result_ex[24] ),
    .Y(net186));
 BUFx3_ASAP7_75t_R _35128_ (.A(\alu_adder_result_ex[25] ),
    .Y(net187));
 BUFx3_ASAP7_75t_R _35129_ (.A(\alu_adder_result_ex[26] ),
    .Y(net188));
 BUFx3_ASAP7_75t_R _35130_ (.A(\alu_adder_result_ex[27] ),
    .Y(net189));
 BUFx3_ASAP7_75t_R _35131_ (.A(\alu_adder_result_ex[28] ),
    .Y(net190));
 BUFx3_ASAP7_75t_R _35132_ (.A(\alu_adder_result_ex[29] ),
    .Y(net191));
 BUFx3_ASAP7_75t_R _35133_ (.A(\alu_adder_result_ex[30] ),
    .Y(net193));
 BUFx3_ASAP7_75t_R _35134_ (.A(net1960),
    .Y(net194));
 BUFx2_ASAP7_75t_R _35135_ (.A(net275),
    .Y(instr_addr_o[0]));
 BUFx2_ASAP7_75t_R _35136_ (.A(net276),
    .Y(instr_addr_o[1]));
 DFFASRHQNx1_ASAP7_75t_R \core_busy_q$_DFF_PN0_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(core_busy_d),
    .QN(_02190_),
    .RESETN(net284),
    .SETN(net1963));
 DLLx1_ASAP7_75t_R \core_clock_gate_i.en_latch$_DLATCH_N_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_00006_),
    .Q(\core_clock_gate_i.en_latch ));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcountinhibit_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02340_),
    .QN(_01396_),
    .RESETN(net285),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcountinhibit_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02341_),
    .QN(_02189_),
    .RESETN(net286),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02342_),
    .QN(_00747_),
    .RESETN(net287),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02343_),
    .QN(_02188_),
    .RESETN(net288),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02344_),
    .QN(_02187_),
    .RESETN(net289),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02345_),
    .QN(_02186_),
    .RESETN(net290),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02346_),
    .QN(_02185_),
    .RESETN(net291),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02347_),
    .QN(_02184_),
    .RESETN(net292),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02348_),
    .QN(_02183_),
    .RESETN(net293),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02349_),
    .QN(_02182_),
    .RESETN(net294),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02350_),
    .QN(_02181_),
    .RESETN(net295),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02351_),
    .QN(_02180_),
    .RESETN(net296),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02352_),
    .QN(_02179_),
    .RESETN(net297),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02353_),
    .QN(_02178_),
    .RESETN(net298),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02354_),
    .QN(_02177_),
    .RESETN(net299),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02355_),
    .QN(_02176_),
    .RESETN(net300),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02356_),
    .QN(_02175_),
    .RESETN(net301),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02357_),
    .QN(_02174_),
    .RESETN(net302),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02358_),
    .QN(_02173_),
    .RESETN(net303),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02359_),
    .QN(_02172_),
    .RESETN(net304),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02360_),
    .QN(_02171_),
    .RESETN(net305),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02361_),
    .QN(_02170_),
    .RESETN(net306),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02362_),
    .QN(_02169_),
    .RESETN(net307),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02363_),
    .QN(_02168_),
    .RESETN(net308),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02364_),
    .QN(_02167_),
    .RESETN(net309),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02365_),
    .QN(_02166_),
    .RESETN(net310),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02366_),
    .QN(_02165_),
    .RESETN(net311),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[32]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02367_),
    .QN(_02164_),
    .RESETN(net312),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[33]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02368_),
    .QN(_02163_),
    .RESETN(net313),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[34]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02369_),
    .QN(_02162_),
    .RESETN(net314),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[35]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02370_),
    .QN(_02161_),
    .RESETN(net315),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[36]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02371_),
    .QN(_02160_),
    .RESETN(net316),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[37]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02372_),
    .QN(_02159_),
    .RESETN(net317),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[38]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02373_),
    .QN(_02158_),
    .RESETN(net318),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[39]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02374_),
    .QN(_02157_),
    .RESETN(net319),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02375_),
    .QN(_02156_),
    .RESETN(net320),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[40]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02376_),
    .QN(_02155_),
    .RESETN(net321),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[41]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02377_),
    .QN(_02154_),
    .RESETN(net322),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[42]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02378_),
    .QN(_02153_),
    .RESETN(net323),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[43]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02379_),
    .QN(_02152_),
    .RESETN(net324),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[44]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02380_),
    .QN(_02151_),
    .RESETN(net325),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[45]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02381_),
    .QN(_02150_),
    .RESETN(net326),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[46]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02382_),
    .QN(_02149_),
    .RESETN(net327),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[47]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02383_),
    .QN(_02148_),
    .RESETN(net328),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[48]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02384_),
    .QN(_02147_),
    .RESETN(net329),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[49]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02385_),
    .QN(_02146_),
    .RESETN(net330),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02386_),
    .QN(_02145_),
    .RESETN(net331),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[50]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02387_),
    .QN(_02144_),
    .RESETN(net332),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[51]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02388_),
    .QN(_02143_),
    .RESETN(net333),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[52]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02389_),
    .QN(_02142_),
    .RESETN(net334),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[53]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02390_),
    .QN(_02141_),
    .RESETN(net335),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[54]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02391_),
    .QN(_02140_),
    .RESETN(net336),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[55]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02392_),
    .QN(_02139_),
    .RESETN(net337),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[56]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02393_),
    .QN(_02138_),
    .RESETN(net338),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[57]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02394_),
    .QN(_02137_),
    .RESETN(net339),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[58]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02395_),
    .QN(_02136_),
    .RESETN(net340),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[59]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02396_),
    .QN(_02135_),
    .RESETN(net341),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02397_),
    .QN(_02134_),
    .RESETN(net342),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[60]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02398_),
    .QN(_02133_),
    .RESETN(net343),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[61]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02399_),
    .QN(_02132_),
    .RESETN(net344),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[62]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02400_),
    .QN(_02131_),
    .RESETN(net345),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[63]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02401_),
    .QN(_02130_),
    .RESETN(net346),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02402_),
    .QN(_02129_),
    .RESETN(net347),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02403_),
    .QN(_02128_),
    .RESETN(net348),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02404_),
    .QN(_02127_),
    .RESETN(net349),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02405_),
    .QN(_02126_),
    .RESETN(net350),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02406_),
    .QN(_00748_),
    .RESETN(net351),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02407_),
    .QN(_02125_),
    .RESETN(net352),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02408_),
    .QN(_02124_),
    .RESETN(net353),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02409_),
    .QN(_02123_),
    .RESETN(net354),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02410_),
    .QN(_02122_),
    .RESETN(net355),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02411_),
    .QN(_02121_),
    .RESETN(net356),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02412_),
    .QN(_02120_),
    .RESETN(net357),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02413_),
    .QN(_02119_),
    .RESETN(net358),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02414_),
    .QN(_02118_),
    .RESETN(net359),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02415_),
    .QN(_02117_),
    .RESETN(net360),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02416_),
    .QN(_02116_),
    .RESETN(net361),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02417_),
    .QN(_02115_),
    .RESETN(net362),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02418_),
    .QN(_02114_),
    .RESETN(net363),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02419_),
    .QN(_02113_),
    .RESETN(net364),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02420_),
    .QN(_02112_),
    .RESETN(net365),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02421_),
    .QN(_02111_),
    .RESETN(net366),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02422_),
    .QN(_02110_),
    .RESETN(net367),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02423_),
    .QN(_02109_),
    .RESETN(net368),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02424_),
    .QN(_02108_),
    .RESETN(net369),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02425_),
    .QN(_02107_),
    .RESETN(net370),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02426_),
    .QN(_02106_),
    .RESETN(net371),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02427_),
    .QN(_02105_),
    .RESETN(net372),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02428_),
    .QN(_02104_),
    .RESETN(net373),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02429_),
    .QN(_02103_),
    .RESETN(net374),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02430_),
    .QN(_02102_),
    .RESETN(net375),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[32]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02431_),
    .QN(_02101_),
    .RESETN(net376),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[33]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02432_),
    .QN(_02100_),
    .RESETN(net377),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[34]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02433_),
    .QN(_02099_),
    .RESETN(net378),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[35]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02434_),
    .QN(_02098_),
    .RESETN(net379),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[36]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02435_),
    .QN(_02097_),
    .RESETN(net380),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[37]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02436_),
    .QN(_02096_),
    .RESETN(net381),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[38]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02437_),
    .QN(_02095_),
    .RESETN(net382),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[39]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02438_),
    .QN(_02094_),
    .RESETN(net383),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02439_),
    .QN(_02093_),
    .RESETN(net384),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[40]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02440_),
    .QN(_02092_),
    .RESETN(net385),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[41]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02441_),
    .QN(_02091_),
    .RESETN(net386),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[42]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02442_),
    .QN(_02090_),
    .RESETN(net387),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[43]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02443_),
    .QN(_02089_),
    .RESETN(net388),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[44]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02444_),
    .QN(_02088_),
    .RESETN(net389),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[45]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02445_),
    .QN(_02087_),
    .RESETN(net390),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[46]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02446_),
    .QN(_02086_),
    .RESETN(net391),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[47]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02447_),
    .QN(_02085_),
    .RESETN(net392),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[48]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02448_),
    .QN(_02084_),
    .RESETN(net393),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[49]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02449_),
    .QN(_02083_),
    .RESETN(net394),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02450_),
    .QN(_02082_),
    .RESETN(net395),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[50]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02451_),
    .QN(_02081_),
    .RESETN(net396),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[51]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02452_),
    .QN(_02080_),
    .RESETN(net397),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[52]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02453_),
    .QN(_02079_),
    .RESETN(net398),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[53]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02454_),
    .QN(_02078_),
    .RESETN(net399),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[54]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02455_),
    .QN(_02077_),
    .RESETN(net400),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[55]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02456_),
    .QN(_02076_),
    .RESETN(net401),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[56]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02457_),
    .QN(_02075_),
    .RESETN(net402),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[57]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02458_),
    .QN(_02074_),
    .RESETN(net403),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[58]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02459_),
    .QN(_02073_),
    .RESETN(net404),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[59]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02460_),
    .QN(_02072_),
    .RESETN(net405),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02461_),
    .QN(_02071_),
    .RESETN(net406),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[60]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02462_),
    .QN(_02070_),
    .RESETN(net407),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[61]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02463_),
    .QN(_02069_),
    .RESETN(net408),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[62]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02464_),
    .QN(_02068_),
    .RESETN(net409),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[63]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02465_),
    .QN(_02067_),
    .RESETN(net410),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02466_),
    .QN(_02066_),
    .RESETN(net411),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02467_),
    .QN(_02065_),
    .RESETN(net412),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02468_),
    .QN(_02064_),
    .RESETN(net413),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_02469_),
    .QN(_02063_),
    .RESETN(net414),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.priv_mode_id_o[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .D(_02470_),
    .QN(_02062_),
    .RESETN(net51),
    .SETN(net415));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.priv_mode_id_o[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .D(_02471_),
    .QN(_18080_),
    .RESETN(net51),
    .SETN(net416));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_1_clk),
    .D(_02472_),
    .QN(_02061_),
    .RESETN(net51),
    .SETN(net417));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02473_),
    .QN(_02060_),
    .RESETN(net418),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02474_),
    .QN(_02059_),
    .RESETN(net419),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02475_),
    .QN(_02058_),
    .RESETN(net420),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02476_),
    .QN(_02057_),
    .RESETN(net421),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_1_clk),
    .D(_02477_),
    .QN(_02056_),
    .RESETN(net51),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02478_),
    .QN(_01398_),
    .RESETN(net423),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02479_),
    .QN(_02055_),
    .RESETN(net424),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02480_),
    .QN(_02054_),
    .RESETN(net425),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02481_),
    .QN(_02053_),
    .RESETN(net426),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02482_),
    .QN(_02052_),
    .RESETN(net427),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02483_),
    .QN(_02051_),
    .RESETN(net428),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02484_),
    .QN(_02050_),
    .RESETN(net429),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02485_),
    .QN(_02049_),
    .RESETN(net430),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02486_),
    .QN(_02048_),
    .RESETN(net431),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02487_),
    .QN(_02047_),
    .RESETN(net432),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02488_),
    .QN(_02046_),
    .RESETN(net433),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02489_),
    .QN(_02045_),
    .RESETN(net434),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02490_),
    .QN(_02044_),
    .RESETN(net435),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02491_),
    .QN(_02043_),
    .RESETN(net436),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02492_),
    .QN(_00749_),
    .RESETN(net437),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02493_),
    .QN(_02042_),
    .RESETN(net438),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02494_),
    .QN(_02041_),
    .RESETN(net439),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02495_),
    .QN(_02040_),
    .RESETN(net440),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02496_),
    .QN(_02039_),
    .RESETN(net441),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02497_),
    .QN(_02038_),
    .RESETN(net442),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02498_),
    .QN(_02037_),
    .RESETN(net443),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02499_),
    .QN(_02036_),
    .RESETN(net444),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02500_),
    .QN(_02035_),
    .RESETN(net445),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02501_),
    .QN(_02034_),
    .RESETN(net446),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02502_),
    .QN(_02033_),
    .RESETN(net447),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02503_),
    .QN(_02032_),
    .RESETN(net448),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02504_),
    .QN(_02031_),
    .RESETN(net449),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02505_),
    .QN(_02030_),
    .RESETN(net450),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02506_),
    .QN(_01399_),
    .RESETN(net451),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02507_),
    .QN(_01400_),
    .RESETN(net452),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02508_),
    .QN(_01401_),
    .RESETN(net453),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02509_),
    .QN(_01402_),
    .RESETN(net454),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02510_),
    .QN(_02029_),
    .RESETN(net455),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02511_),
    .QN(_02028_),
    .RESETN(net456),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02512_),
    .QN(_02027_),
    .RESETN(net457),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02513_),
    .QN(_02026_),
    .RESETN(net458),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02514_),
    .QN(_02025_),
    .RESETN(net459),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02515_),
    .QN(_02024_),
    .RESETN(net460),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02516_),
    .QN(_02023_),
    .RESETN(net461),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02517_),
    .QN(_02022_),
    .RESETN(net462),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02518_),
    .QN(_02021_),
    .RESETN(net463),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02519_),
    .QN(_02020_),
    .RESETN(net464),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02520_),
    .QN(_02019_),
    .RESETN(net465),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02521_),
    .QN(_02018_),
    .RESETN(net466),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02522_),
    .QN(_02017_),
    .RESETN(net467),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02523_),
    .QN(_02016_),
    .RESETN(net468),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02524_),
    .QN(_02015_),
    .RESETN(net469),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02525_),
    .QN(_02014_),
    .RESETN(net470),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02526_),
    .QN(_02013_),
    .RESETN(net471),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02527_),
    .QN(_02012_),
    .RESETN(net472),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02528_),
    .QN(_02011_),
    .RESETN(net473),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02529_),
    .QN(_02010_),
    .RESETN(net474),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02530_),
    .QN(_02009_),
    .RESETN(net475),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02531_),
    .QN(_02008_),
    .RESETN(net476),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02532_),
    .QN(_02007_),
    .RESETN(net477),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02533_),
    .QN(_02006_),
    .RESETN(net478),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02534_),
    .QN(_02005_),
    .RESETN(net479),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02535_),
    .QN(_02004_),
    .RESETN(net480),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02536_),
    .QN(_02003_),
    .RESETN(net481),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02537_),
    .QN(_02002_),
    .RESETN(net482),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02538_),
    .QN(_02001_),
    .RESETN(net483),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02539_),
    .QN(_02000_),
    .RESETN(net484),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02540_),
    .QN(_01999_),
    .RESETN(net485),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02541_),
    .QN(_01998_),
    .RESETN(net486),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02542_),
    .QN(_01997_),
    .RESETN(net487),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02543_),
    .QN(_01996_),
    .RESETN(net488),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02544_),
    .QN(_01995_),
    .RESETN(net489),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02545_),
    .QN(_01994_),
    .RESETN(net490),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02546_),
    .QN(_01993_),
    .RESETN(net491),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02547_),
    .QN(_01992_),
    .RESETN(net492),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02548_),
    .QN(_01991_),
    .RESETN(net493),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02549_),
    .QN(_01990_),
    .RESETN(net494),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02550_),
    .QN(_01989_),
    .RESETN(net495),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02551_),
    .QN(_01988_),
    .RESETN(net496),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02552_),
    .QN(_01987_),
    .RESETN(net497),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02553_),
    .QN(_01986_),
    .RESETN(net498),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02554_),
    .QN(_01985_),
    .RESETN(net499),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02555_),
    .QN(_01984_),
    .RESETN(net500),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02556_),
    .QN(_01983_),
    .RESETN(net501),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02557_),
    .QN(_01982_),
    .RESETN(net502),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02558_),
    .QN(_01981_),
    .RESETN(net503),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02559_),
    .QN(_01980_),
    .RESETN(net504),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02560_),
    .QN(_01979_),
    .RESETN(net505),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02561_),
    .QN(_01978_),
    .RESETN(net506),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02562_),
    .QN(_01977_),
    .RESETN(net507),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02563_),
    .QN(_01976_),
    .RESETN(net508),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02564_),
    .QN(_01975_),
    .RESETN(net509),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02565_),
    .QN(_01974_),
    .RESETN(net510),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02566_),
    .QN(_01973_),
    .RESETN(net511),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02567_),
    .QN(_01972_),
    .RESETN(net512),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02568_),
    .QN(_01971_),
    .RESETN(net513),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02569_),
    .QN(_01970_),
    .RESETN(net514),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02570_),
    .QN(_01969_),
    .RESETN(net515),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02571_),
    .QN(_01968_),
    .RESETN(net516),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02572_),
    .QN(_01967_),
    .RESETN(net517),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02573_),
    .QN(_01966_),
    .RESETN(net518),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02574_),
    .QN(_01965_),
    .RESETN(net519),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02575_),
    .QN(_01964_),
    .RESETN(net520),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02576_),
    .QN(_01963_),
    .RESETN(net521),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02577_),
    .QN(_01962_),
    .RESETN(net522),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02578_),
    .QN(_01961_),
    .RESETN(net523),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02579_),
    .QN(_01960_),
    .RESETN(net524),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02580_),
    .QN(_01959_),
    .RESETN(net525),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02581_),
    .QN(_01958_),
    .RESETN(net526),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02582_),
    .QN(_01957_),
    .RESETN(net527),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02583_),
    .QN(_01956_),
    .RESETN(net528),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02584_),
    .QN(_01955_),
    .RESETN(net529),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02585_),
    .QN(_01954_),
    .RESETN(net530),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02586_),
    .QN(_01953_),
    .RESETN(net531),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02587_),
    .QN(_01952_),
    .RESETN(net532),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02588_),
    .QN(_01951_),
    .RESETN(net533),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02589_),
    .QN(_01950_),
    .RESETN(net534),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02590_),
    .QN(_01949_),
    .RESETN(net535),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02591_),
    .QN(_01948_),
    .RESETN(net536),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02592_),
    .QN(_01947_),
    .RESETN(net537),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02593_),
    .QN(_01946_),
    .RESETN(net538),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02594_),
    .QN(_01945_),
    .RESETN(net539),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02595_),
    .QN(_01944_),
    .RESETN(net540),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02596_),
    .QN(_01943_),
    .RESETN(net541),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02597_),
    .QN(_01942_),
    .RESETN(net542),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02598_),
    .QN(_01941_),
    .RESETN(net543),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02599_),
    .QN(_01940_),
    .RESETN(net544),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02600_),
    .QN(_01939_),
    .RESETN(net545),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02601_),
    .QN(_01938_),
    .RESETN(net546),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02602_),
    .QN(_01937_),
    .RESETN(net547),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02603_),
    .QN(_01936_),
    .RESETN(net548),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02604_),
    .QN(_01935_),
    .RESETN(net549),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02605_),
    .QN(_01934_),
    .RESETN(net550),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02606_),
    .QN(_01933_),
    .RESETN(net551),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02607_),
    .QN(_01932_),
    .RESETN(net552),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02608_),
    .QN(_01931_),
    .RESETN(net553),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02609_),
    .QN(_01930_),
    .RESETN(net554),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02610_),
    .QN(_01929_),
    .RESETN(net555),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02611_),
    .QN(_01928_),
    .RESETN(net556),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02612_),
    .QN(_01927_),
    .RESETN(net557),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02613_),
    .QN(_01926_),
    .RESETN(net558),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02614_),
    .QN(_01925_),
    .RESETN(net559),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02615_),
    .QN(_01924_),
    .RESETN(net560),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02616_),
    .QN(_01923_),
    .RESETN(net561),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02617_),
    .QN(_01922_),
    .RESETN(net562),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02618_),
    .QN(_01921_),
    .RESETN(net563),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02619_),
    .QN(_01920_),
    .RESETN(net564),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02620_),
    .QN(_01919_),
    .RESETN(net565),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02621_),
    .QN(_01918_),
    .RESETN(net566),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02622_),
    .QN(_01917_),
    .RESETN(net567),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02623_),
    .QN(_01916_),
    .RESETN(net568),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02624_),
    .QN(_01915_),
    .RESETN(net569),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02625_),
    .QN(_01914_),
    .RESETN(net570),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02626_),
    .QN(_01913_),
    .RESETN(net571),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02627_),
    .QN(_01912_),
    .RESETN(net572),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02628_),
    .QN(_01911_),
    .RESETN(net573),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02629_),
    .QN(_01910_),
    .RESETN(net574),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02630_),
    .QN(_01909_),
    .RESETN(net575),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02631_),
    .QN(_01908_),
    .RESETN(net576),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02632_),
    .QN(_01907_),
    .RESETN(net577),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02633_),
    .QN(_01906_),
    .RESETN(net578),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02634_),
    .QN(_01905_),
    .RESETN(net579),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02635_),
    .QN(_01904_),
    .RESETN(net580),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02636_),
    .QN(_01903_),
    .RESETN(net581),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02637_),
    .QN(_01902_),
    .RESETN(net582),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02638_),
    .QN(_01901_),
    .RESETN(net583),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02639_),
    .QN(_01900_),
    .RESETN(net584),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02640_),
    .QN(_01899_),
    .RESETN(net585),
    .SETN(net48));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02641_),
    .QN(_01898_),
    .RESETN(net586),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02642_),
    .QN(_01897_),
    .RESETN(net587),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02643_),
    .QN(_01896_),
    .RESETN(net588),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02644_),
    .QN(_01895_),
    .RESETN(net589),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02645_),
    .QN(_01894_),
    .RESETN(net590),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02646_),
    .QN(_01893_),
    .RESETN(net591),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02647_),
    .QN(_01892_),
    .RESETN(net592),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02648_),
    .QN(_01891_),
    .RESETN(net593),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02649_),
    .QN(_01890_),
    .RESETN(net594),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02650_),
    .QN(_01889_),
    .RESETN(net595),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02651_),
    .QN(_01888_),
    .RESETN(net596),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02652_),
    .QN(_01887_),
    .RESETN(net597),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02653_),
    .QN(_01886_),
    .RESETN(net598),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02654_),
    .QN(_01885_),
    .RESETN(net599),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02655_),
    .QN(_01884_),
    .RESETN(net600),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02656_),
    .QN(_01883_),
    .RESETN(net601),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02657_),
    .QN(_01882_),
    .RESETN(net602),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02658_),
    .QN(_01881_),
    .RESETN(net603),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02659_),
    .QN(_01880_),
    .RESETN(net604),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02660_),
    .QN(_01879_),
    .RESETN(net605),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02661_),
    .QN(_01878_),
    .RESETN(net606),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02662_),
    .QN(_01877_),
    .RESETN(net607),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_02663_),
    .QN(_01876_),
    .RESETN(net608),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_02664_),
    .QN(_01875_),
    .RESETN(net609),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02665_),
    .QN(_01874_),
    .RESETN(net610),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02666_),
    .QN(_01873_),
    .RESETN(net611),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02667_),
    .QN(_01872_),
    .RESETN(net612),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02668_),
    .QN(_01871_),
    .RESETN(net613),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02669_),
    .QN(_01870_),
    .RESETN(net614),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02670_),
    .QN(_01869_),
    .RESETN(net615),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rd_data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02671_),
    .QN(_01868_),
    .RESETN(net616),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02672_),
    .QN(_01867_),
    .RESETN(net617),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rd_data_o[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .D(_02673_),
    .QN(_01866_),
    .RESETN(net51),
    .SETN(net618));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02674_),
    .QN(_01865_),
    .RESETN(net619),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02675_),
    .QN(_01864_),
    .RESETN(net620),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02676_),
    .QN(_01863_),
    .RESETN(net621),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02677_),
    .QN(_01862_),
    .RESETN(net622),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02678_),
    .QN(_01861_),
    .RESETN(net623),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02679_),
    .QN(_01860_),
    .RESETN(net624),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02680_),
    .QN(_01859_),
    .RESETN(net625),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02681_),
    .QN(_01858_),
    .RESETN(net626),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02682_),
    .QN(_01857_),
    .RESETN(net627),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02683_),
    .QN(_01856_),
    .RESETN(net628),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02684_),
    .QN(_01855_),
    .RESETN(net629),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02685_),
    .QN(_01854_),
    .RESETN(net630),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02686_),
    .QN(_01853_),
    .RESETN(net631),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02687_),
    .QN(_01852_),
    .RESETN(net632),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02688_),
    .QN(_01851_),
    .RESETN(net633),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02689_),
    .QN(_01850_),
    .RESETN(net634),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02690_),
    .QN(_01849_),
    .RESETN(net635),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02691_),
    .QN(_01848_),
    .RESETN(net636),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02692_),
    .QN(_01847_),
    .RESETN(net637),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02693_),
    .QN(_01846_),
    .RESETN(net638),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02694_),
    .QN(_01845_),
    .RESETN(net639),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02695_),
    .QN(_01844_),
    .RESETN(net640),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02696_),
    .QN(_01843_),
    .RESETN(net641),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02697_),
    .QN(_01842_),
    .RESETN(net642),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02698_),
    .QN(_01841_),
    .RESETN(net643),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02699_),
    .QN(_01840_),
    .RESETN(net644),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02700_),
    .QN(_01839_),
    .RESETN(net645),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02701_),
    .QN(_01838_),
    .RESETN(net646),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02702_),
    .QN(_01837_),
    .RESETN(net647),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02703_),
    .QN(_01836_),
    .RESETN(net648),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02704_),
    .QN(_01835_),
    .RESETN(net649),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02705_),
    .QN(_01834_),
    .RESETN(net650),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02706_),
    .QN(_01833_),
    .RESETN(net651),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02707_),
    .QN(_01832_),
    .RESETN(net652),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_9_clk),
    .D(_02708_),
    .QN(_00331_),
    .RESETN(net653),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .D(_02709_),
    .QN(_00332_),
    .RESETN(net654),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[4]$_DFFE_PN1N_  (.CLK(clknet_leaf_9_clk),
    .D(_02710_),
    .QN(_00333_),
    .RESETN(net51),
    .SETN(net655));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_9_clk),
    .D(_02711_),
    .QN(_00759_),
    .RESETN(net656),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02712_),
    .QN(_01831_),
    .RESETN(net657),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02713_),
    .QN(_01830_),
    .RESETN(net658),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02714_),
    .QN(_01829_),
    .RESETN(net659),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02715_),
    .QN(_01828_),
    .RESETN(net660),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02716_),
    .QN(_01827_),
    .RESETN(net661),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02717_),
    .QN(_01826_),
    .RESETN(net662),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02718_),
    .QN(_01825_),
    .RESETN(net663),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02719_),
    .QN(_01824_),
    .RESETN(net664),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02720_),
    .QN(_01823_),
    .RESETN(net665),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_02721_),
    .QN(_01822_),
    .RESETN(net666),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02722_),
    .QN(_01821_),
    .RESETN(net667),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02723_),
    .QN(_01820_),
    .RESETN(net668),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02724_),
    .QN(_01819_),
    .RESETN(net669),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02725_),
    .QN(_01818_),
    .RESETN(net670),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02726_),
    .QN(_01817_),
    .RESETN(net671),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02727_),
    .QN(_01816_),
    .RESETN(net672),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02728_),
    .QN(_01815_),
    .RESETN(net673),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02729_),
    .QN(_01814_),
    .RESETN(net674),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02730_),
    .QN(_01813_),
    .RESETN(net675),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02731_),
    .QN(_01812_),
    .RESETN(net676),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02732_),
    .QN(_01811_),
    .RESETN(net677),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02733_),
    .QN(_01810_),
    .RESETN(net678),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02734_),
    .QN(_01809_),
    .RESETN(net679),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02735_),
    .QN(_01808_),
    .RESETN(net680),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02736_),
    .QN(_01807_),
    .RESETN(net681),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02737_),
    .QN(_01806_),
    .RESETN(net682),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_02738_),
    .QN(_01805_),
    .RESETN(net683),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02739_),
    .QN(_01804_),
    .RESETN(net684),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02740_),
    .QN(_01803_),
    .RESETN(net685),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_02741_),
    .QN(_01802_),
    .RESETN(net686),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02742_),
    .QN(_01801_),
    .RESETN(net687),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02743_),
    .QN(_01800_),
    .RESETN(net688),
    .SETN(net50));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02744_),
    .QN(_01405_),
    .RESETN(net689),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02745_),
    .QN(_00746_),
    .RESETN(net690),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02746_),
    .QN(_00745_),
    .RESETN(net691),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02747_),
    .QN(_01406_),
    .RESETN(net692),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02748_),
    .QN(_01407_),
    .RESETN(net693),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02749_),
    .QN(_01408_),
    .RESETN(net694),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02750_),
    .QN(_01409_),
    .RESETN(net695),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02751_),
    .QN(_01410_),
    .RESETN(net696),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02752_),
    .QN(_01411_),
    .RESETN(net697),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02753_),
    .QN(_01412_),
    .RESETN(net698),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02754_),
    .QN(_01413_),
    .RESETN(net699),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02755_),
    .QN(_01414_),
    .RESETN(net700),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02756_),
    .QN(_01415_),
    .RESETN(net701),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02757_),
    .QN(_00007_),
    .RESETN(net702),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02758_),
    .QN(_00008_),
    .RESETN(net703),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02759_),
    .QN(_00009_),
    .RESETN(net704),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02760_),
    .QN(_00010_),
    .RESETN(net705),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02761_),
    .QN(_00011_),
    .RESETN(net706),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_02762_),
    .QN(_00012_),
    .RESETN(net707),
    .SETN(net49));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02763_),
    .QN(_00013_),
    .RESETN(net708),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02764_),
    .QN(_00014_),
    .RESETN(net709),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02765_),
    .QN(_00015_),
    .RESETN(net710),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_02766_),
    .QN(_01403_),
    .RESETN(net711),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_02767_),
    .QN(_01404_),
    .RESETN(net712),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02768_),
    .QN(_01799_),
    .RESETN(net713),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02769_),
    .QN(_18083_),
    .RESETN(net714),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02770_),
    .QN(_18084_),
    .RESETN(net715),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02771_),
    .QN(_00026_),
    .RESETN(net716),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02772_),
    .QN(_00027_),
    .RESETN(net717),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02773_),
    .QN(_01394_),
    .RESETN(net718),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1_  (.CLK(clknet_leaf_19_clk),
    .D(_00000_),
    .QN(_02197_),
    .RESETN(net44),
    .SETN(net719));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .D(_00001_),
    .QN(_01397_),
    .RESETN(net720),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .D(_00002_),
    .QN(_02198_),
    .RESETN(net721),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .D(_00003_),
    .QN(_02199_),
    .RESETN(net722),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .D(_00004_),
    .QN(_00752_),
    .RESETN(net723),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .D(_00005_),
    .QN(_01798_),
    .RESETN(net724),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02774_),
    .QN(_00066_),
    .RESETN(net725),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02775_),
    .QN(_00076_),
    .RESETN(net726),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02776_),
    .QN(_00075_),
    .RESETN(net727),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02777_),
    .QN(_00078_),
    .RESETN(net728),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02778_),
    .QN(_00077_),
    .RESETN(net729),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02779_),
    .QN(_00080_),
    .RESETN(net730),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .D(_02780_),
    .QN(_00079_),
    .RESETN(net731),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02781_),
    .QN(_00082_),
    .RESETN(net732),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02782_),
    .QN(_00081_),
    .RESETN(net733),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02783_),
    .QN(_00084_),
    .RESETN(net734),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .D(_02784_),
    .QN(_00083_),
    .RESETN(net735),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .D(_02785_),
    .QN(_00065_),
    .RESETN(net736),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .D(_02786_),
    .QN(_00086_),
    .RESETN(net737),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .D(_02787_),
    .QN(_00085_),
    .RESETN(net738),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .D(_02788_),
    .QN(_00088_),
    .RESETN(net739),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .D(_02789_),
    .QN(_00087_),
    .RESETN(net740),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02790_),
    .QN(_00090_),
    .RESETN(net741),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .D(_02791_),
    .QN(_00089_),
    .RESETN(net742),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02792_),
    .QN(_00092_),
    .RESETN(net743),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .D(_02793_),
    .QN(_00091_),
    .RESETN(net744),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02794_),
    .QN(_00094_),
    .RESETN(net745),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02795_),
    .QN(_00093_),
    .RESETN(net746),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02796_),
    .QN(_00068_),
    .RESETN(net747),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02797_),
    .QN(_00096_),
    .RESETN(net748),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02798_),
    .QN(_00095_),
    .RESETN(net749),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02799_),
    .QN(_00067_),
    .RESETN(net750),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02800_),
    .QN(_00070_),
    .RESETN(net751),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02801_),
    .QN(_00069_),
    .RESETN(net752),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02802_),
    .QN(_00072_),
    .RESETN(net753),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02803_),
    .QN(_00071_),
    .RESETN(net754),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02804_),
    .QN(_00074_),
    .RESETN(net755),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02805_),
    .QN(_00073_),
    .RESETN(net756),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02806_),
    .QN(_00028_),
    .RESETN(net757),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02807_),
    .QN(_00040_),
    .RESETN(net758),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02808_),
    .QN(_00041_),
    .RESETN(net759),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02809_),
    .QN(_00042_),
    .RESETN(net760),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02810_),
    .QN(_00043_),
    .RESETN(net761),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02811_),
    .QN(_00044_),
    .RESETN(net762),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02812_),
    .QN(_00045_),
    .RESETN(net763),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02813_),
    .QN(_00046_),
    .RESETN(net764),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02814_),
    .QN(_00047_),
    .RESETN(net765),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02815_),
    .QN(_00048_),
    .RESETN(net766),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02816_),
    .QN(_00049_),
    .RESETN(net767),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02817_),
    .QN(_00030_),
    .RESETN(net768),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02818_),
    .QN(_00050_),
    .RESETN(net769),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02819_),
    .QN(_00051_),
    .RESETN(net770),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02820_),
    .QN(_00052_),
    .RESETN(net771),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02821_),
    .QN(_00053_),
    .RESETN(net772),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02822_),
    .QN(_00054_),
    .RESETN(net773),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02823_),
    .QN(_00055_),
    .RESETN(net774),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02824_),
    .QN(_00056_),
    .RESETN(net775),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02825_),
    .QN(_00057_),
    .RESETN(net776),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02826_),
    .QN(_00058_),
    .RESETN(net777),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02827_),
    .QN(_00059_),
    .RESETN(net778),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02828_),
    .QN(_00031_),
    .RESETN(net779),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02829_),
    .QN(_00060_),
    .RESETN(net780),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02830_),
    .QN(_00061_),
    .RESETN(net781),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02831_),
    .QN(_00033_),
    .RESETN(net782),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02832_),
    .QN(_00034_),
    .RESETN(net783),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02833_),
    .QN(_00035_),
    .RESETN(net784),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02834_),
    .QN(_00036_),
    .RESETN(net785),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02835_),
    .QN(_00037_),
    .RESETN(net786),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02836_),
    .QN(_00038_),
    .RESETN(net787),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_02837_),
    .QN(_00039_),
    .RESETN(net788),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \fetch_enable_q$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_02838_),
    .QN(_01797_),
    .RESETN(net789),
    .SETN(net1963));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1000]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02839_),
    .QN(_00654_),
    .RESETN(net790),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1001]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_02840_),
    .QN(_00684_),
    .RESETN(net791),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1002]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_02841_),
    .QN(_00714_),
    .RESETN(net792),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1003]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_02842_),
    .QN(_00744_),
    .RESETN(net793),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1004]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_02843_),
    .QN(_00374_),
    .RESETN(net794),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1005]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02844_),
    .QN(_00812_),
    .RESETN(net795),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1006]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02845_),
    .QN(_00844_),
    .RESETN(net796),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1007]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02846_),
    .QN(_00876_),
    .RESETN(net797),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1008]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_02847_),
    .QN(_00908_),
    .RESETN(net798),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1009]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_02848_),
    .QN(_00940_),
    .RESETN(net799),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[100]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02849_),
    .QN(_00506_),
    .RESETN(net800),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1010]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_02850_),
    .QN(_00972_),
    .RESETN(net801),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1011]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_02851_),
    .QN(_01004_),
    .RESETN(net802),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1012]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02852_),
    .QN(_01036_),
    .RESETN(net803),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1013]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02853_),
    .QN(_01068_),
    .RESETN(net804),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1014]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02854_),
    .QN(_01100_),
    .RESETN(net805),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1015]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_02855_),
    .QN(_01132_),
    .RESETN(net806),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1016]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02856_),
    .QN(_01164_),
    .RESETN(net807),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1017]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_02857_),
    .QN(_01196_),
    .RESETN(net808),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1018]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02858_),
    .QN(_01228_),
    .RESETN(net809),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1019]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_02859_),
    .QN(_01260_),
    .RESETN(net810),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[101]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02860_),
    .QN(_00536_),
    .RESETN(net811),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1020]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02861_),
    .QN(_01292_),
    .RESETN(net812),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1021]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_02862_),
    .QN(_01324_),
    .RESETN(net813),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1022]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02863_),
    .QN(_01356_),
    .RESETN(net814),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1023]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_02864_),
    .QN(_01388_),
    .RESETN(net815),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[102]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02865_),
    .QN(_00566_),
    .RESETN(net816),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[103]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02866_),
    .QN(_00596_),
    .RESETN(net817),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[104]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02867_),
    .QN(_00626_),
    .RESETN(net818),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[105]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02868_),
    .QN(_00656_),
    .RESETN(net819),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[106]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02869_),
    .QN(_00686_),
    .RESETN(net820),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[107]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02870_),
    .QN(_00716_),
    .RESETN(net821),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[108]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02871_),
    .QN(_00346_),
    .RESETN(net822),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[109]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02872_),
    .QN(_00784_),
    .RESETN(net823),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[110]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02873_),
    .QN(_00816_),
    .RESETN(net824),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[111]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02874_),
    .QN(_00848_),
    .RESETN(net825),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[112]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02875_),
    .QN(_00880_),
    .RESETN(net826),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[113]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02876_),
    .QN(_00912_),
    .RESETN(net827),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[114]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02877_),
    .QN(_00944_),
    .RESETN(net828),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[115]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02878_),
    .QN(_00976_),
    .RESETN(net829),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[116]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02879_),
    .QN(_01008_),
    .RESETN(net830),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[117]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02880_),
    .QN(_01040_),
    .RESETN(net831),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[118]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_02881_),
    .QN(_01072_),
    .RESETN(net832),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[119]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02882_),
    .QN(_01104_),
    .RESETN(net833),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[120]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_02883_),
    .QN(_01136_),
    .RESETN(net834),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[121]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_02884_),
    .QN(_01168_),
    .RESETN(net835),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[122]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_02885_),
    .QN(_01200_),
    .RESETN(net836),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[123]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_02886_),
    .QN(_01232_),
    .RESETN(net837),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[124]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02887_),
    .QN(_01264_),
    .RESETN(net838),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[125]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02888_),
    .QN(_01296_),
    .RESETN(net839),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[126]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02889_),
    .QN(_01328_),
    .RESETN(net840),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[127]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02890_),
    .QN(_01360_),
    .RESETN(net841),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[128]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02891_),
    .QN(_00383_),
    .RESETN(net842),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[129]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02892_),
    .QN(_00416_),
    .RESETN(net843),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[130]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_02893_),
    .QN(_00447_),
    .RESETN(net844),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[131]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02894_),
    .QN(_00477_),
    .RESETN(net845),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[132]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02895_),
    .QN(_00507_),
    .RESETN(net846),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[133]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02896_),
    .QN(_00537_),
    .RESETN(net847),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[134]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02897_),
    .QN(_00567_),
    .RESETN(net848),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[135]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02898_),
    .QN(_00597_),
    .RESETN(net849),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[136]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02899_),
    .QN(_00627_),
    .RESETN(net850),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[137]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02900_),
    .QN(_00657_),
    .RESETN(net851),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[138]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02901_),
    .QN(_00687_),
    .RESETN(net852),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[139]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_02902_),
    .QN(_00717_),
    .RESETN(net853),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[140]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02903_),
    .QN(_00347_),
    .RESETN(net854),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[141]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_02904_),
    .QN(_00785_),
    .RESETN(net855),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[142]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02905_),
    .QN(_00817_),
    .RESETN(net856),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[143]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02906_),
    .QN(_00849_),
    .RESETN(net857),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[144]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_02907_),
    .QN(_00881_),
    .RESETN(net858),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[145]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02908_),
    .QN(_00913_),
    .RESETN(net859),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[146]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_02909_),
    .QN(_00945_),
    .RESETN(net860),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[147]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02910_),
    .QN(_00977_),
    .RESETN(net861),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[148]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02911_),
    .QN(_01009_),
    .RESETN(net862),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[149]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02912_),
    .QN(_01041_),
    .RESETN(net863),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[150]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02913_),
    .QN(_01073_),
    .RESETN(net864),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[151]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02914_),
    .QN(_01105_),
    .RESETN(net865),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[152]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02915_),
    .QN(_01137_),
    .RESETN(net866),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[153]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_02916_),
    .QN(_01169_),
    .RESETN(net867),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[154]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02917_),
    .QN(_01201_),
    .RESETN(net868),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[155]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02918_),
    .QN(_01233_),
    .RESETN(net869),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[156]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02919_),
    .QN(_01265_),
    .RESETN(net870),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[157]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02920_),
    .QN(_01297_),
    .RESETN(net871),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[158]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02921_),
    .QN(_01329_),
    .RESETN(net872),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[159]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02922_),
    .QN(_01361_),
    .RESETN(net873),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[160]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02923_),
    .QN(_00384_),
    .RESETN(net874),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[161]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02924_),
    .QN(_00417_),
    .RESETN(net875),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[162]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02925_),
    .QN(_00448_),
    .RESETN(net876),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[163]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02926_),
    .QN(_00478_),
    .RESETN(net877),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[164]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02927_),
    .QN(_00508_),
    .RESETN(net878),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[165]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02928_),
    .QN(_00538_),
    .RESETN(net879),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[166]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02929_),
    .QN(_00568_),
    .RESETN(net880),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[167]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02930_),
    .QN(_00598_),
    .RESETN(net881),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[168]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02931_),
    .QN(_00628_),
    .RESETN(net882),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[169]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02932_),
    .QN(_00658_),
    .RESETN(net883),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[170]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_02933_),
    .QN(_00688_),
    .RESETN(net884),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[171]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_02934_),
    .QN(_00718_),
    .RESETN(net885),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[172]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_02935_),
    .QN(_00348_),
    .RESETN(net886),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[173]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_02936_),
    .QN(_00786_),
    .RESETN(net887),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[174]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02937_),
    .QN(_00818_),
    .RESETN(net888),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[175]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02938_),
    .QN(_00850_),
    .RESETN(net889),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[176]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02939_),
    .QN(_00882_),
    .RESETN(net890),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[177]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02940_),
    .QN(_00914_),
    .RESETN(net891),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[178]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02941_),
    .QN(_00946_),
    .RESETN(net892),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[179]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02942_),
    .QN(_00978_),
    .RESETN(net893),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[180]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02943_),
    .QN(_01010_),
    .RESETN(net894),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[181]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02944_),
    .QN(_01042_),
    .RESETN(net895),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[182]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02945_),
    .QN(_01074_),
    .RESETN(net896),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[183]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02946_),
    .QN(_01106_),
    .RESETN(net897),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[184]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02947_),
    .QN(_01138_),
    .RESETN(net898),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[185]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02948_),
    .QN(_01170_),
    .RESETN(net899),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[186]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02949_),
    .QN(_01202_),
    .RESETN(net900),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[187]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02950_),
    .QN(_01234_),
    .RESETN(net901),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[188]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02951_),
    .QN(_01266_),
    .RESETN(net902),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[189]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02952_),
    .QN(_01298_),
    .RESETN(net903),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[190]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02953_),
    .QN(_01330_),
    .RESETN(net904),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[191]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02954_),
    .QN(_01362_),
    .RESETN(net905),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[192]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02955_),
    .QN(_00385_),
    .RESETN(net906),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[193]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02956_),
    .QN(_00418_),
    .RESETN(net907),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[194]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_02957_),
    .QN(_00449_),
    .RESETN(net908),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[195]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02958_),
    .QN(_00479_),
    .RESETN(net909),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[196]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02959_),
    .QN(_00509_),
    .RESETN(net910),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[197]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02960_),
    .QN(_00539_),
    .RESETN(net911),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[198]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02961_),
    .QN(_00569_),
    .RESETN(net912),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[199]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02962_),
    .QN(_00599_),
    .RESETN(net913),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[200]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02963_),
    .QN(_00629_),
    .RESETN(net914),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[201]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02964_),
    .QN(_00659_),
    .RESETN(net915),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[202]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02965_),
    .QN(_00689_),
    .RESETN(net916),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[203]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_02966_),
    .QN(_00719_),
    .RESETN(net917),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[204]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02967_),
    .QN(_00349_),
    .RESETN(net918),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[205]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02968_),
    .QN(_00787_),
    .RESETN(net919),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[206]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02969_),
    .QN(_00819_),
    .RESETN(net920),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[207]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02970_),
    .QN(_00851_),
    .RESETN(net921),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[208]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_02971_),
    .QN(_00883_),
    .RESETN(net922),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[209]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02972_),
    .QN(_00915_),
    .RESETN(net923),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[210]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_02973_),
    .QN(_00947_),
    .RESETN(net924),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[211]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02974_),
    .QN(_00979_),
    .RESETN(net925),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[212]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_02975_),
    .QN(_01011_),
    .RESETN(net926),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[213]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02976_),
    .QN(_01043_),
    .RESETN(net927),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[214]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_02977_),
    .QN(_01075_),
    .RESETN(net928),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[215]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02978_),
    .QN(_01107_),
    .RESETN(net929),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[216]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_02979_),
    .QN(_01139_),
    .RESETN(net930),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[217]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_02980_),
    .QN(_01171_),
    .RESETN(net931),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[218]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02981_),
    .QN(_01203_),
    .RESETN(net932),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[219]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02982_),
    .QN(_01235_),
    .RESETN(net933),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[220]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_02983_),
    .QN(_01267_),
    .RESETN(net934),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[221]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02984_),
    .QN(_01299_),
    .RESETN(net935),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[222]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02985_),
    .QN(_01331_),
    .RESETN(net936),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[223]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02986_),
    .QN(_01363_),
    .RESETN(net937),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[224]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02987_),
    .QN(_00386_),
    .RESETN(net938),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[225]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02988_),
    .QN(_00419_),
    .RESETN(net939),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[226]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02989_),
    .QN(_00450_),
    .RESETN(net940),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[227]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02990_),
    .QN(_00480_),
    .RESETN(net941),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[228]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02991_),
    .QN(_00510_),
    .RESETN(net942),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[229]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02992_),
    .QN(_00540_),
    .RESETN(net943),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[230]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02993_),
    .QN(_00570_),
    .RESETN(net944),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[231]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02994_),
    .QN(_00600_),
    .RESETN(net945),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[232]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02995_),
    .QN(_00630_),
    .RESETN(net946),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[233]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02996_),
    .QN(_00660_),
    .RESETN(net947),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[234]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02997_),
    .QN(_00690_),
    .RESETN(net948),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[235]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_02998_),
    .QN(_00720_),
    .RESETN(net949),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[236]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02999_),
    .QN(_00350_),
    .RESETN(net950),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[237]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03000_),
    .QN(_00788_),
    .RESETN(net951),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[238]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03001_),
    .QN(_00820_),
    .RESETN(net952),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[239]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03002_),
    .QN(_00852_),
    .RESETN(net953),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[240]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03003_),
    .QN(_00884_),
    .RESETN(net954),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[241]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03004_),
    .QN(_00916_),
    .RESETN(net955),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[242]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03005_),
    .QN(_00948_),
    .RESETN(net956),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[243]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03006_),
    .QN(_00980_),
    .RESETN(net957),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[244]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03007_),
    .QN(_01012_),
    .RESETN(net958),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[245]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03008_),
    .QN(_01044_),
    .RESETN(net959),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[246]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03009_),
    .QN(_01076_),
    .RESETN(net960),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[247]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03010_),
    .QN(_01108_),
    .RESETN(net961),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[248]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03011_),
    .QN(_01140_),
    .RESETN(net962),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[249]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03012_),
    .QN(_01172_),
    .RESETN(net963),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[250]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03013_),
    .QN(_01204_),
    .RESETN(net964),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[251]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03014_),
    .QN(_01236_),
    .RESETN(net965),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[252]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03015_),
    .QN(_01268_),
    .RESETN(net966),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[253]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03016_),
    .QN(_01300_),
    .RESETN(net967),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[254]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03017_),
    .QN(_01332_),
    .RESETN(net968),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[255]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03018_),
    .QN(_01364_),
    .RESETN(net969),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[256]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03019_),
    .QN(_00387_),
    .RESETN(net970),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[257]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03020_),
    .QN(_00420_),
    .RESETN(net971),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[258]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03021_),
    .QN(_00451_),
    .RESETN(net972),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[259]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03022_),
    .QN(_00481_),
    .RESETN(net973),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[260]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03023_),
    .QN(_00511_),
    .RESETN(net974),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[261]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03024_),
    .QN(_00541_),
    .RESETN(net975),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[262]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03025_),
    .QN(_00571_),
    .RESETN(net976),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[263]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03026_),
    .QN(_00601_),
    .RESETN(net977),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[264]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03027_),
    .QN(_00631_),
    .RESETN(net978),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[265]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03028_),
    .QN(_00661_),
    .RESETN(net979),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[266]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03029_),
    .QN(_00691_),
    .RESETN(net980),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[267]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03030_),
    .QN(_00721_),
    .RESETN(net981),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[268]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03031_),
    .QN(_00351_),
    .RESETN(net982),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[269]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03032_),
    .QN(_00789_),
    .RESETN(net983),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[270]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03033_),
    .QN(_00821_),
    .RESETN(net984),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[271]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03034_),
    .QN(_00853_),
    .RESETN(net985),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[272]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03035_),
    .QN(_00885_),
    .RESETN(net986),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[273]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03036_),
    .QN(_00917_),
    .RESETN(net987),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[274]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03037_),
    .QN(_00949_),
    .RESETN(net988),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[275]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03038_),
    .QN(_00981_),
    .RESETN(net989),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[276]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03039_),
    .QN(_01013_),
    .RESETN(net990),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[277]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03040_),
    .QN(_01045_),
    .RESETN(net991),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[278]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03041_),
    .QN(_01077_),
    .RESETN(net992),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[279]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03042_),
    .QN(_01109_),
    .RESETN(net993),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[280]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03043_),
    .QN(_01141_),
    .RESETN(net994),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[281]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03044_),
    .QN(_01173_),
    .RESETN(net995),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[282]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03045_),
    .QN(_01205_),
    .RESETN(net996),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[283]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03046_),
    .QN(_01237_),
    .RESETN(net997),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[284]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03047_),
    .QN(_01269_),
    .RESETN(net998),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[285]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03048_),
    .QN(_01301_),
    .RESETN(net999),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[286]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03049_),
    .QN(_01333_),
    .RESETN(net1000),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[287]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03050_),
    .QN(_01365_),
    .RESETN(net1001),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[288]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03051_),
    .QN(_00388_),
    .RESETN(net1002),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[289]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03052_),
    .QN(_00421_),
    .RESETN(net1003),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[290]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03053_),
    .QN(_00452_),
    .RESETN(net1004),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[291]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03054_),
    .QN(_00482_),
    .RESETN(net1005),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[292]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03055_),
    .QN(_00512_),
    .RESETN(net1006),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[293]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03056_),
    .QN(_00542_),
    .RESETN(net1007),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[294]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03057_),
    .QN(_00572_),
    .RESETN(net1008),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[295]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03058_),
    .QN(_00602_),
    .RESETN(net1009),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[296]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03059_),
    .QN(_00632_),
    .RESETN(net1010),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[297]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03060_),
    .QN(_00662_),
    .RESETN(net1011),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[298]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03061_),
    .QN(_00692_),
    .RESETN(net1012),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[299]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03062_),
    .QN(_00722_),
    .RESETN(net1013),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[300]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03063_),
    .QN(_00352_),
    .RESETN(net1014),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[301]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03064_),
    .QN(_00790_),
    .RESETN(net1015),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[302]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03065_),
    .QN(_00822_),
    .RESETN(net1016),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[303]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03066_),
    .QN(_00854_),
    .RESETN(net1017),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[304]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03067_),
    .QN(_00886_),
    .RESETN(net1018),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[305]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03068_),
    .QN(_00918_),
    .RESETN(net1019),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[306]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03069_),
    .QN(_00950_),
    .RESETN(net1020),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[307]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03070_),
    .QN(_00982_),
    .RESETN(net1021),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[308]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03071_),
    .QN(_01014_),
    .RESETN(net1022),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[309]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03072_),
    .QN(_01046_),
    .RESETN(net1023),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[310]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03073_),
    .QN(_01078_),
    .RESETN(net1024),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[311]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03074_),
    .QN(_01110_),
    .RESETN(net1025),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[312]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03075_),
    .QN(_01142_),
    .RESETN(net1026),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[313]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03076_),
    .QN(_01174_),
    .RESETN(net1027),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[314]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03077_),
    .QN(_01206_),
    .RESETN(net1028),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[315]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03078_),
    .QN(_01238_),
    .RESETN(net1029),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[316]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03079_),
    .QN(_01270_),
    .RESETN(net1030),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[317]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03080_),
    .QN(_01302_),
    .RESETN(net1031),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[318]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03081_),
    .QN(_01334_),
    .RESETN(net1032),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[319]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03082_),
    .QN(_01366_),
    .RESETN(net1033),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[320]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03083_),
    .QN(_00389_),
    .RESETN(net1034),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[321]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03084_),
    .QN(_00422_),
    .RESETN(net1035),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[322]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03085_),
    .QN(_00453_),
    .RESETN(net1036),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[323]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03086_),
    .QN(_00483_),
    .RESETN(net1037),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[324]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03087_),
    .QN(_00513_),
    .RESETN(net1038),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[325]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03088_),
    .QN(_00543_),
    .RESETN(net1039),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[326]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03089_),
    .QN(_00573_),
    .RESETN(net1040),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[327]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03090_),
    .QN(_00603_),
    .RESETN(net1041),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[328]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03091_),
    .QN(_00633_),
    .RESETN(net1042),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[329]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03092_),
    .QN(_00663_),
    .RESETN(net1043),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[32]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03093_),
    .QN(_01796_),
    .RESETN(net1044),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[330]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03094_),
    .QN(_00693_),
    .RESETN(net1045),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[331]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03095_),
    .QN(_00723_),
    .RESETN(net1046),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[332]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03096_),
    .QN(_00353_),
    .RESETN(net1047),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[333]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03097_),
    .QN(_00791_),
    .RESETN(net1048),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[334]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03098_),
    .QN(_00823_),
    .RESETN(net1049),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[335]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03099_),
    .QN(_00855_),
    .RESETN(net1050),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[336]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03100_),
    .QN(_00887_),
    .RESETN(net1051),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[337]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03101_),
    .QN(_00919_),
    .RESETN(net1052),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[338]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03102_),
    .QN(_00951_),
    .RESETN(net1053),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[339]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03103_),
    .QN(_00983_),
    .RESETN(net1054),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[33]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03104_),
    .QN(_01795_),
    .RESETN(net1055),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[340]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03105_),
    .QN(_01015_),
    .RESETN(net1056),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[341]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03106_),
    .QN(_01047_),
    .RESETN(net1057),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[342]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03107_),
    .QN(_01079_),
    .RESETN(net1058),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[343]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03108_),
    .QN(_01111_),
    .RESETN(net1059),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[344]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03109_),
    .QN(_01143_),
    .RESETN(net1060),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[345]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03110_),
    .QN(_01175_),
    .RESETN(net1061),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[346]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03111_),
    .QN(_01207_),
    .RESETN(net1062),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[347]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03112_),
    .QN(_01239_),
    .RESETN(net1063),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[348]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03113_),
    .QN(_01271_),
    .RESETN(net1064),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[349]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03114_),
    .QN(_01303_),
    .RESETN(net1065),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[34]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03115_),
    .QN(_01794_),
    .RESETN(net1066),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[350]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03116_),
    .QN(_01335_),
    .RESETN(net1067),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[351]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03117_),
    .QN(_01367_),
    .RESETN(net1068),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[352]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03118_),
    .QN(_00390_),
    .RESETN(net1069),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[353]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03119_),
    .QN(_00423_),
    .RESETN(net1070),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[354]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03120_),
    .QN(_00454_),
    .RESETN(net1071),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[355]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03121_),
    .QN(_00484_),
    .RESETN(net1072),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[356]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03122_),
    .QN(_00514_),
    .RESETN(net1073),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[357]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03123_),
    .QN(_00544_),
    .RESETN(net1074),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[358]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03124_),
    .QN(_00574_),
    .RESETN(net1075),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[359]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03125_),
    .QN(_00604_),
    .RESETN(net1076),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[35]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03126_),
    .QN(_01793_),
    .RESETN(net1077),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[360]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03127_),
    .QN(_00634_),
    .RESETN(net1078),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[361]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03128_),
    .QN(_00664_),
    .RESETN(net1079),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[362]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03129_),
    .QN(_00694_),
    .RESETN(net1080),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[363]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03130_),
    .QN(_00724_),
    .RESETN(net1081),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[364]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03131_),
    .QN(_00354_),
    .RESETN(net1082),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[365]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03132_),
    .QN(_00792_),
    .RESETN(net1083),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[366]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03133_),
    .QN(_00824_),
    .RESETN(net1084),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[367]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03134_),
    .QN(_00856_),
    .RESETN(net1085),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[368]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03135_),
    .QN(_00888_),
    .RESETN(net1086),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[369]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03136_),
    .QN(_00920_),
    .RESETN(net1087),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[36]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03137_),
    .QN(_01792_),
    .RESETN(net1088),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[370]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03138_),
    .QN(_00952_),
    .RESETN(net1089),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[371]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03139_),
    .QN(_00984_),
    .RESETN(net1090),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[372]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03140_),
    .QN(_01016_),
    .RESETN(net1091),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[373]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03141_),
    .QN(_01048_),
    .RESETN(net1092),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[374]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03142_),
    .QN(_01080_),
    .RESETN(net1093),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[375]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03143_),
    .QN(_01112_),
    .RESETN(net1094),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[376]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03144_),
    .QN(_01144_),
    .RESETN(net1095),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[377]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03145_),
    .QN(_01176_),
    .RESETN(net1096),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[378]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03146_),
    .QN(_01208_),
    .RESETN(net1097),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[379]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03147_),
    .QN(_01240_),
    .RESETN(net1098),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[37]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03148_),
    .QN(_01791_),
    .RESETN(net1099),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[380]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03149_),
    .QN(_01272_),
    .RESETN(net1100),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[381]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03150_),
    .QN(_01304_),
    .RESETN(net1101),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[382]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03151_),
    .QN(_01336_),
    .RESETN(net1102),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[383]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03152_),
    .QN(_01368_),
    .RESETN(net1103),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[384]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03153_),
    .QN(_00391_),
    .RESETN(net1104),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[385]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03154_),
    .QN(_00424_),
    .RESETN(net1105),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[386]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03155_),
    .QN(_00455_),
    .RESETN(net1106),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[387]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03156_),
    .QN(_00485_),
    .RESETN(net1107),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[388]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03157_),
    .QN(_00515_),
    .RESETN(net1108),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[389]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03158_),
    .QN(_00545_),
    .RESETN(net1109),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[38]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03159_),
    .QN(_01790_),
    .RESETN(net1110),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[390]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03160_),
    .QN(_00575_),
    .RESETN(net1111),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[391]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03161_),
    .QN(_00605_),
    .RESETN(net1112),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[392]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03162_),
    .QN(_00635_),
    .RESETN(net1113),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[393]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03163_),
    .QN(_00665_),
    .RESETN(net1114),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[394]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03164_),
    .QN(_00695_),
    .RESETN(net1115),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[395]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03165_),
    .QN(_00725_),
    .RESETN(net1116),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[396]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03166_),
    .QN(_00355_),
    .RESETN(net1117),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[397]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03167_),
    .QN(_00793_),
    .RESETN(net1118),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[398]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03168_),
    .QN(_00825_),
    .RESETN(net1119),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[399]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03169_),
    .QN(_00857_),
    .RESETN(net1120),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[39]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03170_),
    .QN(_01789_),
    .RESETN(net1121),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[400]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03171_),
    .QN(_00889_),
    .RESETN(net1122),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[401]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03172_),
    .QN(_00921_),
    .RESETN(net1123),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[402]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03173_),
    .QN(_00953_),
    .RESETN(net1124),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[403]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03174_),
    .QN(_00985_),
    .RESETN(net1125),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[404]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03175_),
    .QN(_01017_),
    .RESETN(net1126),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[405]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03176_),
    .QN(_01049_),
    .RESETN(net1127),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[406]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03177_),
    .QN(_01081_),
    .RESETN(net1128),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[407]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03178_),
    .QN(_01113_),
    .RESETN(net1129),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[408]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03179_),
    .QN(_01145_),
    .RESETN(net1130),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[409]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03180_),
    .QN(_01177_),
    .RESETN(net1131),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[40]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03181_),
    .QN(_01788_),
    .RESETN(net1132),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[410]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03182_),
    .QN(_01209_),
    .RESETN(net1133),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[411]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03183_),
    .QN(_01241_),
    .RESETN(net1134),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[412]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03184_),
    .QN(_01273_),
    .RESETN(net1135),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[413]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03185_),
    .QN(_01305_),
    .RESETN(net1136),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[414]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03186_),
    .QN(_01337_),
    .RESETN(net1137),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[415]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03187_),
    .QN(_01369_),
    .RESETN(net1138),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[416]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03188_),
    .QN(_00392_),
    .RESETN(net1139),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[417]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03189_),
    .QN(_00425_),
    .RESETN(net1140),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[418]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03190_),
    .QN(_00456_),
    .RESETN(net1141),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[419]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03191_),
    .QN(_00486_),
    .RESETN(net1142),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[41]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03192_),
    .QN(_01787_),
    .RESETN(net1143),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[420]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03193_),
    .QN(_00516_),
    .RESETN(net1144),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[421]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03194_),
    .QN(_00546_),
    .RESETN(net1145),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[422]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03195_),
    .QN(_00576_),
    .RESETN(net1146),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[423]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03196_),
    .QN(_00606_),
    .RESETN(net1147),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[424]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03197_),
    .QN(_00636_),
    .RESETN(net1148),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[425]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03198_),
    .QN(_00666_),
    .RESETN(net1149),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[426]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03199_),
    .QN(_00696_),
    .RESETN(net1150),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[427]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03200_),
    .QN(_00726_),
    .RESETN(net1151),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[428]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03201_),
    .QN(_00356_),
    .RESETN(net1152),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[429]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03202_),
    .QN(_00794_),
    .RESETN(net1153),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[42]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03203_),
    .QN(_01786_),
    .RESETN(net1154),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[430]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03204_),
    .QN(_00826_),
    .RESETN(net1155),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[431]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03205_),
    .QN(_00858_),
    .RESETN(net1156),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[432]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03206_),
    .QN(_00890_),
    .RESETN(net1157),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[433]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03207_),
    .QN(_00922_),
    .RESETN(net1158),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[434]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03208_),
    .QN(_00954_),
    .RESETN(net1159),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[435]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03209_),
    .QN(_00986_),
    .RESETN(net1160),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[436]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03210_),
    .QN(_01018_),
    .RESETN(net1161),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[437]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03211_),
    .QN(_01050_),
    .RESETN(net1162),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[438]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03212_),
    .QN(_01082_),
    .RESETN(net1163),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[439]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03213_),
    .QN(_01114_),
    .RESETN(net1164),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[43]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03214_),
    .QN(_01785_),
    .RESETN(net1165),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[440]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03215_),
    .QN(_01146_),
    .RESETN(net1166),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[441]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03216_),
    .QN(_01178_),
    .RESETN(net1167),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[442]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03217_),
    .QN(_01210_),
    .RESETN(net1168),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[443]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03218_),
    .QN(_01242_),
    .RESETN(net1169),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[444]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03219_),
    .QN(_01274_),
    .RESETN(net1170),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[445]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03220_),
    .QN(_01306_),
    .RESETN(net1171),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[446]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03221_),
    .QN(_01338_),
    .RESETN(net1172),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[447]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03222_),
    .QN(_01370_),
    .RESETN(net1173),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[448]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03223_),
    .QN(_00393_),
    .RESETN(net1174),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[449]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03224_),
    .QN(_00426_),
    .RESETN(net1175),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[44]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03225_),
    .QN(_01784_),
    .RESETN(net1176),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[450]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03226_),
    .QN(_00457_),
    .RESETN(net1177),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[451]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03227_),
    .QN(_00487_),
    .RESETN(net1178),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[452]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03228_),
    .QN(_00517_),
    .RESETN(net1179),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[453]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03229_),
    .QN(_00547_),
    .RESETN(net1180),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[454]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03230_),
    .QN(_00577_),
    .RESETN(net1181),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[455]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03231_),
    .QN(_00607_),
    .RESETN(net1182),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[456]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03232_),
    .QN(_00637_),
    .RESETN(net1183),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[457]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03233_),
    .QN(_00667_),
    .RESETN(net1184),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[458]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03234_),
    .QN(_00697_),
    .RESETN(net1185),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[459]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03235_),
    .QN(_00727_),
    .RESETN(net1186),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[45]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03236_),
    .QN(_01783_),
    .RESETN(net1187),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[460]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03237_),
    .QN(_00357_),
    .RESETN(net1188),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[461]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03238_),
    .QN(_00795_),
    .RESETN(net1189),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[462]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03239_),
    .QN(_00827_),
    .RESETN(net1190),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[463]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03240_),
    .QN(_00859_),
    .RESETN(net1191),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[464]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03241_),
    .QN(_00891_),
    .RESETN(net1192),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[465]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03242_),
    .QN(_00923_),
    .RESETN(net1193),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[466]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03243_),
    .QN(_00955_),
    .RESETN(net1194),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[467]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03244_),
    .QN(_00987_),
    .RESETN(net1195),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[468]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03245_),
    .QN(_01019_),
    .RESETN(net1196),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[469]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03246_),
    .QN(_01051_),
    .RESETN(net1197),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[46]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03247_),
    .QN(_01782_),
    .RESETN(net1198),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[470]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03248_),
    .QN(_01083_),
    .RESETN(net1199),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[471]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03249_),
    .QN(_01115_),
    .RESETN(net1200),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[472]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03250_),
    .QN(_01147_),
    .RESETN(net1201),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[473]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03251_),
    .QN(_01179_),
    .RESETN(net1202),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[474]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03252_),
    .QN(_01211_),
    .RESETN(net1203),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[475]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03253_),
    .QN(_01243_),
    .RESETN(net1204),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[476]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03254_),
    .QN(_01275_),
    .RESETN(net1205),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[477]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03255_),
    .QN(_01307_),
    .RESETN(net1206),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[478]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03256_),
    .QN(_01339_),
    .RESETN(net1207),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[479]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03257_),
    .QN(_01371_),
    .RESETN(net1208),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[47]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03258_),
    .QN(_01781_),
    .RESETN(net1209),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[480]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03259_),
    .QN(_00394_),
    .RESETN(net1210),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[481]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03260_),
    .QN(_00427_),
    .RESETN(net1211),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[482]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03261_),
    .QN(_00458_),
    .RESETN(net1212),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[483]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03262_),
    .QN(_00488_),
    .RESETN(net1213),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[484]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03263_),
    .QN(_00518_),
    .RESETN(net1214),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[485]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03264_),
    .QN(_00548_),
    .RESETN(net1215),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[486]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03265_),
    .QN(_00578_),
    .RESETN(net1216),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[487]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03266_),
    .QN(_00608_),
    .RESETN(net1217),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[488]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03267_),
    .QN(_00638_),
    .RESETN(net1218),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[489]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03268_),
    .QN(_00668_),
    .RESETN(net1219),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[48]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03269_),
    .QN(_01780_),
    .RESETN(net1220),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[490]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03270_),
    .QN(_00698_),
    .RESETN(net1221),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[491]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03271_),
    .QN(_00728_),
    .RESETN(net1222),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[492]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03272_),
    .QN(_00358_),
    .RESETN(net1223),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[493]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03273_),
    .QN(_00796_),
    .RESETN(net1224),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[494]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03274_),
    .QN(_00828_),
    .RESETN(net1225),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[495]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03275_),
    .QN(_00860_),
    .RESETN(net1226),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[496]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03276_),
    .QN(_00892_),
    .RESETN(net1227),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[497]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03277_),
    .QN(_00924_),
    .RESETN(net1228),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[498]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03278_),
    .QN(_00956_),
    .RESETN(net1229),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[499]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03279_),
    .QN(_00988_),
    .RESETN(net1230),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[49]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03280_),
    .QN(_01779_),
    .RESETN(net1231),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[500]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03281_),
    .QN(_01020_),
    .RESETN(net1232),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[501]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03282_),
    .QN(_01052_),
    .RESETN(net1233),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[502]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03283_),
    .QN(_01084_),
    .RESETN(net1234),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[503]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03284_),
    .QN(_01116_),
    .RESETN(net1235),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[504]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03285_),
    .QN(_01148_),
    .RESETN(net1236),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[505]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03286_),
    .QN(_01180_),
    .RESETN(net1237),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[506]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03287_),
    .QN(_01212_),
    .RESETN(net1238),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[507]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03288_),
    .QN(_01244_),
    .RESETN(net1239),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[508]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03289_),
    .QN(_01276_),
    .RESETN(net1240),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[509]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03290_),
    .QN(_01308_),
    .RESETN(net1241),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[50]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03291_),
    .QN(_01778_),
    .RESETN(net1242),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[510]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03292_),
    .QN(_01340_),
    .RESETN(net1243),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[511]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03293_),
    .QN(_01372_),
    .RESETN(net1244),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[512]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03294_),
    .QN(_00395_),
    .RESETN(net1245),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[513]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03295_),
    .QN(_00428_),
    .RESETN(net1246),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[514]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03296_),
    .QN(_00459_),
    .RESETN(net1247),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[515]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03297_),
    .QN(_00489_),
    .RESETN(net1248),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[516]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03298_),
    .QN(_00519_),
    .RESETN(net1249),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[517]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03299_),
    .QN(_00549_),
    .RESETN(net1250),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[518]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03300_),
    .QN(_00579_),
    .RESETN(net1251),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[519]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03301_),
    .QN(_00609_),
    .RESETN(net1252),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[51]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03302_),
    .QN(_01777_),
    .RESETN(net1253),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[520]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03303_),
    .QN(_00639_),
    .RESETN(net1254),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[521]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03304_),
    .QN(_00669_),
    .RESETN(net1255),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[522]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03305_),
    .QN(_00699_),
    .RESETN(net1256),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[523]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03306_),
    .QN(_00729_),
    .RESETN(net1257),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[524]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03307_),
    .QN(_00359_),
    .RESETN(net1258),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[525]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03308_),
    .QN(_00797_),
    .RESETN(net1259),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[526]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03309_),
    .QN(_00829_),
    .RESETN(net1260),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[527]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03310_),
    .QN(_00861_),
    .RESETN(net1261),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[528]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03311_),
    .QN(_00893_),
    .RESETN(net1262),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[529]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03312_),
    .QN(_00925_),
    .RESETN(net1263),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[52]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03313_),
    .QN(_01776_),
    .RESETN(net1264),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[530]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03314_),
    .QN(_00957_),
    .RESETN(net1265),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[531]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03315_),
    .QN(_00989_),
    .RESETN(net1266),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[532]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03316_),
    .QN(_01021_),
    .RESETN(net1267),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[533]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03317_),
    .QN(_01053_),
    .RESETN(net1268),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[534]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03318_),
    .QN(_01085_),
    .RESETN(net1269),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[535]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03319_),
    .QN(_01117_),
    .RESETN(net1270),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[536]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03320_),
    .QN(_01149_),
    .RESETN(net1271),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[537]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03321_),
    .QN(_01181_),
    .RESETN(net1272),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[538]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03322_),
    .QN(_01213_),
    .RESETN(net1273),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[539]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03323_),
    .QN(_01245_),
    .RESETN(net1274),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[53]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03324_),
    .QN(_01775_),
    .RESETN(net1275),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[540]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03325_),
    .QN(_01277_),
    .RESETN(net1276),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[541]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03326_),
    .QN(_01309_),
    .RESETN(net1277),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[542]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03327_),
    .QN(_01341_),
    .RESETN(net1278),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[543]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03328_),
    .QN(_01373_),
    .RESETN(net1279),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[544]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03329_),
    .QN(_00396_),
    .RESETN(net1280),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[545]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03330_),
    .QN(_00429_),
    .RESETN(net1281),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[546]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03331_),
    .QN(_00460_),
    .RESETN(net1282),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[547]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03332_),
    .QN(_00490_),
    .RESETN(net1283),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[548]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03333_),
    .QN(_00520_),
    .RESETN(net1284),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[549]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03334_),
    .QN(_00550_),
    .RESETN(net1285),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[54]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03335_),
    .QN(_01774_),
    .RESETN(net1286),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[550]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03336_),
    .QN(_00580_),
    .RESETN(net1287),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[551]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03337_),
    .QN(_00610_),
    .RESETN(net1288),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[552]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03338_),
    .QN(_00640_),
    .RESETN(net1289),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[553]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03339_),
    .QN(_00670_),
    .RESETN(net1290),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[554]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03340_),
    .QN(_00700_),
    .RESETN(net1291),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[555]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03341_),
    .QN(_00730_),
    .RESETN(net1292),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[556]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03342_),
    .QN(_00360_),
    .RESETN(net1293),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[557]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03343_),
    .QN(_00798_),
    .RESETN(net1294),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[558]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03344_),
    .QN(_00830_),
    .RESETN(net1295),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[559]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03345_),
    .QN(_00862_),
    .RESETN(net1296),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[55]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03346_),
    .QN(_01773_),
    .RESETN(net1297),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[560]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03347_),
    .QN(_00894_),
    .RESETN(net1298),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[561]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03348_),
    .QN(_00926_),
    .RESETN(net1299),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[562]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03349_),
    .QN(_00958_),
    .RESETN(net1300),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[563]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03350_),
    .QN(_00990_),
    .RESETN(net1301),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[564]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03351_),
    .QN(_01022_),
    .RESETN(net1302),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[565]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03352_),
    .QN(_01054_),
    .RESETN(net1303),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[566]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03353_),
    .QN(_01086_),
    .RESETN(net1304),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[567]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03354_),
    .QN(_01118_),
    .RESETN(net1305),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[568]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03355_),
    .QN(_01150_),
    .RESETN(net1306),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[569]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03356_),
    .QN(_01182_),
    .RESETN(net1307),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[56]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03357_),
    .QN(_01772_),
    .RESETN(net1308),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[570]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03358_),
    .QN(_01214_),
    .RESETN(net1309),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[571]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03359_),
    .QN(_01246_),
    .RESETN(net1310),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[572]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03360_),
    .QN(_01278_),
    .RESETN(net1311),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[573]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03361_),
    .QN(_01310_),
    .RESETN(net1312),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[574]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03362_),
    .QN(_01342_),
    .RESETN(net1313),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[575]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03363_),
    .QN(_01374_),
    .RESETN(net1314),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[576]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03364_),
    .QN(_00397_),
    .RESETN(net1315),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[577]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03365_),
    .QN(_00430_),
    .RESETN(net1316),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[578]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03366_),
    .QN(_00461_),
    .RESETN(net1317),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[579]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03367_),
    .QN(_00491_),
    .RESETN(net1318),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[57]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03368_),
    .QN(_01771_),
    .RESETN(net1319),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[580]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03369_),
    .QN(_00521_),
    .RESETN(net1320),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[581]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03370_),
    .QN(_00551_),
    .RESETN(net1321),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[582]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03371_),
    .QN(_00581_),
    .RESETN(net1322),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[583]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03372_),
    .QN(_00611_),
    .RESETN(net1323),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[584]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03373_),
    .QN(_00641_),
    .RESETN(net1324),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[585]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03374_),
    .QN(_00671_),
    .RESETN(net1325),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[586]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03375_),
    .QN(_00701_),
    .RESETN(net1326),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[587]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03376_),
    .QN(_00731_),
    .RESETN(net1327),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[588]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03377_),
    .QN(_00361_),
    .RESETN(net1328),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[589]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03378_),
    .QN(_00799_),
    .RESETN(net1329),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[58]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03379_),
    .QN(_01770_),
    .RESETN(net1330),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[590]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03380_),
    .QN(_00831_),
    .RESETN(net1331),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[591]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03381_),
    .QN(_00863_),
    .RESETN(net1332),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[592]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03382_),
    .QN(_00895_),
    .RESETN(net1333),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[593]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03383_),
    .QN(_00927_),
    .RESETN(net1334),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[594]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03384_),
    .QN(_00959_),
    .RESETN(net1335),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[595]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03385_),
    .QN(_00991_),
    .RESETN(net1336),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[596]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03386_),
    .QN(_01023_),
    .RESETN(net1337),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[597]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03387_),
    .QN(_01055_),
    .RESETN(net1338),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[598]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03388_),
    .QN(_01087_),
    .RESETN(net1339),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[599]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03389_),
    .QN(_01119_),
    .RESETN(net1340),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[59]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03390_),
    .QN(_01769_),
    .RESETN(net1341),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[600]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03391_),
    .QN(_01151_),
    .RESETN(net1342),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[601]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03392_),
    .QN(_01183_),
    .RESETN(net1343),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[602]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03393_),
    .QN(_01215_),
    .RESETN(net1344),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[603]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03394_),
    .QN(_01247_),
    .RESETN(net1345),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[604]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03395_),
    .QN(_01279_),
    .RESETN(net1346),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[605]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03396_),
    .QN(_01311_),
    .RESETN(net1347),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[606]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03397_),
    .QN(_01343_),
    .RESETN(net1348),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[607]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03398_),
    .QN(_01375_),
    .RESETN(net1349),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[608]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03399_),
    .QN(_00398_),
    .RESETN(net1350),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[609]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03400_),
    .QN(_00431_),
    .RESETN(net1351),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[60]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03401_),
    .QN(_01768_),
    .RESETN(net1352),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[610]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03402_),
    .QN(_00462_),
    .RESETN(net1353),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[611]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03403_),
    .QN(_00492_),
    .RESETN(net1354),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[612]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03404_),
    .QN(_00522_),
    .RESETN(net1355),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[613]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03405_),
    .QN(_00552_),
    .RESETN(net1356),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[614]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03406_),
    .QN(_00582_),
    .RESETN(net1357),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[615]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03407_),
    .QN(_00612_),
    .RESETN(net1358),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[616]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03408_),
    .QN(_00642_),
    .RESETN(net1359),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[617]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03409_),
    .QN(_00672_),
    .RESETN(net1360),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[618]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03410_),
    .QN(_00702_),
    .RESETN(net1361),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[619]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03411_),
    .QN(_00732_),
    .RESETN(net1362),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[61]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03412_),
    .QN(_01767_),
    .RESETN(net1363),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[620]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03413_),
    .QN(_00362_),
    .RESETN(net1364),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[621]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03414_),
    .QN(_00800_),
    .RESETN(net1365),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[622]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03415_),
    .QN(_00832_),
    .RESETN(net1366),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[623]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03416_),
    .QN(_00864_),
    .RESETN(net1367),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[624]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03417_),
    .QN(_00896_),
    .RESETN(net1368),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[625]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03418_),
    .QN(_00928_),
    .RESETN(net1369),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[626]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03419_),
    .QN(_00960_),
    .RESETN(net1370),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[627]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03420_),
    .QN(_00992_),
    .RESETN(net1371),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[628]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03421_),
    .QN(_01024_),
    .RESETN(net1372),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[629]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03422_),
    .QN(_01056_),
    .RESETN(net1373),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[62]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03423_),
    .QN(_01766_),
    .RESETN(net1374),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[630]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03424_),
    .QN(_01088_),
    .RESETN(net1375),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[631]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03425_),
    .QN(_01120_),
    .RESETN(net1376),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[632]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03426_),
    .QN(_01152_),
    .RESETN(net1377),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[633]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03427_),
    .QN(_01184_),
    .RESETN(net1378),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[634]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03428_),
    .QN(_01216_),
    .RESETN(net1379),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[635]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03429_),
    .QN(_01248_),
    .RESETN(net1380),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[636]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03430_),
    .QN(_01280_),
    .RESETN(net1381),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[637]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03431_),
    .QN(_01312_),
    .RESETN(net1382),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[638]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03432_),
    .QN(_01344_),
    .RESETN(net1383),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[639]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03433_),
    .QN(_01376_),
    .RESETN(net1384),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[63]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03434_),
    .QN(_01765_),
    .RESETN(net1385),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[640]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03435_),
    .QN(_00399_),
    .RESETN(net1386),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[641]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03436_),
    .QN(_00432_),
    .RESETN(net1387),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[642]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03437_),
    .QN(_00463_),
    .RESETN(net1388),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[643]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03438_),
    .QN(_00493_),
    .RESETN(net1389),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[644]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03439_),
    .QN(_00523_),
    .RESETN(net1390),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[645]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03440_),
    .QN(_00553_),
    .RESETN(net1391),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[646]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03441_),
    .QN(_00583_),
    .RESETN(net1392),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[647]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03442_),
    .QN(_00613_),
    .RESETN(net1393),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[648]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03443_),
    .QN(_00643_),
    .RESETN(net1394),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[649]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03444_),
    .QN(_00673_),
    .RESETN(net1395),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[64]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03445_),
    .QN(_00381_),
    .RESETN(net1396),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[650]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03446_),
    .QN(_00703_),
    .RESETN(net1397),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[651]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03447_),
    .QN(_00733_),
    .RESETN(net1398),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[652]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03448_),
    .QN(_00363_),
    .RESETN(net1399),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[653]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03449_),
    .QN(_00801_),
    .RESETN(net1400),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[654]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03450_),
    .QN(_00833_),
    .RESETN(net1401),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[655]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03451_),
    .QN(_00865_),
    .RESETN(net1402),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[656]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03452_),
    .QN(_00897_),
    .RESETN(net1403),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[657]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03453_),
    .QN(_00929_),
    .RESETN(net1404),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[658]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03454_),
    .QN(_00961_),
    .RESETN(net1405),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[659]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03455_),
    .QN(_00993_),
    .RESETN(net1406),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[65]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03456_),
    .QN(_00414_),
    .RESETN(net1407),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[660]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03457_),
    .QN(_01025_),
    .RESETN(net1408),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[661]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03458_),
    .QN(_01057_),
    .RESETN(net1409),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[662]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03459_),
    .QN(_01089_),
    .RESETN(net1410),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[663]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03460_),
    .QN(_01121_),
    .RESETN(net1411),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[664]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03461_),
    .QN(_01153_),
    .RESETN(net1412),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[665]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03462_),
    .QN(_01185_),
    .RESETN(net1413),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[666]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03463_),
    .QN(_01217_),
    .RESETN(net1414),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[667]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03464_),
    .QN(_01249_),
    .RESETN(net1415),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[668]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03465_),
    .QN(_01281_),
    .RESETN(net1416),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[669]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03466_),
    .QN(_01313_),
    .RESETN(net1417),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[66]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03467_),
    .QN(_00445_),
    .RESETN(net1418),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[670]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03468_),
    .QN(_01345_),
    .RESETN(net1419),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[671]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03469_),
    .QN(_01377_),
    .RESETN(net1420),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[672]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03470_),
    .QN(_00400_),
    .RESETN(net1421),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[673]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03471_),
    .QN(_00433_),
    .RESETN(net1422),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[674]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03472_),
    .QN(_00464_),
    .RESETN(net1423),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[675]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03473_),
    .QN(_00494_),
    .RESETN(net1424),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[676]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03474_),
    .QN(_00524_),
    .RESETN(net1425),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[677]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03475_),
    .QN(_00554_),
    .RESETN(net1426),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[678]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03476_),
    .QN(_00584_),
    .RESETN(net1427),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[679]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03477_),
    .QN(_00614_),
    .RESETN(net1428),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[67]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03478_),
    .QN(_00475_),
    .RESETN(net1429),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[680]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03479_),
    .QN(_00644_),
    .RESETN(net1430),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[681]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03480_),
    .QN(_00674_),
    .RESETN(net1431),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[682]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03481_),
    .QN(_00704_),
    .RESETN(net1432),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[683]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03482_),
    .QN(_00734_),
    .RESETN(net1433),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[684]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03483_),
    .QN(_00364_),
    .RESETN(net1434),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[685]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03484_),
    .QN(_00802_),
    .RESETN(net1435),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[686]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03485_),
    .QN(_00834_),
    .RESETN(net1436),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[687]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03486_),
    .QN(_00866_),
    .RESETN(net1437),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[688]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03487_),
    .QN(_00898_),
    .RESETN(net1438),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[689]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03488_),
    .QN(_00930_),
    .RESETN(net1439),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[68]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03489_),
    .QN(_00505_),
    .RESETN(net1440),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[690]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03490_),
    .QN(_00962_),
    .RESETN(net1441),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[691]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03491_),
    .QN(_00994_),
    .RESETN(net1442),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[692]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03492_),
    .QN(_01026_),
    .RESETN(net1443),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[693]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03493_),
    .QN(_01058_),
    .RESETN(net1444),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[694]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03494_),
    .QN(_01090_),
    .RESETN(net1445),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[695]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03495_),
    .QN(_01122_),
    .RESETN(net1446),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[696]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03496_),
    .QN(_01154_),
    .RESETN(net1447),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[697]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03497_),
    .QN(_01186_),
    .RESETN(net1448),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[698]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03498_),
    .QN(_01218_),
    .RESETN(net1449),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[699]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03499_),
    .QN(_01250_),
    .RESETN(net1450),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[69]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03500_),
    .QN(_00535_),
    .RESETN(net1451),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[700]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03501_),
    .QN(_01282_),
    .RESETN(net1452),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[701]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03502_),
    .QN(_01314_),
    .RESETN(net1453),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[702]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03503_),
    .QN(_01346_),
    .RESETN(net1454),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[703]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03504_),
    .QN(_01378_),
    .RESETN(net1455),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[704]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03505_),
    .QN(_00401_),
    .RESETN(net1456),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[705]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03506_),
    .QN(_00434_),
    .RESETN(net1457),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[706]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03507_),
    .QN(_00465_),
    .RESETN(net1458),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[707]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03508_),
    .QN(_00495_),
    .RESETN(net1459),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[708]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03509_),
    .QN(_00525_),
    .RESETN(net1460),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[709]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03510_),
    .QN(_00555_),
    .RESETN(net1461),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[70]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03511_),
    .QN(_00565_),
    .RESETN(net1462),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[710]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03512_),
    .QN(_00585_),
    .RESETN(net1463),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[711]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03513_),
    .QN(_00615_),
    .RESETN(net1464),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[712]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03514_),
    .QN(_00645_),
    .RESETN(net1465),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[713]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03515_),
    .QN(_00675_),
    .RESETN(net1466),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[714]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03516_),
    .QN(_00705_),
    .RESETN(net1467),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[715]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03517_),
    .QN(_00735_),
    .RESETN(net1468),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[716]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03518_),
    .QN(_00365_),
    .RESETN(net1469),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[717]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03519_),
    .QN(_00803_),
    .RESETN(net1470),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[718]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03520_),
    .QN(_00835_),
    .RESETN(net1471),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[719]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03521_),
    .QN(_00867_),
    .RESETN(net1472),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[71]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03522_),
    .QN(_00595_),
    .RESETN(net1473),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[720]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03523_),
    .QN(_00899_),
    .RESETN(net1474),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[721]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03524_),
    .QN(_00931_),
    .RESETN(net1475),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[722]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03525_),
    .QN(_00963_),
    .RESETN(net1476),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[723]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03526_),
    .QN(_00995_),
    .RESETN(net1477),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[724]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03527_),
    .QN(_01027_),
    .RESETN(net1478),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[725]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03528_),
    .QN(_01059_),
    .RESETN(net1479),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[726]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03529_),
    .QN(_01091_),
    .RESETN(net1480),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[727]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03530_),
    .QN(_01123_),
    .RESETN(net1481),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[728]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03531_),
    .QN(_01155_),
    .RESETN(net1482),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[729]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03532_),
    .QN(_01187_),
    .RESETN(net1483),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[72]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03533_),
    .QN(_00625_),
    .RESETN(net1484),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[730]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03534_),
    .QN(_01219_),
    .RESETN(net1485),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[731]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03535_),
    .QN(_01251_),
    .RESETN(net1486),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[732]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03536_),
    .QN(_01283_),
    .RESETN(net1487),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[733]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03537_),
    .QN(_01315_),
    .RESETN(net1488),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[734]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03538_),
    .QN(_01347_),
    .RESETN(net1489),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[735]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03539_),
    .QN(_01379_),
    .RESETN(net1490),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[736]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03540_),
    .QN(_00402_),
    .RESETN(net1491),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[737]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03541_),
    .QN(_00435_),
    .RESETN(net1492),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[738]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03542_),
    .QN(_00466_),
    .RESETN(net1493),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[739]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03543_),
    .QN(_00496_),
    .RESETN(net1494),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[73]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03544_),
    .QN(_00655_),
    .RESETN(net1495),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[740]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03545_),
    .QN(_00526_),
    .RESETN(net1496),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[741]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03546_),
    .QN(_00556_),
    .RESETN(net1497),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[742]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03547_),
    .QN(_00586_),
    .RESETN(net1498),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[743]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03548_),
    .QN(_00616_),
    .RESETN(net1499),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[744]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03549_),
    .QN(_00646_),
    .RESETN(net1500),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[745]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03550_),
    .QN(_00676_),
    .RESETN(net1501),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[746]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03551_),
    .QN(_00706_),
    .RESETN(net1502),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[747]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03552_),
    .QN(_00736_),
    .RESETN(net1503),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[748]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03553_),
    .QN(_00366_),
    .RESETN(net1504),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[749]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03554_),
    .QN(_00804_),
    .RESETN(net1505),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[74]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03555_),
    .QN(_00685_),
    .RESETN(net1506),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[750]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03556_),
    .QN(_00836_),
    .RESETN(net1507),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[751]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03557_),
    .QN(_00868_),
    .RESETN(net1508),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[752]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03558_),
    .QN(_00900_),
    .RESETN(net1509),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[753]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03559_),
    .QN(_00932_),
    .RESETN(net1510),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[754]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03560_),
    .QN(_00964_),
    .RESETN(net1511),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[755]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03561_),
    .QN(_00996_),
    .RESETN(net1512),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[756]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03562_),
    .QN(_01028_),
    .RESETN(net1513),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[757]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03563_),
    .QN(_01060_),
    .RESETN(net1514),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[758]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03564_),
    .QN(_01092_),
    .RESETN(net1515),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[759]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03565_),
    .QN(_01124_),
    .RESETN(net1516),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[75]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03566_),
    .QN(_00715_),
    .RESETN(net1517),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[760]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03567_),
    .QN(_01156_),
    .RESETN(net1518),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[761]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03568_),
    .QN(_01188_),
    .RESETN(net1519),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[762]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03569_),
    .QN(_01220_),
    .RESETN(net1520),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[763]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03570_),
    .QN(_01252_),
    .RESETN(net1521),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[764]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03571_),
    .QN(_01284_),
    .RESETN(net1522),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[765]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03572_),
    .QN(_01316_),
    .RESETN(net1523),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[766]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03573_),
    .QN(_01348_),
    .RESETN(net1524),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[767]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03574_),
    .QN(_01380_),
    .RESETN(net1525),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[768]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03575_),
    .QN(_00403_),
    .RESETN(net1526),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[769]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03576_),
    .QN(_00436_),
    .RESETN(net1527),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[76]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03577_),
    .QN(_00345_),
    .RESETN(net1528),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[770]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03578_),
    .QN(_00467_),
    .RESETN(net1529),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[771]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03579_),
    .QN(_00497_),
    .RESETN(net1530),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[772]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03580_),
    .QN(_00527_),
    .RESETN(net1531),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[773]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03581_),
    .QN(_00557_),
    .RESETN(net1532),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[774]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03582_),
    .QN(_00587_),
    .RESETN(net1533),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[775]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03583_),
    .QN(_00617_),
    .RESETN(net1534),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[776]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03584_),
    .QN(_00647_),
    .RESETN(net1535),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[777]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03585_),
    .QN(_00677_),
    .RESETN(net1536),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[778]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03586_),
    .QN(_00707_),
    .RESETN(net1537),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[779]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03587_),
    .QN(_00737_),
    .RESETN(net1538),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[77]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03588_),
    .QN(_00783_),
    .RESETN(net1539),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[780]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03589_),
    .QN(_00367_),
    .RESETN(net1540),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[781]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03590_),
    .QN(_00805_),
    .RESETN(net1541),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[782]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03591_),
    .QN(_00837_),
    .RESETN(net1542),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[783]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03592_),
    .QN(_00869_),
    .RESETN(net1543),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[784]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03593_),
    .QN(_00901_),
    .RESETN(net1544),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[785]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03594_),
    .QN(_00933_),
    .RESETN(net1545),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[786]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03595_),
    .QN(_00965_),
    .RESETN(net1546),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[787]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03596_),
    .QN(_00997_),
    .RESETN(net1547),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[788]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03597_),
    .QN(_01029_),
    .RESETN(net1548),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[789]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03598_),
    .QN(_01061_),
    .RESETN(net1549),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[78]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03599_),
    .QN(_00815_),
    .RESETN(net1550),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[790]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03600_),
    .QN(_01093_),
    .RESETN(net1551),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[791]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03601_),
    .QN(_01125_),
    .RESETN(net1552),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[792]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03602_),
    .QN(_01157_),
    .RESETN(net1553),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[793]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03603_),
    .QN(_01189_),
    .RESETN(net1554),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[794]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03604_),
    .QN(_01221_),
    .RESETN(net1555),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[795]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03605_),
    .QN(_01253_),
    .RESETN(net1556),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[796]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03606_),
    .QN(_01285_),
    .RESETN(net1557),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[797]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03607_),
    .QN(_01317_),
    .RESETN(net1558),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[798]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03608_),
    .QN(_01349_),
    .RESETN(net1559),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[799]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03609_),
    .QN(_01381_),
    .RESETN(net1560),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[79]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03610_),
    .QN(_00847_),
    .RESETN(net1561),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[800]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03611_),
    .QN(_00404_),
    .RESETN(net1562),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[801]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03612_),
    .QN(_00437_),
    .RESETN(net1563),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[802]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03613_),
    .QN(_00468_),
    .RESETN(net1564),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[803]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03614_),
    .QN(_00498_),
    .RESETN(net1565),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[804]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03615_),
    .QN(_00528_),
    .RESETN(net1566),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[805]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03616_),
    .QN(_00558_),
    .RESETN(net1567),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[806]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03617_),
    .QN(_00588_),
    .RESETN(net1568),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[807]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03618_),
    .QN(_00618_),
    .RESETN(net1569),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[808]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03619_),
    .QN(_00648_),
    .RESETN(net1570),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[809]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03620_),
    .QN(_00678_),
    .RESETN(net1571),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[80]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03621_),
    .QN(_00879_),
    .RESETN(net1572),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[810]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03622_),
    .QN(_00708_),
    .RESETN(net1573),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[811]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03623_),
    .QN(_00738_),
    .RESETN(net1574),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[812]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03624_),
    .QN(_00368_),
    .RESETN(net1575),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[813]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03625_),
    .QN(_00806_),
    .RESETN(net1576),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[814]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03626_),
    .QN(_00838_),
    .RESETN(net1577),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[815]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03627_),
    .QN(_00870_),
    .RESETN(net1578),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[816]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03628_),
    .QN(_00902_),
    .RESETN(net1579),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[817]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03629_),
    .QN(_00934_),
    .RESETN(net1580),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[818]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03630_),
    .QN(_00966_),
    .RESETN(net1581),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[819]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03631_),
    .QN(_00998_),
    .RESETN(net1582),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[81]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03632_),
    .QN(_00911_),
    .RESETN(net1583),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[820]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03633_),
    .QN(_01030_),
    .RESETN(net1584),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[821]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03634_),
    .QN(_01062_),
    .RESETN(net1585),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[822]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03635_),
    .QN(_01094_),
    .RESETN(net1586),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[823]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03636_),
    .QN(_01126_),
    .RESETN(net1587),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[824]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03637_),
    .QN(_01158_),
    .RESETN(net1588),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[825]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03638_),
    .QN(_01190_),
    .RESETN(net1589),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[826]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03639_),
    .QN(_01222_),
    .RESETN(net1590),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[827]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03640_),
    .QN(_01254_),
    .RESETN(net1591),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[828]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03641_),
    .QN(_01286_),
    .RESETN(net1592),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[829]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03642_),
    .QN(_01318_),
    .RESETN(net1593),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[82]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03643_),
    .QN(_00943_),
    .RESETN(net1594),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[830]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03644_),
    .QN(_01350_),
    .RESETN(net1595),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[831]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03645_),
    .QN(_01382_),
    .RESETN(net1596),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[832]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03646_),
    .QN(_00405_),
    .RESETN(net1597),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[833]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03647_),
    .QN(_00438_),
    .RESETN(net1598),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[834]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03648_),
    .QN(_00469_),
    .RESETN(net1599),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[835]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03649_),
    .QN(_00499_),
    .RESETN(net1600),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[836]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03650_),
    .QN(_00529_),
    .RESETN(net1601),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[837]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03651_),
    .QN(_00559_),
    .RESETN(net1602),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[838]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03652_),
    .QN(_00589_),
    .RESETN(net1603),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[839]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03653_),
    .QN(_00619_),
    .RESETN(net1604),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[83]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03654_),
    .QN(_00975_),
    .RESETN(net1605),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[840]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03655_),
    .QN(_00649_),
    .RESETN(net1606),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[841]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03656_),
    .QN(_00679_),
    .RESETN(net1607),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[842]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03657_),
    .QN(_00709_),
    .RESETN(net1608),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[843]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03658_),
    .QN(_00739_),
    .RESETN(net1609),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[844]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03659_),
    .QN(_00369_),
    .RESETN(net1610),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[845]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03660_),
    .QN(_00807_),
    .RESETN(net1611),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[846]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03661_),
    .QN(_00839_),
    .RESETN(net1612),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[847]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03662_),
    .QN(_00871_),
    .RESETN(net1613),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[848]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03663_),
    .QN(_00903_),
    .RESETN(net1614),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[849]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03664_),
    .QN(_00935_),
    .RESETN(net1615),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[84]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03665_),
    .QN(_01007_),
    .RESETN(net1616),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[850]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03666_),
    .QN(_00967_),
    .RESETN(net1617),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[851]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03667_),
    .QN(_00999_),
    .RESETN(net1618),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[852]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03668_),
    .QN(_01031_),
    .RESETN(net1619),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[853]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03669_),
    .QN(_01063_),
    .RESETN(net1620),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[854]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03670_),
    .QN(_01095_),
    .RESETN(net1621),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[855]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03671_),
    .QN(_01127_),
    .RESETN(net1622),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[856]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03672_),
    .QN(_01159_),
    .RESETN(net1623),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[857]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03673_),
    .QN(_01191_),
    .RESETN(net1624),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[858]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03674_),
    .QN(_01223_),
    .RESETN(net1625),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[859]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03675_),
    .QN(_01255_),
    .RESETN(net1626),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[85]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03676_),
    .QN(_01039_),
    .RESETN(net1627),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[860]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03677_),
    .QN(_01287_),
    .RESETN(net1628),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[861]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03678_),
    .QN(_01319_),
    .RESETN(net1629),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[862]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03679_),
    .QN(_01351_),
    .RESETN(net1630),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[863]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03680_),
    .QN(_01383_),
    .RESETN(net1631),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[864]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03681_),
    .QN(_00406_),
    .RESETN(net1632),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[865]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03682_),
    .QN(_00439_),
    .RESETN(net1633),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[866]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03683_),
    .QN(_00470_),
    .RESETN(net1634),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[867]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03684_),
    .QN(_00500_),
    .RESETN(net1635),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[868]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03685_),
    .QN(_00530_),
    .RESETN(net1636),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[869]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03686_),
    .QN(_00560_),
    .RESETN(net1637),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[86]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03687_),
    .QN(_01071_),
    .RESETN(net1638),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[870]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03688_),
    .QN(_00590_),
    .RESETN(net1639),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[871]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03689_),
    .QN(_00620_),
    .RESETN(net1640),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[872]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03690_),
    .QN(_00650_),
    .RESETN(net1641),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[873]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03691_),
    .QN(_00680_),
    .RESETN(net1642),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[874]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03692_),
    .QN(_00710_),
    .RESETN(net1643),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[875]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03693_),
    .QN(_00740_),
    .RESETN(net1644),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[876]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03694_),
    .QN(_00370_),
    .RESETN(net1645),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[877]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03695_),
    .QN(_00808_),
    .RESETN(net1646),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[878]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03696_),
    .QN(_00840_),
    .RESETN(net1647),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[879]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03697_),
    .QN(_00872_),
    .RESETN(net1648),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[87]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03698_),
    .QN(_01103_),
    .RESETN(net1649),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[880]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03699_),
    .QN(_00904_),
    .RESETN(net1650),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[881]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03700_),
    .QN(_00936_),
    .RESETN(net1651),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[882]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03701_),
    .QN(_00968_),
    .RESETN(net1652),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[883]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03702_),
    .QN(_01000_),
    .RESETN(net1653),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[884]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03703_),
    .QN(_01032_),
    .RESETN(net1654),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[885]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03704_),
    .QN(_01064_),
    .RESETN(net1655),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[886]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03705_),
    .QN(_01096_),
    .RESETN(net1656),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[887]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03706_),
    .QN(_01128_),
    .RESETN(net1657),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[888]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03707_),
    .QN(_01160_),
    .RESETN(net1658),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[889]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03708_),
    .QN(_01192_),
    .RESETN(net1659),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[88]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03709_),
    .QN(_01135_),
    .RESETN(net1660),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[890]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03710_),
    .QN(_01224_),
    .RESETN(net1661),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[891]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03711_),
    .QN(_01256_),
    .RESETN(net1662),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[892]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03712_),
    .QN(_01288_),
    .RESETN(net1663),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[893]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03713_),
    .QN(_01320_),
    .RESETN(net1664),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[894]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03714_),
    .QN(_01352_),
    .RESETN(net1665),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[895]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03715_),
    .QN(_01384_),
    .RESETN(net1666),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[896]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03716_),
    .QN(_00407_),
    .RESETN(net1667),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[897]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03717_),
    .QN(_00440_),
    .RESETN(net1668),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[898]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03718_),
    .QN(_00471_),
    .RESETN(net1669),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[899]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03719_),
    .QN(_00501_),
    .RESETN(net1670),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[89]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03720_),
    .QN(_01167_),
    .RESETN(net1671),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[900]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03721_),
    .QN(_00531_),
    .RESETN(net1672),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[901]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03722_),
    .QN(_00561_),
    .RESETN(net1673),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[902]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03723_),
    .QN(_00591_),
    .RESETN(net1674),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[903]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03724_),
    .QN(_00621_),
    .RESETN(net1675),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[904]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03725_),
    .QN(_00651_),
    .RESETN(net1676),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[905]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03726_),
    .QN(_00681_),
    .RESETN(net1677),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[906]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03727_),
    .QN(_00711_),
    .RESETN(net1678),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[907]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03728_),
    .QN(_00741_),
    .RESETN(net1679),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[908]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03729_),
    .QN(_00371_),
    .RESETN(net1680),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[909]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03730_),
    .QN(_00809_),
    .RESETN(net1681),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[90]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03731_),
    .QN(_01199_),
    .RESETN(net1682),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[910]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03732_),
    .QN(_00841_),
    .RESETN(net1683),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[911]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03733_),
    .QN(_00873_),
    .RESETN(net1684),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[912]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03734_),
    .QN(_00905_),
    .RESETN(net1685),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[913]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03735_),
    .QN(_00937_),
    .RESETN(net1686),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[914]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03736_),
    .QN(_00969_),
    .RESETN(net1687),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[915]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03737_),
    .QN(_01001_),
    .RESETN(net1688),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[916]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03738_),
    .QN(_01033_),
    .RESETN(net1689),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[917]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03739_),
    .QN(_01065_),
    .RESETN(net1690),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[918]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03740_),
    .QN(_01097_),
    .RESETN(net1691),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[919]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03741_),
    .QN(_01129_),
    .RESETN(net1692),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[91]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03742_),
    .QN(_01231_),
    .RESETN(net1693),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[920]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03743_),
    .QN(_01161_),
    .RESETN(net1694),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[921]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03744_),
    .QN(_01193_),
    .RESETN(net1695),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[922]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03745_),
    .QN(_01225_),
    .RESETN(net1696),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[923]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03746_),
    .QN(_01257_),
    .RESETN(net1697),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[924]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03747_),
    .QN(_01289_),
    .RESETN(net1698),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[925]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03748_),
    .QN(_01321_),
    .RESETN(net1699),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[926]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03749_),
    .QN(_01353_),
    .RESETN(net1700),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[927]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03750_),
    .QN(_01385_),
    .RESETN(net1701),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[928]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03751_),
    .QN(_00408_),
    .RESETN(net1702),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[929]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03752_),
    .QN(_00441_),
    .RESETN(net1703),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[92]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03753_),
    .QN(_01263_),
    .RESETN(net1704),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[930]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03754_),
    .QN(_00472_),
    .RESETN(net1705),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[931]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03755_),
    .QN(_00502_),
    .RESETN(net1706),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[932]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03756_),
    .QN(_00532_),
    .RESETN(net1707),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[933]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03757_),
    .QN(_00562_),
    .RESETN(net1708),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[934]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03758_),
    .QN(_00592_),
    .RESETN(net1709),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[935]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03759_),
    .QN(_00622_),
    .RESETN(net1710),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[936]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03760_),
    .QN(_00652_),
    .RESETN(net1711),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[937]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03761_),
    .QN(_00682_),
    .RESETN(net1712),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[938]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03762_),
    .QN(_00712_),
    .RESETN(net1713),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[939]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03763_),
    .QN(_00742_),
    .RESETN(net1714),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[93]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03764_),
    .QN(_01295_),
    .RESETN(net1715),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[940]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03765_),
    .QN(_00372_),
    .RESETN(net1716),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[941]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03766_),
    .QN(_00810_),
    .RESETN(net1717),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[942]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03767_),
    .QN(_00842_),
    .RESETN(net1718),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[943]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03768_),
    .QN(_00874_),
    .RESETN(net1719),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[944]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03769_),
    .QN(_00906_),
    .RESETN(net1720),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[945]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03770_),
    .QN(_00938_),
    .RESETN(net1721),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[946]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03771_),
    .QN(_00970_),
    .RESETN(net1722),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[947]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03772_),
    .QN(_01002_),
    .RESETN(net1723),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[948]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03773_),
    .QN(_01034_),
    .RESETN(net1724),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[949]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03774_),
    .QN(_01066_),
    .RESETN(net1725),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[94]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03775_),
    .QN(_01327_),
    .RESETN(net1726),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[950]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03776_),
    .QN(_01098_),
    .RESETN(net1727),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[951]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03777_),
    .QN(_01130_),
    .RESETN(net1728),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[952]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03778_),
    .QN(_01162_),
    .RESETN(net1729),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[953]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03779_),
    .QN(_01194_),
    .RESETN(net1730),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[954]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03780_),
    .QN(_01226_),
    .RESETN(net1731),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[955]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03781_),
    .QN(_01258_),
    .RESETN(net1732),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[956]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03782_),
    .QN(_01290_),
    .RESETN(net1733),
    .SETN(net43));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[957]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03783_),
    .QN(_01322_),
    .RESETN(net1734),
    .SETN(net42));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[958]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03784_),
    .QN(_01354_),
    .RESETN(net1735),
    .SETN(net37));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[959]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03785_),
    .QN(_01386_),
    .RESETN(net1736),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[95]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03786_),
    .QN(_01359_),
    .RESETN(net1737),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[960]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03787_),
    .QN(_00409_),
    .RESETN(net1738),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[961]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03788_),
    .QN(_00442_),
    .RESETN(net1739),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[962]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03789_),
    .QN(_00473_),
    .RESETN(net1740),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[963]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03790_),
    .QN(_00503_),
    .RESETN(net1741),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[964]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03791_),
    .QN(_00533_),
    .RESETN(net1742),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[965]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03792_),
    .QN(_00563_),
    .RESETN(net1743),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[966]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03793_),
    .QN(_00593_),
    .RESETN(net1744),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[967]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03794_),
    .QN(_00623_),
    .RESETN(net1745),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[968]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03795_),
    .QN(_00653_),
    .RESETN(net1746),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[969]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03796_),
    .QN(_00683_),
    .RESETN(net1747),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[96]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03797_),
    .QN(_00382_),
    .RESETN(net1748),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[970]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03798_),
    .QN(_00713_),
    .RESETN(net1749),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[971]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03799_),
    .QN(_00743_),
    .RESETN(net1750),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[972]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03800_),
    .QN(_00373_),
    .RESETN(net1751),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[973]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03801_),
    .QN(_00811_),
    .RESETN(net1752),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[974]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03802_),
    .QN(_00843_),
    .RESETN(net1753),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[975]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03803_),
    .QN(_00875_),
    .RESETN(net1754),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[976]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03804_),
    .QN(_00907_),
    .RESETN(net1755),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[977]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03805_),
    .QN(_00939_),
    .RESETN(net1756),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[978]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03806_),
    .QN(_00971_),
    .RESETN(net1757),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[979]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03807_),
    .QN(_01003_),
    .RESETN(net1758),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[97]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03808_),
    .QN(_00415_),
    .RESETN(net1759),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[980]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03809_),
    .QN(_01035_),
    .RESETN(net1760),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[981]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03810_),
    .QN(_01067_),
    .RESETN(net1761),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[982]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03811_),
    .QN(_01099_),
    .RESETN(net1762),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[983]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03812_),
    .QN(_01131_),
    .RESETN(net1763),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[984]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03813_),
    .QN(_01163_),
    .RESETN(net1764),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[985]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03814_),
    .QN(_01195_),
    .RESETN(net1765),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[986]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03815_),
    .QN(_01227_),
    .RESETN(net1766),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[987]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03816_),
    .QN(_01259_),
    .RESETN(net1767),
    .SETN(net41));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[988]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03817_),
    .QN(_01291_),
    .RESETN(net1768),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[989]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03818_),
    .QN(_01323_),
    .RESETN(net1769),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[98]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03819_),
    .QN(_00446_),
    .RESETN(net1770),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[990]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03820_),
    .QN(_01355_),
    .RESETN(net1771),
    .SETN(net39));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[991]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03821_),
    .QN(_01387_),
    .RESETN(net1772),
    .SETN(net40));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[992]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03822_),
    .QN(_00410_),
    .RESETN(net1773),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[993]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03823_),
    .QN(_00443_),
    .RESETN(net1774),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[994]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03824_),
    .QN(_00474_),
    .RESETN(net1775),
    .SETN(net33));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[995]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03825_),
    .QN(_00504_),
    .RESETN(net1776),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[996]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03826_),
    .QN(_00534_),
    .RESETN(net1777),
    .SETN(net35));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[997]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03827_),
    .QN(_00564_),
    .RESETN(net1778),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[998]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03828_),
    .QN(_00594_),
    .RESETN(net1779),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[999]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03829_),
    .QN(_00624_),
    .RESETN(net1780),
    .SETN(net34));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[99]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03830_),
    .QN(_00476_),
    .RESETN(net1781),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.branch_set$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .D(\id_stage_i.branch_set_d ),
    .QN(_01764_),
    .RESETN(net1782),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_03831_),
    .QN(_01763_),
    .RESETN(net1783),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_03832_),
    .QN(_01762_),
    .RESETN(net1784),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_03833_),
    .QN(_01761_),
    .RESETN(net1785),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_03834_),
    .QN(_01760_),
    .RESETN(net1786),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.debug_mode_o$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_03835_),
    .QN(_00758_),
    .RESETN(net1787),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.exc_req_q$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .D(\id_stage_i.controller_i.exc_req_d ),
    .QN(_02200_),
    .RESETN(net1788),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.illegal_insn_q$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .D(\id_stage_i.controller_i.illegal_insn_d ),
    .QN(_01391_),
    .RESETN(net1789),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.load_err_q$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .D(\id_stage_i.controller_i.load_err_i ),
    .QN(_01759_),
    .RESETN(net1790),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.nmi_mode_o$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_03836_),
    .QN(_00334_),
    .RESETN(net1791),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.store_err_q$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .D(\id_stage_i.controller_i.store_err_i ),
    .QN(_01758_),
    .RESETN(net1792),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.id_fsm_q$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_03837_),
    .QN(_01757_),
    .RESETN(net1793),
    .SETN(net51));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03838_),
    .QN(_01756_),
    .RESETN(net1794),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03839_),
    .QN(_01755_),
    .RESETN(net1795),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03840_),
    .QN(_01754_),
    .RESETN(net1796),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03841_),
    .QN(_01753_),
    .RESETN(net1797),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03842_),
    .QN(_01752_),
    .RESETN(net1798),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03843_),
    .QN(_01751_),
    .RESETN(net1799),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03844_),
    .QN(_01750_),
    .RESETN(net1800),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03845_),
    .QN(_01749_),
    .RESETN(net1801),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03846_),
    .QN(_01748_),
    .RESETN(net1802),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03847_),
    .QN(_01747_),
    .RESETN(net1803),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03848_),
    .QN(_01746_),
    .RESETN(net1804),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03849_),
    .QN(_01745_),
    .RESETN(net1805),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03850_),
    .QN(_01744_),
    .RESETN(net1806),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03851_),
    .QN(_01743_),
    .RESETN(net1807),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03852_),
    .QN(_01742_),
    .RESETN(net1808),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03853_),
    .QN(_01741_),
    .RESETN(net1809),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03854_),
    .QN(_01740_),
    .RESETN(net1810),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03855_),
    .QN(_01739_),
    .RESETN(net1811),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03856_),
    .QN(_01738_),
    .RESETN(net1812),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03857_),
    .QN(_01737_),
    .RESETN(net1813),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03858_),
    .QN(_01736_),
    .RESETN(net1814),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03859_),
    .QN(_01735_),
    .RESETN(net1815),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03860_),
    .QN(_01734_),
    .RESETN(net1816),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03861_),
    .QN(_01733_),
    .RESETN(net1817),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03862_),
    .QN(_01732_),
    .RESETN(net1818),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[34]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03863_),
    .QN(_00062_),
    .RESETN(net1819),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[35]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03864_),
    .QN(_00097_),
    .RESETN(net1820),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[36]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03865_),
    .QN(_00100_),
    .RESETN(net1821),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[37]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03866_),
    .QN(_00104_),
    .RESETN(net1822),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[38]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03867_),
    .QN(_00109_),
    .RESETN(net1823),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[39]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03868_),
    .QN(_00114_),
    .RESETN(net1824),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03869_),
    .QN(_01731_),
    .RESETN(net1825),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[40]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03870_),
    .QN(_00121_),
    .RESETN(net1826),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[41]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03871_),
    .QN(_00128_),
    .RESETN(net1827),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[42]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03872_),
    .QN(_00135_),
    .RESETN(net1828),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[43]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03873_),
    .QN(_00144_),
    .RESETN(net1829),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[44]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03874_),
    .QN(_00152_),
    .RESETN(net1830),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[45]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03875_),
    .QN(_00160_),
    .RESETN(net1831),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[46]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03876_),
    .QN(_00168_),
    .RESETN(net1832),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[47]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03877_),
    .QN(_00175_),
    .RESETN(net1833),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[48]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_03878_),
    .QN(_00180_),
    .RESETN(net1834),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[49]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03879_),
    .QN(_00187_),
    .RESETN(net1835),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03880_),
    .QN(_01730_),
    .RESETN(net1836),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[50]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03881_),
    .QN(_00063_),
    .RESETN(net1837),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[51]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_03882_),
    .QN(_00098_),
    .RESETN(net1838),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[52]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_03883_),
    .QN(_00101_),
    .RESETN(net1839),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[53]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_03884_),
    .QN(_00105_),
    .RESETN(net1840),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[54]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_03885_),
    .QN(_00110_),
    .RESETN(net1841),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[55]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03886_),
    .QN(_00115_),
    .RESETN(net1842),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[56]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03887_),
    .QN(_00122_),
    .RESETN(net1843),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[57]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_03888_),
    .QN(_00129_),
    .RESETN(net1844),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[58]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03889_),
    .QN(_00136_),
    .RESETN(net1845),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[59]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03890_),
    .QN(_00145_),
    .RESETN(net1846),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03891_),
    .QN(_01729_),
    .RESETN(net1847),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[60]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03892_),
    .QN(_00153_),
    .RESETN(net1848),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[61]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03893_),
    .QN(_00161_),
    .RESETN(net1849),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[62]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03894_),
    .QN(_00169_),
    .RESETN(net1850),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[63]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03895_),
    .QN(_00176_),
    .RESETN(net1851),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[64]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03896_),
    .QN(_00181_),
    .RESETN(net1852),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[65]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03897_),
    .QN(_00029_),
    .RESETN(net1853),
    .SETN(net44));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[66]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_03898_),
    .QN(_01728_),
    .RESETN(net1854),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[67]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_03899_),
    .QN(_00205_),
    .RESETN(net1855),
    .SETN(net45));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03900_),
    .QN(_01727_),
    .RESETN(net1856),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03901_),
    .QN(_01726_),
    .RESETN(net1857),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_03902_),
    .QN(_01725_),
    .RESETN(net1858),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_03903_),
    .QN(_02201_),
    .RESETN(net1859),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ),
    .QN(_02202_),
    .RESETN(net1860),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ),
    .QN(_02203_),
    .RESETN(net1861),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .QN(_01724_),
    .RESETN(net1862),
    .SETN(net169));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03904_),
    .QN(_01723_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03905_),
    .QN(_01722_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03906_),
    .QN(_01721_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03907_),
    .QN(_01720_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03908_),
    .QN(_01719_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03909_),
    .QN(_01718_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03910_),
    .QN(_01717_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03911_),
    .QN(_01716_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03912_),
    .QN(_01715_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03913_),
    .QN(_01714_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03914_),
    .QN(_01713_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03915_),
    .QN(_01712_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03916_),
    .QN(_01711_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03917_),
    .QN(_01710_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03918_),
    .QN(_01709_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03919_),
    .QN(_01708_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03920_),
    .QN(_01707_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03921_),
    .QN(_01706_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03922_),
    .QN(_01705_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03923_),
    .QN(_01704_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03924_),
    .QN(_01703_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03925_),
    .QN(_01702_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03926_),
    .QN(_01701_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03927_),
    .QN(_01700_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03928_),
    .QN(_01699_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03929_),
    .QN(_01698_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03930_),
    .QN(_01697_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03931_),
    .QN(_01696_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03932_),
    .QN(_01695_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03933_),
    .QN(_01694_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03934_),
    .QN(_01693_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03935_),
    .QN(_01692_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03936_),
    .QN(_01691_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[0]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03937_),
    .QN(_00750_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[10]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03938_),
    .QN(_01690_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[11]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03939_),
    .QN(_01689_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[12]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03940_),
    .QN(_01688_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[13]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03941_),
    .QN(_01687_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[14]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03942_),
    .QN(_01686_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[15]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03943_),
    .QN(_01685_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[16]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03944_),
    .QN(_01684_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[17]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03945_),
    .QN(_00023_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[18]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03946_),
    .QN(_01683_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[19]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03947_),
    .QN(_01682_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[1]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03948_),
    .QN(_17997_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[20]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03949_),
    .QN(_01681_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[21]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03950_),
    .QN(_01680_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[22]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03951_),
    .QN(_01679_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[23]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03952_),
    .QN(_01678_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[24]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03953_),
    .QN(_01677_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[25]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03954_),
    .QN(_01676_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[26]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03955_),
    .QN(_01675_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[27]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03956_),
    .QN(_01674_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[28]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03957_),
    .QN(_01673_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[29]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03958_),
    .QN(_01672_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03959_),
    .QN(_00021_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[30]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03960_),
    .QN(_01671_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[3]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03961_),
    .QN(_01670_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[4]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03962_),
    .QN(_01669_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[5]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03963_),
    .QN(_01668_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[6]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03964_),
    .QN(_01667_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[7]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03965_),
    .QN(_01666_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[8]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03966_),
    .QN(_01665_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[9]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_03967_),
    .QN(_00022_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03968_),
    .QN(_01664_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03969_),
    .QN(_01663_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03970_),
    .QN(_01662_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03971_),
    .QN(_01661_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03972_),
    .QN(_01660_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03973_),
    .QN(_01659_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03974_),
    .QN(_01658_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03975_),
    .QN(_01657_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03976_),
    .QN(_01656_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03977_),
    .QN(_01655_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03978_),
    .QN(_01654_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03979_),
    .QN(_01653_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03980_),
    .QN(_01652_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03981_),
    .QN(_01651_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03982_),
    .QN(_01650_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03983_),
    .QN(_01649_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03984_),
    .QN(_01648_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03985_),
    .QN(_01647_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03986_),
    .QN(_01646_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03987_),
    .QN(_01645_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03988_),
    .QN(_01644_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03989_),
    .QN(_01643_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03990_),
    .QN(_01642_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03991_),
    .QN(_01641_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03992_),
    .QN(_01640_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03993_),
    .QN(_01639_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03994_),
    .QN(_01638_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03995_),
    .QN(_01637_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03996_),
    .QN(_01636_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03997_),
    .QN(_01635_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03998_),
    .QN(_01634_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03999_),
    .QN(_01633_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04000_),
    .QN(_01632_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04001_),
    .QN(_01631_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04002_),
    .QN(_01630_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04003_),
    .QN(_01629_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04004_),
    .QN(_01628_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04005_),
    .QN(_01627_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04006_),
    .QN(_01626_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04007_),
    .QN(_01625_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04008_),
    .QN(_01624_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04009_),
    .QN(_01623_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04010_),
    .QN(_01622_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04011_),
    .QN(_01621_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04012_),
    .QN(_01620_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04013_),
    .QN(_01619_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04014_),
    .QN(_01618_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04015_),
    .QN(_01617_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04016_),
    .QN(_01616_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04017_),
    .QN(_01615_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04018_),
    .QN(_01614_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04019_),
    .QN(_01613_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04020_),
    .QN(_01612_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04021_),
    .QN(_01611_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04022_),
    .QN(_01610_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04023_),
    .QN(_01609_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04024_),
    .QN(_01608_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04025_),
    .QN(_01607_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04026_),
    .QN(_01606_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04027_),
    .QN(_01605_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04028_),
    .QN(_01604_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04029_),
    .QN(_01603_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04030_),
    .QN(_01602_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04031_),
    .QN(_01601_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04032_),
    .QN(_01600_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04033_),
    .QN(_01599_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04034_),
    .QN(_01598_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04035_),
    .QN(_01597_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04036_),
    .QN(_01596_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04037_),
    .QN(_01595_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04038_),
    .QN(_01594_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04039_),
    .QN(_01593_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04040_),
    .QN(_01592_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04041_),
    .QN(_01591_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04042_),
    .QN(_01590_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04043_),
    .QN(_01589_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04044_),
    .QN(_01588_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04045_),
    .QN(_01587_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04046_),
    .QN(_01586_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04047_),
    .QN(_01585_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04048_),
    .QN(_01584_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04049_),
    .QN(_01583_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04050_),
    .QN(_01582_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04051_),
    .QN(_01581_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04052_),
    .QN(_01580_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04053_),
    .QN(_01579_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04054_),
    .QN(_01578_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04055_),
    .QN(_01577_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04056_),
    .QN(_01576_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04057_),
    .QN(_01575_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04058_),
    .QN(_01574_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04059_),
    .QN(_01573_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04060_),
    .QN(_01572_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04061_),
    .QN(_01571_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04062_),
    .QN(_01570_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04063_),
    .QN(_02204_));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ),
    .QN(_00263_),
    .RESETN(net1863),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ),
    .QN(_00262_),
    .RESETN(net1864),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ),
    .QN(_02205_),
    .RESETN(net1865),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ),
    .QN(_02206_),
    .RESETN(net1866),
    .SETN(net169));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ),
    .QN(_00261_),
    .RESETN(net1867),
    .SETN(net169));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04064_),
    .QN(_01569_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04065_),
    .QN(_01568_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04066_),
    .QN(_01567_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04067_),
    .QN(_01566_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04068_),
    .QN(_01565_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04069_),
    .QN(_01564_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04070_),
    .QN(_01563_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04071_),
    .QN(_01562_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04072_),
    .QN(_01561_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04073_),
    .QN(_01560_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04074_),
    .QN(_01559_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04075_),
    .QN(_01558_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04076_),
    .QN(_01557_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04077_),
    .QN(_01556_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04078_),
    .QN(_01555_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04079_),
    .QN(_01554_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04080_),
    .QN(_01553_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04081_),
    .QN(_01552_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04082_),
    .QN(_01551_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04083_),
    .QN(_01550_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04084_),
    .QN(_01549_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04085_),
    .QN(_01548_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04086_),
    .QN(_01547_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04087_),
    .QN(_01546_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04088_),
    .QN(_01545_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04089_),
    .QN(_01544_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04090_),
    .QN(_01543_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_04091_),
    .QN(_01542_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04092_),
    .QN(_01541_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_04093_),
    .QN(_02207_));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ),
    .QN(_00260_),
    .RESETN(net1868),
    .SETN(net169));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.illegal_c_insn_id_o$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04094_),
    .QN(_01540_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_fetch_err_o$_DFFE_PN_  (.CLK(clknet_leaf_9_clk),
    .D(_04095_),
    .QN(_01539_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_fetch_err_plus2_o$_SDFFCE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .D(_04096_),
    .QN(_01538_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_is_compressed_id_o$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04097_),
    .QN(_00444_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[0]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04098_),
    .QN(_01537_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[10]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04099_),
    .QN(_01536_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[11]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04100_),
    .QN(_01535_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[12]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04101_),
    .QN(_01534_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[13]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04102_),
    .QN(_01533_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[14]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04103_),
    .QN(_01532_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[15]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04104_),
    .QN(_01531_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[1]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04105_),
    .QN(_01530_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[2]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04106_),
    .QN(_01529_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[3]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04107_),
    .QN(_01528_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[4]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04108_),
    .QN(_01527_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[5]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04109_),
    .QN(_01526_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[6]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04110_),
    .QN(_01525_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[7]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04111_),
    .QN(_01524_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[8]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04112_),
    .QN(_01523_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[9]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04113_),
    .QN(_01522_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[0]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04114_),
    .QN(_01521_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[10]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04115_),
    .QN(_01520_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[11]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04116_),
    .QN(_00339_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[12]$_DFFE_PN_  (.CLK(clknet_leaf_18_clk),
    .D(_04117_),
    .QN(_01519_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[13]$_DFFE_PN_  (.CLK(clknet_leaf_18_clk),
    .D(_04118_),
    .QN(_00413_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[14]$_DFFE_PN_  (.CLK(clknet_leaf_18_clk),
    .D(_04119_),
    .QN(_00377_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[15]$_DFFE_PN_  (.CLK(clknet_leaf_21_clk),
    .D(_04120_),
    .QN(_00344_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[16]$_DFFE_PN_  (.CLK(clknet_leaf_21_clk),
    .D(_04121_),
    .QN(_00343_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[17]$_DFFE_PN_  (.CLK(clknet_leaf_21_clk),
    .D(_04122_),
    .QN(_00342_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[18]$_DFFE_PN_  (.CLK(clknet_leaf_21_clk),
    .D(_04123_),
    .QN(_00341_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[19]$_DFFE_PN_  (.CLK(clknet_leaf_21_clk),
    .D(_04124_),
    .QN(_00340_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[1]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04125_),
    .QN(_01518_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[20]$_DFFE_PN_  (.CLK(clknet_leaf_22_clk),
    .D(_04126_),
    .QN(_00380_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[21]$_DFFE_PN_  (.CLK(clknet_leaf_22_clk),
    .D(_04127_),
    .QN(_01517_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[22]$_DFFE_PN_  (.CLK(clknet_leaf_21_clk),
    .D(_04128_),
    .QN(_01516_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[23]$_DFFE_PN_  (.CLK(clknet_leaf_21_clk),
    .D(_04129_),
    .QN(_00379_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[24]$_DFFE_PN_  (.CLK(clknet_leaf_21_clk),
    .D(_04130_),
    .QN(_00378_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[25]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04131_),
    .QN(_01515_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[26]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04132_),
    .QN(_00411_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[27]$_DFFE_PN_  (.CLK(clknet_leaf_1_clk),
    .D(_04133_),
    .QN(_01514_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[28]$_DFFE_PN_  (.CLK(clknet_leaf_1_clk),
    .D(_04134_),
    .QN(_01513_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[29]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04135_),
    .QN(_01512_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[2]$_DFFE_PN_  (.CLK(clknet_leaf_9_clk),
    .D(_04136_),
    .QN(_01511_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[30]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04137_),
    .QN(_01510_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[31]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04138_),
    .QN(_00412_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[3]$_DFFE_PN_  (.CLK(clknet_leaf_9_clk),
    .D(_04139_),
    .QN(_01509_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[4]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04140_),
    .QN(_01508_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[5]$_DFFE_PN_  (.CLK(clknet_leaf_9_clk),
    .D(_04141_),
    .QN(_01507_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[6]$_DFFE_PN_  (.CLK(clknet_leaf_9_clk),
    .D(_04142_),
    .QN(_00376_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[7]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04143_),
    .QN(_01506_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[8]$_DFFE_PN_  (.CLK(clknet_leaf_9_clk),
    .D(_04144_),
    .QN(_01505_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.instr_rdata_id_o[9]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04145_),
    .QN(_02208_));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.instr_valid_id_o$_DFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .D(\if_stage_i.instr_valid_id_d ),
    .QN(_00760_),
    .RESETN(net1869),
    .SETN(net51));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[10]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04146_),
    .QN(_00019_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[11]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04147_),
    .QN(_01504_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[12]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04148_),
    .QN(_01503_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[13]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04149_),
    .QN(_01502_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[14]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04150_),
    .QN(_01501_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[15]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04151_),
    .QN(_01500_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[16]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04152_),
    .QN(_01499_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[17]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04153_),
    .QN(_01498_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[18]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04154_),
    .QN(_00020_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[19]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04155_),
    .QN(_01497_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[1]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04156_),
    .QN(_01496_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[20]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04157_),
    .QN(_01495_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[21]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04158_),
    .QN(_01494_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[22]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04159_),
    .QN(_01493_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[23]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04160_),
    .QN(_01492_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[24]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04161_),
    .QN(_01491_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[25]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04162_),
    .QN(_01490_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[26]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04163_),
    .QN(_01489_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[27]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04164_),
    .QN(_01488_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[28]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04165_),
    .QN(_01487_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[29]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04166_),
    .QN(_01486_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[2]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04167_),
    .QN(_00016_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[30]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04168_),
    .QN(_01485_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[31]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04169_),
    .QN(_01484_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[3]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04170_),
    .QN(_00018_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[4]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04171_),
    .QN(_01483_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[5]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04172_),
    .QN(_01482_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[6]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04173_),
    .QN(_01481_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.pc_id_o[7]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04174_),
    .QN(_01480_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[8]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04175_),
    .QN(_01479_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.pc_id_o[9]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .D(_04176_),
    .QN(_01478_));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04177_),
    .QN(_01477_),
    .RESETN(net1870),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_04178_),
    .QN(_01476_),
    .RESETN(net1871),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_04179_),
    .QN(_01475_),
    .RESETN(net1872),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04180_),
    .QN(_01474_),
    .RESETN(net1873),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04181_),
    .QN(_01473_),
    .RESETN(net1874),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04182_),
    .QN(_01472_),
    .RESETN(net1875),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04183_),
    .QN(_01471_),
    .RESETN(net1876),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04184_),
    .QN(_01470_),
    .RESETN(net1877),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04185_),
    .QN(_01469_),
    .RESETN(net1878),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04186_),
    .QN(_01468_),
    .RESETN(net1879),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04187_),
    .QN(_01467_),
    .RESETN(net1880),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04188_),
    .QN(_01466_),
    .RESETN(net1881),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04189_),
    .QN(_01465_),
    .RESETN(net1882),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04190_),
    .QN(_01464_),
    .RESETN(net1883),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04191_),
    .QN(_01463_),
    .RESETN(net1884),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04192_),
    .QN(_01462_),
    .RESETN(net1885),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04193_),
    .QN(_01461_),
    .RESETN(net1886),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04194_),
    .QN(_01460_),
    .RESETN(net1887),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04195_),
    .QN(_01459_),
    .RESETN(net1888),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04196_),
    .QN(_01458_),
    .RESETN(net1889),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04197_),
    .QN(_01457_),
    .RESETN(net1890),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04198_),
    .QN(_01456_),
    .RESETN(net1891),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_04199_),
    .QN(_01455_),
    .RESETN(net1892),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04200_),
    .QN(_01454_),
    .RESETN(net1893),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04201_),
    .QN(_01453_),
    .RESETN(net1894),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_04202_),
    .QN(_01452_),
    .RESETN(net1895),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04203_),
    .QN(_01451_),
    .RESETN(net1896),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_04204_),
    .QN(_01450_),
    .RESETN(net1897),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04205_),
    .QN(_01449_),
    .RESETN(net1898),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_04206_),
    .QN(_01448_),
    .RESETN(net1899),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_04207_),
    .QN(_01447_),
    .RESETN(net1900),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_04208_),
    .QN(_01446_),
    .RESETN(net1901),
    .SETN(net52));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.data_sign_ext_q$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04209_),
    .QN(_01445_),
    .RESETN(net1902),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.data_we_q$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04210_),
    .QN(_01393_),
    .RESETN(net1903),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.handle_misaligned_q$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_04211_),
    .QN(_18707_),
    .RESETN(net1904),
    .SETN(net38));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_04212_),
    .QN(_01444_),
    .RESETN(net1905),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_04213_),
    .QN(_01443_),
    .RESETN(net1906),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04214_),
    .QN(_00375_),
    .RESETN(net1907),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.lsu_err_q$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04215_),
    .QN(_01442_),
    .RESETN(net1908),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_offset_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04216_),
    .QN(_01441_),
    .RESETN(net1909),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_offset_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04217_),
    .QN(_01440_),
    .RESETN(net1910),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04218_),
    .QN(_01439_),
    .RESETN(net1911),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04219_),
    .QN(_01438_),
    .RESETN(net1912),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04220_),
    .QN(_01437_),
    .RESETN(net1913),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04221_),
    .QN(_01436_),
    .RESETN(net1914),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04222_),
    .QN(_01435_),
    .RESETN(net1915),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04223_),
    .QN(_01434_),
    .RESETN(net1916),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04224_),
    .QN(_01433_),
    .RESETN(net1917),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04225_),
    .QN(_01432_),
    .RESETN(net1918),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04226_),
    .QN(_01431_),
    .RESETN(net1919),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04227_),
    .QN(_01430_),
    .RESETN(net1920),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04228_),
    .QN(_01429_),
    .RESETN(net1921),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04229_),
    .QN(_01428_),
    .RESETN(net1922),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04230_),
    .QN(_01427_),
    .RESETN(net1923),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04231_),
    .QN(_01426_),
    .RESETN(net1924),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04232_),
    .QN(_01425_),
    .RESETN(net1925),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04233_),
    .QN(_01424_),
    .RESETN(net1926),
    .SETN(net36));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04234_),
    .QN(_01423_),
    .RESETN(net1927),
    .SETN(net47));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04235_),
    .QN(_01422_),
    .RESETN(net1928),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04236_),
    .QN(_01421_),
    .RESETN(net1929),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04237_),
    .QN(_01420_),
    .RESETN(net1930),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04238_),
    .QN(_01419_),
    .RESETN(net1931),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04239_),
    .QN(_01418_),
    .RESETN(net1932),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04240_),
    .QN(_01417_),
    .RESETN(net1933),
    .SETN(net46));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_04241_),
    .QN(_01416_),
    .RESETN(net1934),
    .SETN(net46));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_Right_227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_Right_228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_Right_229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_Right_230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_Right_231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_Right_232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_Right_233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_Right_234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_Right_235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_Right_236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_Right_237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_Right_238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_Right_239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_Right_240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_Right_241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_Right_242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_Right_243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_Right_244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_Right_245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_Right_246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_Right_247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_Right_248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_Right_249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_Right_250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_Right_251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_Right_252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_Right_253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_Right_254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_Right_255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_Right_256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_Right_257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_Right_258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_Right_259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_Right_260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_Right_261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_Right_262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_Right_263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_Right_264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_Right_265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_Right_266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_Right_267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_Right_268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_Right_269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_Right_270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_Right_271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_Right_272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_Right_273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_Right_274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_Right_275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_Right_276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_Right_277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Left_333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Left_334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Left_335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Left_336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Left_337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Left_338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Left_339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Left_340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Left_341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Left_342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Left_343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Left_344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Left_345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Left_346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Left_347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Left_348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Left_349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Left_350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Left_351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Left_352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Left_353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Left_354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Left_355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Left_356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Left_357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Left_358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Left_359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Left_360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Left_361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Left_362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Left_363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Left_364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Left_365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Left_366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Left_367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Left_368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Left_369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Left_370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Left_371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Left_372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Left_373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Left_374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Left_375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Left_376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Left_377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Left_378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Left_379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Left_380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Left_381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Left_382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Left_383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Left_384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Left_385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Left_386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Left_387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Left_388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Left_389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Left_390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Left_391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Left_392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Left_393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Left_394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Left_395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Left_396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Left_397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Left_398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Left_399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Left_400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Left_401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Left_402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Left_403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Left_404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Left_405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Left_406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Left_407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Left_408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Left_409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Left_410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Left_411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Left_412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Left_413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Left_414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Left_415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Left_416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Left_417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Left_418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Left_419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Left_420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Left_421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Left_422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Left_423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Left_424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Left_425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Left_426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Left_427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Left_428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Left_429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_Left_430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_Left_431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_Left_432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_Left_433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_Left_434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_Left_435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_Left_436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_Left_437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_Left_438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_Left_439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Left_440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Left_441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Left_442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Left_443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Left_444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Left_445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Left_446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Left_447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Left_448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Left_449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Left_450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Left_451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_Left_452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_Left_453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_Left_454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_Left_455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Left_456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_Left_457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_Left_458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_Left_459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_Left_460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_Left_461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_Left_462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_Left_463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_Left_464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_Left_465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_Left_466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_Left_467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_Left_468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_Left_469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_Left_470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_Left_471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_Left_472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_Left_473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_Left_474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_Left_475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_Left_476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_Left_477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_Left_478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_Left_479 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_Left_480 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_Left_481 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_Left_482 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_Left_483 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_Left_484 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_Left_485 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_Left_486 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_Left_487 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_Left_488 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_Left_489 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_Left_490 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_Left_491 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_Left_492 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_Left_493 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_Left_494 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_Left_495 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_Left_496 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_Left_497 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_Left_498 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_Left_499 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_Left_500 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_Left_501 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_Left_502 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_Left_503 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_Left_504 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_Left_505 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_Left_506 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_Left_507 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_Left_508 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_Left_509 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_Left_510 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_Left_511 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_Left_512 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_Left_513 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_Left_514 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_Left_515 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_Left_516 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_Left_517 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_Left_518 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_Left_519 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_Left_520 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_Left_521 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_Left_522 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_Left_523 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_Left_524 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_Left_525 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_Left_526 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_Left_527 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_Left_528 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_Left_529 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_Left_530 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_Left_531 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_Left_532 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_Left_533 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_Left_534 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_Left_535 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_Left_536 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_Left_537 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_Left_538 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_Left_539 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_Left_540 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_Left_541 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_Left_542 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_Left_543 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_Left_544 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_Left_545 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_Left_546 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_Left_547 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_Left_548 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_Left_549 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_Left_550 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_Left_551 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_Left_552 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_Left_553 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_Left_554 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_Left_555 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_556 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_557 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_558 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_559 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_560 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_561 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_562 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_563 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_564 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_565 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_566 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_567 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_568 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_569 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_570 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_571 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_572 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_573 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_574 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_575 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_576 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_577 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_14_578 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_14_579 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_15_580 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_16_581 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_16_582 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_17_583 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_18_584 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_18_585 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_19_586 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_20_587 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_20_588 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_21_589 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_22_590 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_22_591 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_23_592 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_24_593 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_24_594 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_25_595 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_26_596 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_26_597 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_27_598 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_28_599 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_28_600 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_29_601 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_30_602 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_30_603 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_31_604 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_32_605 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_32_606 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_33_607 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_34_608 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_34_609 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_35_610 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_36_611 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_36_612 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_37_613 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_38_614 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_38_615 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_39_616 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_40_617 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_40_618 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_41_619 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_42_620 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_42_621 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_43_622 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_44_623 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_44_624 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_45_625 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_46_626 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_46_627 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_47_628 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_48_629 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_48_630 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_49_631 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_50_632 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_50_633 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_51_634 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_52_635 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_52_636 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_53_637 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_54_638 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_54_639 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_55_640 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_56_641 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_56_642 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_57_643 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_58_644 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_58_645 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_59_646 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_60_647 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_60_648 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_61_649 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_62_650 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_62_651 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_63_652 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_64_653 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_64_654 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_65_655 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_66_656 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_66_657 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_67_658 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_68_659 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_68_660 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_69_661 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_70_662 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_70_663 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_71_664 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_72_665 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_72_666 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_73_667 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_74_668 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_74_669 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_75_670 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_76_671 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_76_672 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_77_673 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_78_674 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_78_675 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_79_676 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_80_677 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_80_678 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_81_679 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_680 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_681 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_83_682 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_84_683 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_84_684 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_85_685 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_86_686 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_86_687 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_87_688 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_88_689 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_88_690 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_89_691 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_90_692 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_90_693 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_91_694 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_92_695 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_92_696 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_93_697 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_94_698 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_94_699 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_95_700 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_96_701 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_96_702 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_97_703 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_98_704 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_98_705 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_99_706 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_100_707 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_100_708 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_101_709 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_102_710 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_102_711 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_103_712 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_104_713 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_104_714 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_105_715 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_106_716 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_106_717 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_107_718 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_108_719 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_108_720 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_109_721 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_110_722 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_110_723 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_111_724 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_112_725 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_112_726 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_113_727 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_114_728 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_114_729 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_115_730 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_116_731 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_116_732 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_117_733 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_118_734 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_118_735 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_119_736 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_120_737 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_120_738 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_121_739 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_122_740 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_122_741 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_123_742 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_124_743 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_124_744 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_125_745 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_126_746 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_126_747 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_127_748 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_128_749 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_128_750 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_129_751 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_130_752 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_130_753 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_131_754 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_132_755 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_132_756 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_133_757 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_134_758 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_134_759 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_135_760 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_136_761 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_136_762 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_137_763 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_138_764 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_138_765 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_139_766 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_140_767 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_140_768 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_141_769 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_142_770 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_142_771 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_143_772 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_144_773 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_144_774 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_145_775 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_146_776 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_146_777 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_147_778 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_148_779 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_148_780 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_149_781 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_150_782 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_150_783 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_151_784 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_152_785 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_152_786 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_153_787 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_154_788 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_154_789 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_155_790 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_156_791 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_156_792 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_157_793 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_158_794 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_158_795 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_159_796 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_160_797 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_160_798 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_161_799 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_162_800 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_162_801 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_163_802 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_164_803 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_164_804 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_165_805 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_166_806 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_166_807 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_167_808 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_168_809 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_168_810 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_169_811 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_170_812 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_170_813 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_171_814 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_172_815 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_172_816 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_173_817 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_174_818 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_174_819 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_175_820 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_176_821 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_176_822 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_177_823 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_824 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_825 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_826 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_827 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_828 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_829 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_830 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_831 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_832 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_833 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_834 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_835 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_836 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_837 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_838 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_839 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_840 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_841 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_190_842 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_190_843 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_191_844 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_192_845 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_192_846 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_193_847 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_194_848 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_194_849 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_195_850 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_196_851 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_196_852 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_197_853 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_198_854 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_198_855 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_199_856 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_200_857 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_200_858 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_201_859 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_202_860 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_202_861 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_203_862 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_204_863 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_204_864 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_205_865 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_206_866 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_206_867 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_207_868 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_208_869 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_208_870 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_209_871 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_210_872 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_210_873 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_211_874 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_212_875 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_212_876 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_213_877 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_214_878 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_214_879 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_215_880 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_216_881 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_216_882 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_217_883 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_218_884 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_218_885 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_219_886 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_220_887 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_220_888 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_221_889 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_222_890 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_222_891 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_223_892 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_224_893 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_224_894 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_225_895 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_226_896 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_226_897 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_227_898 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_228_899 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_228_900 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_229_901 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_230_902 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_230_903 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_231_904 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_232_905 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_232_906 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_233_907 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_234_908 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_234_909 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_235_910 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_236_911 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_236_912 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_237_913 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_238_914 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_238_915 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_239_916 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_240_917 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_240_918 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_241_919 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_242_920 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_242_921 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_243_922 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_244_923 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_244_924 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_245_925 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_246_926 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_246_927 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_247_928 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_248_929 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_248_930 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_249_931 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_250_932 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_250_933 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_251_934 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_252_935 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_252_936 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_253_937 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_254_938 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_254_939 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_255_940 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_256_941 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_256_942 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_257_943 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_258_944 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_258_945 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_259_946 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_260_947 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_260_948 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_261_949 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_262_950 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_262_951 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_263_952 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_264_953 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_264_954 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_265_955 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_266_956 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_266_957 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_267_958 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_268_959 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_268_960 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_269_961 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_270_962 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_270_963 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_271_964 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_272_965 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_272_966 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_273_967 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_274_968 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_274_969 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_275_970 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_276_971 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_276_972 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_277_973 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_277_974 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_277_975 ();
 BUFx6f_ASAP7_75t_R load_slew32 (.A(_17564_),
    .Y(net32));
 BUFx12f_ASAP7_75t_R load_slew33 (.A(net37),
    .Y(net33));
 BUFx12f_ASAP7_75t_R load_slew34 (.A(net38),
    .Y(net34));
 BUFx12f_ASAP7_75t_R load_slew35 (.A(net38),
    .Y(net35));
 BUFx12f_ASAP7_75t_R load_slew36 (.A(net38),
    .Y(net36));
 BUFx12f_ASAP7_75t_R load_slew37 (.A(net38),
    .Y(net37));
 BUFx12f_ASAP7_75t_R load_slew38 (.A(net44),
    .Y(net38));
 BUFx12f_ASAP7_75t_R load_slew39 (.A(net40),
    .Y(net39));
 BUFx12f_ASAP7_75t_R load_slew40 (.A(net44),
    .Y(net40));
 BUFx12f_ASAP7_75t_R load_slew41 (.A(net42),
    .Y(net41));
 BUFx12f_ASAP7_75t_R load_slew42 (.A(net43),
    .Y(net42));
 BUFx12f_ASAP7_75t_R load_slew43 (.A(net44),
    .Y(net43));
 BUFx12f_ASAP7_75t_R load_slew44 (.A(net52),
    .Y(net44));
 BUFx12f_ASAP7_75t_R load_slew45 (.A(net52),
    .Y(net45));
 BUFx12f_ASAP7_75t_R load_slew46 (.A(net47),
    .Y(net46));
 BUFx12f_ASAP7_75t_R load_slew47 (.A(net50),
    .Y(net47));
 BUFx12f_ASAP7_75t_R load_slew48 (.A(net49),
    .Y(net48));
 BUFx12f_ASAP7_75t_R load_slew49 (.A(net50),
    .Y(net49));
 BUFx12f_ASAP7_75t_R load_slew50 (.A(net1963),
    .Y(net50));
 BUFx12f_ASAP7_75t_R load_slew51 (.A(net169),
    .Y(net51));
 BUFx12f_ASAP7_75t_R max_length52 (.A(net169),
    .Y(net52));
 BUFx3_ASAP7_75t_R input1 (.A(boot_addr_i[10]),
    .Y(net1));
 BUFx3_ASAP7_75t_R input2 (.A(boot_addr_i[11]),
    .Y(net2));
 BUFx3_ASAP7_75t_R input3 (.A(boot_addr_i[12]),
    .Y(net3));
 BUFx3_ASAP7_75t_R input4 (.A(boot_addr_i[13]),
    .Y(net4));
 BUFx3_ASAP7_75t_R input5 (.A(boot_addr_i[14]),
    .Y(net5));
 BUFx3_ASAP7_75t_R input6 (.A(boot_addr_i[15]),
    .Y(net6));
 BUFx3_ASAP7_75t_R input7 (.A(boot_addr_i[16]),
    .Y(net7));
 BUFx3_ASAP7_75t_R input8 (.A(boot_addr_i[17]),
    .Y(net8));
 BUFx3_ASAP7_75t_R input9 (.A(boot_addr_i[18]),
    .Y(net9));
 BUFx3_ASAP7_75t_R input10 (.A(boot_addr_i[19]),
    .Y(net10));
 BUFx3_ASAP7_75t_R input11 (.A(boot_addr_i[20]),
    .Y(net11));
 BUFx3_ASAP7_75t_R input12 (.A(boot_addr_i[21]),
    .Y(net12));
 BUFx3_ASAP7_75t_R input13 (.A(boot_addr_i[22]),
    .Y(net13));
 BUFx3_ASAP7_75t_R input14 (.A(boot_addr_i[23]),
    .Y(net14));
 BUFx3_ASAP7_75t_R input15 (.A(boot_addr_i[24]),
    .Y(net15));
 BUFx3_ASAP7_75t_R input16 (.A(boot_addr_i[25]),
    .Y(net16));
 BUFx3_ASAP7_75t_R input17 (.A(boot_addr_i[26]),
    .Y(net17));
 BUFx3_ASAP7_75t_R input18 (.A(boot_addr_i[27]),
    .Y(net18));
 BUFx3_ASAP7_75t_R input19 (.A(boot_addr_i[28]),
    .Y(net19));
 BUFx3_ASAP7_75t_R input20 (.A(boot_addr_i[29]),
    .Y(net20));
 BUFx3_ASAP7_75t_R input21 (.A(boot_addr_i[30]),
    .Y(net21));
 BUFx3_ASAP7_75t_R input22 (.A(boot_addr_i[31]),
    .Y(net22));
 BUFx3_ASAP7_75t_R input23 (.A(boot_addr_i[8]),
    .Y(net23));
 BUFx3_ASAP7_75t_R input24 (.A(boot_addr_i[9]),
    .Y(net24));
 BUFx3_ASAP7_75t_R input25 (.A(data_err_i),
    .Y(net25));
 BUFx6f_ASAP7_75t_R input26 (.A(data_gnt_i),
    .Y(net26));
 BUFx3_ASAP7_75t_R input27 (.A(data_rdata_i[0]),
    .Y(net27));
 BUFx3_ASAP7_75t_R input28 (.A(data_rdata_i[10]),
    .Y(net28));
 BUFx3_ASAP7_75t_R input29 (.A(data_rdata_i[11]),
    .Y(net29));
 BUFx3_ASAP7_75t_R input30 (.A(data_rdata_i[12]),
    .Y(net30));
 BUFx3_ASAP7_75t_R input31 (.A(data_rdata_i[13]),
    .Y(net31));
 BUFx3_ASAP7_75t_R input32 (.A(data_rdata_i[14]),
    .Y(net53));
 BUFx3_ASAP7_75t_R input33 (.A(data_rdata_i[15]),
    .Y(net54));
 BUFx3_ASAP7_75t_R input34 (.A(data_rdata_i[16]),
    .Y(net55));
 BUFx3_ASAP7_75t_R input35 (.A(data_rdata_i[17]),
    .Y(net56));
 BUFx3_ASAP7_75t_R input36 (.A(data_rdata_i[18]),
    .Y(net57));
 BUFx3_ASAP7_75t_R input37 (.A(data_rdata_i[19]),
    .Y(net58));
 BUFx3_ASAP7_75t_R input38 (.A(data_rdata_i[1]),
    .Y(net59));
 BUFx3_ASAP7_75t_R input39 (.A(data_rdata_i[20]),
    .Y(net60));
 BUFx3_ASAP7_75t_R input40 (.A(data_rdata_i[21]),
    .Y(net61));
 BUFx3_ASAP7_75t_R input41 (.A(data_rdata_i[22]),
    .Y(net62));
 BUFx3_ASAP7_75t_R input42 (.A(data_rdata_i[23]),
    .Y(net63));
 BUFx3_ASAP7_75t_R input43 (.A(data_rdata_i[24]),
    .Y(net64));
 BUFx3_ASAP7_75t_R input44 (.A(data_rdata_i[25]),
    .Y(net65));
 BUFx3_ASAP7_75t_R input45 (.A(data_rdata_i[26]),
    .Y(net66));
 BUFx3_ASAP7_75t_R input46 (.A(data_rdata_i[27]),
    .Y(net67));
 BUFx3_ASAP7_75t_R input47 (.A(data_rdata_i[28]),
    .Y(net68));
 BUFx3_ASAP7_75t_R input48 (.A(data_rdata_i[29]),
    .Y(net69));
 BUFx3_ASAP7_75t_R input49 (.A(data_rdata_i[2]),
    .Y(net70));
 BUFx3_ASAP7_75t_R input50 (.A(data_rdata_i[30]),
    .Y(net71));
 BUFx3_ASAP7_75t_R input51 (.A(data_rdata_i[31]),
    .Y(net72));
 BUFx3_ASAP7_75t_R input52 (.A(data_rdata_i[3]),
    .Y(net73));
 BUFx3_ASAP7_75t_R input53 (.A(data_rdata_i[4]),
    .Y(net74));
 BUFx3_ASAP7_75t_R input54 (.A(data_rdata_i[5]),
    .Y(net75));
 BUFx3_ASAP7_75t_R input55 (.A(data_rdata_i[6]),
    .Y(net76));
 BUFx3_ASAP7_75t_R input56 (.A(data_rdata_i[7]),
    .Y(net77));
 BUFx3_ASAP7_75t_R input57 (.A(data_rdata_i[8]),
    .Y(net78));
 BUFx3_ASAP7_75t_R input58 (.A(data_rdata_i[9]),
    .Y(net79));
 BUFx6f_ASAP7_75t_R input59 (.A(data_rvalid_i),
    .Y(net80));
 BUFx6f_ASAP7_75t_R input60 (.A(debug_req_i),
    .Y(net81));
 BUFx3_ASAP7_75t_R input61 (.A(fetch_enable_i),
    .Y(net82));
 BUFx3_ASAP7_75t_R input62 (.A(hart_id_i[0]),
    .Y(net83));
 BUFx3_ASAP7_75t_R input63 (.A(hart_id_i[10]),
    .Y(net84));
 BUFx3_ASAP7_75t_R input64 (.A(hart_id_i[11]),
    .Y(net85));
 BUFx3_ASAP7_75t_R input65 (.A(hart_id_i[12]),
    .Y(net86));
 BUFx3_ASAP7_75t_R input66 (.A(hart_id_i[13]),
    .Y(net87));
 BUFx3_ASAP7_75t_R input67 (.A(hart_id_i[14]),
    .Y(net88));
 BUFx3_ASAP7_75t_R input68 (.A(hart_id_i[15]),
    .Y(net89));
 BUFx3_ASAP7_75t_R input69 (.A(hart_id_i[16]),
    .Y(net90));
 BUFx3_ASAP7_75t_R input70 (.A(hart_id_i[17]),
    .Y(net91));
 BUFx3_ASAP7_75t_R input71 (.A(hart_id_i[18]),
    .Y(net92));
 BUFx3_ASAP7_75t_R input72 (.A(hart_id_i[19]),
    .Y(net93));
 BUFx3_ASAP7_75t_R input73 (.A(hart_id_i[1]),
    .Y(net94));
 BUFx3_ASAP7_75t_R input74 (.A(hart_id_i[20]),
    .Y(net95));
 BUFx3_ASAP7_75t_R input75 (.A(hart_id_i[21]),
    .Y(net96));
 BUFx3_ASAP7_75t_R input76 (.A(hart_id_i[22]),
    .Y(net97));
 BUFx3_ASAP7_75t_R input77 (.A(hart_id_i[23]),
    .Y(net98));
 BUFx3_ASAP7_75t_R input78 (.A(hart_id_i[24]),
    .Y(net99));
 BUFx3_ASAP7_75t_R input79 (.A(hart_id_i[25]),
    .Y(net100));
 BUFx3_ASAP7_75t_R input80 (.A(hart_id_i[26]),
    .Y(net101));
 BUFx3_ASAP7_75t_R input81 (.A(hart_id_i[27]),
    .Y(net102));
 BUFx3_ASAP7_75t_R input82 (.A(hart_id_i[28]),
    .Y(net103));
 BUFx3_ASAP7_75t_R input83 (.A(hart_id_i[29]),
    .Y(net104));
 BUFx3_ASAP7_75t_R input84 (.A(hart_id_i[2]),
    .Y(net105));
 BUFx3_ASAP7_75t_R input85 (.A(hart_id_i[30]),
    .Y(net106));
 BUFx3_ASAP7_75t_R input86 (.A(hart_id_i[31]),
    .Y(net107));
 BUFx3_ASAP7_75t_R input87 (.A(hart_id_i[3]),
    .Y(net108));
 BUFx3_ASAP7_75t_R input88 (.A(hart_id_i[4]),
    .Y(net109));
 BUFx3_ASAP7_75t_R input89 (.A(hart_id_i[5]),
    .Y(net110));
 BUFx3_ASAP7_75t_R input90 (.A(hart_id_i[6]),
    .Y(net111));
 BUFx3_ASAP7_75t_R input91 (.A(hart_id_i[7]),
    .Y(net112));
 BUFx3_ASAP7_75t_R input92 (.A(hart_id_i[8]),
    .Y(net113));
 BUFx3_ASAP7_75t_R input93 (.A(hart_id_i[9]),
    .Y(net114));
 BUFx3_ASAP7_75t_R input94 (.A(instr_err_i),
    .Y(net115));
 BUFx3_ASAP7_75t_R input95 (.A(instr_gnt_i),
    .Y(net116));
 BUFx3_ASAP7_75t_R input96 (.A(instr_rdata_i[0]),
    .Y(net117));
 BUFx3_ASAP7_75t_R input97 (.A(instr_rdata_i[10]),
    .Y(net118));
 BUFx3_ASAP7_75t_R input98 (.A(instr_rdata_i[11]),
    .Y(net119));
 BUFx3_ASAP7_75t_R input99 (.A(instr_rdata_i[12]),
    .Y(net120));
 BUFx3_ASAP7_75t_R input100 (.A(instr_rdata_i[13]),
    .Y(net121));
 BUFx3_ASAP7_75t_R input101 (.A(instr_rdata_i[14]),
    .Y(net122));
 BUFx3_ASAP7_75t_R input102 (.A(instr_rdata_i[15]),
    .Y(net123));
 BUFx6f_ASAP7_75t_R input103 (.A(instr_rdata_i[16]),
    .Y(net124));
 BUFx6f_ASAP7_75t_R input104 (.A(instr_rdata_i[17]),
    .Y(net125));
 BUFx3_ASAP7_75t_R input105 (.A(instr_rdata_i[18]),
    .Y(net126));
 BUFx3_ASAP7_75t_R input106 (.A(instr_rdata_i[19]),
    .Y(net127));
 BUFx3_ASAP7_75t_R input107 (.A(instr_rdata_i[1]),
    .Y(net128));
 BUFx3_ASAP7_75t_R input108 (.A(instr_rdata_i[20]),
    .Y(net129));
 BUFx3_ASAP7_75t_R input109 (.A(instr_rdata_i[21]),
    .Y(net130));
 BUFx3_ASAP7_75t_R input110 (.A(instr_rdata_i[22]),
    .Y(net131));
 BUFx3_ASAP7_75t_R input111 (.A(instr_rdata_i[23]),
    .Y(net132));
 BUFx3_ASAP7_75t_R input112 (.A(instr_rdata_i[24]),
    .Y(net133));
 BUFx3_ASAP7_75t_R input113 (.A(instr_rdata_i[25]),
    .Y(net134));
 BUFx3_ASAP7_75t_R input114 (.A(instr_rdata_i[26]),
    .Y(net135));
 BUFx3_ASAP7_75t_R input115 (.A(instr_rdata_i[27]),
    .Y(net136));
 BUFx3_ASAP7_75t_R input116 (.A(instr_rdata_i[28]),
    .Y(net137));
 BUFx3_ASAP7_75t_R input117 (.A(instr_rdata_i[29]),
    .Y(net138));
 BUFx3_ASAP7_75t_R input118 (.A(instr_rdata_i[2]),
    .Y(net139));
 BUFx3_ASAP7_75t_R input119 (.A(instr_rdata_i[30]),
    .Y(net140));
 BUFx3_ASAP7_75t_R input120 (.A(instr_rdata_i[31]),
    .Y(net141));
 BUFx3_ASAP7_75t_R input121 (.A(instr_rdata_i[3]),
    .Y(net142));
 BUFx3_ASAP7_75t_R input122 (.A(instr_rdata_i[4]),
    .Y(net143));
 BUFx3_ASAP7_75t_R input123 (.A(instr_rdata_i[5]),
    .Y(net144));
 BUFx3_ASAP7_75t_R input124 (.A(instr_rdata_i[6]),
    .Y(net145));
 BUFx3_ASAP7_75t_R input125 (.A(instr_rdata_i[7]),
    .Y(net146));
 BUFx6f_ASAP7_75t_R input126 (.A(instr_rdata_i[8]),
    .Y(net147));
 BUFx3_ASAP7_75t_R input127 (.A(instr_rdata_i[9]),
    .Y(net148));
 BUFx3_ASAP7_75t_R input128 (.A(instr_rvalid_i),
    .Y(net149));
 BUFx3_ASAP7_75t_R input129 (.A(irq_external_i),
    .Y(net150));
 BUFx3_ASAP7_75t_R input130 (.A(irq_fast_i[0]),
    .Y(net151));
 BUFx3_ASAP7_75t_R input131 (.A(irq_fast_i[10]),
    .Y(net152));
 BUFx3_ASAP7_75t_R input132 (.A(irq_fast_i[11]),
    .Y(net153));
 BUFx3_ASAP7_75t_R input133 (.A(irq_fast_i[12]),
    .Y(net154));
 BUFx3_ASAP7_75t_R input134 (.A(irq_fast_i[13]),
    .Y(net155));
 BUFx3_ASAP7_75t_R input135 (.A(irq_fast_i[14]),
    .Y(net156));
 BUFx3_ASAP7_75t_R input136 (.A(irq_fast_i[1]),
    .Y(net157));
 BUFx3_ASAP7_75t_R input137 (.A(irq_fast_i[2]),
    .Y(net158));
 BUFx3_ASAP7_75t_R input138 (.A(irq_fast_i[3]),
    .Y(net159));
 BUFx3_ASAP7_75t_R input139 (.A(irq_fast_i[4]),
    .Y(net160));
 BUFx3_ASAP7_75t_R input140 (.A(irq_fast_i[5]),
    .Y(net161));
 BUFx3_ASAP7_75t_R input141 (.A(irq_fast_i[6]),
    .Y(net162));
 BUFx3_ASAP7_75t_R input142 (.A(irq_fast_i[7]),
    .Y(net163));
 BUFx3_ASAP7_75t_R input143 (.A(irq_fast_i[8]),
    .Y(net164));
 BUFx3_ASAP7_75t_R input144 (.A(irq_fast_i[9]),
    .Y(net165));
 BUFx6f_ASAP7_75t_R input145 (.A(irq_nm_i),
    .Y(net166));
 BUFx3_ASAP7_75t_R input146 (.A(irq_software_i),
    .Y(net167));
 BUFx3_ASAP7_75t_R input147 (.A(irq_timer_i),
    .Y(net168));
 BUFx6f_ASAP7_75t_R input148 (.A(rst_ni),
    .Y(net169));
 BUFx3_ASAP7_75t_R input149 (.A(test_en_i),
    .Y(net170));
 BUFx3_ASAP7_75t_R output150 (.A(net171),
    .Y(core_sleep_o));
 BUFx3_ASAP7_75t_R output151 (.A(net172),
    .Y(data_addr_o[10]));
 BUFx3_ASAP7_75t_R output152 (.A(net173),
    .Y(data_addr_o[11]));
 BUFx3_ASAP7_75t_R output153 (.A(net174),
    .Y(data_addr_o[12]));
 BUFx3_ASAP7_75t_R output154 (.A(net175),
    .Y(data_addr_o[13]));
 BUFx3_ASAP7_75t_R output155 (.A(net176),
    .Y(data_addr_o[14]));
 BUFx3_ASAP7_75t_R output156 (.A(net177),
    .Y(data_addr_o[15]));
 BUFx3_ASAP7_75t_R output157 (.A(net178),
    .Y(data_addr_o[16]));
 BUFx3_ASAP7_75t_R output158 (.A(net179),
    .Y(data_addr_o[17]));
 BUFx3_ASAP7_75t_R output159 (.A(net180),
    .Y(data_addr_o[18]));
 BUFx3_ASAP7_75t_R output160 (.A(net181),
    .Y(data_addr_o[19]));
 BUFx3_ASAP7_75t_R output161 (.A(net182),
    .Y(data_addr_o[20]));
 BUFx3_ASAP7_75t_R output162 (.A(net183),
    .Y(data_addr_o[21]));
 BUFx3_ASAP7_75t_R output163 (.A(net184),
    .Y(data_addr_o[22]));
 BUFx3_ASAP7_75t_R output164 (.A(net185),
    .Y(data_addr_o[23]));
 BUFx3_ASAP7_75t_R output165 (.A(net186),
    .Y(data_addr_o[24]));
 BUFx3_ASAP7_75t_R output166 (.A(net187),
    .Y(data_addr_o[25]));
 BUFx3_ASAP7_75t_R output167 (.A(net188),
    .Y(data_addr_o[26]));
 BUFx3_ASAP7_75t_R output168 (.A(net189),
    .Y(data_addr_o[27]));
 BUFx3_ASAP7_75t_R output169 (.A(net190),
    .Y(data_addr_o[28]));
 BUFx3_ASAP7_75t_R output170 (.A(net191),
    .Y(data_addr_o[29]));
 BUFx3_ASAP7_75t_R output171 (.A(net192),
    .Y(data_addr_o[2]));
 BUFx3_ASAP7_75t_R output172 (.A(net193),
    .Y(data_addr_o[30]));
 BUFx3_ASAP7_75t_R output173 (.A(net194),
    .Y(data_addr_o[31]));
 BUFx3_ASAP7_75t_R output174 (.A(net195),
    .Y(data_addr_o[3]));
 BUFx3_ASAP7_75t_R output175 (.A(net196),
    .Y(data_addr_o[4]));
 BUFx3_ASAP7_75t_R output176 (.A(net197),
    .Y(data_addr_o[5]));
 BUFx3_ASAP7_75t_R output177 (.A(net198),
    .Y(data_addr_o[6]));
 BUFx3_ASAP7_75t_R output178 (.A(net199),
    .Y(data_addr_o[7]));
 BUFx3_ASAP7_75t_R output179 (.A(net200),
    .Y(data_addr_o[8]));
 BUFx3_ASAP7_75t_R output180 (.A(net201),
    .Y(data_addr_o[9]));
 BUFx3_ASAP7_75t_R output181 (.A(net202),
    .Y(data_be_o[0]));
 BUFx3_ASAP7_75t_R output182 (.A(net203),
    .Y(data_be_o[1]));
 BUFx3_ASAP7_75t_R output183 (.A(net204),
    .Y(data_be_o[2]));
 BUFx3_ASAP7_75t_R output184 (.A(net205),
    .Y(data_be_o[3]));
 BUFx3_ASAP7_75t_R output185 (.A(net206),
    .Y(data_req_o));
 BUFx3_ASAP7_75t_R output186 (.A(net207),
    .Y(data_wdata_o[0]));
 BUFx3_ASAP7_75t_R output187 (.A(net208),
    .Y(data_wdata_o[10]));
 BUFx3_ASAP7_75t_R output188 (.A(net209),
    .Y(data_wdata_o[11]));
 BUFx3_ASAP7_75t_R output189 (.A(net210),
    .Y(data_wdata_o[12]));
 BUFx3_ASAP7_75t_R output190 (.A(net211),
    .Y(data_wdata_o[13]));
 BUFx3_ASAP7_75t_R output191 (.A(net212),
    .Y(data_wdata_o[14]));
 BUFx3_ASAP7_75t_R output192 (.A(net213),
    .Y(data_wdata_o[15]));
 BUFx3_ASAP7_75t_R output193 (.A(net214),
    .Y(data_wdata_o[16]));
 BUFx3_ASAP7_75t_R output194 (.A(net215),
    .Y(data_wdata_o[17]));
 BUFx3_ASAP7_75t_R output195 (.A(net216),
    .Y(data_wdata_o[18]));
 BUFx3_ASAP7_75t_R output196 (.A(net217),
    .Y(data_wdata_o[19]));
 BUFx3_ASAP7_75t_R output197 (.A(net218),
    .Y(data_wdata_o[1]));
 BUFx3_ASAP7_75t_R output198 (.A(net219),
    .Y(data_wdata_o[20]));
 BUFx3_ASAP7_75t_R output199 (.A(net220),
    .Y(data_wdata_o[21]));
 BUFx3_ASAP7_75t_R output200 (.A(net221),
    .Y(data_wdata_o[22]));
 BUFx3_ASAP7_75t_R output201 (.A(net222),
    .Y(data_wdata_o[23]));
 BUFx3_ASAP7_75t_R output202 (.A(net223),
    .Y(data_wdata_o[24]));
 BUFx3_ASAP7_75t_R output203 (.A(net224),
    .Y(data_wdata_o[25]));
 BUFx3_ASAP7_75t_R output204 (.A(net225),
    .Y(data_wdata_o[26]));
 BUFx3_ASAP7_75t_R output205 (.A(net226),
    .Y(data_wdata_o[27]));
 BUFx3_ASAP7_75t_R output206 (.A(net227),
    .Y(data_wdata_o[28]));
 BUFx3_ASAP7_75t_R output207 (.A(net228),
    .Y(data_wdata_o[29]));
 BUFx3_ASAP7_75t_R output208 (.A(net229),
    .Y(data_wdata_o[2]));
 BUFx3_ASAP7_75t_R output209 (.A(net230),
    .Y(data_wdata_o[30]));
 BUFx3_ASAP7_75t_R output210 (.A(net231),
    .Y(data_wdata_o[31]));
 BUFx3_ASAP7_75t_R output211 (.A(net232),
    .Y(data_wdata_o[3]));
 BUFx3_ASAP7_75t_R output212 (.A(net233),
    .Y(data_wdata_o[4]));
 BUFx3_ASAP7_75t_R output213 (.A(net234),
    .Y(data_wdata_o[5]));
 BUFx3_ASAP7_75t_R output214 (.A(net235),
    .Y(data_wdata_o[6]));
 BUFx3_ASAP7_75t_R output215 (.A(net236),
    .Y(data_wdata_o[7]));
 BUFx3_ASAP7_75t_R output216 (.A(net237),
    .Y(data_wdata_o[8]));
 BUFx3_ASAP7_75t_R output217 (.A(net238),
    .Y(data_wdata_o[9]));
 BUFx3_ASAP7_75t_R output218 (.A(net239),
    .Y(data_we_o));
 BUFx3_ASAP7_75t_R output219 (.A(net240),
    .Y(instr_addr_o[10]));
 BUFx3_ASAP7_75t_R output220 (.A(net241),
    .Y(instr_addr_o[11]));
 BUFx3_ASAP7_75t_R output221 (.A(net242),
    .Y(instr_addr_o[12]));
 BUFx3_ASAP7_75t_R output222 (.A(net243),
    .Y(instr_addr_o[13]));
 BUFx3_ASAP7_75t_R output223 (.A(net244),
    .Y(instr_addr_o[14]));
 BUFx3_ASAP7_75t_R output224 (.A(net245),
    .Y(instr_addr_o[15]));
 BUFx3_ASAP7_75t_R output225 (.A(net246),
    .Y(instr_addr_o[16]));
 BUFx3_ASAP7_75t_R output226 (.A(net247),
    .Y(instr_addr_o[17]));
 BUFx3_ASAP7_75t_R output227 (.A(net248),
    .Y(instr_addr_o[18]));
 BUFx3_ASAP7_75t_R output228 (.A(net249),
    .Y(instr_addr_o[19]));
 BUFx3_ASAP7_75t_R output229 (.A(net250),
    .Y(instr_addr_o[20]));
 BUFx3_ASAP7_75t_R output230 (.A(net251),
    .Y(instr_addr_o[21]));
 BUFx3_ASAP7_75t_R output231 (.A(net252),
    .Y(instr_addr_o[22]));
 BUFx3_ASAP7_75t_R output232 (.A(net253),
    .Y(instr_addr_o[23]));
 BUFx3_ASAP7_75t_R output233 (.A(net254),
    .Y(instr_addr_o[24]));
 BUFx3_ASAP7_75t_R output234 (.A(net255),
    .Y(instr_addr_o[25]));
 BUFx3_ASAP7_75t_R output235 (.A(net256),
    .Y(instr_addr_o[26]));
 BUFx3_ASAP7_75t_R output236 (.A(net257),
    .Y(instr_addr_o[27]));
 BUFx3_ASAP7_75t_R output237 (.A(net258),
    .Y(instr_addr_o[28]));
 BUFx3_ASAP7_75t_R output238 (.A(net259),
    .Y(instr_addr_o[29]));
 BUFx3_ASAP7_75t_R output239 (.A(net260),
    .Y(instr_addr_o[2]));
 BUFx3_ASAP7_75t_R output240 (.A(net261),
    .Y(instr_addr_o[30]));
 BUFx3_ASAP7_75t_R output241 (.A(net262),
    .Y(instr_addr_o[31]));
 BUFx3_ASAP7_75t_R output242 (.A(net263),
    .Y(instr_addr_o[3]));
 BUFx3_ASAP7_75t_R output243 (.A(net264),
    .Y(instr_addr_o[4]));
 BUFx3_ASAP7_75t_R output244 (.A(net265),
    .Y(instr_addr_o[5]));
 BUFx3_ASAP7_75t_R output245 (.A(net266),
    .Y(instr_addr_o[6]));
 BUFx3_ASAP7_75t_R output246 (.A(net267),
    .Y(instr_addr_o[7]));
 BUFx3_ASAP7_75t_R output247 (.A(net268),
    .Y(instr_addr_o[8]));
 BUFx3_ASAP7_75t_R output248 (.A(net269),
    .Y(instr_addr_o[9]));
 BUFx3_ASAP7_75t_R output249 (.A(net270),
    .Y(instr_req_o));
 TIELOx1_ASAP7_75t_R _35101__250 (.L(net271));
 TIELOx1_ASAP7_75t_R _35102__251 (.L(net272));
 TIELOx1_ASAP7_75t_R _35103__252 (.L(net273));
 TIELOx1_ASAP7_75t_R _35104__253 (.L(net274));
 TIELOx1_ASAP7_75t_R _35135__254 (.L(net275));
 TIELOx1_ASAP7_75t_R _35136__255 (.L(net276));
 TIEHIx1_ASAP7_75t_R _35093__257 (.H(net278));
 TIEHIx1_ASAP7_75t_R _35094__258 (.H(net279));
 TIEHIx1_ASAP7_75t_R _35095__259 (.H(net280));
 TIEHIx1_ASAP7_75t_R _35096__260 (.H(net281));
 TIEHIx1_ASAP7_75t_R _35097__261 (.H(net282));
 TIEHIx1_ASAP7_75t_R _35098__262 (.H(net283));
 TIEHIx1_ASAP7_75t_R \core_busy_q$_DFF_PN0__263  (.H(net284));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcountinhibit_q[0]$_DFFE_PN0P__264  (.H(net285));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcountinhibit_q[2]$_DFFE_PN0P__265  (.H(net286));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[0]$_DFFE_PN0P__266  (.H(net287));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[10]$_DFFE_PN0P__267  (.H(net288));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[11]$_DFFE_PN0P__268  (.H(net289));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[12]$_DFFE_PN0P__269  (.H(net290));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[13]$_DFFE_PN0P__270  (.H(net291));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[14]$_DFFE_PN0P__271  (.H(net292));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[15]$_DFFE_PN0P__272  (.H(net293));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[16]$_DFFE_PN0P__273  (.H(net294));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[17]$_DFFE_PN0P__274  (.H(net295));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[18]$_DFFE_PN0P__275  (.H(net296));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[19]$_DFFE_PN0P__276  (.H(net297));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[1]$_DFFE_PN0P__277  (.H(net298));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[20]$_DFFE_PN0P__278  (.H(net299));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[21]$_DFFE_PN0P__279  (.H(net300));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[22]$_DFFE_PN0P__280  (.H(net301));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[23]$_DFFE_PN0P__281  (.H(net302));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[24]$_DFFE_PN0P__282  (.H(net303));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[25]$_DFFE_PN0P__283  (.H(net304));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[26]$_DFFE_PN0P__284  (.H(net305));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[27]$_DFFE_PN0P__285  (.H(net306));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[28]$_DFFE_PN0P__286  (.H(net307));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[29]$_DFFE_PN0P__287  (.H(net308));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[2]$_DFFE_PN0P__288  (.H(net309));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[30]$_DFFE_PN0P__289  (.H(net310));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[31]$_DFFE_PN0P__290  (.H(net311));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[32]$_DFFE_PN0P__291  (.H(net312));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[33]$_DFFE_PN0P__292  (.H(net313));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[34]$_DFFE_PN0P__293  (.H(net314));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[35]$_DFFE_PN0P__294  (.H(net315));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[36]$_DFFE_PN0P__295  (.H(net316));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[37]$_DFFE_PN0P__296  (.H(net317));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[38]$_DFFE_PN0P__297  (.H(net318));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[39]$_DFFE_PN0P__298  (.H(net319));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[3]$_DFFE_PN0P__299  (.H(net320));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[40]$_DFFE_PN0P__300  (.H(net321));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[41]$_DFFE_PN0P__301  (.H(net322));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[42]$_DFFE_PN0P__302  (.H(net323));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[43]$_DFFE_PN0P__303  (.H(net324));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[44]$_DFFE_PN0P__304  (.H(net325));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[45]$_DFFE_PN0P__305  (.H(net326));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[46]$_DFFE_PN0P__306  (.H(net327));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[47]$_DFFE_PN0P__307  (.H(net328));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[48]$_DFFE_PN0P__308  (.H(net329));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[49]$_DFFE_PN0P__309  (.H(net330));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[4]$_DFFE_PN0P__310  (.H(net331));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[50]$_DFFE_PN0P__311  (.H(net332));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[51]$_DFFE_PN0P__312  (.H(net333));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[52]$_DFFE_PN0P__313  (.H(net334));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[53]$_DFFE_PN0P__314  (.H(net335));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[54]$_DFFE_PN0P__315  (.H(net336));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[55]$_DFFE_PN0P__316  (.H(net337));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[56]$_DFFE_PN0P__317  (.H(net338));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[57]$_DFFE_PN0P__318  (.H(net339));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[58]$_DFFE_PN0P__319  (.H(net340));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[59]$_DFFE_PN0P__320  (.H(net341));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[5]$_DFFE_PN0P__321  (.H(net342));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[60]$_DFFE_PN0P__322  (.H(net343));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[61]$_DFFE_PN0P__323  (.H(net344));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[62]$_DFFE_PN0P__324  (.H(net345));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[63]$_DFFE_PN0P__325  (.H(net346));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[6]$_DFFE_PN0P__326  (.H(net347));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[7]$_DFFE_PN0P__327  (.H(net348));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[8]$_DFFE_PN0P__328  (.H(net349));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_val_o[9]$_DFFE_PN0P__329  (.H(net350));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[0]$_DFFE_PN0P__330  (.H(net351));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[10]$_DFFE_PN0P__331  (.H(net352));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[11]$_DFFE_PN0P__332  (.H(net353));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[12]$_DFFE_PN0P__333  (.H(net354));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[13]$_DFFE_PN0P__334  (.H(net355));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[14]$_DFFE_PN0P__335  (.H(net356));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[15]$_DFFE_PN0P__336  (.H(net357));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[16]$_DFFE_PN0P__337  (.H(net358));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[17]$_DFFE_PN0P__338  (.H(net359));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[18]$_DFFE_PN0P__339  (.H(net360));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[19]$_DFFE_PN0P__340  (.H(net361));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[1]$_DFFE_PN0P__341  (.H(net362));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[20]$_DFFE_PN0P__342  (.H(net363));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[21]$_DFFE_PN0P__343  (.H(net364));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[22]$_DFFE_PN0P__344  (.H(net365));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[23]$_DFFE_PN0P__345  (.H(net366));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[24]$_DFFE_PN0P__346  (.H(net367));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[25]$_DFFE_PN0P__347  (.H(net368));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[26]$_DFFE_PN0P__348  (.H(net369));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[27]$_DFFE_PN0P__349  (.H(net370));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[28]$_DFFE_PN0P__350  (.H(net371));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[29]$_DFFE_PN0P__351  (.H(net372));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[2]$_DFFE_PN0P__352  (.H(net373));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[30]$_DFFE_PN0P__353  (.H(net374));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[31]$_DFFE_PN0P__354  (.H(net375));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[32]$_DFFE_PN0P__355  (.H(net376));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[33]$_DFFE_PN0P__356  (.H(net377));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[34]$_DFFE_PN0P__357  (.H(net378));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[35]$_DFFE_PN0P__358  (.H(net379));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[36]$_DFFE_PN0P__359  (.H(net380));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[37]$_DFFE_PN0P__360  (.H(net381));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[38]$_DFFE_PN0P__361  (.H(net382));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[39]$_DFFE_PN0P__362  (.H(net383));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[3]$_DFFE_PN0P__363  (.H(net384));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[40]$_DFFE_PN0P__364  (.H(net385));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[41]$_DFFE_PN0P__365  (.H(net386));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[42]$_DFFE_PN0P__366  (.H(net387));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[43]$_DFFE_PN0P__367  (.H(net388));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[44]$_DFFE_PN0P__368  (.H(net389));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[45]$_DFFE_PN0P__369  (.H(net390));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[46]$_DFFE_PN0P__370  (.H(net391));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[47]$_DFFE_PN0P__371  (.H(net392));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[48]$_DFFE_PN0P__372  (.H(net393));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[49]$_DFFE_PN0P__373  (.H(net394));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[4]$_DFFE_PN0P__374  (.H(net395));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[50]$_DFFE_PN0P__375  (.H(net396));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[51]$_DFFE_PN0P__376  (.H(net397));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[52]$_DFFE_PN0P__377  (.H(net398));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[53]$_DFFE_PN0P__378  (.H(net399));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[54]$_DFFE_PN0P__379  (.H(net400));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[55]$_DFFE_PN0P__380  (.H(net401));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[56]$_DFFE_PN0P__381  (.H(net402));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[57]$_DFFE_PN0P__382  (.H(net403));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[58]$_DFFE_PN0P__383  (.H(net404));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[59]$_DFFE_PN0P__384  (.H(net405));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[5]$_DFFE_PN0P__385  (.H(net406));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[60]$_DFFE_PN0P__386  (.H(net407));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[61]$_DFFE_PN0P__387  (.H(net408));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[62]$_DFFE_PN0P__388  (.H(net409));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[63]$_DFFE_PN0P__389  (.H(net410));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[6]$_DFFE_PN0P__390  (.H(net411));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[7]$_DFFE_PN0P__391  (.H(net412));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[8]$_DFFE_PN0P__392  (.H(net413));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_val_o[9]$_DFFE_PN0P__393  (.H(net414));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.priv_mode_id_o[0]$_DFFE_PN1P__394  (.H(net415));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.priv_mode_id_o[1]$_DFFE_PN1P__395  (.H(net416));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[0]$_DFFE_PN1P__396  (.H(net417));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[11]$_DFFE_PN0P__397  (.H(net418));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[12]$_DFFE_PN0P__398  (.H(net419));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[13]$_DFFE_PN0P__399  (.H(net420));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[15]$_DFFE_PN0P__400  (.H(net421));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[1]$_DFFE_PN1P__401  (.H(net422));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[2]$_DFFE_PN0P__402  (.H(net423));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[6]$_DFFE_PN0P__403  (.H(net424));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[7]$_DFFE_PN0P__404  (.H(net425));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rd_data_o[8]$_DFFE_PN0P__405  (.H(net426));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[10]$_DFFE_PN0P__406  (.H(net427));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[11]$_DFFE_PN0P__407  (.H(net428));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[12]$_DFFE_PN0P__408  (.H(net429));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[13]$_DFFE_PN0P__409  (.H(net430));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[14]$_DFFE_PN0P__410  (.H(net431));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[15]$_DFFE_PN0P__411  (.H(net432));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[16]$_DFFE_PN0P__412  (.H(net433));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[17]$_DFFE_PN0P__413  (.H(net434));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[18]$_DFFE_PN0P__414  (.H(net435));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[19]$_DFFE_PN0P__415  (.H(net436));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[1]$_DFFE_PN0P__416  (.H(net437));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[20]$_DFFE_PN0P__417  (.H(net438));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[21]$_DFFE_PN0P__418  (.H(net439));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[22]$_DFFE_PN0P__419  (.H(net440));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[23]$_DFFE_PN0P__420  (.H(net441));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[24]$_DFFE_PN0P__421  (.H(net442));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[25]$_DFFE_PN0P__422  (.H(net443));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[26]$_DFFE_PN0P__423  (.H(net444));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[27]$_DFFE_PN0P__424  (.H(net445));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[28]$_DFFE_PN0P__425  (.H(net446));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[29]$_DFFE_PN0P__426  (.H(net447));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[2]$_DFFE_PN0P__427  (.H(net448));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[30]$_DFFE_PN0P__428  (.H(net449));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[31]$_DFFE_PN0P__429  (.H(net450));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[3]$_DFFE_PN0P__430  (.H(net451));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[4]$_DFFE_PN0P__431  (.H(net452));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[5]$_DFFE_PN0P__432  (.H(net453));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[6]$_DFFE_PN0P__433  (.H(net454));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[7]$_DFFE_PN0P__434  (.H(net455));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[8]$_DFFE_PN0P__435  (.H(net456));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rd_data_o[9]$_DFFE_PN0P__436  (.H(net457));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[0]$_DFFE_PN0P__437  (.H(net458));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[10]$_DFFE_PN0P__438  (.H(net459));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[11]$_DFFE_PN0P__439  (.H(net460));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[12]$_DFFE_PN0P__440  (.H(net461));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[13]$_DFFE_PN0P__441  (.H(net462));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[14]$_DFFE_PN0P__442  (.H(net463));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[15]$_DFFE_PN0P__443  (.H(net464));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[16]$_DFFE_PN0P__444  (.H(net465));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[17]$_DFFE_PN0P__445  (.H(net466));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[18]$_DFFE_PN0P__446  (.H(net467));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[19]$_DFFE_PN0P__447  (.H(net468));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[1]$_DFFE_PN0P__448  (.H(net469));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[20]$_DFFE_PN0P__449  (.H(net470));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[21]$_DFFE_PN0P__450  (.H(net471));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[22]$_DFFE_PN0P__451  (.H(net472));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[23]$_DFFE_PN0P__452  (.H(net473));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[24]$_DFFE_PN0P__453  (.H(net474));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[25]$_DFFE_PN0P__454  (.H(net475));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[26]$_DFFE_PN0P__455  (.H(net476));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[27]$_DFFE_PN0P__456  (.H(net477));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[28]$_DFFE_PN0P__457  (.H(net478));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[29]$_DFFE_PN0P__458  (.H(net479));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[2]$_DFFE_PN0P__459  (.H(net480));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[30]$_DFFE_PN0P__460  (.H(net481));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[31]$_DFFE_PN0P__461  (.H(net482));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[3]$_DFFE_PN0P__462  (.H(net483));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[4]$_DFFE_PN0P__463  (.H(net484));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[5]$_DFFE_PN0P__464  (.H(net485));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[6]$_DFFE_PN0P__465  (.H(net486));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[7]$_DFFE_PN0P__466  (.H(net487));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[8]$_DFFE_PN0P__467  (.H(net488));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rd_data_o[9]$_DFFE_PN0P__468  (.H(net489));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[0]$_DFFE_PN0P__469  (.H(net490));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[10]$_DFFE_PN0P__470  (.H(net491));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[11]$_DFFE_PN0P__471  (.H(net492));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[12]$_DFFE_PN0P__472  (.H(net493));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[13]$_DFFE_PN0P__473  (.H(net494));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[14]$_DFFE_PN0P__474  (.H(net495));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[15]$_DFFE_PN0P__475  (.H(net496));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[16]$_DFFE_PN0P__476  (.H(net497));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[17]$_DFFE_PN0P__477  (.H(net498));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[18]$_DFFE_PN0P__478  (.H(net499));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[19]$_DFFE_PN0P__479  (.H(net500));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[1]$_DFFE_PN0P__480  (.H(net501));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[20]$_DFFE_PN0P__481  (.H(net502));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[21]$_DFFE_PN0P__482  (.H(net503));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[22]$_DFFE_PN0P__483  (.H(net504));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[23]$_DFFE_PN0P__484  (.H(net505));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[24]$_DFFE_PN0P__485  (.H(net506));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[25]$_DFFE_PN0P__486  (.H(net507));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[26]$_DFFE_PN0P__487  (.H(net508));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[27]$_DFFE_PN0P__488  (.H(net509));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[28]$_DFFE_PN0P__489  (.H(net510));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[29]$_DFFE_PN0P__490  (.H(net511));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[2]$_DFFE_PN0P__491  (.H(net512));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[30]$_DFFE_PN0P__492  (.H(net513));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[31]$_DFFE_PN0P__493  (.H(net514));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[3]$_DFFE_PN0P__494  (.H(net515));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[4]$_DFFE_PN0P__495  (.H(net516));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[5]$_DFFE_PN0P__496  (.H(net517));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[6]$_DFFE_PN0P__497  (.H(net518));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[7]$_DFFE_PN0P__498  (.H(net519));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[8]$_DFFE_PN0P__499  (.H(net520));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rd_data_o[9]$_DFFE_PN0P__500  (.H(net521));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[0]$_DFFE_PN0P__501  (.H(net522));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[1]$_DFFE_PN0P__502  (.H(net523));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[2]$_DFFE_PN0P__503  (.H(net524));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[3]$_DFFE_PN0P__504  (.H(net525));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[4]$_DFFE_PN0P__505  (.H(net526));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rd_data_o[5]$_DFFE_PN0P__506  (.H(net527));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[0]$_DFFE_PN0P__507  (.H(net528));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[10]$_DFFE_PN0P__508  (.H(net529));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[11]$_DFFE_PN0P__509  (.H(net530));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[12]$_DFFE_PN0P__510  (.H(net531));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[13]$_DFFE_PN0P__511  (.H(net532));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[14]$_DFFE_PN0P__512  (.H(net533));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[15]$_DFFE_PN0P__513  (.H(net534));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[16]$_DFFE_PN0P__514  (.H(net535));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[17]$_DFFE_PN0P__515  (.H(net536));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[18]$_DFFE_PN0P__516  (.H(net537));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[19]$_DFFE_PN0P__517  (.H(net538));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[1]$_DFFE_PN0P__518  (.H(net539));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[20]$_DFFE_PN0P__519  (.H(net540));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[21]$_DFFE_PN0P__520  (.H(net541));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[22]$_DFFE_PN0P__521  (.H(net542));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[23]$_DFFE_PN0P__522  (.H(net543));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[24]$_DFFE_PN0P__523  (.H(net544));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[25]$_DFFE_PN0P__524  (.H(net545));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[26]$_DFFE_PN0P__525  (.H(net546));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[27]$_DFFE_PN0P__526  (.H(net547));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[28]$_DFFE_PN0P__527  (.H(net548));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[29]$_DFFE_PN0P__528  (.H(net549));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[2]$_DFFE_PN0P__529  (.H(net550));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[30]$_DFFE_PN0P__530  (.H(net551));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[31]$_DFFE_PN0P__531  (.H(net552));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[3]$_DFFE_PN0P__532  (.H(net553));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[4]$_DFFE_PN0P__533  (.H(net554));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[5]$_DFFE_PN0P__534  (.H(net555));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[6]$_DFFE_PN0P__535  (.H(net556));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[7]$_DFFE_PN0P__536  (.H(net557));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[8]$_DFFE_PN0P__537  (.H(net558));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rd_data_o[9]$_DFFE_PN0P__538  (.H(net559));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[0]$_DFFE_PN0P__539  (.H(net560));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[10]$_DFFE_PN0P__540  (.H(net561));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[11]$_DFFE_PN0P__541  (.H(net562));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[12]$_DFFE_PN0P__542  (.H(net563));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[13]$_DFFE_PN0P__543  (.H(net564));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[14]$_DFFE_PN0P__544  (.H(net565));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[15]$_DFFE_PN0P__545  (.H(net566));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[16]$_DFFE_PN0P__546  (.H(net567));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[17]$_DFFE_PN0P__547  (.H(net568));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[1]$_DFFE_PN0P__548  (.H(net569));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[2]$_DFFE_PN0P__549  (.H(net570));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[3]$_DFFE_PN0P__550  (.H(net571));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[4]$_DFFE_PN0P__551  (.H(net572));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[5]$_DFFE_PN0P__552  (.H(net573));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[6]$_DFFE_PN0P__553  (.H(net574));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[7]$_DFFE_PN0P__554  (.H(net575));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[8]$_DFFE_PN0P__555  (.H(net576));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rd_data_o[9]$_DFFE_PN0P__556  (.H(net577));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[0]$_DFFE_PN0P__557  (.H(net578));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[10]$_DFFE_PN0P__558  (.H(net579));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[11]$_DFFE_PN0P__559  (.H(net580));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[12]$_DFFE_PN0P__560  (.H(net581));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[13]$_DFFE_PN0P__561  (.H(net582));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[14]$_DFFE_PN0P__562  (.H(net583));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[15]$_DFFE_PN0P__563  (.H(net584));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[16]$_DFFE_PN0P__564  (.H(net585));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[17]$_DFFE_PN0P__565  (.H(net586));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[18]$_DFFE_PN0P__566  (.H(net587));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[19]$_DFFE_PN0P__567  (.H(net588));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[1]$_DFFE_PN0P__568  (.H(net589));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[20]$_DFFE_PN0P__569  (.H(net590));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[21]$_DFFE_PN0P__570  (.H(net591));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[22]$_DFFE_PN0P__571  (.H(net592));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[23]$_DFFE_PN0P__572  (.H(net593));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[24]$_DFFE_PN0P__573  (.H(net594));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[25]$_DFFE_PN0P__574  (.H(net595));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[26]$_DFFE_PN0P__575  (.H(net596));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[27]$_DFFE_PN0P__576  (.H(net597));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[28]$_DFFE_PN0P__577  (.H(net598));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[29]$_DFFE_PN0P__578  (.H(net599));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[2]$_DFFE_PN0P__579  (.H(net600));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[30]$_DFFE_PN0P__580  (.H(net601));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[31]$_DFFE_PN0P__581  (.H(net602));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[3]$_DFFE_PN0P__582  (.H(net603));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[4]$_DFFE_PN0P__583  (.H(net604));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[5]$_DFFE_PN0P__584  (.H(net605));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[6]$_DFFE_PN0P__585  (.H(net606));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[7]$_DFFE_PN0P__586  (.H(net607));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[8]$_DFFE_PN0P__587  (.H(net608));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rd_data_o[9]$_DFFE_PN0P__588  (.H(net609));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[0]$_DFFE_PN0P__589  (.H(net610));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[1]$_DFFE_PN0P__590  (.H(net611));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[2]$_DFFE_PN0P__591  (.H(net612));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[3]$_DFFE_PN0P__592  (.H(net613));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[4]$_DFFE_PN0P__593  (.H(net614));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rd_data_o[5]$_DFFE_PN0P__594  (.H(net615));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rd_data_o[0]$_DFFE_PN0P__595  (.H(net616));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rd_data_o[1]$_DFFE_PN0P__596  (.H(net617));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rd_data_o[2]$_DFFE_PN1P__597  (.H(net618));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[0]$_DFFE_PN0P__598  (.H(net619));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[10]$_DFFE_PN0P__599  (.H(net620));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[11]$_DFFE_PN0P__600  (.H(net621));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[12]$_DFFE_PN0P__601  (.H(net622));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[13]$_DFFE_PN0P__602  (.H(net623));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[14]$_DFFE_PN0P__603  (.H(net624));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[15]$_DFFE_PN0P__604  (.H(net625));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[16]$_DFFE_PN0P__605  (.H(net626));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[17]$_DFFE_PN0P__606  (.H(net627));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[18]$_DFFE_PN0P__607  (.H(net628));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[19]$_DFFE_PN0P__608  (.H(net629));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[1]$_DFFE_PN0P__609  (.H(net630));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[20]$_DFFE_PN0P__610  (.H(net631));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[21]$_DFFE_PN0P__611  (.H(net632));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[22]$_DFFE_PN0P__612  (.H(net633));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[23]$_DFFE_PN0P__613  (.H(net634));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[24]$_DFFE_PN0P__614  (.H(net635));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[25]$_DFFE_PN0P__615  (.H(net636));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[26]$_DFFE_PN0P__616  (.H(net637));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[27]$_DFFE_PN0P__617  (.H(net638));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[28]$_DFFE_PN0P__618  (.H(net639));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[29]$_DFFE_PN0P__619  (.H(net640));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[2]$_DFFE_PN0P__620  (.H(net641));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[30]$_DFFE_PN0P__621  (.H(net642));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[31]$_DFFE_PN0P__622  (.H(net643));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[3]$_DFFE_PN0P__623  (.H(net644));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[4]$_DFFE_PN0P__624  (.H(net645));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[5]$_DFFE_PN0P__625  (.H(net646));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[6]$_DFFE_PN0P__626  (.H(net647));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[7]$_DFFE_PN0P__627  (.H(net648));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[8]$_DFFE_PN0P__628  (.H(net649));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rd_data_o[9]$_DFFE_PN0P__629  (.H(net650));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[0]$_DFFE_PN0P__630  (.H(net651));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[1]$_DFFE_PN0P__631  (.H(net652));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[2]$_DFFE_PN0N__632  (.H(net653));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[3]$_DFFE_PN0N__633  (.H(net654));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[4]$_DFFE_PN1N__634  (.H(net655));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rd_data_o[5]$_DFFE_PN0N__635  (.H(net656));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[0]$_DFFE_PN0P__636  (.H(net657));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[10]$_DFFE_PN0P__637  (.H(net658));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[11]$_DFFE_PN0P__638  (.H(net659));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[12]$_DFFE_PN0P__639  (.H(net660));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[13]$_DFFE_PN0P__640  (.H(net661));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[14]$_DFFE_PN0P__641  (.H(net662));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[15]$_DFFE_PN0P__642  (.H(net663));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[16]$_DFFE_PN0P__643  (.H(net664));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[17]$_DFFE_PN0P__644  (.H(net665));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[18]$_DFFE_PN0P__645  (.H(net666));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[19]$_DFFE_PN0P__646  (.H(net667));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[1]$_DFFE_PN0P__647  (.H(net668));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[20]$_DFFE_PN0P__648  (.H(net669));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[21]$_DFFE_PN0P__649  (.H(net670));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[22]$_DFFE_PN0P__650  (.H(net671));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[23]$_DFFE_PN0P__651  (.H(net672));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[24]$_DFFE_PN0P__652  (.H(net673));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[25]$_DFFE_PN0P__653  (.H(net674));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[26]$_DFFE_PN0P__654  (.H(net675));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[27]$_DFFE_PN0P__655  (.H(net676));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[28]$_DFFE_PN0P__656  (.H(net677));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[29]$_DFFE_PN0P__657  (.H(net678));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[2]$_DFFE_PN0P__658  (.H(net679));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[30]$_DFFE_PN0P__659  (.H(net680));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[31]$_DFFE_PN0P__660  (.H(net681));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[3]$_DFFE_PN0P__661  (.H(net682));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[4]$_DFFE_PN0P__662  (.H(net683));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[5]$_DFFE_PN0P__663  (.H(net684));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[6]$_DFFE_PN0P__664  (.H(net685));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[7]$_DFFE_PN0P__665  (.H(net686));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[8]$_DFFE_PN0P__666  (.H(net687));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rd_data_o[9]$_DFFE_PN0P__667  (.H(net688));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[10]$_DFFE_PN0P__668  (.H(net689));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[11]$_DFFE_PN0P__669  (.H(net690));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[12]$_DFFE_PN0P__670  (.H(net691));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[13]$_DFFE_PN0P__671  (.H(net692));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[14]$_DFFE_PN0P__672  (.H(net693));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[15]$_DFFE_PN0P__673  (.H(net694));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[16]$_DFFE_PN0P__674  (.H(net695));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[17]$_DFFE_PN0P__675  (.H(net696));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[18]$_DFFE_PN0P__676  (.H(net697));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[19]$_DFFE_PN0P__677  (.H(net698));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[20]$_DFFE_PN0P__678  (.H(net699));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[21]$_DFFE_PN0P__679  (.H(net700));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[22]$_DFFE_PN0P__680  (.H(net701));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[23]$_DFFE_PN0P__681  (.H(net702));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[24]$_DFFE_PN0P__682  (.H(net703));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[25]$_DFFE_PN0P__683  (.H(net704));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[26]$_DFFE_PN0P__684  (.H(net705));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[27]$_DFFE_PN0P__685  (.H(net706));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[28]$_DFFE_PN0P__686  (.H(net707));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[29]$_DFFE_PN0P__687  (.H(net708));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[30]$_DFFE_PN0P__688  (.H(net709));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[31]$_DFFE_PN0P__689  (.H(net710));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[8]$_DFFE_PN0P__690  (.H(net711));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rd_data_o[9]$_DFFE_PN0P__691  (.H(net712));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P__692  (.H(net713));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P__693  (.H(net714));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P__694  (.H(net715));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P__695  (.H(net716));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P__696  (.H(net717));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P__697  (.H(net718));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1__698  (.H(net719));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0__699  (.H(net720));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0__700  (.H(net721));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0__701  (.H(net722));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0__702  (.H(net723));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0__703  (.H(net724));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P__704  (.H(net725));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P__705  (.H(net726));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P__706  (.H(net727));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P__707  (.H(net728));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P__708  (.H(net729));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P__709  (.H(net730));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P__710  (.H(net731));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P__711  (.H(net732));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P__712  (.H(net733));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P__713  (.H(net734));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P__714  (.H(net735));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P__715  (.H(net736));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P__716  (.H(net737));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P__717  (.H(net738));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P__718  (.H(net739));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P__719  (.H(net740));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P__720  (.H(net741));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P__721  (.H(net742));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P__722  (.H(net743));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P__723  (.H(net744));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P__724  (.H(net745));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P__725  (.H(net746));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P__726  (.H(net747));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P__727  (.H(net748));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P__728  (.H(net749));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P__729  (.H(net750));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P__730  (.H(net751));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P__731  (.H(net752));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P__732  (.H(net753));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P__733  (.H(net754));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P__734  (.H(net755));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P__735  (.H(net756));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P__736  (.H(net757));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P__737  (.H(net758));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P__738  (.H(net759));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P__739  (.H(net760));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P__740  (.H(net761));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P__741  (.H(net762));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P__742  (.H(net763));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P__743  (.H(net764));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P__744  (.H(net765));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P__745  (.H(net766));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P__746  (.H(net767));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P__747  (.H(net768));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P__748  (.H(net769));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P__749  (.H(net770));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P__750  (.H(net771));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P__751  (.H(net772));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P__752  (.H(net773));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P__753  (.H(net774));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P__754  (.H(net775));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P__755  (.H(net776));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P__756  (.H(net777));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P__757  (.H(net778));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P__758  (.H(net779));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P__759  (.H(net780));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P__760  (.H(net781));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P__761  (.H(net782));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P__762  (.H(net783));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P__763  (.H(net784));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P__764  (.H(net785));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P__765  (.H(net786));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P__766  (.H(net787));
 TIEHIx1_ASAP7_75t_R \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P__767  (.H(net788));
 TIEHIx1_ASAP7_75t_R \fetch_enable_q$_DFFE_PN0P__768  (.H(net789));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1000]$_DFFE_PN0P__769  (.H(net790));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1001]$_DFFE_PN0P__770  (.H(net791));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1002]$_DFFE_PN0P__771  (.H(net792));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1003]$_DFFE_PN0P__772  (.H(net793));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1004]$_DFFE_PN0P__773  (.H(net794));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1005]$_DFFE_PN0P__774  (.H(net795));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1006]$_DFFE_PN0P__775  (.H(net796));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1007]$_DFFE_PN0P__776  (.H(net797));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1008]$_DFFE_PN0P__777  (.H(net798));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1009]$_DFFE_PN0P__778  (.H(net799));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[100]$_DFFE_PN0P__779  (.H(net800));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1010]$_DFFE_PN0P__780  (.H(net801));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1011]$_DFFE_PN0P__781  (.H(net802));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1012]$_DFFE_PN0P__782  (.H(net803));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1013]$_DFFE_PN0P__783  (.H(net804));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1014]$_DFFE_PN0P__784  (.H(net805));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1015]$_DFFE_PN0P__785  (.H(net806));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1016]$_DFFE_PN0P__786  (.H(net807));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1017]$_DFFE_PN0P__787  (.H(net808));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1018]$_DFFE_PN0P__788  (.H(net809));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1019]$_DFFE_PN0P__789  (.H(net810));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[101]$_DFFE_PN0P__790  (.H(net811));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1020]$_DFFE_PN0P__791  (.H(net812));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1021]$_DFFE_PN0P__792  (.H(net813));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1022]$_DFFE_PN0P__793  (.H(net814));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[1023]$_DFFE_PN0P__794  (.H(net815));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[102]$_DFFE_PN0P__795  (.H(net816));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[103]$_DFFE_PN0P__796  (.H(net817));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[104]$_DFFE_PN0P__797  (.H(net818));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[105]$_DFFE_PN0P__798  (.H(net819));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[106]$_DFFE_PN0P__799  (.H(net820));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[107]$_DFFE_PN0P__800  (.H(net821));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[108]$_DFFE_PN0P__801  (.H(net822));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[109]$_DFFE_PN0P__802  (.H(net823));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[110]$_DFFE_PN0P__803  (.H(net824));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[111]$_DFFE_PN0P__804  (.H(net825));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[112]$_DFFE_PN0P__805  (.H(net826));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[113]$_DFFE_PN0P__806  (.H(net827));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[114]$_DFFE_PN0P__807  (.H(net828));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[115]$_DFFE_PN0P__808  (.H(net829));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[116]$_DFFE_PN0P__809  (.H(net830));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[117]$_DFFE_PN0P__810  (.H(net831));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[118]$_DFFE_PN0P__811  (.H(net832));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[119]$_DFFE_PN0P__812  (.H(net833));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[120]$_DFFE_PN0P__813  (.H(net834));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[121]$_DFFE_PN0P__814  (.H(net835));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[122]$_DFFE_PN0P__815  (.H(net836));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[123]$_DFFE_PN0P__816  (.H(net837));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[124]$_DFFE_PN0P__817  (.H(net838));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[125]$_DFFE_PN0P__818  (.H(net839));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[126]$_DFFE_PN0P__819  (.H(net840));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[127]$_DFFE_PN0P__820  (.H(net841));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[128]$_DFFE_PN0P__821  (.H(net842));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[129]$_DFFE_PN0P__822  (.H(net843));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[130]$_DFFE_PN0P__823  (.H(net844));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[131]$_DFFE_PN0P__824  (.H(net845));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[132]$_DFFE_PN0P__825  (.H(net846));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[133]$_DFFE_PN0P__826  (.H(net847));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[134]$_DFFE_PN0P__827  (.H(net848));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[135]$_DFFE_PN0P__828  (.H(net849));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[136]$_DFFE_PN0P__829  (.H(net850));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[137]$_DFFE_PN0P__830  (.H(net851));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[138]$_DFFE_PN0P__831  (.H(net852));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[139]$_DFFE_PN0P__832  (.H(net853));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[140]$_DFFE_PN0P__833  (.H(net854));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[141]$_DFFE_PN0P__834  (.H(net855));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[142]$_DFFE_PN0P__835  (.H(net856));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[143]$_DFFE_PN0P__836  (.H(net857));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[144]$_DFFE_PN0P__837  (.H(net858));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[145]$_DFFE_PN0P__838  (.H(net859));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[146]$_DFFE_PN0P__839  (.H(net860));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[147]$_DFFE_PN0P__840  (.H(net861));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[148]$_DFFE_PN0P__841  (.H(net862));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[149]$_DFFE_PN0P__842  (.H(net863));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[150]$_DFFE_PN0P__843  (.H(net864));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[151]$_DFFE_PN0P__844  (.H(net865));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[152]$_DFFE_PN0P__845  (.H(net866));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[153]$_DFFE_PN0P__846  (.H(net867));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[154]$_DFFE_PN0P__847  (.H(net868));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[155]$_DFFE_PN0P__848  (.H(net869));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[156]$_DFFE_PN0P__849  (.H(net870));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[157]$_DFFE_PN0P__850  (.H(net871));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[158]$_DFFE_PN0P__851  (.H(net872));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[159]$_DFFE_PN0P__852  (.H(net873));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[160]$_DFFE_PN0P__853  (.H(net874));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[161]$_DFFE_PN0P__854  (.H(net875));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[162]$_DFFE_PN0P__855  (.H(net876));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[163]$_DFFE_PN0P__856  (.H(net877));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[164]$_DFFE_PN0P__857  (.H(net878));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[165]$_DFFE_PN0P__858  (.H(net879));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[166]$_DFFE_PN0P__859  (.H(net880));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[167]$_DFFE_PN0P__860  (.H(net881));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[168]$_DFFE_PN0P__861  (.H(net882));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[169]$_DFFE_PN0P__862  (.H(net883));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[170]$_DFFE_PN0P__863  (.H(net884));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[171]$_DFFE_PN0P__864  (.H(net885));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[172]$_DFFE_PN0P__865  (.H(net886));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[173]$_DFFE_PN0P__866  (.H(net887));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[174]$_DFFE_PN0P__867  (.H(net888));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[175]$_DFFE_PN0P__868  (.H(net889));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[176]$_DFFE_PN0P__869  (.H(net890));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[177]$_DFFE_PN0P__870  (.H(net891));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[178]$_DFFE_PN0P__871  (.H(net892));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[179]$_DFFE_PN0P__872  (.H(net893));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[180]$_DFFE_PN0P__873  (.H(net894));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[181]$_DFFE_PN0P__874  (.H(net895));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[182]$_DFFE_PN0P__875  (.H(net896));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[183]$_DFFE_PN0P__876  (.H(net897));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[184]$_DFFE_PN0P__877  (.H(net898));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[185]$_DFFE_PN0P__878  (.H(net899));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[186]$_DFFE_PN0P__879  (.H(net900));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[187]$_DFFE_PN0P__880  (.H(net901));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[188]$_DFFE_PN0P__881  (.H(net902));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[189]$_DFFE_PN0P__882  (.H(net903));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[190]$_DFFE_PN0P__883  (.H(net904));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[191]$_DFFE_PN0P__884  (.H(net905));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[192]$_DFFE_PN0P__885  (.H(net906));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[193]$_DFFE_PN0P__886  (.H(net907));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[194]$_DFFE_PN0P__887  (.H(net908));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[195]$_DFFE_PN0P__888  (.H(net909));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[196]$_DFFE_PN0P__889  (.H(net910));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[197]$_DFFE_PN0P__890  (.H(net911));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[198]$_DFFE_PN0P__891  (.H(net912));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[199]$_DFFE_PN0P__892  (.H(net913));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[200]$_DFFE_PN0P__893  (.H(net914));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[201]$_DFFE_PN0P__894  (.H(net915));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[202]$_DFFE_PN0P__895  (.H(net916));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[203]$_DFFE_PN0P__896  (.H(net917));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[204]$_DFFE_PN0P__897  (.H(net918));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[205]$_DFFE_PN0P__898  (.H(net919));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[206]$_DFFE_PN0P__899  (.H(net920));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[207]$_DFFE_PN0P__900  (.H(net921));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[208]$_DFFE_PN0P__901  (.H(net922));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[209]$_DFFE_PN0P__902  (.H(net923));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[210]$_DFFE_PN0P__903  (.H(net924));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[211]$_DFFE_PN0P__904  (.H(net925));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[212]$_DFFE_PN0P__905  (.H(net926));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[213]$_DFFE_PN0P__906  (.H(net927));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[214]$_DFFE_PN0P__907  (.H(net928));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[215]$_DFFE_PN0P__908  (.H(net929));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[216]$_DFFE_PN0P__909  (.H(net930));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[217]$_DFFE_PN0P__910  (.H(net931));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[218]$_DFFE_PN0P__911  (.H(net932));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[219]$_DFFE_PN0P__912  (.H(net933));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[220]$_DFFE_PN0P__913  (.H(net934));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[221]$_DFFE_PN0P__914  (.H(net935));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[222]$_DFFE_PN0P__915  (.H(net936));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[223]$_DFFE_PN0P__916  (.H(net937));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[224]$_DFFE_PN0P__917  (.H(net938));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[225]$_DFFE_PN0P__918  (.H(net939));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[226]$_DFFE_PN0P__919  (.H(net940));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[227]$_DFFE_PN0P__920  (.H(net941));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[228]$_DFFE_PN0P__921  (.H(net942));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[229]$_DFFE_PN0P__922  (.H(net943));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[230]$_DFFE_PN0P__923  (.H(net944));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[231]$_DFFE_PN0P__924  (.H(net945));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[232]$_DFFE_PN0P__925  (.H(net946));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[233]$_DFFE_PN0P__926  (.H(net947));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[234]$_DFFE_PN0P__927  (.H(net948));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[235]$_DFFE_PN0P__928  (.H(net949));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[236]$_DFFE_PN0P__929  (.H(net950));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[237]$_DFFE_PN0P__930  (.H(net951));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[238]$_DFFE_PN0P__931  (.H(net952));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[239]$_DFFE_PN0P__932  (.H(net953));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[240]$_DFFE_PN0P__933  (.H(net954));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[241]$_DFFE_PN0P__934  (.H(net955));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[242]$_DFFE_PN0P__935  (.H(net956));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[243]$_DFFE_PN0P__936  (.H(net957));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[244]$_DFFE_PN0P__937  (.H(net958));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[245]$_DFFE_PN0P__938  (.H(net959));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[246]$_DFFE_PN0P__939  (.H(net960));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[247]$_DFFE_PN0P__940  (.H(net961));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[248]$_DFFE_PN0P__941  (.H(net962));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[249]$_DFFE_PN0P__942  (.H(net963));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[250]$_DFFE_PN0P__943  (.H(net964));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[251]$_DFFE_PN0P__944  (.H(net965));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[252]$_DFFE_PN0P__945  (.H(net966));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[253]$_DFFE_PN0P__946  (.H(net967));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[254]$_DFFE_PN0P__947  (.H(net968));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[255]$_DFFE_PN0P__948  (.H(net969));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[256]$_DFFE_PN0P__949  (.H(net970));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[257]$_DFFE_PN0P__950  (.H(net971));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[258]$_DFFE_PN0P__951  (.H(net972));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[259]$_DFFE_PN0P__952  (.H(net973));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[260]$_DFFE_PN0P__953  (.H(net974));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[261]$_DFFE_PN0P__954  (.H(net975));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[262]$_DFFE_PN0P__955  (.H(net976));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[263]$_DFFE_PN0P__956  (.H(net977));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[264]$_DFFE_PN0P__957  (.H(net978));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[265]$_DFFE_PN0P__958  (.H(net979));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[266]$_DFFE_PN0P__959  (.H(net980));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[267]$_DFFE_PN0P__960  (.H(net981));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[268]$_DFFE_PN0P__961  (.H(net982));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[269]$_DFFE_PN0P__962  (.H(net983));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[270]$_DFFE_PN0P__963  (.H(net984));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[271]$_DFFE_PN0P__964  (.H(net985));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[272]$_DFFE_PN0P__965  (.H(net986));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[273]$_DFFE_PN0P__966  (.H(net987));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[274]$_DFFE_PN0P__967  (.H(net988));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[275]$_DFFE_PN0P__968  (.H(net989));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[276]$_DFFE_PN0P__969  (.H(net990));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[277]$_DFFE_PN0P__970  (.H(net991));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[278]$_DFFE_PN0P__971  (.H(net992));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[279]$_DFFE_PN0P__972  (.H(net993));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[280]$_DFFE_PN0P__973  (.H(net994));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[281]$_DFFE_PN0P__974  (.H(net995));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[282]$_DFFE_PN0P__975  (.H(net996));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[283]$_DFFE_PN0P__976  (.H(net997));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[284]$_DFFE_PN0P__977  (.H(net998));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[285]$_DFFE_PN0P__978  (.H(net999));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[286]$_DFFE_PN0P__979  (.H(net1000));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[287]$_DFFE_PN0P__980  (.H(net1001));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[288]$_DFFE_PN0P__981  (.H(net1002));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[289]$_DFFE_PN0P__982  (.H(net1003));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[290]$_DFFE_PN0P__983  (.H(net1004));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[291]$_DFFE_PN0P__984  (.H(net1005));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[292]$_DFFE_PN0P__985  (.H(net1006));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[293]$_DFFE_PN0P__986  (.H(net1007));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[294]$_DFFE_PN0P__987  (.H(net1008));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[295]$_DFFE_PN0P__988  (.H(net1009));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[296]$_DFFE_PN0P__989  (.H(net1010));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[297]$_DFFE_PN0P__990  (.H(net1011));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[298]$_DFFE_PN0P__991  (.H(net1012));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[299]$_DFFE_PN0P__992  (.H(net1013));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[300]$_DFFE_PN0P__993  (.H(net1014));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[301]$_DFFE_PN0P__994  (.H(net1015));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[302]$_DFFE_PN0P__995  (.H(net1016));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[303]$_DFFE_PN0P__996  (.H(net1017));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[304]$_DFFE_PN0P__997  (.H(net1018));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[305]$_DFFE_PN0P__998  (.H(net1019));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[306]$_DFFE_PN0P__999  (.H(net1020));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[307]$_DFFE_PN0P__1000  (.H(net1021));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[308]$_DFFE_PN0P__1001  (.H(net1022));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[309]$_DFFE_PN0P__1002  (.H(net1023));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[310]$_DFFE_PN0P__1003  (.H(net1024));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[311]$_DFFE_PN0P__1004  (.H(net1025));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[312]$_DFFE_PN0P__1005  (.H(net1026));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[313]$_DFFE_PN0P__1006  (.H(net1027));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[314]$_DFFE_PN0P__1007  (.H(net1028));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[315]$_DFFE_PN0P__1008  (.H(net1029));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[316]$_DFFE_PN0P__1009  (.H(net1030));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[317]$_DFFE_PN0P__1010  (.H(net1031));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[318]$_DFFE_PN0P__1011  (.H(net1032));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[319]$_DFFE_PN0P__1012  (.H(net1033));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[320]$_DFFE_PN0P__1013  (.H(net1034));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[321]$_DFFE_PN0P__1014  (.H(net1035));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[322]$_DFFE_PN0P__1015  (.H(net1036));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[323]$_DFFE_PN0P__1016  (.H(net1037));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[324]$_DFFE_PN0P__1017  (.H(net1038));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[325]$_DFFE_PN0P__1018  (.H(net1039));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[326]$_DFFE_PN0P__1019  (.H(net1040));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[327]$_DFFE_PN0P__1020  (.H(net1041));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[328]$_DFFE_PN0P__1021  (.H(net1042));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[329]$_DFFE_PN0P__1022  (.H(net1043));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[32]$_DFFE_PN0P__1023  (.H(net1044));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[330]$_DFFE_PN0P__1024  (.H(net1045));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[331]$_DFFE_PN0P__1025  (.H(net1046));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[332]$_DFFE_PN0P__1026  (.H(net1047));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[333]$_DFFE_PN0P__1027  (.H(net1048));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[334]$_DFFE_PN0P__1028  (.H(net1049));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[335]$_DFFE_PN0P__1029  (.H(net1050));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[336]$_DFFE_PN0P__1030  (.H(net1051));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[337]$_DFFE_PN0P__1031  (.H(net1052));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[338]$_DFFE_PN0P__1032  (.H(net1053));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[339]$_DFFE_PN0P__1033  (.H(net1054));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[33]$_DFFE_PN0P__1034  (.H(net1055));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[340]$_DFFE_PN0P__1035  (.H(net1056));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[341]$_DFFE_PN0P__1036  (.H(net1057));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[342]$_DFFE_PN0P__1037  (.H(net1058));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[343]$_DFFE_PN0P__1038  (.H(net1059));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[344]$_DFFE_PN0P__1039  (.H(net1060));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[345]$_DFFE_PN0P__1040  (.H(net1061));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[346]$_DFFE_PN0P__1041  (.H(net1062));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[347]$_DFFE_PN0P__1042  (.H(net1063));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[348]$_DFFE_PN0P__1043  (.H(net1064));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[349]$_DFFE_PN0P__1044  (.H(net1065));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[34]$_DFFE_PN0P__1045  (.H(net1066));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[350]$_DFFE_PN0P__1046  (.H(net1067));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[351]$_DFFE_PN0P__1047  (.H(net1068));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[352]$_DFFE_PN0P__1048  (.H(net1069));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[353]$_DFFE_PN0P__1049  (.H(net1070));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[354]$_DFFE_PN0P__1050  (.H(net1071));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[355]$_DFFE_PN0P__1051  (.H(net1072));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[356]$_DFFE_PN0P__1052  (.H(net1073));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[357]$_DFFE_PN0P__1053  (.H(net1074));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[358]$_DFFE_PN0P__1054  (.H(net1075));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[359]$_DFFE_PN0P__1055  (.H(net1076));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[35]$_DFFE_PN0P__1056  (.H(net1077));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[360]$_DFFE_PN0P__1057  (.H(net1078));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[361]$_DFFE_PN0P__1058  (.H(net1079));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[362]$_DFFE_PN0P__1059  (.H(net1080));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[363]$_DFFE_PN0P__1060  (.H(net1081));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[364]$_DFFE_PN0P__1061  (.H(net1082));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[365]$_DFFE_PN0P__1062  (.H(net1083));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[366]$_DFFE_PN0P__1063  (.H(net1084));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[367]$_DFFE_PN0P__1064  (.H(net1085));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[368]$_DFFE_PN0P__1065  (.H(net1086));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[369]$_DFFE_PN0P__1066  (.H(net1087));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[36]$_DFFE_PN0P__1067  (.H(net1088));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[370]$_DFFE_PN0P__1068  (.H(net1089));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[371]$_DFFE_PN0P__1069  (.H(net1090));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[372]$_DFFE_PN0P__1070  (.H(net1091));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[373]$_DFFE_PN0P__1071  (.H(net1092));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[374]$_DFFE_PN0P__1072  (.H(net1093));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[375]$_DFFE_PN0P__1073  (.H(net1094));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[376]$_DFFE_PN0P__1074  (.H(net1095));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[377]$_DFFE_PN0P__1075  (.H(net1096));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[378]$_DFFE_PN0P__1076  (.H(net1097));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[379]$_DFFE_PN0P__1077  (.H(net1098));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[37]$_DFFE_PN0P__1078  (.H(net1099));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[380]$_DFFE_PN0P__1079  (.H(net1100));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[381]$_DFFE_PN0P__1080  (.H(net1101));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[382]$_DFFE_PN0P__1081  (.H(net1102));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[383]$_DFFE_PN0P__1082  (.H(net1103));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[384]$_DFFE_PN0P__1083  (.H(net1104));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[385]$_DFFE_PN0P__1084  (.H(net1105));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[386]$_DFFE_PN0P__1085  (.H(net1106));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[387]$_DFFE_PN0P__1086  (.H(net1107));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[388]$_DFFE_PN0P__1087  (.H(net1108));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[389]$_DFFE_PN0P__1088  (.H(net1109));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[38]$_DFFE_PN0P__1089  (.H(net1110));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[390]$_DFFE_PN0P__1090  (.H(net1111));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[391]$_DFFE_PN0P__1091  (.H(net1112));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[392]$_DFFE_PN0P__1092  (.H(net1113));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[393]$_DFFE_PN0P__1093  (.H(net1114));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[394]$_DFFE_PN0P__1094  (.H(net1115));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[395]$_DFFE_PN0P__1095  (.H(net1116));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[396]$_DFFE_PN0P__1096  (.H(net1117));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[397]$_DFFE_PN0P__1097  (.H(net1118));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[398]$_DFFE_PN0P__1098  (.H(net1119));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[399]$_DFFE_PN0P__1099  (.H(net1120));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[39]$_DFFE_PN0P__1100  (.H(net1121));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[400]$_DFFE_PN0P__1101  (.H(net1122));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[401]$_DFFE_PN0P__1102  (.H(net1123));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[402]$_DFFE_PN0P__1103  (.H(net1124));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[403]$_DFFE_PN0P__1104  (.H(net1125));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[404]$_DFFE_PN0P__1105  (.H(net1126));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[405]$_DFFE_PN0P__1106  (.H(net1127));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[406]$_DFFE_PN0P__1107  (.H(net1128));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[407]$_DFFE_PN0P__1108  (.H(net1129));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[408]$_DFFE_PN0P__1109  (.H(net1130));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[409]$_DFFE_PN0P__1110  (.H(net1131));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[40]$_DFFE_PN0P__1111  (.H(net1132));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[410]$_DFFE_PN0P__1112  (.H(net1133));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[411]$_DFFE_PN0P__1113  (.H(net1134));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[412]$_DFFE_PN0P__1114  (.H(net1135));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[413]$_DFFE_PN0P__1115  (.H(net1136));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[414]$_DFFE_PN0P__1116  (.H(net1137));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[415]$_DFFE_PN0P__1117  (.H(net1138));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[416]$_DFFE_PN0P__1118  (.H(net1139));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[417]$_DFFE_PN0P__1119  (.H(net1140));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[418]$_DFFE_PN0P__1120  (.H(net1141));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[419]$_DFFE_PN0P__1121  (.H(net1142));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[41]$_DFFE_PN0P__1122  (.H(net1143));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[420]$_DFFE_PN0P__1123  (.H(net1144));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[421]$_DFFE_PN0P__1124  (.H(net1145));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[422]$_DFFE_PN0P__1125  (.H(net1146));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[423]$_DFFE_PN0P__1126  (.H(net1147));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[424]$_DFFE_PN0P__1127  (.H(net1148));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[425]$_DFFE_PN0P__1128  (.H(net1149));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[426]$_DFFE_PN0P__1129  (.H(net1150));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[427]$_DFFE_PN0P__1130  (.H(net1151));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[428]$_DFFE_PN0P__1131  (.H(net1152));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[429]$_DFFE_PN0P__1132  (.H(net1153));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[42]$_DFFE_PN0P__1133  (.H(net1154));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[430]$_DFFE_PN0P__1134  (.H(net1155));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[431]$_DFFE_PN0P__1135  (.H(net1156));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[432]$_DFFE_PN0P__1136  (.H(net1157));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[433]$_DFFE_PN0P__1137  (.H(net1158));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[434]$_DFFE_PN0P__1138  (.H(net1159));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[435]$_DFFE_PN0P__1139  (.H(net1160));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[436]$_DFFE_PN0P__1140  (.H(net1161));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[437]$_DFFE_PN0P__1141  (.H(net1162));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[438]$_DFFE_PN0P__1142  (.H(net1163));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[439]$_DFFE_PN0P__1143  (.H(net1164));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[43]$_DFFE_PN0P__1144  (.H(net1165));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[440]$_DFFE_PN0P__1145  (.H(net1166));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[441]$_DFFE_PN0P__1146  (.H(net1167));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[442]$_DFFE_PN0P__1147  (.H(net1168));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[443]$_DFFE_PN0P__1148  (.H(net1169));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[444]$_DFFE_PN0P__1149  (.H(net1170));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[445]$_DFFE_PN0P__1150  (.H(net1171));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[446]$_DFFE_PN0P__1151  (.H(net1172));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[447]$_DFFE_PN0P__1152  (.H(net1173));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[448]$_DFFE_PN0P__1153  (.H(net1174));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[449]$_DFFE_PN0P__1154  (.H(net1175));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[44]$_DFFE_PN0P__1155  (.H(net1176));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[450]$_DFFE_PN0P__1156  (.H(net1177));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[451]$_DFFE_PN0P__1157  (.H(net1178));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[452]$_DFFE_PN0P__1158  (.H(net1179));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[453]$_DFFE_PN0P__1159  (.H(net1180));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[454]$_DFFE_PN0P__1160  (.H(net1181));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[455]$_DFFE_PN0P__1161  (.H(net1182));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[456]$_DFFE_PN0P__1162  (.H(net1183));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[457]$_DFFE_PN0P__1163  (.H(net1184));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[458]$_DFFE_PN0P__1164  (.H(net1185));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[459]$_DFFE_PN0P__1165  (.H(net1186));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[45]$_DFFE_PN0P__1166  (.H(net1187));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[460]$_DFFE_PN0P__1167  (.H(net1188));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[461]$_DFFE_PN0P__1168  (.H(net1189));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[462]$_DFFE_PN0P__1169  (.H(net1190));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[463]$_DFFE_PN0P__1170  (.H(net1191));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[464]$_DFFE_PN0P__1171  (.H(net1192));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[465]$_DFFE_PN0P__1172  (.H(net1193));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[466]$_DFFE_PN0P__1173  (.H(net1194));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[467]$_DFFE_PN0P__1174  (.H(net1195));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[468]$_DFFE_PN0P__1175  (.H(net1196));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[469]$_DFFE_PN0P__1176  (.H(net1197));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[46]$_DFFE_PN0P__1177  (.H(net1198));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[470]$_DFFE_PN0P__1178  (.H(net1199));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[471]$_DFFE_PN0P__1179  (.H(net1200));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[472]$_DFFE_PN0P__1180  (.H(net1201));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[473]$_DFFE_PN0P__1181  (.H(net1202));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[474]$_DFFE_PN0P__1182  (.H(net1203));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[475]$_DFFE_PN0P__1183  (.H(net1204));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[476]$_DFFE_PN0P__1184  (.H(net1205));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[477]$_DFFE_PN0P__1185  (.H(net1206));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[478]$_DFFE_PN0P__1186  (.H(net1207));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[479]$_DFFE_PN0P__1187  (.H(net1208));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[47]$_DFFE_PN0P__1188  (.H(net1209));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[480]$_DFFE_PN0P__1189  (.H(net1210));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[481]$_DFFE_PN0P__1190  (.H(net1211));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[482]$_DFFE_PN0P__1191  (.H(net1212));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[483]$_DFFE_PN0P__1192  (.H(net1213));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[484]$_DFFE_PN0P__1193  (.H(net1214));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[485]$_DFFE_PN0P__1194  (.H(net1215));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[486]$_DFFE_PN0P__1195  (.H(net1216));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[487]$_DFFE_PN0P__1196  (.H(net1217));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[488]$_DFFE_PN0P__1197  (.H(net1218));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[489]$_DFFE_PN0P__1198  (.H(net1219));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[48]$_DFFE_PN0P__1199  (.H(net1220));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[490]$_DFFE_PN0P__1200  (.H(net1221));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[491]$_DFFE_PN0P__1201  (.H(net1222));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[492]$_DFFE_PN0P__1202  (.H(net1223));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[493]$_DFFE_PN0P__1203  (.H(net1224));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[494]$_DFFE_PN0P__1204  (.H(net1225));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[495]$_DFFE_PN0P__1205  (.H(net1226));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[496]$_DFFE_PN0P__1206  (.H(net1227));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[497]$_DFFE_PN0P__1207  (.H(net1228));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[498]$_DFFE_PN0P__1208  (.H(net1229));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[499]$_DFFE_PN0P__1209  (.H(net1230));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[49]$_DFFE_PN0P__1210  (.H(net1231));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[500]$_DFFE_PN0P__1211  (.H(net1232));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[501]$_DFFE_PN0P__1212  (.H(net1233));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[502]$_DFFE_PN0P__1213  (.H(net1234));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[503]$_DFFE_PN0P__1214  (.H(net1235));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[504]$_DFFE_PN0P__1215  (.H(net1236));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[505]$_DFFE_PN0P__1216  (.H(net1237));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[506]$_DFFE_PN0P__1217  (.H(net1238));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[507]$_DFFE_PN0P__1218  (.H(net1239));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[508]$_DFFE_PN0P__1219  (.H(net1240));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[509]$_DFFE_PN0P__1220  (.H(net1241));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[50]$_DFFE_PN0P__1221  (.H(net1242));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[510]$_DFFE_PN0P__1222  (.H(net1243));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[511]$_DFFE_PN0P__1223  (.H(net1244));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[512]$_DFFE_PN0P__1224  (.H(net1245));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[513]$_DFFE_PN0P__1225  (.H(net1246));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[514]$_DFFE_PN0P__1226  (.H(net1247));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[515]$_DFFE_PN0P__1227  (.H(net1248));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[516]$_DFFE_PN0P__1228  (.H(net1249));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[517]$_DFFE_PN0P__1229  (.H(net1250));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[518]$_DFFE_PN0P__1230  (.H(net1251));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[519]$_DFFE_PN0P__1231  (.H(net1252));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[51]$_DFFE_PN0P__1232  (.H(net1253));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[520]$_DFFE_PN0P__1233  (.H(net1254));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[521]$_DFFE_PN0P__1234  (.H(net1255));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[522]$_DFFE_PN0P__1235  (.H(net1256));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[523]$_DFFE_PN0P__1236  (.H(net1257));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[524]$_DFFE_PN0P__1237  (.H(net1258));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[525]$_DFFE_PN0P__1238  (.H(net1259));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[526]$_DFFE_PN0P__1239  (.H(net1260));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[527]$_DFFE_PN0P__1240  (.H(net1261));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[528]$_DFFE_PN0P__1241  (.H(net1262));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[529]$_DFFE_PN0P__1242  (.H(net1263));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[52]$_DFFE_PN0P__1243  (.H(net1264));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[530]$_DFFE_PN0P__1244  (.H(net1265));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[531]$_DFFE_PN0P__1245  (.H(net1266));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[532]$_DFFE_PN0P__1246  (.H(net1267));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[533]$_DFFE_PN0P__1247  (.H(net1268));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[534]$_DFFE_PN0P__1248  (.H(net1269));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[535]$_DFFE_PN0P__1249  (.H(net1270));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[536]$_DFFE_PN0P__1250  (.H(net1271));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[537]$_DFFE_PN0P__1251  (.H(net1272));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[538]$_DFFE_PN0P__1252  (.H(net1273));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[539]$_DFFE_PN0P__1253  (.H(net1274));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[53]$_DFFE_PN0P__1254  (.H(net1275));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[540]$_DFFE_PN0P__1255  (.H(net1276));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[541]$_DFFE_PN0P__1256  (.H(net1277));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[542]$_DFFE_PN0P__1257  (.H(net1278));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[543]$_DFFE_PN0P__1258  (.H(net1279));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[544]$_DFFE_PN0P__1259  (.H(net1280));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[545]$_DFFE_PN0P__1260  (.H(net1281));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[546]$_DFFE_PN0P__1261  (.H(net1282));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[547]$_DFFE_PN0P__1262  (.H(net1283));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[548]$_DFFE_PN0P__1263  (.H(net1284));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[549]$_DFFE_PN0P__1264  (.H(net1285));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[54]$_DFFE_PN0P__1265  (.H(net1286));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[550]$_DFFE_PN0P__1266  (.H(net1287));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[551]$_DFFE_PN0P__1267  (.H(net1288));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[552]$_DFFE_PN0P__1268  (.H(net1289));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[553]$_DFFE_PN0P__1269  (.H(net1290));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[554]$_DFFE_PN0P__1270  (.H(net1291));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[555]$_DFFE_PN0P__1271  (.H(net1292));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[556]$_DFFE_PN0P__1272  (.H(net1293));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[557]$_DFFE_PN0P__1273  (.H(net1294));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[558]$_DFFE_PN0P__1274  (.H(net1295));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[559]$_DFFE_PN0P__1275  (.H(net1296));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[55]$_DFFE_PN0P__1276  (.H(net1297));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[560]$_DFFE_PN0P__1277  (.H(net1298));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[561]$_DFFE_PN0P__1278  (.H(net1299));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[562]$_DFFE_PN0P__1279  (.H(net1300));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[563]$_DFFE_PN0P__1280  (.H(net1301));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[564]$_DFFE_PN0P__1281  (.H(net1302));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[565]$_DFFE_PN0P__1282  (.H(net1303));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[566]$_DFFE_PN0P__1283  (.H(net1304));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[567]$_DFFE_PN0P__1284  (.H(net1305));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[568]$_DFFE_PN0P__1285  (.H(net1306));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[569]$_DFFE_PN0P__1286  (.H(net1307));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[56]$_DFFE_PN0P__1287  (.H(net1308));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[570]$_DFFE_PN0P__1288  (.H(net1309));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[571]$_DFFE_PN0P__1289  (.H(net1310));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[572]$_DFFE_PN0P__1290  (.H(net1311));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[573]$_DFFE_PN0P__1291  (.H(net1312));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[574]$_DFFE_PN0P__1292  (.H(net1313));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[575]$_DFFE_PN0P__1293  (.H(net1314));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[576]$_DFFE_PN0P__1294  (.H(net1315));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[577]$_DFFE_PN0P__1295  (.H(net1316));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[578]$_DFFE_PN0P__1296  (.H(net1317));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[579]$_DFFE_PN0P__1297  (.H(net1318));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[57]$_DFFE_PN0P__1298  (.H(net1319));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[580]$_DFFE_PN0P__1299  (.H(net1320));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[581]$_DFFE_PN0P__1300  (.H(net1321));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[582]$_DFFE_PN0P__1301  (.H(net1322));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[583]$_DFFE_PN0P__1302  (.H(net1323));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[584]$_DFFE_PN0P__1303  (.H(net1324));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[585]$_DFFE_PN0P__1304  (.H(net1325));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[586]$_DFFE_PN0P__1305  (.H(net1326));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[587]$_DFFE_PN0P__1306  (.H(net1327));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[588]$_DFFE_PN0P__1307  (.H(net1328));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[589]$_DFFE_PN0P__1308  (.H(net1329));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[58]$_DFFE_PN0P__1309  (.H(net1330));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[590]$_DFFE_PN0P__1310  (.H(net1331));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[591]$_DFFE_PN0P__1311  (.H(net1332));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[592]$_DFFE_PN0P__1312  (.H(net1333));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[593]$_DFFE_PN0P__1313  (.H(net1334));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[594]$_DFFE_PN0P__1314  (.H(net1335));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[595]$_DFFE_PN0P__1315  (.H(net1336));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[596]$_DFFE_PN0P__1316  (.H(net1337));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[597]$_DFFE_PN0P__1317  (.H(net1338));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[598]$_DFFE_PN0P__1318  (.H(net1339));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[599]$_DFFE_PN0P__1319  (.H(net1340));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[59]$_DFFE_PN0P__1320  (.H(net1341));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[600]$_DFFE_PN0P__1321  (.H(net1342));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[601]$_DFFE_PN0P__1322  (.H(net1343));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[602]$_DFFE_PN0P__1323  (.H(net1344));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[603]$_DFFE_PN0P__1324  (.H(net1345));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[604]$_DFFE_PN0P__1325  (.H(net1346));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[605]$_DFFE_PN0P__1326  (.H(net1347));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[606]$_DFFE_PN0P__1327  (.H(net1348));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[607]$_DFFE_PN0P__1328  (.H(net1349));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[608]$_DFFE_PN0P__1329  (.H(net1350));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[609]$_DFFE_PN0P__1330  (.H(net1351));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[60]$_DFFE_PN0P__1331  (.H(net1352));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[610]$_DFFE_PN0P__1332  (.H(net1353));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[611]$_DFFE_PN0P__1333  (.H(net1354));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[612]$_DFFE_PN0P__1334  (.H(net1355));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[613]$_DFFE_PN0P__1335  (.H(net1356));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[614]$_DFFE_PN0P__1336  (.H(net1357));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[615]$_DFFE_PN0P__1337  (.H(net1358));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[616]$_DFFE_PN0P__1338  (.H(net1359));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[617]$_DFFE_PN0P__1339  (.H(net1360));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[618]$_DFFE_PN0P__1340  (.H(net1361));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[619]$_DFFE_PN0P__1341  (.H(net1362));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[61]$_DFFE_PN0P__1342  (.H(net1363));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[620]$_DFFE_PN0P__1343  (.H(net1364));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[621]$_DFFE_PN0P__1344  (.H(net1365));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[622]$_DFFE_PN0P__1345  (.H(net1366));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[623]$_DFFE_PN0P__1346  (.H(net1367));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[624]$_DFFE_PN0P__1347  (.H(net1368));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[625]$_DFFE_PN0P__1348  (.H(net1369));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[626]$_DFFE_PN0P__1349  (.H(net1370));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[627]$_DFFE_PN0P__1350  (.H(net1371));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[628]$_DFFE_PN0P__1351  (.H(net1372));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[629]$_DFFE_PN0P__1352  (.H(net1373));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[62]$_DFFE_PN0P__1353  (.H(net1374));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[630]$_DFFE_PN0P__1354  (.H(net1375));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[631]$_DFFE_PN0P__1355  (.H(net1376));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[632]$_DFFE_PN0P__1356  (.H(net1377));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[633]$_DFFE_PN0P__1357  (.H(net1378));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[634]$_DFFE_PN0P__1358  (.H(net1379));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[635]$_DFFE_PN0P__1359  (.H(net1380));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[636]$_DFFE_PN0P__1360  (.H(net1381));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[637]$_DFFE_PN0P__1361  (.H(net1382));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[638]$_DFFE_PN0P__1362  (.H(net1383));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[639]$_DFFE_PN0P__1363  (.H(net1384));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[63]$_DFFE_PN0P__1364  (.H(net1385));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[640]$_DFFE_PN0P__1365  (.H(net1386));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[641]$_DFFE_PN0P__1366  (.H(net1387));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[642]$_DFFE_PN0P__1367  (.H(net1388));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[643]$_DFFE_PN0P__1368  (.H(net1389));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[644]$_DFFE_PN0P__1369  (.H(net1390));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[645]$_DFFE_PN0P__1370  (.H(net1391));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[646]$_DFFE_PN0P__1371  (.H(net1392));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[647]$_DFFE_PN0P__1372  (.H(net1393));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[648]$_DFFE_PN0P__1373  (.H(net1394));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[649]$_DFFE_PN0P__1374  (.H(net1395));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[64]$_DFFE_PN0P__1375  (.H(net1396));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[650]$_DFFE_PN0P__1376  (.H(net1397));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[651]$_DFFE_PN0P__1377  (.H(net1398));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[652]$_DFFE_PN0P__1378  (.H(net1399));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[653]$_DFFE_PN0P__1379  (.H(net1400));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[654]$_DFFE_PN0P__1380  (.H(net1401));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[655]$_DFFE_PN0P__1381  (.H(net1402));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[656]$_DFFE_PN0P__1382  (.H(net1403));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[657]$_DFFE_PN0P__1383  (.H(net1404));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[658]$_DFFE_PN0P__1384  (.H(net1405));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[659]$_DFFE_PN0P__1385  (.H(net1406));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[65]$_DFFE_PN0P__1386  (.H(net1407));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[660]$_DFFE_PN0P__1387  (.H(net1408));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[661]$_DFFE_PN0P__1388  (.H(net1409));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[662]$_DFFE_PN0P__1389  (.H(net1410));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[663]$_DFFE_PN0P__1390  (.H(net1411));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[664]$_DFFE_PN0P__1391  (.H(net1412));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[665]$_DFFE_PN0P__1392  (.H(net1413));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[666]$_DFFE_PN0P__1393  (.H(net1414));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[667]$_DFFE_PN0P__1394  (.H(net1415));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[668]$_DFFE_PN0P__1395  (.H(net1416));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[669]$_DFFE_PN0P__1396  (.H(net1417));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[66]$_DFFE_PN0P__1397  (.H(net1418));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[670]$_DFFE_PN0P__1398  (.H(net1419));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[671]$_DFFE_PN0P__1399  (.H(net1420));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[672]$_DFFE_PN0P__1400  (.H(net1421));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[673]$_DFFE_PN0P__1401  (.H(net1422));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[674]$_DFFE_PN0P__1402  (.H(net1423));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[675]$_DFFE_PN0P__1403  (.H(net1424));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[676]$_DFFE_PN0P__1404  (.H(net1425));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[677]$_DFFE_PN0P__1405  (.H(net1426));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[678]$_DFFE_PN0P__1406  (.H(net1427));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[679]$_DFFE_PN0P__1407  (.H(net1428));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[67]$_DFFE_PN0P__1408  (.H(net1429));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[680]$_DFFE_PN0P__1409  (.H(net1430));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[681]$_DFFE_PN0P__1410  (.H(net1431));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[682]$_DFFE_PN0P__1411  (.H(net1432));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[683]$_DFFE_PN0P__1412  (.H(net1433));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[684]$_DFFE_PN0P__1413  (.H(net1434));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[685]$_DFFE_PN0P__1414  (.H(net1435));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[686]$_DFFE_PN0P__1415  (.H(net1436));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[687]$_DFFE_PN0P__1416  (.H(net1437));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[688]$_DFFE_PN0P__1417  (.H(net1438));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[689]$_DFFE_PN0P__1418  (.H(net1439));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[68]$_DFFE_PN0P__1419  (.H(net1440));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[690]$_DFFE_PN0P__1420  (.H(net1441));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[691]$_DFFE_PN0P__1421  (.H(net1442));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[692]$_DFFE_PN0P__1422  (.H(net1443));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[693]$_DFFE_PN0P__1423  (.H(net1444));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[694]$_DFFE_PN0P__1424  (.H(net1445));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[695]$_DFFE_PN0P__1425  (.H(net1446));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[696]$_DFFE_PN0P__1426  (.H(net1447));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[697]$_DFFE_PN0P__1427  (.H(net1448));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[698]$_DFFE_PN0P__1428  (.H(net1449));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[699]$_DFFE_PN0P__1429  (.H(net1450));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[69]$_DFFE_PN0P__1430  (.H(net1451));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[700]$_DFFE_PN0P__1431  (.H(net1452));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[701]$_DFFE_PN0P__1432  (.H(net1453));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[702]$_DFFE_PN0P__1433  (.H(net1454));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[703]$_DFFE_PN0P__1434  (.H(net1455));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[704]$_DFFE_PN0P__1435  (.H(net1456));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[705]$_DFFE_PN0P__1436  (.H(net1457));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[706]$_DFFE_PN0P__1437  (.H(net1458));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[707]$_DFFE_PN0P__1438  (.H(net1459));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[708]$_DFFE_PN0P__1439  (.H(net1460));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[709]$_DFFE_PN0P__1440  (.H(net1461));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[70]$_DFFE_PN0P__1441  (.H(net1462));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[710]$_DFFE_PN0P__1442  (.H(net1463));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[711]$_DFFE_PN0P__1443  (.H(net1464));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[712]$_DFFE_PN0P__1444  (.H(net1465));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[713]$_DFFE_PN0P__1445  (.H(net1466));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[714]$_DFFE_PN0P__1446  (.H(net1467));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[715]$_DFFE_PN0P__1447  (.H(net1468));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[716]$_DFFE_PN0P__1448  (.H(net1469));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[717]$_DFFE_PN0P__1449  (.H(net1470));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[718]$_DFFE_PN0P__1450  (.H(net1471));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[719]$_DFFE_PN0P__1451  (.H(net1472));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[71]$_DFFE_PN0P__1452  (.H(net1473));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[720]$_DFFE_PN0P__1453  (.H(net1474));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[721]$_DFFE_PN0P__1454  (.H(net1475));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[722]$_DFFE_PN0P__1455  (.H(net1476));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[723]$_DFFE_PN0P__1456  (.H(net1477));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[724]$_DFFE_PN0P__1457  (.H(net1478));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[725]$_DFFE_PN0P__1458  (.H(net1479));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[726]$_DFFE_PN0P__1459  (.H(net1480));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[727]$_DFFE_PN0P__1460  (.H(net1481));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[728]$_DFFE_PN0P__1461  (.H(net1482));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[729]$_DFFE_PN0P__1462  (.H(net1483));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[72]$_DFFE_PN0P__1463  (.H(net1484));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[730]$_DFFE_PN0P__1464  (.H(net1485));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[731]$_DFFE_PN0P__1465  (.H(net1486));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[732]$_DFFE_PN0P__1466  (.H(net1487));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[733]$_DFFE_PN0P__1467  (.H(net1488));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[734]$_DFFE_PN0P__1468  (.H(net1489));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[735]$_DFFE_PN0P__1469  (.H(net1490));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[736]$_DFFE_PN0P__1470  (.H(net1491));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[737]$_DFFE_PN0P__1471  (.H(net1492));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[738]$_DFFE_PN0P__1472  (.H(net1493));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[739]$_DFFE_PN0P__1473  (.H(net1494));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[73]$_DFFE_PN0P__1474  (.H(net1495));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[740]$_DFFE_PN0P__1475  (.H(net1496));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[741]$_DFFE_PN0P__1476  (.H(net1497));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[742]$_DFFE_PN0P__1477  (.H(net1498));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[743]$_DFFE_PN0P__1478  (.H(net1499));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[744]$_DFFE_PN0P__1479  (.H(net1500));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[745]$_DFFE_PN0P__1480  (.H(net1501));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[746]$_DFFE_PN0P__1481  (.H(net1502));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[747]$_DFFE_PN0P__1482  (.H(net1503));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[748]$_DFFE_PN0P__1483  (.H(net1504));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[749]$_DFFE_PN0P__1484  (.H(net1505));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[74]$_DFFE_PN0P__1485  (.H(net1506));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[750]$_DFFE_PN0P__1486  (.H(net1507));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[751]$_DFFE_PN0P__1487  (.H(net1508));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[752]$_DFFE_PN0P__1488  (.H(net1509));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[753]$_DFFE_PN0P__1489  (.H(net1510));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[754]$_DFFE_PN0P__1490  (.H(net1511));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[755]$_DFFE_PN0P__1491  (.H(net1512));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[756]$_DFFE_PN0P__1492  (.H(net1513));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[757]$_DFFE_PN0P__1493  (.H(net1514));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[758]$_DFFE_PN0P__1494  (.H(net1515));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[759]$_DFFE_PN0P__1495  (.H(net1516));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[75]$_DFFE_PN0P__1496  (.H(net1517));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[760]$_DFFE_PN0P__1497  (.H(net1518));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[761]$_DFFE_PN0P__1498  (.H(net1519));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[762]$_DFFE_PN0P__1499  (.H(net1520));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[763]$_DFFE_PN0P__1500  (.H(net1521));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[764]$_DFFE_PN0P__1501  (.H(net1522));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[765]$_DFFE_PN0P__1502  (.H(net1523));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[766]$_DFFE_PN0P__1503  (.H(net1524));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[767]$_DFFE_PN0P__1504  (.H(net1525));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[768]$_DFFE_PN0P__1505  (.H(net1526));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[769]$_DFFE_PN0P__1506  (.H(net1527));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[76]$_DFFE_PN0P__1507  (.H(net1528));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[770]$_DFFE_PN0P__1508  (.H(net1529));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[771]$_DFFE_PN0P__1509  (.H(net1530));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[772]$_DFFE_PN0P__1510  (.H(net1531));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[773]$_DFFE_PN0P__1511  (.H(net1532));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[774]$_DFFE_PN0P__1512  (.H(net1533));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[775]$_DFFE_PN0P__1513  (.H(net1534));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[776]$_DFFE_PN0P__1514  (.H(net1535));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[777]$_DFFE_PN0P__1515  (.H(net1536));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[778]$_DFFE_PN0P__1516  (.H(net1537));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[779]$_DFFE_PN0P__1517  (.H(net1538));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[77]$_DFFE_PN0P__1518  (.H(net1539));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[780]$_DFFE_PN0P__1519  (.H(net1540));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[781]$_DFFE_PN0P__1520  (.H(net1541));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[782]$_DFFE_PN0P__1521  (.H(net1542));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[783]$_DFFE_PN0P__1522  (.H(net1543));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[784]$_DFFE_PN0P__1523  (.H(net1544));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[785]$_DFFE_PN0P__1524  (.H(net1545));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[786]$_DFFE_PN0P__1525  (.H(net1546));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[787]$_DFFE_PN0P__1526  (.H(net1547));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[788]$_DFFE_PN0P__1527  (.H(net1548));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[789]$_DFFE_PN0P__1528  (.H(net1549));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[78]$_DFFE_PN0P__1529  (.H(net1550));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[790]$_DFFE_PN0P__1530  (.H(net1551));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[791]$_DFFE_PN0P__1531  (.H(net1552));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[792]$_DFFE_PN0P__1532  (.H(net1553));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[793]$_DFFE_PN0P__1533  (.H(net1554));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[794]$_DFFE_PN0P__1534  (.H(net1555));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[795]$_DFFE_PN0P__1535  (.H(net1556));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[796]$_DFFE_PN0P__1536  (.H(net1557));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[797]$_DFFE_PN0P__1537  (.H(net1558));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[798]$_DFFE_PN0P__1538  (.H(net1559));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[799]$_DFFE_PN0P__1539  (.H(net1560));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[79]$_DFFE_PN0P__1540  (.H(net1561));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[800]$_DFFE_PN0P__1541  (.H(net1562));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[801]$_DFFE_PN0P__1542  (.H(net1563));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[802]$_DFFE_PN0P__1543  (.H(net1564));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[803]$_DFFE_PN0P__1544  (.H(net1565));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[804]$_DFFE_PN0P__1545  (.H(net1566));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[805]$_DFFE_PN0P__1546  (.H(net1567));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[806]$_DFFE_PN0P__1547  (.H(net1568));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[807]$_DFFE_PN0P__1548  (.H(net1569));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[808]$_DFFE_PN0P__1549  (.H(net1570));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[809]$_DFFE_PN0P__1550  (.H(net1571));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[80]$_DFFE_PN0P__1551  (.H(net1572));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[810]$_DFFE_PN0P__1552  (.H(net1573));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[811]$_DFFE_PN0P__1553  (.H(net1574));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[812]$_DFFE_PN0P__1554  (.H(net1575));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[813]$_DFFE_PN0P__1555  (.H(net1576));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[814]$_DFFE_PN0P__1556  (.H(net1577));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[815]$_DFFE_PN0P__1557  (.H(net1578));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[816]$_DFFE_PN0P__1558  (.H(net1579));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[817]$_DFFE_PN0P__1559  (.H(net1580));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[818]$_DFFE_PN0P__1560  (.H(net1581));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[819]$_DFFE_PN0P__1561  (.H(net1582));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[81]$_DFFE_PN0P__1562  (.H(net1583));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[820]$_DFFE_PN0P__1563  (.H(net1584));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[821]$_DFFE_PN0P__1564  (.H(net1585));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[822]$_DFFE_PN0P__1565  (.H(net1586));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[823]$_DFFE_PN0P__1566  (.H(net1587));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[824]$_DFFE_PN0P__1567  (.H(net1588));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[825]$_DFFE_PN0P__1568  (.H(net1589));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[826]$_DFFE_PN0P__1569  (.H(net1590));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[827]$_DFFE_PN0P__1570  (.H(net1591));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[828]$_DFFE_PN0P__1571  (.H(net1592));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[829]$_DFFE_PN0P__1572  (.H(net1593));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[82]$_DFFE_PN0P__1573  (.H(net1594));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[830]$_DFFE_PN0P__1574  (.H(net1595));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[831]$_DFFE_PN0P__1575  (.H(net1596));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[832]$_DFFE_PN0P__1576  (.H(net1597));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[833]$_DFFE_PN0P__1577  (.H(net1598));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[834]$_DFFE_PN0P__1578  (.H(net1599));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[835]$_DFFE_PN0P__1579  (.H(net1600));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[836]$_DFFE_PN0P__1580  (.H(net1601));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[837]$_DFFE_PN0P__1581  (.H(net1602));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[838]$_DFFE_PN0P__1582  (.H(net1603));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[839]$_DFFE_PN0P__1583  (.H(net1604));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[83]$_DFFE_PN0P__1584  (.H(net1605));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[840]$_DFFE_PN0P__1585  (.H(net1606));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[841]$_DFFE_PN0P__1586  (.H(net1607));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[842]$_DFFE_PN0P__1587  (.H(net1608));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[843]$_DFFE_PN0P__1588  (.H(net1609));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[844]$_DFFE_PN0P__1589  (.H(net1610));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[845]$_DFFE_PN0P__1590  (.H(net1611));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[846]$_DFFE_PN0P__1591  (.H(net1612));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[847]$_DFFE_PN0P__1592  (.H(net1613));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[848]$_DFFE_PN0P__1593  (.H(net1614));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[849]$_DFFE_PN0P__1594  (.H(net1615));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[84]$_DFFE_PN0P__1595  (.H(net1616));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[850]$_DFFE_PN0P__1596  (.H(net1617));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[851]$_DFFE_PN0P__1597  (.H(net1618));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[852]$_DFFE_PN0P__1598  (.H(net1619));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[853]$_DFFE_PN0P__1599  (.H(net1620));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[854]$_DFFE_PN0P__1600  (.H(net1621));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[855]$_DFFE_PN0P__1601  (.H(net1622));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[856]$_DFFE_PN0P__1602  (.H(net1623));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[857]$_DFFE_PN0P__1603  (.H(net1624));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[858]$_DFFE_PN0P__1604  (.H(net1625));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[859]$_DFFE_PN0P__1605  (.H(net1626));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[85]$_DFFE_PN0P__1606  (.H(net1627));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[860]$_DFFE_PN0P__1607  (.H(net1628));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[861]$_DFFE_PN0P__1608  (.H(net1629));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[862]$_DFFE_PN0P__1609  (.H(net1630));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[863]$_DFFE_PN0P__1610  (.H(net1631));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[864]$_DFFE_PN0P__1611  (.H(net1632));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[865]$_DFFE_PN0P__1612  (.H(net1633));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[866]$_DFFE_PN0P__1613  (.H(net1634));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[867]$_DFFE_PN0P__1614  (.H(net1635));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[868]$_DFFE_PN0P__1615  (.H(net1636));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[869]$_DFFE_PN0P__1616  (.H(net1637));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[86]$_DFFE_PN0P__1617  (.H(net1638));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[870]$_DFFE_PN0P__1618  (.H(net1639));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[871]$_DFFE_PN0P__1619  (.H(net1640));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[872]$_DFFE_PN0P__1620  (.H(net1641));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[873]$_DFFE_PN0P__1621  (.H(net1642));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[874]$_DFFE_PN0P__1622  (.H(net1643));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[875]$_DFFE_PN0P__1623  (.H(net1644));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[876]$_DFFE_PN0P__1624  (.H(net1645));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[877]$_DFFE_PN0P__1625  (.H(net1646));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[878]$_DFFE_PN0P__1626  (.H(net1647));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[879]$_DFFE_PN0P__1627  (.H(net1648));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[87]$_DFFE_PN0P__1628  (.H(net1649));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[880]$_DFFE_PN0P__1629  (.H(net1650));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[881]$_DFFE_PN0P__1630  (.H(net1651));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[882]$_DFFE_PN0P__1631  (.H(net1652));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[883]$_DFFE_PN0P__1632  (.H(net1653));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[884]$_DFFE_PN0P__1633  (.H(net1654));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[885]$_DFFE_PN0P__1634  (.H(net1655));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[886]$_DFFE_PN0P__1635  (.H(net1656));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[887]$_DFFE_PN0P__1636  (.H(net1657));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[888]$_DFFE_PN0P__1637  (.H(net1658));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[889]$_DFFE_PN0P__1638  (.H(net1659));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[88]$_DFFE_PN0P__1639  (.H(net1660));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[890]$_DFFE_PN0P__1640  (.H(net1661));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[891]$_DFFE_PN0P__1641  (.H(net1662));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[892]$_DFFE_PN0P__1642  (.H(net1663));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[893]$_DFFE_PN0P__1643  (.H(net1664));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[894]$_DFFE_PN0P__1644  (.H(net1665));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[895]$_DFFE_PN0P__1645  (.H(net1666));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[896]$_DFFE_PN0P__1646  (.H(net1667));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[897]$_DFFE_PN0P__1647  (.H(net1668));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[898]$_DFFE_PN0P__1648  (.H(net1669));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[899]$_DFFE_PN0P__1649  (.H(net1670));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[89]$_DFFE_PN0P__1650  (.H(net1671));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[900]$_DFFE_PN0P__1651  (.H(net1672));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[901]$_DFFE_PN0P__1652  (.H(net1673));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[902]$_DFFE_PN0P__1653  (.H(net1674));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[903]$_DFFE_PN0P__1654  (.H(net1675));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[904]$_DFFE_PN0P__1655  (.H(net1676));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[905]$_DFFE_PN0P__1656  (.H(net1677));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[906]$_DFFE_PN0P__1657  (.H(net1678));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[907]$_DFFE_PN0P__1658  (.H(net1679));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[908]$_DFFE_PN0P__1659  (.H(net1680));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[909]$_DFFE_PN0P__1660  (.H(net1681));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[90]$_DFFE_PN0P__1661  (.H(net1682));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[910]$_DFFE_PN0P__1662  (.H(net1683));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[911]$_DFFE_PN0P__1663  (.H(net1684));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[912]$_DFFE_PN0P__1664  (.H(net1685));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[913]$_DFFE_PN0P__1665  (.H(net1686));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[914]$_DFFE_PN0P__1666  (.H(net1687));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[915]$_DFFE_PN0P__1667  (.H(net1688));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[916]$_DFFE_PN0P__1668  (.H(net1689));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[917]$_DFFE_PN0P__1669  (.H(net1690));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[918]$_DFFE_PN0P__1670  (.H(net1691));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[919]$_DFFE_PN0P__1671  (.H(net1692));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[91]$_DFFE_PN0P__1672  (.H(net1693));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[920]$_DFFE_PN0P__1673  (.H(net1694));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[921]$_DFFE_PN0P__1674  (.H(net1695));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[922]$_DFFE_PN0P__1675  (.H(net1696));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[923]$_DFFE_PN0P__1676  (.H(net1697));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[924]$_DFFE_PN0P__1677  (.H(net1698));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[925]$_DFFE_PN0P__1678  (.H(net1699));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[926]$_DFFE_PN0P__1679  (.H(net1700));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[927]$_DFFE_PN0P__1680  (.H(net1701));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[928]$_DFFE_PN0P__1681  (.H(net1702));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[929]$_DFFE_PN0P__1682  (.H(net1703));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[92]$_DFFE_PN0P__1683  (.H(net1704));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[930]$_DFFE_PN0P__1684  (.H(net1705));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[931]$_DFFE_PN0P__1685  (.H(net1706));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[932]$_DFFE_PN0P__1686  (.H(net1707));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[933]$_DFFE_PN0P__1687  (.H(net1708));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[934]$_DFFE_PN0P__1688  (.H(net1709));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[935]$_DFFE_PN0P__1689  (.H(net1710));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[936]$_DFFE_PN0P__1690  (.H(net1711));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[937]$_DFFE_PN0P__1691  (.H(net1712));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[938]$_DFFE_PN0P__1692  (.H(net1713));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[939]$_DFFE_PN0P__1693  (.H(net1714));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[93]$_DFFE_PN0P__1694  (.H(net1715));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[940]$_DFFE_PN0P__1695  (.H(net1716));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[941]$_DFFE_PN0P__1696  (.H(net1717));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[942]$_DFFE_PN0P__1697  (.H(net1718));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[943]$_DFFE_PN0P__1698  (.H(net1719));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[944]$_DFFE_PN0P__1699  (.H(net1720));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[945]$_DFFE_PN0P__1700  (.H(net1721));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[946]$_DFFE_PN0P__1701  (.H(net1722));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[947]$_DFFE_PN0P__1702  (.H(net1723));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[948]$_DFFE_PN0P__1703  (.H(net1724));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[949]$_DFFE_PN0P__1704  (.H(net1725));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[94]$_DFFE_PN0P__1705  (.H(net1726));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[950]$_DFFE_PN0P__1706  (.H(net1727));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[951]$_DFFE_PN0P__1707  (.H(net1728));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[952]$_DFFE_PN0P__1708  (.H(net1729));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[953]$_DFFE_PN0P__1709  (.H(net1730));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[954]$_DFFE_PN0P__1710  (.H(net1731));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[955]$_DFFE_PN0P__1711  (.H(net1732));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[956]$_DFFE_PN0P__1712  (.H(net1733));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[957]$_DFFE_PN0P__1713  (.H(net1734));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[958]$_DFFE_PN0P__1714  (.H(net1735));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[959]$_DFFE_PN0P__1715  (.H(net1736));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[95]$_DFFE_PN0P__1716  (.H(net1737));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[960]$_DFFE_PN0P__1717  (.H(net1738));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[961]$_DFFE_PN0P__1718  (.H(net1739));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[962]$_DFFE_PN0P__1719  (.H(net1740));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[963]$_DFFE_PN0P__1720  (.H(net1741));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[964]$_DFFE_PN0P__1721  (.H(net1742));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[965]$_DFFE_PN0P__1722  (.H(net1743));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[966]$_DFFE_PN0P__1723  (.H(net1744));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[967]$_DFFE_PN0P__1724  (.H(net1745));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[968]$_DFFE_PN0P__1725  (.H(net1746));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[969]$_DFFE_PN0P__1726  (.H(net1747));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[96]$_DFFE_PN0P__1727  (.H(net1748));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[970]$_DFFE_PN0P__1728  (.H(net1749));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[971]$_DFFE_PN0P__1729  (.H(net1750));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[972]$_DFFE_PN0P__1730  (.H(net1751));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[973]$_DFFE_PN0P__1731  (.H(net1752));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[974]$_DFFE_PN0P__1732  (.H(net1753));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[975]$_DFFE_PN0P__1733  (.H(net1754));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[976]$_DFFE_PN0P__1734  (.H(net1755));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[977]$_DFFE_PN0P__1735  (.H(net1756));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[978]$_DFFE_PN0P__1736  (.H(net1757));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[979]$_DFFE_PN0P__1737  (.H(net1758));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[97]$_DFFE_PN0P__1738  (.H(net1759));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[980]$_DFFE_PN0P__1739  (.H(net1760));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[981]$_DFFE_PN0P__1740  (.H(net1761));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[982]$_DFFE_PN0P__1741  (.H(net1762));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[983]$_DFFE_PN0P__1742  (.H(net1763));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[984]$_DFFE_PN0P__1743  (.H(net1764));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[985]$_DFFE_PN0P__1744  (.H(net1765));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[986]$_DFFE_PN0P__1745  (.H(net1766));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[987]$_DFFE_PN0P__1746  (.H(net1767));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[988]$_DFFE_PN0P__1747  (.H(net1768));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[989]$_DFFE_PN0P__1748  (.H(net1769));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[98]$_DFFE_PN0P__1749  (.H(net1770));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[990]$_DFFE_PN0P__1750  (.H(net1771));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[991]$_DFFE_PN0P__1751  (.H(net1772));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[992]$_DFFE_PN0P__1752  (.H(net1773));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[993]$_DFFE_PN0P__1753  (.H(net1774));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[994]$_DFFE_PN0P__1754  (.H(net1775));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[995]$_DFFE_PN0P__1755  (.H(net1776));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[996]$_DFFE_PN0P__1756  (.H(net1777));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[997]$_DFFE_PN0P__1757  (.H(net1778));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[998]$_DFFE_PN0P__1758  (.H(net1779));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[999]$_DFFE_PN0P__1759  (.H(net1780));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg[99]$_DFFE_PN0P__1760  (.H(net1781));
 TIEHIx1_ASAP7_75t_R \id_stage_i.branch_set$_DFF_PN0__1761  (.H(net1782));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFFE_PN0P__1762  (.H(net1783));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[1]$_DFFE_PN0P__1763  (.H(net1784));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[2]$_DFFE_PN0P__1764  (.H(net1785));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[3]$_DFFE_PN0P__1765  (.H(net1786));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.debug_mode_o$_DFFE_PN0P__1766  (.H(net1787));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.exc_req_q$_DFF_PN0__1767  (.H(net1788));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.illegal_insn_q$_DFF_PN0__1768  (.H(net1789));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.load_err_q$_DFF_PN0__1769  (.H(net1790));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.nmi_mode_o$_DFFE_PN0P__1770  (.H(net1791));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.store_err_q$_DFF_PN0__1771  (.H(net1792));
 TIEHIx1_ASAP7_75t_R \id_stage_i.id_fsm_q$_DFFE_PN0P__1772  (.H(net1793));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[0]$_DFFE_PN0P__1773  (.H(net1794));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[10]$_DFFE_PN0P__1774  (.H(net1795));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[11]$_DFFE_PN0P__1775  (.H(net1796));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[12]$_DFFE_PN0P__1776  (.H(net1797));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[13]$_DFFE_PN0P__1777  (.H(net1798));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[14]$_DFFE_PN0P__1778  (.H(net1799));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[15]$_DFFE_PN0P__1779  (.H(net1800));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[16]$_DFFE_PN0P__1780  (.H(net1801));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[17]$_DFFE_PN0P__1781  (.H(net1802));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[18]$_DFFE_PN0P__1782  (.H(net1803));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[19]$_DFFE_PN0P__1783  (.H(net1804));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[1]$_DFFE_PN0P__1784  (.H(net1805));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[20]$_DFFE_PN0P__1785  (.H(net1806));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[21]$_DFFE_PN0P__1786  (.H(net1807));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[22]$_DFFE_PN0P__1787  (.H(net1808));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[23]$_DFFE_PN0P__1788  (.H(net1809));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[24]$_DFFE_PN0P__1789  (.H(net1810));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[25]$_DFFE_PN0P__1790  (.H(net1811));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[26]$_DFFE_PN0P__1791  (.H(net1812));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[27]$_DFFE_PN0P__1792  (.H(net1813));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[28]$_DFFE_PN0P__1793  (.H(net1814));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[29]$_DFFE_PN0P__1794  (.H(net1815));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[2]$_DFFE_PN0P__1795  (.H(net1816));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[30]$_DFFE_PN0P__1796  (.H(net1817));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[31]$_DFFE_PN0P__1797  (.H(net1818));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[34]$_DFFE_PN0P__1798  (.H(net1819));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[35]$_DFFE_PN0P__1799  (.H(net1820));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[36]$_DFFE_PN0P__1800  (.H(net1821));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[37]$_DFFE_PN0P__1801  (.H(net1822));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[38]$_DFFE_PN0P__1802  (.H(net1823));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[39]$_DFFE_PN0P__1803  (.H(net1824));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[3]$_DFFE_PN0P__1804  (.H(net1825));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[40]$_DFFE_PN0P__1805  (.H(net1826));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[41]$_DFFE_PN0P__1806  (.H(net1827));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[42]$_DFFE_PN0P__1807  (.H(net1828));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[43]$_DFFE_PN0P__1808  (.H(net1829));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[44]$_DFFE_PN0P__1809  (.H(net1830));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[45]$_DFFE_PN0P__1810  (.H(net1831));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[46]$_DFFE_PN0P__1811  (.H(net1832));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[47]$_DFFE_PN0P__1812  (.H(net1833));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[48]$_DFFE_PN0P__1813  (.H(net1834));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[49]$_DFFE_PN0P__1814  (.H(net1835));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[4]$_DFFE_PN0P__1815  (.H(net1836));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[50]$_DFFE_PN0P__1816  (.H(net1837));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[51]$_DFFE_PN0P__1817  (.H(net1838));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[52]$_DFFE_PN0P__1818  (.H(net1839));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[53]$_DFFE_PN0P__1819  (.H(net1840));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[54]$_DFFE_PN0P__1820  (.H(net1841));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[55]$_DFFE_PN0P__1821  (.H(net1842));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[56]$_DFFE_PN0P__1822  (.H(net1843));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[57]$_DFFE_PN0P__1823  (.H(net1844));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[58]$_DFFE_PN0P__1824  (.H(net1845));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[59]$_DFFE_PN0P__1825  (.H(net1846));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[5]$_DFFE_PN0P__1826  (.H(net1847));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[60]$_DFFE_PN0P__1827  (.H(net1848));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[61]$_DFFE_PN0P__1828  (.H(net1849));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[62]$_DFFE_PN0P__1829  (.H(net1850));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[63]$_DFFE_PN0P__1830  (.H(net1851));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[64]$_DFFE_PN0P__1831  (.H(net1852));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[65]$_DFFE_PN0P__1832  (.H(net1853));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[66]$_DFFE_PN0P__1833  (.H(net1854));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[67]$_DFFE_PN0P__1834  (.H(net1855));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[6]$_DFFE_PN0P__1835  (.H(net1856));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[7]$_DFFE_PN0P__1836  (.H(net1857));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[8]$_DFFE_PN0P__1837  (.H(net1858));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q_ex_o[9]$_DFFE_PN0P__1838  (.H(net1859));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0__1839  (.H(net1860));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0__1840  (.H(net1861));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0__1841  (.H(net1862));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0__1842  (.H(net1863));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0__1843  (.H(net1864));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0__1844  (.H(net1865));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0__1845  (.H(net1866));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0__1846  (.H(net1867));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0__1847  (.H(net1868));
 TIEHIx1_ASAP7_75t_R \if_stage_i.instr_valid_id_o$_DFF_PN0__1848  (.H(net1869));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[0]$_DFFE_PN0P__1849  (.H(net1870));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[10]$_DFFE_PN0P__1850  (.H(net1871));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[11]$_DFFE_PN0P__1851  (.H(net1872));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[12]$_DFFE_PN0P__1852  (.H(net1873));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[13]$_DFFE_PN0P__1853  (.H(net1874));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[14]$_DFFE_PN0P__1854  (.H(net1875));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[15]$_DFFE_PN0P__1855  (.H(net1876));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[16]$_DFFE_PN0P__1856  (.H(net1877));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[17]$_DFFE_PN0P__1857  (.H(net1878));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[18]$_DFFE_PN0P__1858  (.H(net1879));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[19]$_DFFE_PN0P__1859  (.H(net1880));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[1]$_DFFE_PN0P__1860  (.H(net1881));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[20]$_DFFE_PN0P__1861  (.H(net1882));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[21]$_DFFE_PN0P__1862  (.H(net1883));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[22]$_DFFE_PN0P__1863  (.H(net1884));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[23]$_DFFE_PN0P__1864  (.H(net1885));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[24]$_DFFE_PN0P__1865  (.H(net1886));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[25]$_DFFE_PN0P__1866  (.H(net1887));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[26]$_DFFE_PN0P__1867  (.H(net1888));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[27]$_DFFE_PN0P__1868  (.H(net1889));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[28]$_DFFE_PN0P__1869  (.H(net1890));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[29]$_DFFE_PN0P__1870  (.H(net1891));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[2]$_DFFE_PN0P__1871  (.H(net1892));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[30]$_DFFE_PN0P__1872  (.H(net1893));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[31]$_DFFE_PN0P__1873  (.H(net1894));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[3]$_DFFE_PN0P__1874  (.H(net1895));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[4]$_DFFE_PN0P__1875  (.H(net1896));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[5]$_DFFE_PN0P__1876  (.H(net1897));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[6]$_DFFE_PN0P__1877  (.H(net1898));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[7]$_DFFE_PN0P__1878  (.H(net1899));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[8]$_DFFE_PN0P__1879  (.H(net1900));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_o[9]$_DFFE_PN0P__1880  (.H(net1901));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.data_sign_ext_q$_DFFE_PN0P__1881  (.H(net1902));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.data_we_q$_DFFE_PN0P__1882  (.H(net1903));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.handle_misaligned_q$_DFFE_PN0P__1883  (.H(net1904));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[0]$_DFFE_PN0P__1884  (.H(net1905));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[1]$_DFFE_PN0P__1885  (.H(net1906));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[2]$_DFFE_PN0P__1886  (.H(net1907));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.lsu_err_q$_DFFE_PN0P__1887  (.H(net1908));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_offset_q[0]$_DFFE_PN0P__1888  (.H(net1909));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_offset_q[1]$_DFFE_PN0P__1889  (.H(net1910));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[0]$_DFFE_PN0P__1890  (.H(net1911));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[10]$_DFFE_PN0P__1891  (.H(net1912));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[11]$_DFFE_PN0P__1892  (.H(net1913));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[12]$_DFFE_PN0P__1893  (.H(net1914));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[13]$_DFFE_PN0P__1894  (.H(net1915));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[14]$_DFFE_PN0P__1895  (.H(net1916));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[15]$_DFFE_PN0P__1896  (.H(net1917));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[16]$_DFFE_PN0P__1897  (.H(net1918));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[17]$_DFFE_PN0P__1898  (.H(net1919));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[18]$_DFFE_PN0P__1899  (.H(net1920));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[19]$_DFFE_PN0P__1900  (.H(net1921));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[1]$_DFFE_PN0P__1901  (.H(net1922));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[20]$_DFFE_PN0P__1902  (.H(net1923));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[21]$_DFFE_PN0P__1903  (.H(net1924));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[22]$_DFFE_PN0P__1904  (.H(net1925));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[23]$_DFFE_PN0P__1905  (.H(net1926));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[2]$_DFFE_PN0P__1906  (.H(net1927));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[3]$_DFFE_PN0P__1907  (.H(net1928));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[4]$_DFFE_PN0P__1908  (.H(net1929));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[5]$_DFFE_PN0P__1909  (.H(net1930));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[6]$_DFFE_PN0P__1910  (.H(net1931));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[7]$_DFFE_PN0P__1911  (.H(net1932));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[8]$_DFFE_PN0P__1912  (.H(net1933));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[9]$_DFFE_PN0P__1913  (.H(net1934));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk_i (.A(clk_i),
    .Y(clknet_0_clk_i));
 BUFx16f_ASAP7_75t_R clkbuf_1_0__f_clk_i (.A(clknet_0_clk_i),
    .Y(clknet_1_0__leaf_clk_i));
 BUFx24_ASAP7_75t_R clkbuf_leaf_0_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_0_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_1_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_1_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_2_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_2_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_3_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_3_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_4_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_4_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_5_clk_i_regs (.A(clknet_1_1__leaf_clk_i_regs),
    .Y(clknet_leaf_5_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_6_clk_i_regs (.A(clknet_1_1__leaf_clk_i_regs),
    .Y(clknet_leaf_6_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_7_clk_i_regs (.A(clknet_1_1__leaf_clk_i_regs),
    .Y(clknet_leaf_7_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_8_clk_i_regs (.A(clknet_1_1__leaf_clk_i_regs),
    .Y(clknet_leaf_8_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_9_clk_i_regs (.A(clknet_1_1__leaf_clk_i_regs),
    .Y(clknet_leaf_9_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_10_clk_i_regs (.A(clknet_1_1__leaf_clk_i_regs),
    .Y(clknet_leaf_10_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_11_clk_i_regs (.A(clknet_1_1__leaf_clk_i_regs),
    .Y(clknet_leaf_11_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_12_clk_i_regs (.A(clknet_1_1__leaf_clk_i_regs),
    .Y(clknet_leaf_12_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_13_clk_i_regs (.A(clknet_1_1__leaf_clk_i_regs),
    .Y(clknet_leaf_13_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_14_clk_i_regs (.A(clknet_1_1__leaf_clk_i_regs),
    .Y(clknet_leaf_14_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_15_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_15_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_16_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_16_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_17_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_17_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_18_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_18_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_19_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_19_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_20_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_20_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_21_clk_i_regs (.A(clknet_1_0__leaf_clk_i_regs),
    .Y(clknet_leaf_21_clk_i_regs));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk_i_regs (.A(clk_i_regs),
    .Y(clknet_0_clk_i_regs));
 BUFx16f_ASAP7_75t_R clkbuf_1_0__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Y(clknet_1_0__leaf_clk_i_regs));
 BUFx16f_ASAP7_75t_R clkbuf_1_1__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Y(clknet_1_1__leaf_clk_i_regs));
 INVx8_ASAP7_75t_R clkload0 (.A(clknet_1_1__leaf_clk_i_regs));
 CKINVDCx20_ASAP7_75t_R clkload1 (.A(clknet_leaf_15_clk_i_regs));
 CKINVDCx8_ASAP7_75t_R clkload2 (.A(clknet_leaf_16_clk_i_regs));
 INVx13_ASAP7_75t_R clkload3 (.A(clknet_leaf_21_clk_i_regs));
 CKINVDCx5p33_ASAP7_75t_R clkload4 (.A(clknet_leaf_5_clk_i_regs));
 CKINVDCx16_ASAP7_75t_R clkload5 (.A(clknet_leaf_6_clk_i_regs));
 INVxp67_ASAP7_75t_R clkload6 (.A(clknet_leaf_14_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_0_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_1_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_1_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_2_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_2_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_3_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_3_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_4_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_4_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_5_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_5_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_6_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_6_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_7_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_7_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_8_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_8_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_9_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_9_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_10_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_10_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_11_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_11_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_12_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_12_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_13_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_13_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_14_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_14_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_15_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_15_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_16_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_16_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_17_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_17_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_18_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_18_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_19_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_19_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_20_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_20_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_21_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_21_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_22_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_22_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_23_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_23_clk));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx16f_ASAP7_75t_R clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_1_0__leaf_clk));
 BUFx16f_ASAP7_75t_R clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_1_1__leaf_clk));
 INVx8_ASAP7_75t_R clkload7 (.A(clknet_1_0__leaf_clk));
 CKINVDCx16_ASAP7_75t_R clkload8 (.A(clknet_leaf_10_clk));
 INVxp33_ASAP7_75t_R clkload9 (.A(clknet_leaf_11_clk));
 INVxp33_ASAP7_75t_R clkload10 (.A(clknet_leaf_13_clk));
 BUFx12_ASAP7_75t_R clkload11 (.A(clknet_leaf_14_clk));
 INVxp33_ASAP7_75t_R clkload12 (.A(clknet_leaf_15_clk));
 INVxp67_ASAP7_75t_R clkload13 (.A(clknet_leaf_16_clk));
 INVx3_ASAP7_75t_R clkload14 (.A(clknet_leaf_17_clk));
 CKINVDCx14_ASAP7_75t_R clkload15 (.A(clknet_leaf_18_clk));
 CKINVDCx10_ASAP7_75t_R clkload16 (.A(clknet_leaf_19_clk));
 CKINVDCx20_ASAP7_75t_R clkload17 (.A(clknet_leaf_20_clk));
 CKINVDCx14_ASAP7_75t_R clkload18 (.A(clknet_leaf_0_clk));
 INVxp33_ASAP7_75t_R clkload19 (.A(clknet_leaf_2_clk));
 CKINVDCx16_ASAP7_75t_R clkload20 (.A(clknet_leaf_3_clk));
 CKINVDCx10_ASAP7_75t_R clkload21 (.A(clknet_leaf_4_clk));
 INVxp33_ASAP7_75t_R clkload22 (.A(clknet_leaf_5_clk));
 INVxp33_ASAP7_75t_R clkload23 (.A(clknet_leaf_6_clk));
 INVxp33_ASAP7_75t_R clkload24 (.A(clknet_leaf_7_clk));
 INVxp33_ASAP7_75t_R clkload25 (.A(clknet_leaf_8_clk));
 CKINVDCx11_ASAP7_75t_R clkload26 (.A(clknet_leaf_9_clk));
 CKINVDCx20_ASAP7_75t_R clkload27 (.A(clknet_leaf_21_clk));
 CKINVDCx20_ASAP7_75t_R clkload28 (.A(clknet_leaf_22_clk));
 CKINVDCx16_ASAP7_75t_R clkload29 (.A(clknet_leaf_23_clk));
 BUFx16f_ASAP7_75t_R delaybuf_0_core_clock (.A(delaynet_0_core_clock),
    .Y(delaynet_1_core_clock));
 BUFx16f_ASAP7_75t_R delaybuf_1_core_clock (.A(delaynet_1_core_clock),
    .Y(delaynet_2_core_clock));
 BUFx16f_ASAP7_75t_R delaybuf_2_core_clock (.A(delaynet_2_core_clock),
    .Y(clk_i_regs));
 BUFx3_ASAP7_75t_R rebuffer1 (.A(_00845_),
    .Y(net1935));
 BUFx3_ASAP7_75t_R rebuffer2 (.A(net1935),
    .Y(net1936));
 BUFx3_ASAP7_75t_R rebuffer3 (.A(_00813_),
    .Y(net1937));
 BUFx3_ASAP7_75t_R rebuffer4 (.A(_00781_),
    .Y(net1938));
 BUFx3_ASAP7_75t_R rebuffer5 (.A(net1938),
    .Y(net1939));
 BUFx3_ASAP7_75t_R rebuffer6 (.A(_00941_),
    .Y(net1940));
 BUFx3_ASAP7_75t_R rebuffer7 (.A(_00877_),
    .Y(net1941));
 BUFx3_ASAP7_75t_R rebuffer8 (.A(_00777_),
    .Y(net1942));
 BUFx3_ASAP7_75t_R rebuffer9 (.A(net1942),
    .Y(net1943));
 BUFx3_ASAP7_75t_R rebuffer10 (.A(_00779_),
    .Y(net1944));
 BUFx3_ASAP7_75t_R rebuffer11 (.A(net1944),
    .Y(net1945));
 BUFx3_ASAP7_75t_R rebuffer12 (.A(_15646_),
    .Y(net1946));
 BUFx3_ASAP7_75t_R rebuffer13 (.A(_15646_),
    .Y(net1947));
 BUFx3_ASAP7_75t_R rebuffer14 (.A(_00773_),
    .Y(net1948));
 BUFx3_ASAP7_75t_R rebuffer15 (.A(net1948),
    .Y(net1949));
 BUFx3_ASAP7_75t_R rebuffer16 (.A(_00775_),
    .Y(net1950));
 BUFx3_ASAP7_75t_R rebuffer17 (.A(_01005_),
    .Y(net1951));
 BUFx3_ASAP7_75t_R rebuffer18 (.A(_04971_),
    .Y(net1952));
 BUFx3_ASAP7_75t_R rebuffer19 (.A(_14619_),
    .Y(net1953));
 BUFx3_ASAP7_75t_R rebuffer20 (.A(_16502_),
    .Y(net1954));
 BUFx3_ASAP7_75t_R rebuffer21 (.A(_00814_),
    .Y(net1955));
 BUFx3_ASAP7_75t_R rebuffer22 (.A(_16006_),
    .Y(net1956));
 BUFx3_ASAP7_75t_R rebuffer23 (.A(_15261_),
    .Y(net1957));
 BUFx3_ASAP7_75t_R rebuffer24 (.A(net1968),
    .Y(net1958));
 BUFx3_ASAP7_75t_R rebuffer25 (.A(net1976),
    .Y(net1959));
 BUFx3_ASAP7_75t_R rebuffer26 (.A(\alu_adder_result_ex[31] ),
    .Y(net1960));
 BUFx3_ASAP7_75t_R rebuffer27 (.A(\alu_adder_result_ex[31] ),
    .Y(net1961));
 BUFx3_ASAP7_75t_R rebuffer28 (.A(_17737_),
    .Y(net1962));
 BUFx16f_ASAP7_75t_R load_slew1 (.A(net169),
    .Y(net1963));
 BUFx3_ASAP7_75t_R rebuffer29 (.A(_11694_),
    .Y(net1964));
 BUFx3_ASAP7_75t_R rebuffer30 (.A(_16131_),
    .Y(net1965));
 BUFx3_ASAP7_75t_R rebuffer31 (.A(_16131_),
    .Y(net1966));
 BUFx3_ASAP7_75t_R rebuffer32 (.A(_00185_),
    .Y(net1967));
 BUFx4_ASAP7_75t_R clone33 (.A(_15258_),
    .Y(net1968));
 BUFx3_ASAP7_75t_R rebuffer34 (.A(_15299_),
    .Y(net1969));
 BUFx3_ASAP7_75t_R rebuffer35 (.A(_15502_),
    .Y(net1970));
 BUFx4_ASAP7_75t_R clone36 (.A(_15258_),
    .Y(net1971));
 BUFx6f_ASAP7_75t_R rebuffer37 (.A(_15256_),
    .Y(net1972));
 BUFx3_ASAP7_75t_R rebuffer38 (.A(_15256_),
    .Y(net1973));
 BUFx3_ASAP7_75t_R rebuffer39 (.A(_02221_),
    .Y(net1974));
 BUFx3_ASAP7_75t_R rebuffer41 (.A(_01517_),
    .Y(net1976));
 BUFx3_ASAP7_75t_R rebuffer42 (.A(_13362_),
    .Y(net1977));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_662 ();
 DECAPx2_ASAP7_75t_R FILLER_0_684 ();
 FILLER_ASAP7_75t_R FILLER_0_690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886 ();
 DECAPx6_ASAP7_75t_R FILLER_0_908 ();
 FILLER_ASAP7_75t_R FILLER_0_922 ();
 DECAPx10_ASAP7_75t_R FILLER_0_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1004 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1095 ();
 FILLER_ASAP7_75t_R FILLER_0_1102 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1174 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_1_112 ();
 DECAPx10_ASAP7_75t_R FILLER_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_1_156 ();
 DECAPx10_ASAP7_75t_R FILLER_1_178 ();
 DECAPx10_ASAP7_75t_R FILLER_1_200 ();
 DECAPx10_ASAP7_75t_R FILLER_1_222 ();
 DECAPx10_ASAP7_75t_R FILLER_1_244 ();
 DECAPx10_ASAP7_75t_R FILLER_1_266 ();
 DECAPx10_ASAP7_75t_R FILLER_1_288 ();
 DECAPx10_ASAP7_75t_R FILLER_1_310 ();
 DECAPx10_ASAP7_75t_R FILLER_1_332 ();
 DECAPx10_ASAP7_75t_R FILLER_1_354 ();
 DECAPx10_ASAP7_75t_R FILLER_1_376 ();
 DECAPx10_ASAP7_75t_R FILLER_1_398 ();
 DECAPx10_ASAP7_75t_R FILLER_1_420 ();
 DECAPx10_ASAP7_75t_R FILLER_1_442 ();
 DECAPx10_ASAP7_75t_R FILLER_1_464 ();
 DECAPx10_ASAP7_75t_R FILLER_1_486 ();
 DECAPx10_ASAP7_75t_R FILLER_1_508 ();
 DECAPx10_ASAP7_75t_R FILLER_1_530 ();
 DECAPx10_ASAP7_75t_R FILLER_1_552 ();
 DECAPx10_ASAP7_75t_R FILLER_1_574 ();
 DECAPx10_ASAP7_75t_R FILLER_1_596 ();
 DECAPx10_ASAP7_75t_R FILLER_1_618 ();
 DECAPx10_ASAP7_75t_R FILLER_1_640 ();
 DECAPx10_ASAP7_75t_R FILLER_1_662 ();
 DECAPx4_ASAP7_75t_R FILLER_1_684 ();
 DECAPx6_ASAP7_75t_R FILLER_1_706 ();
 FILLER_ASAP7_75t_R FILLER_1_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_722 ();
 DECAPx2_ASAP7_75t_R FILLER_1_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_743 ();
 DECAPx10_ASAP7_75t_R FILLER_1_747 ();
 DECAPx4_ASAP7_75t_R FILLER_1_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_802 ();
 DECAPx10_ASAP7_75t_R FILLER_1_820 ();
 DECAPx10_ASAP7_75t_R FILLER_1_842 ();
 DECAPx10_ASAP7_75t_R FILLER_1_864 ();
 DECAPx10_ASAP7_75t_R FILLER_1_886 ();
 DECAPx6_ASAP7_75t_R FILLER_1_908 ();
 FILLER_ASAP7_75t_R FILLER_1_922 ();
 DECAPx10_ASAP7_75t_R FILLER_1_926 ();
 DECAPx10_ASAP7_75t_R FILLER_1_948 ();
 DECAPx2_ASAP7_75t_R FILLER_1_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_976 ();
 DECAPx10_ASAP7_75t_R FILLER_1_983 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_1_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1070 ();
 DECAPx4_ASAP7_75t_R FILLER_1_1092 ();
 FILLER_ASAP7_75t_R FILLER_1_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_1_1111 ();
 FILLER_ASAP7_75t_R FILLER_1_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_1_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_1_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_1_1182 ();
 FILLER_ASAP7_75t_R FILLER_1_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1358 ();
 DECAPx4_ASAP7_75t_R FILLER_1_1380 ();
 FILLER_ASAP7_75t_R FILLER_1_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_2_112 ();
 DECAPx10_ASAP7_75t_R FILLER_2_134 ();
 DECAPx10_ASAP7_75t_R FILLER_2_156 ();
 DECAPx10_ASAP7_75t_R FILLER_2_178 ();
 DECAPx10_ASAP7_75t_R FILLER_2_200 ();
 DECAPx10_ASAP7_75t_R FILLER_2_222 ();
 DECAPx10_ASAP7_75t_R FILLER_2_244 ();
 DECAPx10_ASAP7_75t_R FILLER_2_266 ();
 DECAPx10_ASAP7_75t_R FILLER_2_288 ();
 DECAPx10_ASAP7_75t_R FILLER_2_310 ();
 DECAPx10_ASAP7_75t_R FILLER_2_332 ();
 DECAPx10_ASAP7_75t_R FILLER_2_354 ();
 DECAPx10_ASAP7_75t_R FILLER_2_376 ();
 DECAPx10_ASAP7_75t_R FILLER_2_398 ();
 DECAPx10_ASAP7_75t_R FILLER_2_420 ();
 DECAPx6_ASAP7_75t_R FILLER_2_442 ();
 DECAPx2_ASAP7_75t_R FILLER_2_456 ();
 DECAPx10_ASAP7_75t_R FILLER_2_464 ();
 DECAPx10_ASAP7_75t_R FILLER_2_486 ();
 DECAPx10_ASAP7_75t_R FILLER_2_508 ();
 DECAPx10_ASAP7_75t_R FILLER_2_530 ();
 DECAPx10_ASAP7_75t_R FILLER_2_552 ();
 DECAPx10_ASAP7_75t_R FILLER_2_574 ();
 DECAPx10_ASAP7_75t_R FILLER_2_596 ();
 DECAPx10_ASAP7_75t_R FILLER_2_618 ();
 DECAPx10_ASAP7_75t_R FILLER_2_640 ();
 DECAPx10_ASAP7_75t_R FILLER_2_662 ();
 DECAPx10_ASAP7_75t_R FILLER_2_684 ();
 DECAPx4_ASAP7_75t_R FILLER_2_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_729 ();
 DECAPx6_ASAP7_75t_R FILLER_2_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_779 ();
 FILLER_ASAP7_75t_R FILLER_2_800 ();
 DECAPx4_ASAP7_75t_R FILLER_2_822 ();
 FILLER_ASAP7_75t_R FILLER_2_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_834 ();
 DECAPx10_ASAP7_75t_R FILLER_2_841 ();
 DECAPx10_ASAP7_75t_R FILLER_2_863 ();
 DECAPx10_ASAP7_75t_R FILLER_2_885 ();
 DECAPx10_ASAP7_75t_R FILLER_2_907 ();
 DECAPx10_ASAP7_75t_R FILLER_2_929 ();
 DECAPx10_ASAP7_75t_R FILLER_2_951 ();
 DECAPx10_ASAP7_75t_R FILLER_2_973 ();
 DECAPx10_ASAP7_75t_R FILLER_2_995 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_2_1039 ();
 FILLER_ASAP7_75t_R FILLER_2_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1350 ();
 DECAPx6_ASAP7_75t_R FILLER_2_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_2_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_3_112 ();
 DECAPx10_ASAP7_75t_R FILLER_3_134 ();
 DECAPx10_ASAP7_75t_R FILLER_3_156 ();
 DECAPx10_ASAP7_75t_R FILLER_3_178 ();
 DECAPx10_ASAP7_75t_R FILLER_3_200 ();
 DECAPx10_ASAP7_75t_R FILLER_3_222 ();
 DECAPx10_ASAP7_75t_R FILLER_3_244 ();
 DECAPx10_ASAP7_75t_R FILLER_3_266 ();
 DECAPx10_ASAP7_75t_R FILLER_3_288 ();
 DECAPx10_ASAP7_75t_R FILLER_3_310 ();
 DECAPx10_ASAP7_75t_R FILLER_3_332 ();
 DECAPx10_ASAP7_75t_R FILLER_3_354 ();
 DECAPx10_ASAP7_75t_R FILLER_3_376 ();
 DECAPx10_ASAP7_75t_R FILLER_3_398 ();
 DECAPx10_ASAP7_75t_R FILLER_3_420 ();
 DECAPx10_ASAP7_75t_R FILLER_3_442 ();
 DECAPx10_ASAP7_75t_R FILLER_3_464 ();
 DECAPx10_ASAP7_75t_R FILLER_3_486 ();
 DECAPx10_ASAP7_75t_R FILLER_3_508 ();
 DECAPx10_ASAP7_75t_R FILLER_3_530 ();
 DECAPx10_ASAP7_75t_R FILLER_3_552 ();
 DECAPx10_ASAP7_75t_R FILLER_3_574 ();
 DECAPx10_ASAP7_75t_R FILLER_3_596 ();
 DECAPx10_ASAP7_75t_R FILLER_3_618 ();
 DECAPx10_ASAP7_75t_R FILLER_3_640 ();
 DECAPx10_ASAP7_75t_R FILLER_3_662 ();
 DECAPx10_ASAP7_75t_R FILLER_3_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_706 ();
 DECAPx4_ASAP7_75t_R FILLER_3_742 ();
 FILLER_ASAP7_75t_R FILLER_3_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_758 ();
 FILLER_ASAP7_75t_R FILLER_3_774 ();
 DECAPx1_ASAP7_75t_R FILLER_3_805 ();
 FILLER_ASAP7_75t_R FILLER_3_840 ();
 DECAPx10_ASAP7_75t_R FILLER_3_862 ();
 DECAPx10_ASAP7_75t_R FILLER_3_884 ();
 DECAPx6_ASAP7_75t_R FILLER_3_906 ();
 DECAPx1_ASAP7_75t_R FILLER_3_920 ();
 DECAPx10_ASAP7_75t_R FILLER_3_926 ();
 DECAPx10_ASAP7_75t_R FILLER_3_948 ();
 DECAPx10_ASAP7_75t_R FILLER_3_970 ();
 DECAPx10_ASAP7_75t_R FILLER_3_992 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_3_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_4_112 ();
 DECAPx10_ASAP7_75t_R FILLER_4_134 ();
 DECAPx10_ASAP7_75t_R FILLER_4_156 ();
 DECAPx10_ASAP7_75t_R FILLER_4_178 ();
 DECAPx10_ASAP7_75t_R FILLER_4_200 ();
 DECAPx10_ASAP7_75t_R FILLER_4_222 ();
 DECAPx10_ASAP7_75t_R FILLER_4_244 ();
 DECAPx10_ASAP7_75t_R FILLER_4_266 ();
 DECAPx10_ASAP7_75t_R FILLER_4_288 ();
 DECAPx10_ASAP7_75t_R FILLER_4_310 ();
 DECAPx10_ASAP7_75t_R FILLER_4_332 ();
 DECAPx10_ASAP7_75t_R FILLER_4_354 ();
 DECAPx10_ASAP7_75t_R FILLER_4_376 ();
 DECAPx10_ASAP7_75t_R FILLER_4_398 ();
 DECAPx10_ASAP7_75t_R FILLER_4_420 ();
 DECAPx6_ASAP7_75t_R FILLER_4_442 ();
 DECAPx2_ASAP7_75t_R FILLER_4_456 ();
 DECAPx10_ASAP7_75t_R FILLER_4_464 ();
 DECAPx10_ASAP7_75t_R FILLER_4_486 ();
 DECAPx10_ASAP7_75t_R FILLER_4_508 ();
 DECAPx10_ASAP7_75t_R FILLER_4_530 ();
 DECAPx10_ASAP7_75t_R FILLER_4_552 ();
 DECAPx10_ASAP7_75t_R FILLER_4_574 ();
 DECAPx10_ASAP7_75t_R FILLER_4_596 ();
 DECAPx10_ASAP7_75t_R FILLER_4_618 ();
 DECAPx10_ASAP7_75t_R FILLER_4_640 ();
 DECAPx10_ASAP7_75t_R FILLER_4_662 ();
 DECAPx1_ASAP7_75t_R FILLER_4_684 ();
 FILLER_ASAP7_75t_R FILLER_4_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_724 ();
 DECAPx2_ASAP7_75t_R FILLER_4_731 ();
 FILLER_ASAP7_75t_R FILLER_4_754 ();
 DECAPx1_ASAP7_75t_R FILLER_4_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_774 ();
 DECAPx4_ASAP7_75t_R FILLER_4_792 ();
 FILLER_ASAP7_75t_R FILLER_4_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_822 ();
 DECAPx1_ASAP7_75t_R FILLER_4_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_850 ();
 DECAPx10_ASAP7_75t_R FILLER_4_874 ();
 DECAPx10_ASAP7_75t_R FILLER_4_896 ();
 DECAPx10_ASAP7_75t_R FILLER_4_918 ();
 DECAPx10_ASAP7_75t_R FILLER_4_940 ();
 DECAPx10_ASAP7_75t_R FILLER_4_962 ();
 DECAPx10_ASAP7_75t_R FILLER_4_984 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_4_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_4_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_5_68 ();
 DECAPx10_ASAP7_75t_R FILLER_5_90 ();
 DECAPx10_ASAP7_75t_R FILLER_5_112 ();
 DECAPx10_ASAP7_75t_R FILLER_5_134 ();
 DECAPx10_ASAP7_75t_R FILLER_5_156 ();
 DECAPx10_ASAP7_75t_R FILLER_5_178 ();
 DECAPx10_ASAP7_75t_R FILLER_5_200 ();
 DECAPx10_ASAP7_75t_R FILLER_5_222 ();
 DECAPx10_ASAP7_75t_R FILLER_5_244 ();
 DECAPx10_ASAP7_75t_R FILLER_5_266 ();
 DECAPx10_ASAP7_75t_R FILLER_5_288 ();
 DECAPx10_ASAP7_75t_R FILLER_5_310 ();
 DECAPx10_ASAP7_75t_R FILLER_5_332 ();
 DECAPx10_ASAP7_75t_R FILLER_5_354 ();
 DECAPx10_ASAP7_75t_R FILLER_5_376 ();
 DECAPx10_ASAP7_75t_R FILLER_5_398 ();
 DECAPx10_ASAP7_75t_R FILLER_5_420 ();
 DECAPx10_ASAP7_75t_R FILLER_5_442 ();
 DECAPx10_ASAP7_75t_R FILLER_5_464 ();
 DECAPx10_ASAP7_75t_R FILLER_5_486 ();
 DECAPx10_ASAP7_75t_R FILLER_5_508 ();
 DECAPx10_ASAP7_75t_R FILLER_5_530 ();
 DECAPx10_ASAP7_75t_R FILLER_5_552 ();
 DECAPx10_ASAP7_75t_R FILLER_5_574 ();
 DECAPx10_ASAP7_75t_R FILLER_5_596 ();
 DECAPx10_ASAP7_75t_R FILLER_5_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_640 ();
 DECAPx2_ASAP7_75t_R FILLER_5_651 ();
 DECAPx6_ASAP7_75t_R FILLER_5_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_707 ();
 DECAPx10_ASAP7_75t_R FILLER_5_728 ();
 DECAPx2_ASAP7_75t_R FILLER_5_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_756 ();
 DECAPx6_ASAP7_75t_R FILLER_5_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_792 ();
 DECAPx6_ASAP7_75t_R FILLER_5_796 ();
 FILLER_ASAP7_75t_R FILLER_5_827 ();
 FILLER_ASAP7_75t_R FILLER_5_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_849 ();
 FILLER_ASAP7_75t_R FILLER_5_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_855 ();
 DECAPx10_ASAP7_75t_R FILLER_5_873 ();
 DECAPx10_ASAP7_75t_R FILLER_5_895 ();
 DECAPx2_ASAP7_75t_R FILLER_5_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_923 ();
 DECAPx10_ASAP7_75t_R FILLER_5_926 ();
 DECAPx10_ASAP7_75t_R FILLER_5_948 ();
 DECAPx10_ASAP7_75t_R FILLER_5_970 ();
 DECAPx10_ASAP7_75t_R FILLER_5_992 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_5_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_6_68 ();
 DECAPx10_ASAP7_75t_R FILLER_6_90 ();
 DECAPx10_ASAP7_75t_R FILLER_6_112 ();
 DECAPx10_ASAP7_75t_R FILLER_6_134 ();
 DECAPx10_ASAP7_75t_R FILLER_6_156 ();
 DECAPx10_ASAP7_75t_R FILLER_6_178 ();
 DECAPx10_ASAP7_75t_R FILLER_6_200 ();
 DECAPx10_ASAP7_75t_R FILLER_6_222 ();
 DECAPx10_ASAP7_75t_R FILLER_6_244 ();
 DECAPx10_ASAP7_75t_R FILLER_6_266 ();
 DECAPx10_ASAP7_75t_R FILLER_6_288 ();
 DECAPx10_ASAP7_75t_R FILLER_6_310 ();
 DECAPx10_ASAP7_75t_R FILLER_6_332 ();
 DECAPx10_ASAP7_75t_R FILLER_6_354 ();
 DECAPx10_ASAP7_75t_R FILLER_6_376 ();
 DECAPx10_ASAP7_75t_R FILLER_6_398 ();
 DECAPx10_ASAP7_75t_R FILLER_6_420 ();
 DECAPx6_ASAP7_75t_R FILLER_6_442 ();
 DECAPx2_ASAP7_75t_R FILLER_6_456 ();
 DECAPx10_ASAP7_75t_R FILLER_6_464 ();
 DECAPx10_ASAP7_75t_R FILLER_6_486 ();
 DECAPx10_ASAP7_75t_R FILLER_6_508 ();
 DECAPx10_ASAP7_75t_R FILLER_6_530 ();
 DECAPx10_ASAP7_75t_R FILLER_6_552 ();
 DECAPx10_ASAP7_75t_R FILLER_6_574 ();
 DECAPx10_ASAP7_75t_R FILLER_6_596 ();
 DECAPx6_ASAP7_75t_R FILLER_6_618 ();
 DECAPx2_ASAP7_75t_R FILLER_6_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_657 ();
 DECAPx2_ASAP7_75t_R FILLER_6_667 ();
 FILLER_ASAP7_75t_R FILLER_6_673 ();
 DECAPx1_ASAP7_75t_R FILLER_6_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_697 ();
 DECAPx2_ASAP7_75t_R FILLER_6_708 ();
 FILLER_ASAP7_75t_R FILLER_6_714 ();
 FILLER_ASAP7_75t_R FILLER_6_722 ();
 DECAPx2_ASAP7_75t_R FILLER_6_727 ();
 FILLER_ASAP7_75t_R FILLER_6_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_735 ();
 DECAPx1_ASAP7_75t_R FILLER_6_742 ();
 DECAPx10_ASAP7_75t_R FILLER_6_749 ();
 DECAPx6_ASAP7_75t_R FILLER_6_771 ();
 DECAPx2_ASAP7_75t_R FILLER_6_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_791 ();
 FILLER_ASAP7_75t_R FILLER_6_806 ();
 FILLER_ASAP7_75t_R FILLER_6_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_813 ();
 DECAPx6_ASAP7_75t_R FILLER_6_817 ();
 FILLER_ASAP7_75t_R FILLER_6_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_833 ();
 FILLER_ASAP7_75t_R FILLER_6_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_842 ();
 DECAPx6_ASAP7_75t_R FILLER_6_846 ();
 DECAPx10_ASAP7_75t_R FILLER_6_869 ();
 DECAPx10_ASAP7_75t_R FILLER_6_891 ();
 DECAPx10_ASAP7_75t_R FILLER_6_913 ();
 DECAPx10_ASAP7_75t_R FILLER_6_935 ();
 DECAPx10_ASAP7_75t_R FILLER_6_957 ();
 DECAPx10_ASAP7_75t_R FILLER_6_979 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1353 ();
 DECAPx4_ASAP7_75t_R FILLER_6_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_6_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_7_90 ();
 DECAPx10_ASAP7_75t_R FILLER_7_112 ();
 DECAPx10_ASAP7_75t_R FILLER_7_134 ();
 DECAPx10_ASAP7_75t_R FILLER_7_156 ();
 DECAPx10_ASAP7_75t_R FILLER_7_178 ();
 DECAPx10_ASAP7_75t_R FILLER_7_200 ();
 DECAPx10_ASAP7_75t_R FILLER_7_222 ();
 DECAPx10_ASAP7_75t_R FILLER_7_244 ();
 DECAPx10_ASAP7_75t_R FILLER_7_266 ();
 DECAPx10_ASAP7_75t_R FILLER_7_288 ();
 DECAPx10_ASAP7_75t_R FILLER_7_310 ();
 DECAPx10_ASAP7_75t_R FILLER_7_332 ();
 DECAPx10_ASAP7_75t_R FILLER_7_354 ();
 DECAPx10_ASAP7_75t_R FILLER_7_376 ();
 DECAPx10_ASAP7_75t_R FILLER_7_398 ();
 DECAPx10_ASAP7_75t_R FILLER_7_420 ();
 DECAPx10_ASAP7_75t_R FILLER_7_442 ();
 DECAPx10_ASAP7_75t_R FILLER_7_464 ();
 DECAPx10_ASAP7_75t_R FILLER_7_486 ();
 DECAPx10_ASAP7_75t_R FILLER_7_508 ();
 DECAPx10_ASAP7_75t_R FILLER_7_530 ();
 DECAPx10_ASAP7_75t_R FILLER_7_552 ();
 DECAPx10_ASAP7_75t_R FILLER_7_574 ();
 DECAPx10_ASAP7_75t_R FILLER_7_596 ();
 DECAPx6_ASAP7_75t_R FILLER_7_618 ();
 DECAPx2_ASAP7_75t_R FILLER_7_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_638 ();
 FILLER_ASAP7_75t_R FILLER_7_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_651 ();
 DECAPx4_ASAP7_75t_R FILLER_7_658 ();
 DECAPx2_ASAP7_75t_R FILLER_7_671 ();
 FILLER_ASAP7_75t_R FILLER_7_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_693 ();
 DECAPx10_ASAP7_75t_R FILLER_7_712 ();
 FILLER_ASAP7_75t_R FILLER_7_748 ();
 DECAPx1_ASAP7_75t_R FILLER_7_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_771 ();
 DECAPx2_ASAP7_75t_R FILLER_7_800 ();
 DECAPx2_ASAP7_75t_R FILLER_7_826 ();
 DECAPx4_ASAP7_75t_R FILLER_7_842 ();
 DECAPx10_ASAP7_75t_R FILLER_7_866 ();
 DECAPx10_ASAP7_75t_R FILLER_7_888 ();
 DECAPx6_ASAP7_75t_R FILLER_7_910 ();
 DECAPx10_ASAP7_75t_R FILLER_7_926 ();
 DECAPx10_ASAP7_75t_R FILLER_7_948 ();
 DECAPx10_ASAP7_75t_R FILLER_7_970 ();
 DECAPx10_ASAP7_75t_R FILLER_7_992 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_7_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_8_112 ();
 DECAPx10_ASAP7_75t_R FILLER_8_134 ();
 DECAPx10_ASAP7_75t_R FILLER_8_156 ();
 DECAPx10_ASAP7_75t_R FILLER_8_178 ();
 DECAPx10_ASAP7_75t_R FILLER_8_200 ();
 DECAPx10_ASAP7_75t_R FILLER_8_222 ();
 DECAPx10_ASAP7_75t_R FILLER_8_244 ();
 DECAPx10_ASAP7_75t_R FILLER_8_266 ();
 DECAPx10_ASAP7_75t_R FILLER_8_288 ();
 DECAPx10_ASAP7_75t_R FILLER_8_310 ();
 DECAPx10_ASAP7_75t_R FILLER_8_332 ();
 DECAPx10_ASAP7_75t_R FILLER_8_354 ();
 DECAPx10_ASAP7_75t_R FILLER_8_376 ();
 DECAPx10_ASAP7_75t_R FILLER_8_398 ();
 DECAPx10_ASAP7_75t_R FILLER_8_420 ();
 DECAPx6_ASAP7_75t_R FILLER_8_442 ();
 DECAPx2_ASAP7_75t_R FILLER_8_456 ();
 DECAPx10_ASAP7_75t_R FILLER_8_464 ();
 DECAPx10_ASAP7_75t_R FILLER_8_486 ();
 DECAPx10_ASAP7_75t_R FILLER_8_508 ();
 DECAPx10_ASAP7_75t_R FILLER_8_530 ();
 DECAPx10_ASAP7_75t_R FILLER_8_552 ();
 DECAPx10_ASAP7_75t_R FILLER_8_574 ();
 FILLER_ASAP7_75t_R FILLER_8_596 ();
 DECAPx1_ASAP7_75t_R FILLER_8_616 ();
 DECAPx2_ASAP7_75t_R FILLER_8_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_644 ();
 DECAPx2_ASAP7_75t_R FILLER_8_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_657 ();
 DECAPx2_ASAP7_75t_R FILLER_8_664 ();
 FILLER_ASAP7_75t_R FILLER_8_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_672 ();
 FILLER_ASAP7_75t_R FILLER_8_679 ();
 DECAPx2_ASAP7_75t_R FILLER_8_684 ();
 FILLER_ASAP7_75t_R FILLER_8_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_695 ();
 DECAPx6_ASAP7_75t_R FILLER_8_713 ();
 DECAPx1_ASAP7_75t_R FILLER_8_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_731 ();
 DECAPx1_ASAP7_75t_R FILLER_8_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_788 ();
 FILLER_ASAP7_75t_R FILLER_8_799 ();
 DECAPx2_ASAP7_75t_R FILLER_8_821 ();
 DECAPx1_ASAP7_75t_R FILLER_8_847 ();
 DECAPx2_ASAP7_75t_R FILLER_8_857 ();
 FILLER_ASAP7_75t_R FILLER_8_863 ();
 DECAPx10_ASAP7_75t_R FILLER_8_868 ();
 DECAPx10_ASAP7_75t_R FILLER_8_890 ();
 DECAPx10_ASAP7_75t_R FILLER_8_912 ();
 DECAPx10_ASAP7_75t_R FILLER_8_934 ();
 DECAPx10_ASAP7_75t_R FILLER_8_956 ();
 DECAPx10_ASAP7_75t_R FILLER_8_978 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1022 ();
 DECAPx6_ASAP7_75t_R FILLER_8_1044 ();
 DECAPx1_ASAP7_75t_R FILLER_8_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1353 ();
 DECAPx4_ASAP7_75t_R FILLER_8_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_8_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_9_68 ();
 DECAPx10_ASAP7_75t_R FILLER_9_90 ();
 DECAPx10_ASAP7_75t_R FILLER_9_112 ();
 DECAPx10_ASAP7_75t_R FILLER_9_134 ();
 DECAPx10_ASAP7_75t_R FILLER_9_156 ();
 DECAPx10_ASAP7_75t_R FILLER_9_178 ();
 DECAPx10_ASAP7_75t_R FILLER_9_200 ();
 DECAPx10_ASAP7_75t_R FILLER_9_222 ();
 DECAPx10_ASAP7_75t_R FILLER_9_244 ();
 DECAPx10_ASAP7_75t_R FILLER_9_266 ();
 DECAPx10_ASAP7_75t_R FILLER_9_288 ();
 DECAPx10_ASAP7_75t_R FILLER_9_310 ();
 DECAPx10_ASAP7_75t_R FILLER_9_332 ();
 DECAPx10_ASAP7_75t_R FILLER_9_354 ();
 DECAPx10_ASAP7_75t_R FILLER_9_376 ();
 DECAPx10_ASAP7_75t_R FILLER_9_398 ();
 DECAPx10_ASAP7_75t_R FILLER_9_420 ();
 DECAPx10_ASAP7_75t_R FILLER_9_442 ();
 DECAPx10_ASAP7_75t_R FILLER_9_464 ();
 DECAPx10_ASAP7_75t_R FILLER_9_486 ();
 DECAPx10_ASAP7_75t_R FILLER_9_508 ();
 DECAPx10_ASAP7_75t_R FILLER_9_530 ();
 DECAPx10_ASAP7_75t_R FILLER_9_552 ();
 DECAPx10_ASAP7_75t_R FILLER_9_574 ();
 DECAPx10_ASAP7_75t_R FILLER_9_596 ();
 DECAPx1_ASAP7_75t_R FILLER_9_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_622 ();
 DECAPx2_ASAP7_75t_R FILLER_9_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_647 ();
 DECAPx6_ASAP7_75t_R FILLER_9_680 ();
 DECAPx1_ASAP7_75t_R FILLER_9_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_698 ();
 DECAPx2_ASAP7_75t_R FILLER_9_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_711 ();
 DECAPx6_ASAP7_75t_R FILLER_9_730 ();
 DECAPx1_ASAP7_75t_R FILLER_9_744 ();
 DECAPx2_ASAP7_75t_R FILLER_9_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_770 ();
 DECAPx2_ASAP7_75t_R FILLER_9_774 ();
 DECAPx1_ASAP7_75t_R FILLER_9_783 ();
 FILLER_ASAP7_75t_R FILLER_9_796 ();
 DECAPx2_ASAP7_75t_R FILLER_9_801 ();
 DECAPx6_ASAP7_75t_R FILLER_9_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_831 ();
 FILLER_ASAP7_75t_R FILLER_9_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_854 ();
 FILLER_ASAP7_75t_R FILLER_9_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_860 ();
 DECAPx10_ASAP7_75t_R FILLER_9_870 ();
 DECAPx10_ASAP7_75t_R FILLER_9_892 ();
 DECAPx4_ASAP7_75t_R FILLER_9_914 ();
 DECAPx10_ASAP7_75t_R FILLER_9_926 ();
 DECAPx10_ASAP7_75t_R FILLER_9_948 ();
 DECAPx10_ASAP7_75t_R FILLER_9_970 ();
 DECAPx10_ASAP7_75t_R FILLER_9_992 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_9_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_9_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1358 ();
 DECAPx4_ASAP7_75t_R FILLER_9_1380 ();
 FILLER_ASAP7_75t_R FILLER_9_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_10_112 ();
 DECAPx10_ASAP7_75t_R FILLER_10_134 ();
 DECAPx10_ASAP7_75t_R FILLER_10_156 ();
 DECAPx10_ASAP7_75t_R FILLER_10_178 ();
 DECAPx10_ASAP7_75t_R FILLER_10_200 ();
 DECAPx10_ASAP7_75t_R FILLER_10_222 ();
 DECAPx10_ASAP7_75t_R FILLER_10_244 ();
 DECAPx10_ASAP7_75t_R FILLER_10_266 ();
 DECAPx10_ASAP7_75t_R FILLER_10_288 ();
 DECAPx10_ASAP7_75t_R FILLER_10_310 ();
 DECAPx10_ASAP7_75t_R FILLER_10_332 ();
 DECAPx10_ASAP7_75t_R FILLER_10_354 ();
 DECAPx10_ASAP7_75t_R FILLER_10_376 ();
 DECAPx10_ASAP7_75t_R FILLER_10_398 ();
 DECAPx10_ASAP7_75t_R FILLER_10_420 ();
 DECAPx6_ASAP7_75t_R FILLER_10_442 ();
 DECAPx2_ASAP7_75t_R FILLER_10_456 ();
 DECAPx10_ASAP7_75t_R FILLER_10_464 ();
 DECAPx10_ASAP7_75t_R FILLER_10_486 ();
 DECAPx10_ASAP7_75t_R FILLER_10_508 ();
 DECAPx10_ASAP7_75t_R FILLER_10_530 ();
 DECAPx10_ASAP7_75t_R FILLER_10_552 ();
 DECAPx10_ASAP7_75t_R FILLER_10_574 ();
 DECAPx10_ASAP7_75t_R FILLER_10_596 ();
 DECAPx1_ASAP7_75t_R FILLER_10_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_622 ();
 DECAPx1_ASAP7_75t_R FILLER_10_651 ();
 FILLER_ASAP7_75t_R FILLER_10_664 ();
 FILLER_ASAP7_75t_R FILLER_10_669 ();
 DECAPx2_ASAP7_75t_R FILLER_10_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_691 ();
 DECAPx2_ASAP7_75t_R FILLER_10_706 ();
 FILLER_ASAP7_75t_R FILLER_10_712 ();
 DECAPx1_ASAP7_75t_R FILLER_10_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_738 ();
 DECAPx2_ASAP7_75t_R FILLER_10_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_751 ();
 DECAPx1_ASAP7_75t_R FILLER_10_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_766 ();
 DECAPx1_ASAP7_75t_R FILLER_10_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_780 ();
 DECAPx6_ASAP7_75t_R FILLER_10_790 ();
 DECAPx2_ASAP7_75t_R FILLER_10_804 ();
 FILLER_ASAP7_75t_R FILLER_10_813 ();
 DECAPx4_ASAP7_75t_R FILLER_10_818 ();
 FILLER_ASAP7_75t_R FILLER_10_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_830 ();
 DECAPx2_ASAP7_75t_R FILLER_10_834 ();
 FILLER_ASAP7_75t_R FILLER_10_846 ();
 DECAPx10_ASAP7_75t_R FILLER_10_879 ();
 DECAPx10_ASAP7_75t_R FILLER_10_901 ();
 DECAPx10_ASAP7_75t_R FILLER_10_923 ();
 DECAPx10_ASAP7_75t_R FILLER_10_945 ();
 DECAPx10_ASAP7_75t_R FILLER_10_967 ();
 DECAPx10_ASAP7_75t_R FILLER_10_989 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1011 ();
 DECAPx6_ASAP7_75t_R FILLER_10_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_10_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_11_24 ();
 DECAPx10_ASAP7_75t_R FILLER_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_11_68 ();
 DECAPx10_ASAP7_75t_R FILLER_11_90 ();
 DECAPx10_ASAP7_75t_R FILLER_11_112 ();
 DECAPx10_ASAP7_75t_R FILLER_11_134 ();
 DECAPx10_ASAP7_75t_R FILLER_11_156 ();
 DECAPx10_ASAP7_75t_R FILLER_11_178 ();
 DECAPx10_ASAP7_75t_R FILLER_11_200 ();
 DECAPx10_ASAP7_75t_R FILLER_11_222 ();
 DECAPx10_ASAP7_75t_R FILLER_11_244 ();
 DECAPx10_ASAP7_75t_R FILLER_11_266 ();
 DECAPx10_ASAP7_75t_R FILLER_11_288 ();
 DECAPx10_ASAP7_75t_R FILLER_11_310 ();
 DECAPx10_ASAP7_75t_R FILLER_11_332 ();
 DECAPx10_ASAP7_75t_R FILLER_11_354 ();
 DECAPx10_ASAP7_75t_R FILLER_11_376 ();
 DECAPx10_ASAP7_75t_R FILLER_11_398 ();
 DECAPx10_ASAP7_75t_R FILLER_11_420 ();
 DECAPx10_ASAP7_75t_R FILLER_11_442 ();
 DECAPx10_ASAP7_75t_R FILLER_11_464 ();
 DECAPx10_ASAP7_75t_R FILLER_11_486 ();
 DECAPx10_ASAP7_75t_R FILLER_11_508 ();
 DECAPx10_ASAP7_75t_R FILLER_11_530 ();
 DECAPx6_ASAP7_75t_R FILLER_11_552 ();
 DECAPx2_ASAP7_75t_R FILLER_11_566 ();
 DECAPx2_ASAP7_75t_R FILLER_11_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_614 ();
 DECAPx1_ASAP7_75t_R FILLER_11_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_629 ();
 DECAPx6_ASAP7_75t_R FILLER_11_651 ();
 DECAPx2_ASAP7_75t_R FILLER_11_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_671 ();
 FILLER_ASAP7_75t_R FILLER_11_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_677 ();
 DECAPx2_ASAP7_75t_R FILLER_11_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_687 ();
 DECAPx4_ASAP7_75t_R FILLER_11_694 ();
 DECAPx2_ASAP7_75t_R FILLER_11_713 ();
 DECAPx1_ASAP7_75t_R FILLER_11_728 ();
 FILLER_ASAP7_75t_R FILLER_11_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_737 ();
 DECAPx2_ASAP7_75t_R FILLER_11_750 ();
 FILLER_ASAP7_75t_R FILLER_11_756 ();
 DECAPx2_ASAP7_75t_R FILLER_11_772 ();
 FILLER_ASAP7_75t_R FILLER_11_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_780 ();
 DECAPx2_ASAP7_75t_R FILLER_11_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_807 ();
 DECAPx4_ASAP7_75t_R FILLER_11_822 ();
 DECAPx1_ASAP7_75t_R FILLER_11_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_860 ();
 DECAPx10_ASAP7_75t_R FILLER_11_881 ();
 DECAPx6_ASAP7_75t_R FILLER_11_903 ();
 DECAPx2_ASAP7_75t_R FILLER_11_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_923 ();
 DECAPx10_ASAP7_75t_R FILLER_11_926 ();
 DECAPx10_ASAP7_75t_R FILLER_11_948 ();
 DECAPx10_ASAP7_75t_R FILLER_11_970 ();
 DECAPx10_ASAP7_75t_R FILLER_11_992 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1354 ();
 DECAPx6_ASAP7_75t_R FILLER_11_1376 ();
 FILLER_ASAP7_75t_R FILLER_11_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_12_24 ();
 DECAPx10_ASAP7_75t_R FILLER_12_46 ();
 DECAPx10_ASAP7_75t_R FILLER_12_68 ();
 DECAPx10_ASAP7_75t_R FILLER_12_90 ();
 DECAPx10_ASAP7_75t_R FILLER_12_112 ();
 DECAPx10_ASAP7_75t_R FILLER_12_134 ();
 DECAPx10_ASAP7_75t_R FILLER_12_156 ();
 DECAPx10_ASAP7_75t_R FILLER_12_178 ();
 DECAPx10_ASAP7_75t_R FILLER_12_200 ();
 DECAPx10_ASAP7_75t_R FILLER_12_222 ();
 DECAPx10_ASAP7_75t_R FILLER_12_244 ();
 DECAPx10_ASAP7_75t_R FILLER_12_266 ();
 DECAPx10_ASAP7_75t_R FILLER_12_288 ();
 DECAPx10_ASAP7_75t_R FILLER_12_310 ();
 DECAPx10_ASAP7_75t_R FILLER_12_332 ();
 DECAPx10_ASAP7_75t_R FILLER_12_354 ();
 DECAPx10_ASAP7_75t_R FILLER_12_376 ();
 DECAPx10_ASAP7_75t_R FILLER_12_398 ();
 DECAPx10_ASAP7_75t_R FILLER_12_420 ();
 DECAPx6_ASAP7_75t_R FILLER_12_442 ();
 DECAPx2_ASAP7_75t_R FILLER_12_456 ();
 DECAPx10_ASAP7_75t_R FILLER_12_464 ();
 DECAPx10_ASAP7_75t_R FILLER_12_486 ();
 DECAPx10_ASAP7_75t_R FILLER_12_508 ();
 DECAPx10_ASAP7_75t_R FILLER_12_530 ();
 DECAPx10_ASAP7_75t_R FILLER_12_552 ();
 DECAPx10_ASAP7_75t_R FILLER_12_574 ();
 FILLER_ASAP7_75t_R FILLER_12_596 ();
 FILLER_ASAP7_75t_R FILLER_12_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_646 ();
 DECAPx2_ASAP7_75t_R FILLER_12_650 ();
 FILLER_ASAP7_75t_R FILLER_12_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_665 ();
 DECAPx2_ASAP7_75t_R FILLER_12_680 ();
 FILLER_ASAP7_75t_R FILLER_12_700 ();
 DECAPx1_ASAP7_75t_R FILLER_12_712 ();
 DECAPx1_ASAP7_75t_R FILLER_12_719 ();
 DECAPx2_ASAP7_75t_R FILLER_12_765 ();
 FILLER_ASAP7_75t_R FILLER_12_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_773 ();
 DECAPx2_ASAP7_75t_R FILLER_12_780 ();
 DECAPx1_ASAP7_75t_R FILLER_12_792 ();
 DECAPx1_ASAP7_75t_R FILLER_12_822 ();
 DECAPx10_ASAP7_75t_R FILLER_12_846 ();
 FILLER_ASAP7_75t_R FILLER_12_868 ();
 DECAPx10_ASAP7_75t_R FILLER_12_876 ();
 DECAPx10_ASAP7_75t_R FILLER_12_898 ();
 DECAPx10_ASAP7_75t_R FILLER_12_920 ();
 DECAPx10_ASAP7_75t_R FILLER_12_942 ();
 DECAPx10_ASAP7_75t_R FILLER_12_964 ();
 DECAPx10_ASAP7_75t_R FILLER_12_986 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_12_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_12_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_13_24 ();
 DECAPx10_ASAP7_75t_R FILLER_13_46 ();
 DECAPx10_ASAP7_75t_R FILLER_13_68 ();
 DECAPx10_ASAP7_75t_R FILLER_13_90 ();
 DECAPx10_ASAP7_75t_R FILLER_13_112 ();
 DECAPx10_ASAP7_75t_R FILLER_13_134 ();
 DECAPx10_ASAP7_75t_R FILLER_13_156 ();
 DECAPx10_ASAP7_75t_R FILLER_13_178 ();
 DECAPx10_ASAP7_75t_R FILLER_13_200 ();
 DECAPx10_ASAP7_75t_R FILLER_13_222 ();
 DECAPx10_ASAP7_75t_R FILLER_13_244 ();
 DECAPx10_ASAP7_75t_R FILLER_13_266 ();
 DECAPx10_ASAP7_75t_R FILLER_13_288 ();
 DECAPx10_ASAP7_75t_R FILLER_13_310 ();
 DECAPx10_ASAP7_75t_R FILLER_13_332 ();
 DECAPx10_ASAP7_75t_R FILLER_13_354 ();
 DECAPx10_ASAP7_75t_R FILLER_13_376 ();
 DECAPx10_ASAP7_75t_R FILLER_13_398 ();
 DECAPx10_ASAP7_75t_R FILLER_13_420 ();
 DECAPx10_ASAP7_75t_R FILLER_13_442 ();
 DECAPx10_ASAP7_75t_R FILLER_13_464 ();
 DECAPx10_ASAP7_75t_R FILLER_13_486 ();
 DECAPx10_ASAP7_75t_R FILLER_13_508 ();
 DECAPx10_ASAP7_75t_R FILLER_13_530 ();
 DECAPx10_ASAP7_75t_R FILLER_13_552 ();
 DECAPx10_ASAP7_75t_R FILLER_13_574 ();
 DECAPx6_ASAP7_75t_R FILLER_13_596 ();
 DECAPx1_ASAP7_75t_R FILLER_13_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_614 ();
 DECAPx4_ASAP7_75t_R FILLER_13_627 ();
 FILLER_ASAP7_75t_R FILLER_13_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_639 ();
 DECAPx2_ASAP7_75t_R FILLER_13_643 ();
 FILLER_ASAP7_75t_R FILLER_13_649 ();
 FILLER_ASAP7_75t_R FILLER_13_671 ();
 DECAPx1_ASAP7_75t_R FILLER_13_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_680 ();
 DECAPx1_ASAP7_75t_R FILLER_13_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_698 ();
 DECAPx6_ASAP7_75t_R FILLER_13_719 ();
 DECAPx1_ASAP7_75t_R FILLER_13_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_741 ();
 DECAPx2_ASAP7_75t_R FILLER_13_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_751 ();
 DECAPx4_ASAP7_75t_R FILLER_13_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_765 ();
 FILLER_ASAP7_75t_R FILLER_13_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_771 ();
 DECAPx4_ASAP7_75t_R FILLER_13_789 ();
 DECAPx1_ASAP7_75t_R FILLER_13_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_809 ();
 DECAPx6_ASAP7_75t_R FILLER_13_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_830 ();
 FILLER_ASAP7_75t_R FILLER_13_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_839 ();
 DECAPx2_ASAP7_75t_R FILLER_13_843 ();
 FILLER_ASAP7_75t_R FILLER_13_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_851 ();
 DECAPx10_ASAP7_75t_R FILLER_13_855 ();
 FILLER_ASAP7_75t_R FILLER_13_877 ();
 DECAPx10_ASAP7_75t_R FILLER_13_888 ();
 DECAPx6_ASAP7_75t_R FILLER_13_910 ();
 DECAPx10_ASAP7_75t_R FILLER_13_926 ();
 DECAPx10_ASAP7_75t_R FILLER_13_948 ();
 DECAPx10_ASAP7_75t_R FILLER_13_970 ();
 DECAPx10_ASAP7_75t_R FILLER_13_992 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_13_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_14_2 ();
 DECAPx10_ASAP7_75t_R FILLER_14_24 ();
 DECAPx10_ASAP7_75t_R FILLER_14_46 ();
 DECAPx10_ASAP7_75t_R FILLER_14_68 ();
 DECAPx10_ASAP7_75t_R FILLER_14_90 ();
 DECAPx10_ASAP7_75t_R FILLER_14_112 ();
 DECAPx10_ASAP7_75t_R FILLER_14_134 ();
 DECAPx10_ASAP7_75t_R FILLER_14_156 ();
 DECAPx10_ASAP7_75t_R FILLER_14_178 ();
 DECAPx10_ASAP7_75t_R FILLER_14_200 ();
 DECAPx10_ASAP7_75t_R FILLER_14_222 ();
 DECAPx10_ASAP7_75t_R FILLER_14_244 ();
 DECAPx10_ASAP7_75t_R FILLER_14_266 ();
 DECAPx10_ASAP7_75t_R FILLER_14_288 ();
 DECAPx10_ASAP7_75t_R FILLER_14_310 ();
 DECAPx10_ASAP7_75t_R FILLER_14_332 ();
 DECAPx10_ASAP7_75t_R FILLER_14_354 ();
 DECAPx10_ASAP7_75t_R FILLER_14_376 ();
 DECAPx10_ASAP7_75t_R FILLER_14_398 ();
 DECAPx10_ASAP7_75t_R FILLER_14_420 ();
 DECAPx6_ASAP7_75t_R FILLER_14_442 ();
 DECAPx2_ASAP7_75t_R FILLER_14_456 ();
 DECAPx10_ASAP7_75t_R FILLER_14_464 ();
 DECAPx10_ASAP7_75t_R FILLER_14_486 ();
 DECAPx10_ASAP7_75t_R FILLER_14_508 ();
 DECAPx10_ASAP7_75t_R FILLER_14_530 ();
 DECAPx10_ASAP7_75t_R FILLER_14_552 ();
 DECAPx10_ASAP7_75t_R FILLER_14_574 ();
 DECAPx4_ASAP7_75t_R FILLER_14_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_606 ();
 DECAPx4_ASAP7_75t_R FILLER_14_623 ();
 FILLER_ASAP7_75t_R FILLER_14_633 ();
 DECAPx4_ASAP7_75t_R FILLER_14_645 ();
 FILLER_ASAP7_75t_R FILLER_14_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_657 ();
 DECAPx6_ASAP7_75t_R FILLER_14_668 ();
 DECAPx1_ASAP7_75t_R FILLER_14_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_686 ();
 DECAPx6_ASAP7_75t_R FILLER_14_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_710 ();
 DECAPx2_ASAP7_75t_R FILLER_14_714 ();
 FILLER_ASAP7_75t_R FILLER_14_720 ();
 FILLER_ASAP7_75t_R FILLER_14_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_727 ();
 DECAPx10_ASAP7_75t_R FILLER_14_742 ();
 FILLER_ASAP7_75t_R FILLER_14_764 ();
 DECAPx2_ASAP7_75t_R FILLER_14_780 ();
 DECAPx4_ASAP7_75t_R FILLER_14_789 ();
 FILLER_ASAP7_75t_R FILLER_14_799 ();
 FILLER_ASAP7_75t_R FILLER_14_810 ();
 DECAPx2_ASAP7_75t_R FILLER_14_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_832 ();
 DECAPx1_ASAP7_75t_R FILLER_14_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_869 ();
 DECAPx10_ASAP7_75t_R FILLER_14_876 ();
 DECAPx10_ASAP7_75t_R FILLER_14_898 ();
 DECAPx10_ASAP7_75t_R FILLER_14_920 ();
 DECAPx10_ASAP7_75t_R FILLER_14_942 ();
 DECAPx10_ASAP7_75t_R FILLER_14_964 ();
 DECAPx10_ASAP7_75t_R FILLER_14_986 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_14_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_14_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_15_2 ();
 DECAPx10_ASAP7_75t_R FILLER_15_24 ();
 DECAPx10_ASAP7_75t_R FILLER_15_46 ();
 DECAPx10_ASAP7_75t_R FILLER_15_68 ();
 DECAPx10_ASAP7_75t_R FILLER_15_90 ();
 DECAPx10_ASAP7_75t_R FILLER_15_112 ();
 DECAPx10_ASAP7_75t_R FILLER_15_134 ();
 DECAPx10_ASAP7_75t_R FILLER_15_156 ();
 DECAPx10_ASAP7_75t_R FILLER_15_178 ();
 DECAPx10_ASAP7_75t_R FILLER_15_200 ();
 DECAPx10_ASAP7_75t_R FILLER_15_222 ();
 DECAPx10_ASAP7_75t_R FILLER_15_244 ();
 DECAPx10_ASAP7_75t_R FILLER_15_266 ();
 DECAPx10_ASAP7_75t_R FILLER_15_288 ();
 DECAPx10_ASAP7_75t_R FILLER_15_310 ();
 DECAPx10_ASAP7_75t_R FILLER_15_332 ();
 DECAPx10_ASAP7_75t_R FILLER_15_354 ();
 DECAPx10_ASAP7_75t_R FILLER_15_376 ();
 DECAPx10_ASAP7_75t_R FILLER_15_398 ();
 DECAPx10_ASAP7_75t_R FILLER_15_420 ();
 DECAPx10_ASAP7_75t_R FILLER_15_442 ();
 DECAPx10_ASAP7_75t_R FILLER_15_464 ();
 DECAPx10_ASAP7_75t_R FILLER_15_486 ();
 DECAPx10_ASAP7_75t_R FILLER_15_508 ();
 DECAPx10_ASAP7_75t_R FILLER_15_530 ();
 DECAPx10_ASAP7_75t_R FILLER_15_552 ();
 DECAPx10_ASAP7_75t_R FILLER_15_574 ();
 DECAPx4_ASAP7_75t_R FILLER_15_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_606 ();
 FILLER_ASAP7_75t_R FILLER_15_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_625 ();
 DECAPx4_ASAP7_75t_R FILLER_15_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_670 ();
 DECAPx6_ASAP7_75t_R FILLER_15_681 ();
 DECAPx1_ASAP7_75t_R FILLER_15_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_714 ();
 FILLER_ASAP7_75t_R FILLER_15_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_731 ();
 FILLER_ASAP7_75t_R FILLER_15_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_754 ();
 DECAPx2_ASAP7_75t_R FILLER_15_792 ();
 DECAPx2_ASAP7_75t_R FILLER_15_801 ();
 FILLER_ASAP7_75t_R FILLER_15_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_809 ();
 DECAPx4_ASAP7_75t_R FILLER_15_819 ();
 DECAPx2_ASAP7_75t_R FILLER_15_849 ();
 DECAPx1_ASAP7_75t_R FILLER_15_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_878 ();
 DECAPx10_ASAP7_75t_R FILLER_15_882 ();
 DECAPx6_ASAP7_75t_R FILLER_15_904 ();
 DECAPx2_ASAP7_75t_R FILLER_15_918 ();
 DECAPx10_ASAP7_75t_R FILLER_15_926 ();
 DECAPx10_ASAP7_75t_R FILLER_15_948 ();
 DECAPx10_ASAP7_75t_R FILLER_15_970 ();
 DECAPx10_ASAP7_75t_R FILLER_15_992 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_15_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_16_2 ();
 DECAPx10_ASAP7_75t_R FILLER_16_24 ();
 DECAPx10_ASAP7_75t_R FILLER_16_46 ();
 DECAPx10_ASAP7_75t_R FILLER_16_68 ();
 DECAPx10_ASAP7_75t_R FILLER_16_90 ();
 DECAPx10_ASAP7_75t_R FILLER_16_112 ();
 DECAPx10_ASAP7_75t_R FILLER_16_134 ();
 DECAPx10_ASAP7_75t_R FILLER_16_156 ();
 DECAPx10_ASAP7_75t_R FILLER_16_178 ();
 DECAPx10_ASAP7_75t_R FILLER_16_200 ();
 DECAPx10_ASAP7_75t_R FILLER_16_222 ();
 DECAPx10_ASAP7_75t_R FILLER_16_244 ();
 DECAPx10_ASAP7_75t_R FILLER_16_266 ();
 DECAPx10_ASAP7_75t_R FILLER_16_288 ();
 DECAPx10_ASAP7_75t_R FILLER_16_310 ();
 DECAPx10_ASAP7_75t_R FILLER_16_332 ();
 DECAPx10_ASAP7_75t_R FILLER_16_354 ();
 DECAPx10_ASAP7_75t_R FILLER_16_376 ();
 DECAPx10_ASAP7_75t_R FILLER_16_398 ();
 DECAPx10_ASAP7_75t_R FILLER_16_420 ();
 DECAPx6_ASAP7_75t_R FILLER_16_442 ();
 DECAPx2_ASAP7_75t_R FILLER_16_456 ();
 DECAPx10_ASAP7_75t_R FILLER_16_464 ();
 DECAPx10_ASAP7_75t_R FILLER_16_486 ();
 DECAPx10_ASAP7_75t_R FILLER_16_508 ();
 DECAPx10_ASAP7_75t_R FILLER_16_530 ();
 DECAPx10_ASAP7_75t_R FILLER_16_552 ();
 DECAPx10_ASAP7_75t_R FILLER_16_574 ();
 DECAPx4_ASAP7_75t_R FILLER_16_596 ();
 FILLER_ASAP7_75t_R FILLER_16_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_634 ();
 DECAPx4_ASAP7_75t_R FILLER_16_641 ();
 FILLER_ASAP7_75t_R FILLER_16_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_653 ();
 DECAPx1_ASAP7_75t_R FILLER_16_660 ();
 DECAPx1_ASAP7_75t_R FILLER_16_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_696 ();
 DECAPx1_ASAP7_75t_R FILLER_16_713 ();
 DECAPx4_ASAP7_75t_R FILLER_16_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_736 ();
 DECAPx4_ASAP7_75t_R FILLER_16_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_750 ();
 DECAPx2_ASAP7_75t_R FILLER_16_771 ();
 DECAPx6_ASAP7_75t_R FILLER_16_780 ();
 FILLER_ASAP7_75t_R FILLER_16_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_796 ();
 DECAPx4_ASAP7_75t_R FILLER_16_803 ();
 FILLER_ASAP7_75t_R FILLER_16_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_815 ();
 DECAPx4_ASAP7_75t_R FILLER_16_825 ();
 DECAPx6_ASAP7_75t_R FILLER_16_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_878 ();
 DECAPx10_ASAP7_75t_R FILLER_16_891 ();
 DECAPx10_ASAP7_75t_R FILLER_16_913 ();
 DECAPx10_ASAP7_75t_R FILLER_16_935 ();
 DECAPx10_ASAP7_75t_R FILLER_16_957 ();
 DECAPx10_ASAP7_75t_R FILLER_16_979 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1353 ();
 DECAPx4_ASAP7_75t_R FILLER_16_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_16_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_17_2 ();
 DECAPx10_ASAP7_75t_R FILLER_17_24 ();
 DECAPx10_ASAP7_75t_R FILLER_17_46 ();
 DECAPx10_ASAP7_75t_R FILLER_17_68 ();
 DECAPx10_ASAP7_75t_R FILLER_17_90 ();
 DECAPx10_ASAP7_75t_R FILLER_17_112 ();
 DECAPx10_ASAP7_75t_R FILLER_17_134 ();
 DECAPx10_ASAP7_75t_R FILLER_17_156 ();
 DECAPx10_ASAP7_75t_R FILLER_17_178 ();
 DECAPx10_ASAP7_75t_R FILLER_17_200 ();
 DECAPx10_ASAP7_75t_R FILLER_17_222 ();
 DECAPx10_ASAP7_75t_R FILLER_17_244 ();
 DECAPx10_ASAP7_75t_R FILLER_17_266 ();
 DECAPx10_ASAP7_75t_R FILLER_17_288 ();
 DECAPx10_ASAP7_75t_R FILLER_17_310 ();
 DECAPx10_ASAP7_75t_R FILLER_17_332 ();
 DECAPx10_ASAP7_75t_R FILLER_17_354 ();
 DECAPx10_ASAP7_75t_R FILLER_17_376 ();
 DECAPx10_ASAP7_75t_R FILLER_17_398 ();
 DECAPx10_ASAP7_75t_R FILLER_17_420 ();
 DECAPx10_ASAP7_75t_R FILLER_17_442 ();
 DECAPx10_ASAP7_75t_R FILLER_17_464 ();
 DECAPx10_ASAP7_75t_R FILLER_17_486 ();
 DECAPx10_ASAP7_75t_R FILLER_17_508 ();
 DECAPx10_ASAP7_75t_R FILLER_17_530 ();
 DECAPx10_ASAP7_75t_R FILLER_17_552 ();
 DECAPx10_ASAP7_75t_R FILLER_17_574 ();
 DECAPx4_ASAP7_75t_R FILLER_17_596 ();
 FILLER_ASAP7_75t_R FILLER_17_606 ();
 DECAPx10_ASAP7_75t_R FILLER_17_618 ();
 DECAPx4_ASAP7_75t_R FILLER_17_640 ();
 FILLER_ASAP7_75t_R FILLER_17_650 ();
 DECAPx2_ASAP7_75t_R FILLER_17_662 ();
 FILLER_ASAP7_75t_R FILLER_17_668 ();
 DECAPx4_ASAP7_75t_R FILLER_17_676 ();
 FILLER_ASAP7_75t_R FILLER_17_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_694 ();
 DECAPx1_ASAP7_75t_R FILLER_17_701 ();
 FILLER_ASAP7_75t_R FILLER_17_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_713 ();
 DECAPx1_ASAP7_75t_R FILLER_17_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_721 ();
 DECAPx2_ASAP7_75t_R FILLER_17_725 ();
 FILLER_ASAP7_75t_R FILLER_17_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_733 ();
 DECAPx6_ASAP7_75t_R FILLER_17_748 ();
 FILLER_ASAP7_75t_R FILLER_17_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_764 ();
 DECAPx1_ASAP7_75t_R FILLER_17_774 ();
 DECAPx4_ASAP7_75t_R FILLER_17_781 ();
 FILLER_ASAP7_75t_R FILLER_17_791 ();
 DECAPx4_ASAP7_75t_R FILLER_17_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_812 ();
 DECAPx6_ASAP7_75t_R FILLER_17_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_847 ();
 FILLER_ASAP7_75t_R FILLER_17_854 ();
 DECAPx4_ASAP7_75t_R FILLER_17_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_884 ();
 DECAPx10_ASAP7_75t_R FILLER_17_894 ();
 DECAPx2_ASAP7_75t_R FILLER_17_916 ();
 FILLER_ASAP7_75t_R FILLER_17_922 ();
 DECAPx10_ASAP7_75t_R FILLER_17_926 ();
 DECAPx10_ASAP7_75t_R FILLER_17_948 ();
 DECAPx10_ASAP7_75t_R FILLER_17_970 ();
 DECAPx10_ASAP7_75t_R FILLER_17_992 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_17_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_18_2 ();
 DECAPx10_ASAP7_75t_R FILLER_18_24 ();
 DECAPx10_ASAP7_75t_R FILLER_18_46 ();
 DECAPx10_ASAP7_75t_R FILLER_18_68 ();
 DECAPx10_ASAP7_75t_R FILLER_18_90 ();
 DECAPx10_ASAP7_75t_R FILLER_18_112 ();
 DECAPx10_ASAP7_75t_R FILLER_18_134 ();
 DECAPx10_ASAP7_75t_R FILLER_18_156 ();
 DECAPx10_ASAP7_75t_R FILLER_18_178 ();
 DECAPx10_ASAP7_75t_R FILLER_18_200 ();
 DECAPx10_ASAP7_75t_R FILLER_18_222 ();
 DECAPx10_ASAP7_75t_R FILLER_18_244 ();
 DECAPx10_ASAP7_75t_R FILLER_18_266 ();
 DECAPx10_ASAP7_75t_R FILLER_18_288 ();
 DECAPx10_ASAP7_75t_R FILLER_18_310 ();
 DECAPx10_ASAP7_75t_R FILLER_18_332 ();
 DECAPx10_ASAP7_75t_R FILLER_18_354 ();
 DECAPx10_ASAP7_75t_R FILLER_18_376 ();
 DECAPx10_ASAP7_75t_R FILLER_18_398 ();
 DECAPx10_ASAP7_75t_R FILLER_18_420 ();
 DECAPx6_ASAP7_75t_R FILLER_18_442 ();
 DECAPx2_ASAP7_75t_R FILLER_18_456 ();
 DECAPx10_ASAP7_75t_R FILLER_18_464 ();
 DECAPx10_ASAP7_75t_R FILLER_18_486 ();
 DECAPx10_ASAP7_75t_R FILLER_18_508 ();
 DECAPx10_ASAP7_75t_R FILLER_18_530 ();
 DECAPx10_ASAP7_75t_R FILLER_18_552 ();
 DECAPx6_ASAP7_75t_R FILLER_18_574 ();
 DECAPx1_ASAP7_75t_R FILLER_18_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_592 ();
 FILLER_ASAP7_75t_R FILLER_18_605 ();
 FILLER_ASAP7_75t_R FILLER_18_621 ();
 DECAPx4_ASAP7_75t_R FILLER_18_629 ();
 FILLER_ASAP7_75t_R FILLER_18_639 ();
 DECAPx2_ASAP7_75t_R FILLER_18_647 ();
 DECAPx6_ASAP7_75t_R FILLER_18_665 ();
 FILLER_ASAP7_75t_R FILLER_18_679 ();
 DECAPx6_ASAP7_75t_R FILLER_18_687 ();
 DECAPx2_ASAP7_75t_R FILLER_18_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_707 ();
 DECAPx2_ASAP7_75t_R FILLER_18_717 ();
 FILLER_ASAP7_75t_R FILLER_18_723 ();
 DECAPx2_ASAP7_75t_R FILLER_18_734 ();
 FILLER_ASAP7_75t_R FILLER_18_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_742 ();
 DECAPx2_ASAP7_75t_R FILLER_18_746 ();
 FILLER_ASAP7_75t_R FILLER_18_752 ();
 FILLER_ASAP7_75t_R FILLER_18_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_768 ();
 DECAPx1_ASAP7_75t_R FILLER_18_783 ();
 FILLER_ASAP7_75t_R FILLER_18_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_813 ();
 DECAPx2_ASAP7_75t_R FILLER_18_826 ();
 FILLER_ASAP7_75t_R FILLER_18_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_865 ();
 DECAPx2_ASAP7_75t_R FILLER_18_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_875 ();
 DECAPx10_ASAP7_75t_R FILLER_18_889 ();
 DECAPx10_ASAP7_75t_R FILLER_18_911 ();
 DECAPx10_ASAP7_75t_R FILLER_18_933 ();
 DECAPx10_ASAP7_75t_R FILLER_18_955 ();
 DECAPx10_ASAP7_75t_R FILLER_18_977 ();
 DECAPx10_ASAP7_75t_R FILLER_18_999 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1351 ();
 DECAPx4_ASAP7_75t_R FILLER_18_1373 ();
 FILLER_ASAP7_75t_R FILLER_18_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_18_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_19_2 ();
 DECAPx10_ASAP7_75t_R FILLER_19_24 ();
 DECAPx10_ASAP7_75t_R FILLER_19_46 ();
 DECAPx10_ASAP7_75t_R FILLER_19_68 ();
 DECAPx10_ASAP7_75t_R FILLER_19_90 ();
 DECAPx10_ASAP7_75t_R FILLER_19_112 ();
 DECAPx10_ASAP7_75t_R FILLER_19_134 ();
 DECAPx10_ASAP7_75t_R FILLER_19_156 ();
 DECAPx10_ASAP7_75t_R FILLER_19_178 ();
 DECAPx10_ASAP7_75t_R FILLER_19_200 ();
 DECAPx10_ASAP7_75t_R FILLER_19_222 ();
 DECAPx10_ASAP7_75t_R FILLER_19_244 ();
 DECAPx10_ASAP7_75t_R FILLER_19_266 ();
 DECAPx10_ASAP7_75t_R FILLER_19_288 ();
 DECAPx10_ASAP7_75t_R FILLER_19_310 ();
 DECAPx10_ASAP7_75t_R FILLER_19_332 ();
 DECAPx10_ASAP7_75t_R FILLER_19_354 ();
 DECAPx10_ASAP7_75t_R FILLER_19_376 ();
 DECAPx10_ASAP7_75t_R FILLER_19_398 ();
 DECAPx10_ASAP7_75t_R FILLER_19_420 ();
 DECAPx10_ASAP7_75t_R FILLER_19_442 ();
 DECAPx10_ASAP7_75t_R FILLER_19_464 ();
 DECAPx10_ASAP7_75t_R FILLER_19_486 ();
 DECAPx10_ASAP7_75t_R FILLER_19_508 ();
 DECAPx10_ASAP7_75t_R FILLER_19_530 ();
 DECAPx10_ASAP7_75t_R FILLER_19_552 ();
 DECAPx2_ASAP7_75t_R FILLER_19_574 ();
 FILLER_ASAP7_75t_R FILLER_19_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_582 ();
 DECAPx1_ASAP7_75t_R FILLER_19_589 ();
 FILLER_ASAP7_75t_R FILLER_19_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_612 ();
 FILLER_ASAP7_75t_R FILLER_19_630 ();
 DECAPx1_ASAP7_75t_R FILLER_19_652 ();
 DECAPx2_ASAP7_75t_R FILLER_19_670 ();
 FILLER_ASAP7_75t_R FILLER_19_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_705 ();
 DECAPx4_ASAP7_75t_R FILLER_19_709 ();
 FILLER_ASAP7_75t_R FILLER_19_719 ();
 FILLER_ASAP7_75t_R FILLER_19_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_726 ();
 FILLER_ASAP7_75t_R FILLER_19_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_758 ();
 DECAPx2_ASAP7_75t_R FILLER_19_776 ();
 FILLER_ASAP7_75t_R FILLER_19_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_818 ();
 FILLER_ASAP7_75t_R FILLER_19_840 ();
 DECAPx6_ASAP7_75t_R FILLER_19_856 ();
 DECAPx2_ASAP7_75t_R FILLER_19_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_876 ();
 DECAPx10_ASAP7_75t_R FILLER_19_899 ();
 FILLER_ASAP7_75t_R FILLER_19_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_923 ();
 DECAPx10_ASAP7_75t_R FILLER_19_926 ();
 DECAPx10_ASAP7_75t_R FILLER_19_948 ();
 DECAPx10_ASAP7_75t_R FILLER_19_970 ();
 DECAPx10_ASAP7_75t_R FILLER_19_992 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_19_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_20_2 ();
 DECAPx10_ASAP7_75t_R FILLER_20_24 ();
 DECAPx10_ASAP7_75t_R FILLER_20_46 ();
 DECAPx10_ASAP7_75t_R FILLER_20_68 ();
 DECAPx10_ASAP7_75t_R FILLER_20_90 ();
 DECAPx10_ASAP7_75t_R FILLER_20_112 ();
 DECAPx10_ASAP7_75t_R FILLER_20_134 ();
 DECAPx10_ASAP7_75t_R FILLER_20_156 ();
 DECAPx10_ASAP7_75t_R FILLER_20_178 ();
 DECAPx10_ASAP7_75t_R FILLER_20_200 ();
 DECAPx10_ASAP7_75t_R FILLER_20_222 ();
 DECAPx10_ASAP7_75t_R FILLER_20_244 ();
 DECAPx10_ASAP7_75t_R FILLER_20_266 ();
 DECAPx10_ASAP7_75t_R FILLER_20_288 ();
 DECAPx10_ASAP7_75t_R FILLER_20_310 ();
 DECAPx10_ASAP7_75t_R FILLER_20_332 ();
 DECAPx10_ASAP7_75t_R FILLER_20_354 ();
 DECAPx10_ASAP7_75t_R FILLER_20_376 ();
 DECAPx10_ASAP7_75t_R FILLER_20_398 ();
 DECAPx10_ASAP7_75t_R FILLER_20_420 ();
 DECAPx6_ASAP7_75t_R FILLER_20_442 ();
 DECAPx2_ASAP7_75t_R FILLER_20_456 ();
 DECAPx10_ASAP7_75t_R FILLER_20_464 ();
 DECAPx10_ASAP7_75t_R FILLER_20_486 ();
 DECAPx10_ASAP7_75t_R FILLER_20_508 ();
 DECAPx10_ASAP7_75t_R FILLER_20_530 ();
 DECAPx4_ASAP7_75t_R FILLER_20_552 ();
 FILLER_ASAP7_75t_R FILLER_20_562 ();
 DECAPx4_ASAP7_75t_R FILLER_20_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_596 ();
 DECAPx6_ASAP7_75t_R FILLER_20_603 ();
 DECAPx2_ASAP7_75t_R FILLER_20_629 ();
 FILLER_ASAP7_75t_R FILLER_20_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_637 ();
 FILLER_ASAP7_75t_R FILLER_20_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_667 ();
 FILLER_ASAP7_75t_R FILLER_20_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_673 ();
 FILLER_ASAP7_75t_R FILLER_20_705 ();
 DECAPx2_ASAP7_75t_R FILLER_20_721 ();
 DECAPx4_ASAP7_75t_R FILLER_20_747 ();
 FILLER_ASAP7_75t_R FILLER_20_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_759 ();
 DECAPx6_ASAP7_75t_R FILLER_20_766 ();
 DECAPx2_ASAP7_75t_R FILLER_20_780 ();
 DECAPx1_ASAP7_75t_R FILLER_20_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_811 ();
 DECAPx1_ASAP7_75t_R FILLER_20_830 ();
 DECAPx4_ASAP7_75t_R FILLER_20_850 ();
 FILLER_ASAP7_75t_R FILLER_20_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_862 ();
 DECAPx1_ASAP7_75t_R FILLER_20_875 ();
 DECAPx10_ASAP7_75t_R FILLER_20_897 ();
 DECAPx10_ASAP7_75t_R FILLER_20_919 ();
 DECAPx10_ASAP7_75t_R FILLER_20_941 ();
 DECAPx10_ASAP7_75t_R FILLER_20_963 ();
 DECAPx10_ASAP7_75t_R FILLER_20_985 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_20_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_20_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_21_2 ();
 DECAPx10_ASAP7_75t_R FILLER_21_24 ();
 DECAPx10_ASAP7_75t_R FILLER_21_46 ();
 DECAPx10_ASAP7_75t_R FILLER_21_68 ();
 DECAPx10_ASAP7_75t_R FILLER_21_90 ();
 DECAPx10_ASAP7_75t_R FILLER_21_112 ();
 DECAPx10_ASAP7_75t_R FILLER_21_134 ();
 DECAPx10_ASAP7_75t_R FILLER_21_156 ();
 DECAPx10_ASAP7_75t_R FILLER_21_178 ();
 DECAPx10_ASAP7_75t_R FILLER_21_200 ();
 DECAPx10_ASAP7_75t_R FILLER_21_222 ();
 DECAPx10_ASAP7_75t_R FILLER_21_244 ();
 DECAPx10_ASAP7_75t_R FILLER_21_266 ();
 DECAPx10_ASAP7_75t_R FILLER_21_288 ();
 DECAPx10_ASAP7_75t_R FILLER_21_310 ();
 DECAPx10_ASAP7_75t_R FILLER_21_332 ();
 DECAPx10_ASAP7_75t_R FILLER_21_354 ();
 DECAPx10_ASAP7_75t_R FILLER_21_376 ();
 DECAPx10_ASAP7_75t_R FILLER_21_398 ();
 DECAPx10_ASAP7_75t_R FILLER_21_420 ();
 DECAPx10_ASAP7_75t_R FILLER_21_442 ();
 DECAPx10_ASAP7_75t_R FILLER_21_464 ();
 DECAPx10_ASAP7_75t_R FILLER_21_486 ();
 DECAPx10_ASAP7_75t_R FILLER_21_508 ();
 DECAPx10_ASAP7_75t_R FILLER_21_530 ();
 DECAPx1_ASAP7_75t_R FILLER_21_552 ();
 DECAPx2_ASAP7_75t_R FILLER_21_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_580 ();
 DECAPx10_ASAP7_75t_R FILLER_21_598 ();
 FILLER_ASAP7_75t_R FILLER_21_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_622 ();
 FILLER_ASAP7_75t_R FILLER_21_626 ();
 DECAPx4_ASAP7_75t_R FILLER_21_631 ();
 DECAPx4_ASAP7_75t_R FILLER_21_644 ();
 DECAPx2_ASAP7_75t_R FILLER_21_682 ();
 FILLER_ASAP7_75t_R FILLER_21_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_690 ();
 DECAPx1_ASAP7_75t_R FILLER_21_697 ();
 FILLER_ASAP7_75t_R FILLER_21_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_709 ();
 FILLER_ASAP7_75t_R FILLER_21_727 ();
 DECAPx2_ASAP7_75t_R FILLER_21_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_755 ();
 FILLER_ASAP7_75t_R FILLER_21_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_775 ();
 DECAPx2_ASAP7_75t_R FILLER_21_785 ();
 FILLER_ASAP7_75t_R FILLER_21_791 ();
 DECAPx2_ASAP7_75t_R FILLER_21_805 ();
 FILLER_ASAP7_75t_R FILLER_21_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_813 ();
 DECAPx2_ASAP7_75t_R FILLER_21_820 ();
 FILLER_ASAP7_75t_R FILLER_21_826 ();
 FILLER_ASAP7_75t_R FILLER_21_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_850 ();
 DECAPx10_ASAP7_75t_R FILLER_21_854 ();
 FILLER_ASAP7_75t_R FILLER_21_876 ();
 DECAPx10_ASAP7_75t_R FILLER_21_895 ();
 DECAPx2_ASAP7_75t_R FILLER_21_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_923 ();
 DECAPx10_ASAP7_75t_R FILLER_21_926 ();
 DECAPx10_ASAP7_75t_R FILLER_21_948 ();
 DECAPx10_ASAP7_75t_R FILLER_21_970 ();
 DECAPx10_ASAP7_75t_R FILLER_21_992 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_21_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_22_2 ();
 DECAPx10_ASAP7_75t_R FILLER_22_24 ();
 DECAPx10_ASAP7_75t_R FILLER_22_46 ();
 DECAPx10_ASAP7_75t_R FILLER_22_68 ();
 DECAPx10_ASAP7_75t_R FILLER_22_90 ();
 DECAPx10_ASAP7_75t_R FILLER_22_112 ();
 DECAPx10_ASAP7_75t_R FILLER_22_134 ();
 DECAPx10_ASAP7_75t_R FILLER_22_156 ();
 DECAPx10_ASAP7_75t_R FILLER_22_178 ();
 DECAPx10_ASAP7_75t_R FILLER_22_200 ();
 DECAPx10_ASAP7_75t_R FILLER_22_222 ();
 DECAPx10_ASAP7_75t_R FILLER_22_244 ();
 DECAPx10_ASAP7_75t_R FILLER_22_266 ();
 DECAPx10_ASAP7_75t_R FILLER_22_288 ();
 DECAPx10_ASAP7_75t_R FILLER_22_310 ();
 DECAPx10_ASAP7_75t_R FILLER_22_332 ();
 DECAPx10_ASAP7_75t_R FILLER_22_354 ();
 DECAPx10_ASAP7_75t_R FILLER_22_376 ();
 DECAPx10_ASAP7_75t_R FILLER_22_398 ();
 DECAPx10_ASAP7_75t_R FILLER_22_420 ();
 DECAPx6_ASAP7_75t_R FILLER_22_442 ();
 DECAPx2_ASAP7_75t_R FILLER_22_456 ();
 DECAPx10_ASAP7_75t_R FILLER_22_464 ();
 DECAPx10_ASAP7_75t_R FILLER_22_486 ();
 DECAPx10_ASAP7_75t_R FILLER_22_508 ();
 DECAPx10_ASAP7_75t_R FILLER_22_530 ();
 DECAPx10_ASAP7_75t_R FILLER_22_552 ();
 DECAPx2_ASAP7_75t_R FILLER_22_574 ();
 FILLER_ASAP7_75t_R FILLER_22_580 ();
 DECAPx1_ASAP7_75t_R FILLER_22_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_589 ();
 DECAPx6_ASAP7_75t_R FILLER_22_593 ();
 DECAPx1_ASAP7_75t_R FILLER_22_607 ();
 FILLER_ASAP7_75t_R FILLER_22_617 ();
 DECAPx6_ASAP7_75t_R FILLER_22_653 ();
 FILLER_ASAP7_75t_R FILLER_22_667 ();
 DECAPx6_ASAP7_75t_R FILLER_22_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_692 ();
 DECAPx4_ASAP7_75t_R FILLER_22_702 ();
 FILLER_ASAP7_75t_R FILLER_22_712 ();
 DECAPx1_ASAP7_75t_R FILLER_22_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_732 ();
 DECAPx4_ASAP7_75t_R FILLER_22_736 ();
 FILLER_ASAP7_75t_R FILLER_22_746 ();
 DECAPx6_ASAP7_75t_R FILLER_22_765 ();
 DECAPx1_ASAP7_75t_R FILLER_22_790 ();
 DECAPx4_ASAP7_75t_R FILLER_22_800 ();
 FILLER_ASAP7_75t_R FILLER_22_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_829 ();
 DECAPx1_ASAP7_75t_R FILLER_22_836 ();
 DECAPx4_ASAP7_75t_R FILLER_22_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_864 ();
 DECAPx2_ASAP7_75t_R FILLER_22_868 ();
 FILLER_ASAP7_75t_R FILLER_22_883 ();
 DECAPx10_ASAP7_75t_R FILLER_22_898 ();
 DECAPx10_ASAP7_75t_R FILLER_22_920 ();
 DECAPx10_ASAP7_75t_R FILLER_22_942 ();
 DECAPx10_ASAP7_75t_R FILLER_22_964 ();
 DECAPx10_ASAP7_75t_R FILLER_22_986 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_22_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_22_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_23_2 ();
 DECAPx10_ASAP7_75t_R FILLER_23_24 ();
 DECAPx10_ASAP7_75t_R FILLER_23_46 ();
 DECAPx10_ASAP7_75t_R FILLER_23_68 ();
 DECAPx10_ASAP7_75t_R FILLER_23_90 ();
 DECAPx10_ASAP7_75t_R FILLER_23_112 ();
 DECAPx10_ASAP7_75t_R FILLER_23_134 ();
 DECAPx10_ASAP7_75t_R FILLER_23_156 ();
 DECAPx10_ASAP7_75t_R FILLER_23_178 ();
 DECAPx10_ASAP7_75t_R FILLER_23_200 ();
 DECAPx10_ASAP7_75t_R FILLER_23_222 ();
 DECAPx10_ASAP7_75t_R FILLER_23_244 ();
 DECAPx10_ASAP7_75t_R FILLER_23_266 ();
 DECAPx10_ASAP7_75t_R FILLER_23_288 ();
 DECAPx10_ASAP7_75t_R FILLER_23_310 ();
 DECAPx10_ASAP7_75t_R FILLER_23_332 ();
 DECAPx10_ASAP7_75t_R FILLER_23_354 ();
 DECAPx10_ASAP7_75t_R FILLER_23_376 ();
 DECAPx10_ASAP7_75t_R FILLER_23_398 ();
 DECAPx10_ASAP7_75t_R FILLER_23_420 ();
 DECAPx10_ASAP7_75t_R FILLER_23_442 ();
 DECAPx10_ASAP7_75t_R FILLER_23_464 ();
 DECAPx10_ASAP7_75t_R FILLER_23_486 ();
 DECAPx10_ASAP7_75t_R FILLER_23_508 ();
 DECAPx10_ASAP7_75t_R FILLER_23_530 ();
 DECAPx6_ASAP7_75t_R FILLER_23_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_573 ();
 FILLER_ASAP7_75t_R FILLER_23_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_588 ();
 DECAPx1_ASAP7_75t_R FILLER_23_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_607 ();
 FILLER_ASAP7_75t_R FILLER_23_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_624 ();
 FILLER_ASAP7_75t_R FILLER_23_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_630 ();
 DECAPx2_ASAP7_75t_R FILLER_23_651 ();
 DECAPx2_ASAP7_75t_R FILLER_23_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_672 ();
 DECAPx2_ASAP7_75t_R FILLER_23_676 ();
 DECAPx2_ASAP7_75t_R FILLER_23_702 ();
 FILLER_ASAP7_75t_R FILLER_23_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_717 ();
 DECAPx1_ASAP7_75t_R FILLER_23_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_725 ();
 DECAPx4_ASAP7_75t_R FILLER_23_732 ();
 FILLER_ASAP7_75t_R FILLER_23_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_758 ();
 FILLER_ASAP7_75t_R FILLER_23_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_764 ();
 DECAPx1_ASAP7_75t_R FILLER_23_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_775 ();
 DECAPx10_ASAP7_75t_R FILLER_23_779 ();
 FILLER_ASAP7_75t_R FILLER_23_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_809 ();
 DECAPx10_ASAP7_75t_R FILLER_23_819 ();
 DECAPx2_ASAP7_75t_R FILLER_23_841 ();
 FILLER_ASAP7_75t_R FILLER_23_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_849 ();
 DECAPx1_ASAP7_75t_R FILLER_23_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_857 ();
 DECAPx1_ASAP7_75t_R FILLER_23_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_875 ();
 DECAPx10_ASAP7_75t_R FILLER_23_895 ();
 DECAPx2_ASAP7_75t_R FILLER_23_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_923 ();
 DECAPx10_ASAP7_75t_R FILLER_23_926 ();
 DECAPx10_ASAP7_75t_R FILLER_23_948 ();
 DECAPx10_ASAP7_75t_R FILLER_23_970 ();
 DECAPx10_ASAP7_75t_R FILLER_23_992 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_23_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_24_2 ();
 DECAPx10_ASAP7_75t_R FILLER_24_24 ();
 DECAPx10_ASAP7_75t_R FILLER_24_46 ();
 DECAPx10_ASAP7_75t_R FILLER_24_68 ();
 DECAPx10_ASAP7_75t_R FILLER_24_90 ();
 DECAPx10_ASAP7_75t_R FILLER_24_112 ();
 DECAPx10_ASAP7_75t_R FILLER_24_134 ();
 DECAPx10_ASAP7_75t_R FILLER_24_156 ();
 DECAPx10_ASAP7_75t_R FILLER_24_178 ();
 DECAPx10_ASAP7_75t_R FILLER_24_200 ();
 DECAPx10_ASAP7_75t_R FILLER_24_222 ();
 DECAPx10_ASAP7_75t_R FILLER_24_244 ();
 DECAPx10_ASAP7_75t_R FILLER_24_266 ();
 DECAPx10_ASAP7_75t_R FILLER_24_288 ();
 DECAPx10_ASAP7_75t_R FILLER_24_310 ();
 DECAPx10_ASAP7_75t_R FILLER_24_332 ();
 DECAPx10_ASAP7_75t_R FILLER_24_354 ();
 DECAPx10_ASAP7_75t_R FILLER_24_376 ();
 DECAPx10_ASAP7_75t_R FILLER_24_398 ();
 DECAPx10_ASAP7_75t_R FILLER_24_420 ();
 DECAPx6_ASAP7_75t_R FILLER_24_442 ();
 DECAPx2_ASAP7_75t_R FILLER_24_456 ();
 DECAPx10_ASAP7_75t_R FILLER_24_464 ();
 DECAPx10_ASAP7_75t_R FILLER_24_486 ();
 DECAPx10_ASAP7_75t_R FILLER_24_508 ();
 DECAPx10_ASAP7_75t_R FILLER_24_530 ();
 FILLER_ASAP7_75t_R FILLER_24_552 ();
 DECAPx1_ASAP7_75t_R FILLER_24_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_578 ();
 FILLER_ASAP7_75t_R FILLER_24_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_587 ();
 DECAPx1_ASAP7_75t_R FILLER_24_631 ();
 FILLER_ASAP7_75t_R FILLER_24_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_643 ();
 DECAPx6_ASAP7_75t_R FILLER_24_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_667 ();
 DECAPx1_ASAP7_75t_R FILLER_24_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_704 ();
 DECAPx1_ASAP7_75t_R FILLER_24_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_728 ();
 DECAPx2_ASAP7_75t_R FILLER_24_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_752 ();
 FILLER_ASAP7_75t_R FILLER_24_756 ();
 DECAPx1_ASAP7_75t_R FILLER_24_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_776 ();
 DECAPx2_ASAP7_75t_R FILLER_24_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_795 ();
 DECAPx4_ASAP7_75t_R FILLER_24_816 ();
 FILLER_ASAP7_75t_R FILLER_24_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_828 ();
 DECAPx1_ASAP7_75t_R FILLER_24_869 ();
 FILLER_ASAP7_75t_R FILLER_24_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_881 ();
 DECAPx10_ASAP7_75t_R FILLER_24_891 ();
 DECAPx10_ASAP7_75t_R FILLER_24_913 ();
 DECAPx10_ASAP7_75t_R FILLER_24_935 ();
 DECAPx10_ASAP7_75t_R FILLER_24_957 ();
 DECAPx10_ASAP7_75t_R FILLER_24_979 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1353 ();
 DECAPx4_ASAP7_75t_R FILLER_24_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_24_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_25_2 ();
 DECAPx10_ASAP7_75t_R FILLER_25_24 ();
 DECAPx10_ASAP7_75t_R FILLER_25_46 ();
 DECAPx10_ASAP7_75t_R FILLER_25_68 ();
 DECAPx10_ASAP7_75t_R FILLER_25_90 ();
 DECAPx10_ASAP7_75t_R FILLER_25_112 ();
 DECAPx10_ASAP7_75t_R FILLER_25_134 ();
 DECAPx10_ASAP7_75t_R FILLER_25_156 ();
 DECAPx10_ASAP7_75t_R FILLER_25_178 ();
 DECAPx10_ASAP7_75t_R FILLER_25_200 ();
 DECAPx10_ASAP7_75t_R FILLER_25_222 ();
 DECAPx10_ASAP7_75t_R FILLER_25_244 ();
 DECAPx10_ASAP7_75t_R FILLER_25_266 ();
 DECAPx10_ASAP7_75t_R FILLER_25_288 ();
 DECAPx10_ASAP7_75t_R FILLER_25_310 ();
 DECAPx10_ASAP7_75t_R FILLER_25_332 ();
 DECAPx10_ASAP7_75t_R FILLER_25_354 ();
 DECAPx10_ASAP7_75t_R FILLER_25_376 ();
 DECAPx10_ASAP7_75t_R FILLER_25_398 ();
 DECAPx10_ASAP7_75t_R FILLER_25_420 ();
 DECAPx10_ASAP7_75t_R FILLER_25_442 ();
 DECAPx10_ASAP7_75t_R FILLER_25_464 ();
 DECAPx10_ASAP7_75t_R FILLER_25_486 ();
 DECAPx10_ASAP7_75t_R FILLER_25_508 ();
 DECAPx6_ASAP7_75t_R FILLER_25_530 ();
 DECAPx2_ASAP7_75t_R FILLER_25_544 ();
 DECAPx1_ASAP7_75t_R FILLER_25_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_572 ();
 DECAPx4_ASAP7_75t_R FILLER_25_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_597 ();
 FILLER_ASAP7_75t_R FILLER_25_608 ();
 DECAPx2_ASAP7_75t_R FILLER_25_616 ();
 FILLER_ASAP7_75t_R FILLER_25_631 ();
 DECAPx2_ASAP7_75t_R FILLER_25_636 ();
 FILLER_ASAP7_75t_R FILLER_25_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_644 ();
 DECAPx2_ASAP7_75t_R FILLER_25_651 ();
 DECAPx1_ASAP7_75t_R FILLER_25_660 ();
 FILLER_ASAP7_75t_R FILLER_25_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_684 ();
 DECAPx1_ASAP7_75t_R FILLER_25_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_695 ();
 DECAPx2_ASAP7_75t_R FILLER_25_699 ();
 FILLER_ASAP7_75t_R FILLER_25_705 ();
 DECAPx6_ASAP7_75t_R FILLER_25_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_735 ();
 DECAPx1_ASAP7_75t_R FILLER_25_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_746 ();
 FILLER_ASAP7_75t_R FILLER_25_750 ();
 DECAPx2_ASAP7_75t_R FILLER_25_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_761 ();
 DECAPx2_ASAP7_75t_R FILLER_25_765 ();
 DECAPx4_ASAP7_75t_R FILLER_25_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_798 ();
 DECAPx2_ASAP7_75t_R FILLER_25_811 ();
 DECAPx1_ASAP7_75t_R FILLER_25_840 ();
 DECAPx1_ASAP7_75t_R FILLER_25_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_865 ();
 DECAPx1_ASAP7_75t_R FILLER_25_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_873 ();
 FILLER_ASAP7_75t_R FILLER_25_883 ();
 DECAPx10_ASAP7_75t_R FILLER_25_892 ();
 DECAPx4_ASAP7_75t_R FILLER_25_914 ();
 DECAPx10_ASAP7_75t_R FILLER_25_926 ();
 DECAPx10_ASAP7_75t_R FILLER_25_948 ();
 DECAPx10_ASAP7_75t_R FILLER_25_970 ();
 DECAPx10_ASAP7_75t_R FILLER_25_992 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_26_2 ();
 DECAPx10_ASAP7_75t_R FILLER_26_24 ();
 DECAPx10_ASAP7_75t_R FILLER_26_46 ();
 DECAPx10_ASAP7_75t_R FILLER_26_68 ();
 DECAPx10_ASAP7_75t_R FILLER_26_90 ();
 DECAPx10_ASAP7_75t_R FILLER_26_112 ();
 DECAPx10_ASAP7_75t_R FILLER_26_134 ();
 DECAPx10_ASAP7_75t_R FILLER_26_156 ();
 DECAPx10_ASAP7_75t_R FILLER_26_178 ();
 DECAPx10_ASAP7_75t_R FILLER_26_200 ();
 DECAPx10_ASAP7_75t_R FILLER_26_222 ();
 DECAPx10_ASAP7_75t_R FILLER_26_244 ();
 DECAPx10_ASAP7_75t_R FILLER_26_266 ();
 DECAPx10_ASAP7_75t_R FILLER_26_288 ();
 DECAPx10_ASAP7_75t_R FILLER_26_310 ();
 DECAPx10_ASAP7_75t_R FILLER_26_332 ();
 DECAPx10_ASAP7_75t_R FILLER_26_354 ();
 DECAPx10_ASAP7_75t_R FILLER_26_376 ();
 DECAPx10_ASAP7_75t_R FILLER_26_398 ();
 DECAPx10_ASAP7_75t_R FILLER_26_420 ();
 DECAPx6_ASAP7_75t_R FILLER_26_442 ();
 DECAPx2_ASAP7_75t_R FILLER_26_456 ();
 DECAPx10_ASAP7_75t_R FILLER_26_464 ();
 DECAPx10_ASAP7_75t_R FILLER_26_486 ();
 DECAPx10_ASAP7_75t_R FILLER_26_508 ();
 DECAPx10_ASAP7_75t_R FILLER_26_530 ();
 DECAPx2_ASAP7_75t_R FILLER_26_552 ();
 DECAPx2_ASAP7_75t_R FILLER_26_573 ();
 FILLER_ASAP7_75t_R FILLER_26_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_581 ();
 DECAPx10_ASAP7_75t_R FILLER_26_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_607 ();
 DECAPx6_ASAP7_75t_R FILLER_26_611 ();
 FILLER_ASAP7_75t_R FILLER_26_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_627 ();
 DECAPx1_ASAP7_75t_R FILLER_26_631 ();
 FILLER_ASAP7_75t_R FILLER_26_655 ();
 DECAPx10_ASAP7_75t_R FILLER_26_671 ();
 FILLER_ASAP7_75t_R FILLER_26_693 ();
 DECAPx1_ASAP7_75t_R FILLER_26_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_705 ();
 DECAPx4_ASAP7_75t_R FILLER_26_709 ();
 FILLER_ASAP7_75t_R FILLER_26_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_721 ();
 FILLER_ASAP7_75t_R FILLER_26_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_755 ();
 DECAPx6_ASAP7_75t_R FILLER_26_759 ();
 FILLER_ASAP7_75t_R FILLER_26_773 ();
 DECAPx6_ASAP7_75t_R FILLER_26_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_813 ();
 DECAPx4_ASAP7_75t_R FILLER_26_817 ();
 FILLER_ASAP7_75t_R FILLER_26_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_850 ();
 DECAPx2_ASAP7_75t_R FILLER_26_854 ();
 FILLER_ASAP7_75t_R FILLER_26_860 ();
 DECAPx1_ASAP7_75t_R FILLER_26_871 ();
 FILLER_ASAP7_75t_R FILLER_26_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_880 ();
 DECAPx10_ASAP7_75t_R FILLER_26_893 ();
 DECAPx10_ASAP7_75t_R FILLER_26_915 ();
 DECAPx10_ASAP7_75t_R FILLER_26_937 ();
 DECAPx10_ASAP7_75t_R FILLER_26_959 ();
 DECAPx10_ASAP7_75t_R FILLER_26_981 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_26_1377 ();
 FILLER_ASAP7_75t_R FILLER_26_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_26_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_27_2 ();
 DECAPx10_ASAP7_75t_R FILLER_27_24 ();
 DECAPx10_ASAP7_75t_R FILLER_27_46 ();
 DECAPx10_ASAP7_75t_R FILLER_27_68 ();
 DECAPx10_ASAP7_75t_R FILLER_27_90 ();
 DECAPx10_ASAP7_75t_R FILLER_27_112 ();
 DECAPx10_ASAP7_75t_R FILLER_27_134 ();
 DECAPx10_ASAP7_75t_R FILLER_27_156 ();
 DECAPx10_ASAP7_75t_R FILLER_27_178 ();
 DECAPx10_ASAP7_75t_R FILLER_27_200 ();
 DECAPx10_ASAP7_75t_R FILLER_27_222 ();
 DECAPx10_ASAP7_75t_R FILLER_27_244 ();
 DECAPx10_ASAP7_75t_R FILLER_27_266 ();
 DECAPx10_ASAP7_75t_R FILLER_27_288 ();
 DECAPx10_ASAP7_75t_R FILLER_27_310 ();
 DECAPx10_ASAP7_75t_R FILLER_27_332 ();
 DECAPx10_ASAP7_75t_R FILLER_27_354 ();
 DECAPx10_ASAP7_75t_R FILLER_27_376 ();
 DECAPx10_ASAP7_75t_R FILLER_27_398 ();
 DECAPx10_ASAP7_75t_R FILLER_27_420 ();
 DECAPx10_ASAP7_75t_R FILLER_27_442 ();
 DECAPx10_ASAP7_75t_R FILLER_27_464 ();
 DECAPx10_ASAP7_75t_R FILLER_27_486 ();
 DECAPx10_ASAP7_75t_R FILLER_27_508 ();
 DECAPx10_ASAP7_75t_R FILLER_27_530 ();
 DECAPx4_ASAP7_75t_R FILLER_27_552 ();
 DECAPx2_ASAP7_75t_R FILLER_27_565 ();
 FILLER_ASAP7_75t_R FILLER_27_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_573 ();
 FILLER_ASAP7_75t_R FILLER_27_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_579 ();
 FILLER_ASAP7_75t_R FILLER_27_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_596 ();
 FILLER_ASAP7_75t_R FILLER_27_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_618 ();
 DECAPx1_ASAP7_75t_R FILLER_27_639 ();
 FILLER_ASAP7_75t_R FILLER_27_657 ();
 DECAPx4_ASAP7_75t_R FILLER_27_673 ();
 DECAPx1_ASAP7_75t_R FILLER_27_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_693 ();
 DECAPx2_ASAP7_75t_R FILLER_27_708 ();
 DECAPx4_ASAP7_75t_R FILLER_27_723 ();
 DECAPx10_ASAP7_75t_R FILLER_27_736 ();
 DECAPx10_ASAP7_75t_R FILLER_27_772 ();
 DECAPx2_ASAP7_75t_R FILLER_27_800 ();
 FILLER_ASAP7_75t_R FILLER_27_806 ();
 DECAPx6_ASAP7_75t_R FILLER_27_811 ();
 DECAPx1_ASAP7_75t_R FILLER_27_825 ();
 DECAPx10_ASAP7_75t_R FILLER_27_832 ();
 FILLER_ASAP7_75t_R FILLER_27_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_859 ();
 DECAPx6_ASAP7_75t_R FILLER_27_863 ();
 DECAPx1_ASAP7_75t_R FILLER_27_877 ();
 DECAPx10_ASAP7_75t_R FILLER_27_888 ();
 DECAPx6_ASAP7_75t_R FILLER_27_910 ();
 DECAPx10_ASAP7_75t_R FILLER_27_926 ();
 DECAPx10_ASAP7_75t_R FILLER_27_948 ();
 DECAPx10_ASAP7_75t_R FILLER_27_970 ();
 DECAPx10_ASAP7_75t_R FILLER_27_992 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_27_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_28_24 ();
 DECAPx10_ASAP7_75t_R FILLER_28_46 ();
 DECAPx10_ASAP7_75t_R FILLER_28_68 ();
 DECAPx10_ASAP7_75t_R FILLER_28_90 ();
 DECAPx10_ASAP7_75t_R FILLER_28_112 ();
 DECAPx10_ASAP7_75t_R FILLER_28_134 ();
 DECAPx10_ASAP7_75t_R FILLER_28_156 ();
 DECAPx10_ASAP7_75t_R FILLER_28_178 ();
 DECAPx10_ASAP7_75t_R FILLER_28_200 ();
 DECAPx10_ASAP7_75t_R FILLER_28_222 ();
 DECAPx10_ASAP7_75t_R FILLER_28_244 ();
 DECAPx10_ASAP7_75t_R FILLER_28_266 ();
 DECAPx10_ASAP7_75t_R FILLER_28_288 ();
 DECAPx10_ASAP7_75t_R FILLER_28_310 ();
 DECAPx10_ASAP7_75t_R FILLER_28_332 ();
 DECAPx10_ASAP7_75t_R FILLER_28_354 ();
 DECAPx10_ASAP7_75t_R FILLER_28_376 ();
 DECAPx10_ASAP7_75t_R FILLER_28_398 ();
 DECAPx10_ASAP7_75t_R FILLER_28_420 ();
 DECAPx6_ASAP7_75t_R FILLER_28_442 ();
 DECAPx2_ASAP7_75t_R FILLER_28_456 ();
 DECAPx10_ASAP7_75t_R FILLER_28_464 ();
 DECAPx10_ASAP7_75t_R FILLER_28_486 ();
 DECAPx10_ASAP7_75t_R FILLER_28_508 ();
 DECAPx4_ASAP7_75t_R FILLER_28_530 ();
 FILLER_ASAP7_75t_R FILLER_28_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_542 ();
 DECAPx10_ASAP7_75t_R FILLER_28_563 ();
 DECAPx1_ASAP7_75t_R FILLER_28_585 ();
 DECAPx4_ASAP7_75t_R FILLER_28_609 ();
 FILLER_ASAP7_75t_R FILLER_28_619 ();
 DECAPx10_ASAP7_75t_R FILLER_28_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_653 ();
 DECAPx4_ASAP7_75t_R FILLER_28_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_667 ();
 DECAPx4_ASAP7_75t_R FILLER_28_671 ();
 FILLER_ASAP7_75t_R FILLER_28_681 ();
 FILLER_ASAP7_75t_R FILLER_28_701 ();
 DECAPx1_ASAP7_75t_R FILLER_28_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_742 ();
 DECAPx6_ASAP7_75t_R FILLER_28_769 ();
 DECAPx2_ASAP7_75t_R FILLER_28_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_789 ();
 DECAPx4_ASAP7_75t_R FILLER_28_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_815 ();
 DECAPx2_ASAP7_75t_R FILLER_28_834 ();
 DECAPx4_ASAP7_75t_R FILLER_28_857 ();
 FILLER_ASAP7_75t_R FILLER_28_867 ();
 DECAPx10_ASAP7_75t_R FILLER_28_895 ();
 DECAPx10_ASAP7_75t_R FILLER_28_917 ();
 DECAPx10_ASAP7_75t_R FILLER_28_939 ();
 DECAPx10_ASAP7_75t_R FILLER_28_961 ();
 DECAPx10_ASAP7_75t_R FILLER_28_983 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_28_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_29_2 ();
 DECAPx10_ASAP7_75t_R FILLER_29_24 ();
 DECAPx10_ASAP7_75t_R FILLER_29_46 ();
 DECAPx10_ASAP7_75t_R FILLER_29_68 ();
 DECAPx10_ASAP7_75t_R FILLER_29_90 ();
 DECAPx10_ASAP7_75t_R FILLER_29_112 ();
 DECAPx10_ASAP7_75t_R FILLER_29_134 ();
 DECAPx10_ASAP7_75t_R FILLER_29_156 ();
 DECAPx10_ASAP7_75t_R FILLER_29_178 ();
 DECAPx10_ASAP7_75t_R FILLER_29_200 ();
 DECAPx10_ASAP7_75t_R FILLER_29_222 ();
 DECAPx10_ASAP7_75t_R FILLER_29_244 ();
 DECAPx10_ASAP7_75t_R FILLER_29_266 ();
 DECAPx10_ASAP7_75t_R FILLER_29_288 ();
 DECAPx10_ASAP7_75t_R FILLER_29_310 ();
 DECAPx10_ASAP7_75t_R FILLER_29_332 ();
 DECAPx10_ASAP7_75t_R FILLER_29_354 ();
 DECAPx10_ASAP7_75t_R FILLER_29_376 ();
 DECAPx10_ASAP7_75t_R FILLER_29_398 ();
 DECAPx10_ASAP7_75t_R FILLER_29_420 ();
 DECAPx10_ASAP7_75t_R FILLER_29_442 ();
 DECAPx10_ASAP7_75t_R FILLER_29_464 ();
 DECAPx10_ASAP7_75t_R FILLER_29_486 ();
 DECAPx10_ASAP7_75t_R FILLER_29_508 ();
 DECAPx4_ASAP7_75t_R FILLER_29_530 ();
 FILLER_ASAP7_75t_R FILLER_29_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_542 ();
 DECAPx2_ASAP7_75t_R FILLER_29_561 ();
 DECAPx2_ASAP7_75t_R FILLER_29_599 ();
 FILLER_ASAP7_75t_R FILLER_29_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_607 ();
 FILLER_ASAP7_75t_R FILLER_29_621 ();
 DECAPx4_ASAP7_75t_R FILLER_29_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_647 ();
 DECAPx6_ASAP7_75t_R FILLER_29_654 ();
 DECAPx1_ASAP7_75t_R FILLER_29_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_672 ();
 FILLER_ASAP7_75t_R FILLER_29_691 ();
 DECAPx2_ASAP7_75t_R FILLER_29_713 ();
 DECAPx1_ASAP7_75t_R FILLER_29_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_726 ();
 FILLER_ASAP7_75t_R FILLER_29_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_732 ();
 DECAPx10_ASAP7_75t_R FILLER_29_736 ();
 DECAPx1_ASAP7_75t_R FILLER_29_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_825 ();
 DECAPx2_ASAP7_75t_R FILLER_29_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_846 ();
 DECAPx2_ASAP7_75t_R FILLER_29_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_873 ();
 DECAPx10_ASAP7_75t_R FILLER_29_889 ();
 DECAPx4_ASAP7_75t_R FILLER_29_911 ();
 FILLER_ASAP7_75t_R FILLER_29_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_923 ();
 DECAPx10_ASAP7_75t_R FILLER_29_926 ();
 DECAPx10_ASAP7_75t_R FILLER_29_948 ();
 DECAPx10_ASAP7_75t_R FILLER_29_970 ();
 DECAPx10_ASAP7_75t_R FILLER_29_992 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_29_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1347 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_30_2 ();
 DECAPx10_ASAP7_75t_R FILLER_30_24 ();
 DECAPx10_ASAP7_75t_R FILLER_30_46 ();
 DECAPx10_ASAP7_75t_R FILLER_30_68 ();
 DECAPx10_ASAP7_75t_R FILLER_30_90 ();
 DECAPx10_ASAP7_75t_R FILLER_30_112 ();
 DECAPx10_ASAP7_75t_R FILLER_30_134 ();
 DECAPx10_ASAP7_75t_R FILLER_30_156 ();
 DECAPx10_ASAP7_75t_R FILLER_30_178 ();
 DECAPx10_ASAP7_75t_R FILLER_30_200 ();
 DECAPx10_ASAP7_75t_R FILLER_30_222 ();
 DECAPx10_ASAP7_75t_R FILLER_30_244 ();
 DECAPx10_ASAP7_75t_R FILLER_30_266 ();
 DECAPx10_ASAP7_75t_R FILLER_30_288 ();
 DECAPx10_ASAP7_75t_R FILLER_30_310 ();
 DECAPx10_ASAP7_75t_R FILLER_30_332 ();
 DECAPx10_ASAP7_75t_R FILLER_30_354 ();
 DECAPx10_ASAP7_75t_R FILLER_30_376 ();
 DECAPx10_ASAP7_75t_R FILLER_30_398 ();
 DECAPx10_ASAP7_75t_R FILLER_30_420 ();
 DECAPx6_ASAP7_75t_R FILLER_30_442 ();
 DECAPx2_ASAP7_75t_R FILLER_30_456 ();
 DECAPx10_ASAP7_75t_R FILLER_30_464 ();
 DECAPx10_ASAP7_75t_R FILLER_30_486 ();
 DECAPx10_ASAP7_75t_R FILLER_30_508 ();
 DECAPx6_ASAP7_75t_R FILLER_30_530 ();
 FILLER_ASAP7_75t_R FILLER_30_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_546 ();
 DECAPx2_ASAP7_75t_R FILLER_30_579 ();
 FILLER_ASAP7_75t_R FILLER_30_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_587 ();
 DECAPx1_ASAP7_75t_R FILLER_30_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_601 ();
 FILLER_ASAP7_75t_R FILLER_30_616 ();
 FILLER_ASAP7_75t_R FILLER_30_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_623 ();
 DECAPx1_ASAP7_75t_R FILLER_30_648 ();
 DECAPx1_ASAP7_75t_R FILLER_30_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_674 ();
 DECAPx4_ASAP7_75t_R FILLER_30_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_703 ();
 DECAPx2_ASAP7_75t_R FILLER_30_707 ();
 FILLER_ASAP7_75t_R FILLER_30_713 ();
 DECAPx2_ASAP7_75t_R FILLER_30_743 ();
 FILLER_ASAP7_75t_R FILLER_30_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_751 ();
 DECAPx1_ASAP7_75t_R FILLER_30_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_765 ();
 DECAPx10_ASAP7_75t_R FILLER_30_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_811 ();
 DECAPx1_ASAP7_75t_R FILLER_30_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_833 ();
 DECAPx1_ASAP7_75t_R FILLER_30_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_845 ();
 FILLER_ASAP7_75t_R FILLER_30_858 ();
 DECAPx6_ASAP7_75t_R FILLER_30_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_897 ();
 DECAPx1_ASAP7_75t_R FILLER_30_904 ();
 DECAPx1_ASAP7_75t_R FILLER_30_911 ();
 DECAPx10_ASAP7_75t_R FILLER_30_959 ();
 DECAPx10_ASAP7_75t_R FILLER_30_981 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1135 ();
 DECAPx6_ASAP7_75t_R FILLER_30_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_30_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_30_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_30_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_30_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_31_2 ();
 DECAPx10_ASAP7_75t_R FILLER_31_24 ();
 DECAPx10_ASAP7_75t_R FILLER_31_46 ();
 DECAPx10_ASAP7_75t_R FILLER_31_68 ();
 DECAPx10_ASAP7_75t_R FILLER_31_90 ();
 DECAPx10_ASAP7_75t_R FILLER_31_112 ();
 DECAPx10_ASAP7_75t_R FILLER_31_134 ();
 DECAPx10_ASAP7_75t_R FILLER_31_156 ();
 DECAPx10_ASAP7_75t_R FILLER_31_178 ();
 DECAPx10_ASAP7_75t_R FILLER_31_200 ();
 DECAPx10_ASAP7_75t_R FILLER_31_222 ();
 DECAPx10_ASAP7_75t_R FILLER_31_244 ();
 DECAPx10_ASAP7_75t_R FILLER_31_266 ();
 DECAPx10_ASAP7_75t_R FILLER_31_288 ();
 DECAPx10_ASAP7_75t_R FILLER_31_310 ();
 DECAPx10_ASAP7_75t_R FILLER_31_332 ();
 DECAPx10_ASAP7_75t_R FILLER_31_354 ();
 DECAPx10_ASAP7_75t_R FILLER_31_376 ();
 DECAPx10_ASAP7_75t_R FILLER_31_398 ();
 DECAPx10_ASAP7_75t_R FILLER_31_420 ();
 DECAPx10_ASAP7_75t_R FILLER_31_442 ();
 DECAPx10_ASAP7_75t_R FILLER_31_464 ();
 DECAPx10_ASAP7_75t_R FILLER_31_486 ();
 DECAPx10_ASAP7_75t_R FILLER_31_508 ();
 DECAPx10_ASAP7_75t_R FILLER_31_530 ();
 DECAPx2_ASAP7_75t_R FILLER_31_552 ();
 DECAPx1_ASAP7_75t_R FILLER_31_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_565 ();
 DECAPx2_ASAP7_75t_R FILLER_31_576 ();
 FILLER_ASAP7_75t_R FILLER_31_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_584 ();
 DECAPx4_ASAP7_75t_R FILLER_31_588 ();
 FILLER_ASAP7_75t_R FILLER_31_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_600 ();
 DECAPx10_ASAP7_75t_R FILLER_31_604 ();
 DECAPx1_ASAP7_75t_R FILLER_31_626 ();
 DECAPx1_ASAP7_75t_R FILLER_31_633 ();
 DECAPx10_ASAP7_75t_R FILLER_31_640 ();
 DECAPx1_ASAP7_75t_R FILLER_31_662 ();
 FILLER_ASAP7_75t_R FILLER_31_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_671 ();
 DECAPx2_ASAP7_75t_R FILLER_31_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_695 ();
 DECAPx4_ASAP7_75t_R FILLER_31_699 ();
 FILLER_ASAP7_75t_R FILLER_31_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_711 ();
 DECAPx10_ASAP7_75t_R FILLER_31_726 ();
 DECAPx2_ASAP7_75t_R FILLER_31_748 ();
 FILLER_ASAP7_75t_R FILLER_31_754 ();
 FILLER_ASAP7_75t_R FILLER_31_777 ();
 DECAPx6_ASAP7_75t_R FILLER_31_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_799 ();
 DECAPx4_ASAP7_75t_R FILLER_31_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_826 ();
 FILLER_ASAP7_75t_R FILLER_31_830 ();
 FILLER_ASAP7_75t_R FILLER_31_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_843 ();
 FILLER_ASAP7_75t_R FILLER_31_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_849 ();
 DECAPx2_ASAP7_75t_R FILLER_31_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_865 ();
 DECAPx10_ASAP7_75t_R FILLER_31_869 ();
 FILLER_ASAP7_75t_R FILLER_31_891 ();
 DECAPx1_ASAP7_75t_R FILLER_31_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_923 ();
 DECAPx4_ASAP7_75t_R FILLER_31_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_954 ();
 DECAPx10_ASAP7_75t_R FILLER_31_958 ();
 DECAPx10_ASAP7_75t_R FILLER_31_980 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1112 ();
 FILLER_ASAP7_75t_R FILLER_31_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1127 ();
 FILLER_ASAP7_75t_R FILLER_31_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1383 ();
 FILLER_ASAP7_75t_R FILLER_31_1389 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_32_2 ();
 DECAPx10_ASAP7_75t_R FILLER_32_24 ();
 DECAPx10_ASAP7_75t_R FILLER_32_46 ();
 DECAPx10_ASAP7_75t_R FILLER_32_68 ();
 DECAPx10_ASAP7_75t_R FILLER_32_90 ();
 DECAPx10_ASAP7_75t_R FILLER_32_112 ();
 DECAPx10_ASAP7_75t_R FILLER_32_134 ();
 DECAPx10_ASAP7_75t_R FILLER_32_156 ();
 DECAPx10_ASAP7_75t_R FILLER_32_178 ();
 DECAPx10_ASAP7_75t_R FILLER_32_200 ();
 DECAPx10_ASAP7_75t_R FILLER_32_222 ();
 DECAPx10_ASAP7_75t_R FILLER_32_244 ();
 DECAPx10_ASAP7_75t_R FILLER_32_266 ();
 DECAPx10_ASAP7_75t_R FILLER_32_288 ();
 DECAPx10_ASAP7_75t_R FILLER_32_310 ();
 DECAPx10_ASAP7_75t_R FILLER_32_332 ();
 DECAPx10_ASAP7_75t_R FILLER_32_354 ();
 DECAPx10_ASAP7_75t_R FILLER_32_376 ();
 DECAPx10_ASAP7_75t_R FILLER_32_398 ();
 DECAPx10_ASAP7_75t_R FILLER_32_420 ();
 DECAPx6_ASAP7_75t_R FILLER_32_442 ();
 DECAPx2_ASAP7_75t_R FILLER_32_456 ();
 DECAPx10_ASAP7_75t_R FILLER_32_464 ();
 DECAPx10_ASAP7_75t_R FILLER_32_486 ();
 DECAPx6_ASAP7_75t_R FILLER_32_508 ();
 DECAPx2_ASAP7_75t_R FILLER_32_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_539 ();
 DECAPx2_ASAP7_75t_R FILLER_32_558 ();
 FILLER_ASAP7_75t_R FILLER_32_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_566 ();
 DECAPx6_ASAP7_75t_R FILLER_32_573 ();
 FILLER_ASAP7_75t_R FILLER_32_587 ();
 DECAPx2_ASAP7_75t_R FILLER_32_598 ();
 FILLER_ASAP7_75t_R FILLER_32_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_606 ();
 DECAPx1_ASAP7_75t_R FILLER_32_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_614 ();
 DECAPx4_ASAP7_75t_R FILLER_32_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_628 ();
 DECAPx4_ASAP7_75t_R FILLER_32_635 ();
 FILLER_ASAP7_75t_R FILLER_32_648 ();
 DECAPx2_ASAP7_75t_R FILLER_32_662 ();
 FILLER_ASAP7_75t_R FILLER_32_668 ();
 DECAPx2_ASAP7_75t_R FILLER_32_679 ();
 FILLER_ASAP7_75t_R FILLER_32_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_687 ();
 DECAPx4_ASAP7_75t_R FILLER_32_702 ();
 FILLER_ASAP7_75t_R FILLER_32_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_727 ();
 DECAPx1_ASAP7_75t_R FILLER_32_731 ();
 DECAPx4_ASAP7_75t_R FILLER_32_749 ();
 FILLER_ASAP7_75t_R FILLER_32_759 ();
 DECAPx1_ASAP7_75t_R FILLER_32_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_782 ();
 DECAPx6_ASAP7_75t_R FILLER_32_818 ();
 DECAPx1_ASAP7_75t_R FILLER_32_832 ();
 DECAPx2_ASAP7_75t_R FILLER_32_839 ();
 FILLER_ASAP7_75t_R FILLER_32_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_847 ();
 DECAPx4_ASAP7_75t_R FILLER_32_857 ();
 FILLER_ASAP7_75t_R FILLER_32_867 ();
 FILLER_ASAP7_75t_R FILLER_32_875 ();
 DECAPx1_ASAP7_75t_R FILLER_32_880 ();
 DECAPx2_ASAP7_75t_R FILLER_32_910 ();
 FILLER_ASAP7_75t_R FILLER_32_916 ();
 FILLER_ASAP7_75t_R FILLER_32_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_933 ();
 DECAPx10_ASAP7_75t_R FILLER_32_966 ();
 DECAPx10_ASAP7_75t_R FILLER_32_988 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1054 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1090 ();
 FILLER_ASAP7_75t_R FILLER_32_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1111 ();
 DECAPx4_ASAP7_75t_R FILLER_32_1132 ();
 FILLER_ASAP7_75t_R FILLER_32_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1144 ();
 FILLER_ASAP7_75t_R FILLER_32_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1206 ();
 FILLER_ASAP7_75t_R FILLER_32_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1214 ();
 DECAPx4_ASAP7_75t_R FILLER_32_1228 ();
 FILLER_ASAP7_75t_R FILLER_32_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_32_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_32_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_33_2 ();
 DECAPx10_ASAP7_75t_R FILLER_33_24 ();
 DECAPx10_ASAP7_75t_R FILLER_33_46 ();
 DECAPx10_ASAP7_75t_R FILLER_33_68 ();
 DECAPx10_ASAP7_75t_R FILLER_33_90 ();
 DECAPx10_ASAP7_75t_R FILLER_33_112 ();
 DECAPx10_ASAP7_75t_R FILLER_33_134 ();
 DECAPx10_ASAP7_75t_R FILLER_33_156 ();
 DECAPx10_ASAP7_75t_R FILLER_33_178 ();
 DECAPx10_ASAP7_75t_R FILLER_33_200 ();
 DECAPx10_ASAP7_75t_R FILLER_33_222 ();
 DECAPx10_ASAP7_75t_R FILLER_33_244 ();
 DECAPx10_ASAP7_75t_R FILLER_33_266 ();
 DECAPx10_ASAP7_75t_R FILLER_33_288 ();
 DECAPx10_ASAP7_75t_R FILLER_33_310 ();
 DECAPx10_ASAP7_75t_R FILLER_33_332 ();
 DECAPx10_ASAP7_75t_R FILLER_33_354 ();
 DECAPx10_ASAP7_75t_R FILLER_33_376 ();
 DECAPx10_ASAP7_75t_R FILLER_33_398 ();
 DECAPx10_ASAP7_75t_R FILLER_33_420 ();
 DECAPx10_ASAP7_75t_R FILLER_33_442 ();
 DECAPx10_ASAP7_75t_R FILLER_33_464 ();
 DECAPx10_ASAP7_75t_R FILLER_33_486 ();
 DECAPx10_ASAP7_75t_R FILLER_33_508 ();
 DECAPx6_ASAP7_75t_R FILLER_33_530 ();
 DECAPx2_ASAP7_75t_R FILLER_33_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_570 ();
 DECAPx1_ASAP7_75t_R FILLER_33_580 ();
 FILLER_ASAP7_75t_R FILLER_33_607 ();
 DECAPx2_ASAP7_75t_R FILLER_33_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_664 ();
 DECAPx2_ASAP7_75t_R FILLER_33_679 ();
 FILLER_ASAP7_75t_R FILLER_33_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_687 ();
 DECAPx2_ASAP7_75t_R FILLER_33_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_700 ();
 DECAPx4_ASAP7_75t_R FILLER_33_704 ();
 FILLER_ASAP7_75t_R FILLER_33_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_736 ();
 DECAPx6_ASAP7_75t_R FILLER_33_765 ();
 FILLER_ASAP7_75t_R FILLER_33_779 ();
 DECAPx1_ASAP7_75t_R FILLER_33_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_813 ();
 FILLER_ASAP7_75t_R FILLER_33_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_825 ();
 DECAPx1_ASAP7_75t_R FILLER_33_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_843 ();
 DECAPx1_ASAP7_75t_R FILLER_33_847 ();
 DECAPx2_ASAP7_75t_R FILLER_33_854 ();
 FILLER_ASAP7_75t_R FILLER_33_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_888 ();
 DECAPx6_ASAP7_75t_R FILLER_33_906 ();
 DECAPx1_ASAP7_75t_R FILLER_33_920 ();
 DECAPx2_ASAP7_75t_R FILLER_33_926 ();
 FILLER_ASAP7_75t_R FILLER_33_932 ();
 DECAPx2_ASAP7_75t_R FILLER_33_951 ();
 FILLER_ASAP7_75t_R FILLER_33_957 ();
 DECAPx10_ASAP7_75t_R FILLER_33_962 ();
 DECAPx10_ASAP7_75t_R FILLER_33_984 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_33_1050 ();
 DECAPx6_ASAP7_75t_R FILLER_33_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_33_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1156 ();
 FILLER_ASAP7_75t_R FILLER_33_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1164 ();
 DECAPx6_ASAP7_75t_R FILLER_33_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1192 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1383 ();
 FILLER_ASAP7_75t_R FILLER_33_1389 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_34_2 ();
 DECAPx10_ASAP7_75t_R FILLER_34_24 ();
 DECAPx10_ASAP7_75t_R FILLER_34_46 ();
 DECAPx10_ASAP7_75t_R FILLER_34_68 ();
 DECAPx10_ASAP7_75t_R FILLER_34_90 ();
 DECAPx10_ASAP7_75t_R FILLER_34_112 ();
 DECAPx10_ASAP7_75t_R FILLER_34_134 ();
 DECAPx10_ASAP7_75t_R FILLER_34_156 ();
 DECAPx10_ASAP7_75t_R FILLER_34_178 ();
 DECAPx10_ASAP7_75t_R FILLER_34_200 ();
 DECAPx10_ASAP7_75t_R FILLER_34_222 ();
 DECAPx10_ASAP7_75t_R FILLER_34_244 ();
 DECAPx10_ASAP7_75t_R FILLER_34_266 ();
 DECAPx10_ASAP7_75t_R FILLER_34_288 ();
 DECAPx10_ASAP7_75t_R FILLER_34_310 ();
 DECAPx10_ASAP7_75t_R FILLER_34_332 ();
 DECAPx10_ASAP7_75t_R FILLER_34_354 ();
 DECAPx10_ASAP7_75t_R FILLER_34_376 ();
 DECAPx10_ASAP7_75t_R FILLER_34_398 ();
 DECAPx10_ASAP7_75t_R FILLER_34_420 ();
 DECAPx6_ASAP7_75t_R FILLER_34_442 ();
 DECAPx2_ASAP7_75t_R FILLER_34_456 ();
 DECAPx10_ASAP7_75t_R FILLER_34_464 ();
 DECAPx10_ASAP7_75t_R FILLER_34_486 ();
 DECAPx6_ASAP7_75t_R FILLER_34_508 ();
 DECAPx2_ASAP7_75t_R FILLER_34_522 ();
 DECAPx1_ASAP7_75t_R FILLER_34_546 ();
 DECAPx1_ASAP7_75t_R FILLER_34_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_588 ();
 DECAPx1_ASAP7_75t_R FILLER_34_603 ();
 FILLER_ASAP7_75t_R FILLER_34_621 ();
 DECAPx2_ASAP7_75t_R FILLER_34_640 ();
 FILLER_ASAP7_75t_R FILLER_34_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_648 ();
 DECAPx2_ASAP7_75t_R FILLER_34_663 ();
 FILLER_ASAP7_75t_R FILLER_34_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_712 ();
 DECAPx6_ASAP7_75t_R FILLER_34_719 ();
 DECAPx1_ASAP7_75t_R FILLER_34_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_737 ();
 DECAPx1_ASAP7_75t_R FILLER_34_744 ();
 DECAPx2_ASAP7_75t_R FILLER_34_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_760 ();
 DECAPx10_ASAP7_75t_R FILLER_34_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_796 ();
 DECAPx6_ASAP7_75t_R FILLER_34_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_814 ();
 FILLER_ASAP7_75t_R FILLER_34_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_829 ();
 FILLER_ASAP7_75t_R FILLER_34_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_835 ();
 DECAPx4_ASAP7_75t_R FILLER_34_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_855 ();
 DECAPx6_ASAP7_75t_R FILLER_34_882 ();
 FILLER_ASAP7_75t_R FILLER_34_896 ();
 FILLER_ASAP7_75t_R FILLER_34_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_903 ();
 FILLER_ASAP7_75t_R FILLER_34_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_920 ();
 DECAPx10_ASAP7_75t_R FILLER_34_971 ();
 DECAPx10_ASAP7_75t_R FILLER_34_993 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_34_1037 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1077 ();
 FILLER_ASAP7_75t_R FILLER_34_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1110 ();
 FILLER_ASAP7_75t_R FILLER_34_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1118 ();
 DECAPx1_ASAP7_75t_R FILLER_34_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1136 ();
 FILLER_ASAP7_75t_R FILLER_34_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1178 ();
 DECAPx4_ASAP7_75t_R FILLER_34_1205 ();
 FILLER_ASAP7_75t_R FILLER_34_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_34_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_34_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_35_2 ();
 DECAPx10_ASAP7_75t_R FILLER_35_24 ();
 DECAPx10_ASAP7_75t_R FILLER_35_46 ();
 DECAPx10_ASAP7_75t_R FILLER_35_68 ();
 DECAPx10_ASAP7_75t_R FILLER_35_90 ();
 DECAPx10_ASAP7_75t_R FILLER_35_112 ();
 DECAPx10_ASAP7_75t_R FILLER_35_134 ();
 DECAPx10_ASAP7_75t_R FILLER_35_156 ();
 DECAPx10_ASAP7_75t_R FILLER_35_178 ();
 DECAPx10_ASAP7_75t_R FILLER_35_200 ();
 DECAPx10_ASAP7_75t_R FILLER_35_222 ();
 DECAPx10_ASAP7_75t_R FILLER_35_244 ();
 DECAPx10_ASAP7_75t_R FILLER_35_266 ();
 DECAPx10_ASAP7_75t_R FILLER_35_288 ();
 DECAPx10_ASAP7_75t_R FILLER_35_310 ();
 DECAPx10_ASAP7_75t_R FILLER_35_332 ();
 DECAPx10_ASAP7_75t_R FILLER_35_354 ();
 DECAPx10_ASAP7_75t_R FILLER_35_376 ();
 DECAPx10_ASAP7_75t_R FILLER_35_398 ();
 DECAPx10_ASAP7_75t_R FILLER_35_420 ();
 DECAPx10_ASAP7_75t_R FILLER_35_442 ();
 DECAPx10_ASAP7_75t_R FILLER_35_464 ();
 DECAPx10_ASAP7_75t_R FILLER_35_486 ();
 DECAPx10_ASAP7_75t_R FILLER_35_508 ();
 DECAPx6_ASAP7_75t_R FILLER_35_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_544 ();
 DECAPx4_ASAP7_75t_R FILLER_35_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_571 ();
 DECAPx1_ASAP7_75t_R FILLER_35_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_590 ();
 DECAPx4_ASAP7_75t_R FILLER_35_597 ();
 FILLER_ASAP7_75t_R FILLER_35_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_609 ();
 DECAPx2_ASAP7_75t_R FILLER_35_613 ();
 DECAPx2_ASAP7_75t_R FILLER_35_622 ();
 DECAPx4_ASAP7_75t_R FILLER_35_642 ();
 FILLER_ASAP7_75t_R FILLER_35_652 ();
 DECAPx2_ASAP7_75t_R FILLER_35_657 ();
 FILLER_ASAP7_75t_R FILLER_35_663 ();
 DECAPx6_ASAP7_75t_R FILLER_35_668 ();
 FILLER_ASAP7_75t_R FILLER_35_682 ();
 DECAPx2_ASAP7_75t_R FILLER_35_696 ();
 DECAPx2_ASAP7_75t_R FILLER_35_716 ();
 FILLER_ASAP7_75t_R FILLER_35_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_734 ();
 DECAPx2_ASAP7_75t_R FILLER_35_752 ();
 FILLER_ASAP7_75t_R FILLER_35_772 ();
 FILLER_ASAP7_75t_R FILLER_35_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_785 ();
 DECAPx2_ASAP7_75t_R FILLER_35_800 ();
 FILLER_ASAP7_75t_R FILLER_35_806 ();
 DECAPx4_ASAP7_75t_R FILLER_35_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_821 ();
 FILLER_ASAP7_75t_R FILLER_35_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_837 ();
 DECAPx2_ASAP7_75t_R FILLER_35_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_870 ();
 DECAPx2_ASAP7_75t_R FILLER_35_878 ();
 FILLER_ASAP7_75t_R FILLER_35_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_897 ();
 DECAPx2_ASAP7_75t_R FILLER_35_926 ();
 FILLER_ASAP7_75t_R FILLER_35_932 ();
 FILLER_ASAP7_75t_R FILLER_35_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_943 ();
 DECAPx10_ASAP7_75t_R FILLER_35_970 ();
 DECAPx10_ASAP7_75t_R FILLER_35_992 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1014 ();
 DECAPx1_ASAP7_75t_R FILLER_35_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1066 ();
 DECAPx4_ASAP7_75t_R FILLER_35_1074 ();
 FILLER_ASAP7_75t_R FILLER_35_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_35_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1105 ();
 FILLER_ASAP7_75t_R FILLER_35_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1113 ();
 FILLER_ASAP7_75t_R FILLER_35_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1126 ();
 FILLER_ASAP7_75t_R FILLER_35_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1157 ();
 FILLER_ASAP7_75t_R FILLER_35_1163 ();
 FILLER_ASAP7_75t_R FILLER_35_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_35_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1340 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1384 ();
 FILLER_ASAP7_75t_R FILLER_35_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_36_2 ();
 DECAPx10_ASAP7_75t_R FILLER_36_24 ();
 DECAPx10_ASAP7_75t_R FILLER_36_46 ();
 DECAPx10_ASAP7_75t_R FILLER_36_68 ();
 DECAPx10_ASAP7_75t_R FILLER_36_90 ();
 DECAPx10_ASAP7_75t_R FILLER_36_112 ();
 DECAPx10_ASAP7_75t_R FILLER_36_134 ();
 DECAPx10_ASAP7_75t_R FILLER_36_156 ();
 DECAPx10_ASAP7_75t_R FILLER_36_178 ();
 DECAPx10_ASAP7_75t_R FILLER_36_200 ();
 DECAPx10_ASAP7_75t_R FILLER_36_222 ();
 DECAPx10_ASAP7_75t_R FILLER_36_244 ();
 DECAPx10_ASAP7_75t_R FILLER_36_266 ();
 DECAPx10_ASAP7_75t_R FILLER_36_288 ();
 DECAPx10_ASAP7_75t_R FILLER_36_310 ();
 DECAPx10_ASAP7_75t_R FILLER_36_332 ();
 DECAPx10_ASAP7_75t_R FILLER_36_354 ();
 DECAPx10_ASAP7_75t_R FILLER_36_376 ();
 DECAPx10_ASAP7_75t_R FILLER_36_398 ();
 DECAPx10_ASAP7_75t_R FILLER_36_420 ();
 DECAPx6_ASAP7_75t_R FILLER_36_442 ();
 DECAPx2_ASAP7_75t_R FILLER_36_456 ();
 DECAPx10_ASAP7_75t_R FILLER_36_464 ();
 DECAPx10_ASAP7_75t_R FILLER_36_486 ();
 DECAPx10_ASAP7_75t_R FILLER_36_508 ();
 DECAPx10_ASAP7_75t_R FILLER_36_542 ();
 DECAPx2_ASAP7_75t_R FILLER_36_564 ();
 FILLER_ASAP7_75t_R FILLER_36_579 ();
 DECAPx2_ASAP7_75t_R FILLER_36_584 ();
 FILLER_ASAP7_75t_R FILLER_36_590 ();
 FILLER_ASAP7_75t_R FILLER_36_595 ();
 DECAPx2_ASAP7_75t_R FILLER_36_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_606 ();
 FILLER_ASAP7_75t_R FILLER_36_619 ();
 DECAPx6_ASAP7_75t_R FILLER_36_624 ();
 DECAPx1_ASAP7_75t_R FILLER_36_638 ();
 DECAPx2_ASAP7_75t_R FILLER_36_645 ();
 DECAPx1_ASAP7_75t_R FILLER_36_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_658 ();
 DECAPx2_ASAP7_75t_R FILLER_36_662 ();
 DECAPx6_ASAP7_75t_R FILLER_36_682 ();
 DECAPx2_ASAP7_75t_R FILLER_36_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_702 ();
 DECAPx6_ASAP7_75t_R FILLER_36_709 ();
 DECAPx1_ASAP7_75t_R FILLER_36_723 ();
 FILLER_ASAP7_75t_R FILLER_36_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_753 ();
 FILLER_ASAP7_75t_R FILLER_36_766 ();
 FILLER_ASAP7_75t_R FILLER_36_782 ();
 DECAPx1_ASAP7_75t_R FILLER_36_794 ();
 FILLER_ASAP7_75t_R FILLER_36_810 ();
 FILLER_ASAP7_75t_R FILLER_36_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_817 ();
 DECAPx2_ASAP7_75t_R FILLER_36_857 ();
 DECAPx2_ASAP7_75t_R FILLER_36_879 ();
 DECAPx10_ASAP7_75t_R FILLER_36_911 ();
 DECAPx1_ASAP7_75t_R FILLER_36_933 ();
 DECAPx4_ASAP7_75t_R FILLER_36_947 ();
 FILLER_ASAP7_75t_R FILLER_36_957 ();
 DECAPx10_ASAP7_75t_R FILLER_36_962 ();
 DECAPx10_ASAP7_75t_R FILLER_36_984 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_36_1028 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_36_1062 ();
 DECAPx1_ASAP7_75t_R FILLER_36_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1112 ();
 DECAPx1_ASAP7_75t_R FILLER_36_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1138 ();
 DECAPx6_ASAP7_75t_R FILLER_36_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1174 ();
 DECAPx6_ASAP7_75t_R FILLER_36_1186 ();
 FILLER_ASAP7_75t_R FILLER_36_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1209 ();
 FILLER_ASAP7_75t_R FILLER_36_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_36_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_37_2 ();
 DECAPx10_ASAP7_75t_R FILLER_37_24 ();
 DECAPx10_ASAP7_75t_R FILLER_37_46 ();
 DECAPx10_ASAP7_75t_R FILLER_37_68 ();
 DECAPx10_ASAP7_75t_R FILLER_37_90 ();
 DECAPx10_ASAP7_75t_R FILLER_37_112 ();
 DECAPx10_ASAP7_75t_R FILLER_37_134 ();
 DECAPx10_ASAP7_75t_R FILLER_37_156 ();
 DECAPx10_ASAP7_75t_R FILLER_37_178 ();
 DECAPx10_ASAP7_75t_R FILLER_37_200 ();
 DECAPx10_ASAP7_75t_R FILLER_37_222 ();
 DECAPx10_ASAP7_75t_R FILLER_37_244 ();
 DECAPx10_ASAP7_75t_R FILLER_37_266 ();
 DECAPx10_ASAP7_75t_R FILLER_37_288 ();
 DECAPx10_ASAP7_75t_R FILLER_37_310 ();
 DECAPx10_ASAP7_75t_R FILLER_37_332 ();
 DECAPx10_ASAP7_75t_R FILLER_37_354 ();
 DECAPx10_ASAP7_75t_R FILLER_37_376 ();
 DECAPx10_ASAP7_75t_R FILLER_37_398 ();
 DECAPx10_ASAP7_75t_R FILLER_37_420 ();
 DECAPx10_ASAP7_75t_R FILLER_37_442 ();
 DECAPx10_ASAP7_75t_R FILLER_37_464 ();
 DECAPx10_ASAP7_75t_R FILLER_37_486 ();
 DECAPx6_ASAP7_75t_R FILLER_37_508 ();
 DECAPx2_ASAP7_75t_R FILLER_37_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_528 ();
 DECAPx1_ASAP7_75t_R FILLER_37_547 ();
 FILLER_ASAP7_75t_R FILLER_37_555 ();
 FILLER_ASAP7_75t_R FILLER_37_589 ();
 FILLER_ASAP7_75t_R FILLER_37_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_607 ();
 DECAPx4_ASAP7_75t_R FILLER_37_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_632 ();
 DECAPx2_ASAP7_75t_R FILLER_37_636 ();
 FILLER_ASAP7_75t_R FILLER_37_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_644 ();
 FILLER_ASAP7_75t_R FILLER_37_662 ();
 DECAPx1_ASAP7_75t_R FILLER_37_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_695 ();
 DECAPx4_ASAP7_75t_R FILLER_37_713 ();
 DECAPx10_ASAP7_75t_R FILLER_37_726 ();
 DECAPx1_ASAP7_75t_R FILLER_37_748 ();
 FILLER_ASAP7_75t_R FILLER_37_772 ();
 DECAPx2_ASAP7_75t_R FILLER_37_780 ();
 DECAPx1_ASAP7_75t_R FILLER_37_792 ();
 DECAPx1_ASAP7_75t_R FILLER_37_799 ();
 DECAPx10_ASAP7_75t_R FILLER_37_812 ();
 DECAPx10_ASAP7_75t_R FILLER_37_834 ();
 DECAPx6_ASAP7_75t_R FILLER_37_856 ();
 FILLER_ASAP7_75t_R FILLER_37_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_899 ();
 DECAPx6_ASAP7_75t_R FILLER_37_903 ();
 DECAPx2_ASAP7_75t_R FILLER_37_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_923 ();
 DECAPx2_ASAP7_75t_R FILLER_37_926 ();
 FILLER_ASAP7_75t_R FILLER_37_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_934 ();
 DECAPx2_ASAP7_75t_R FILLER_37_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_951 ();
 DECAPx10_ASAP7_75t_R FILLER_37_955 ();
 DECAPx10_ASAP7_75t_R FILLER_37_977 ();
 DECAPx10_ASAP7_75t_R FILLER_37_999 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1021 ();
 DECAPx4_ASAP7_75t_R FILLER_37_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1115 ();
 DECAPx6_ASAP7_75t_R FILLER_37_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1143 ();
 FILLER_ASAP7_75t_R FILLER_37_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1205 ();
 FILLER_ASAP7_75t_R FILLER_37_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1358 ();
 DECAPx10_ASAP7_75t_R FILLER_38_2 ();
 DECAPx10_ASAP7_75t_R FILLER_38_24 ();
 DECAPx10_ASAP7_75t_R FILLER_38_46 ();
 DECAPx10_ASAP7_75t_R FILLER_38_68 ();
 DECAPx10_ASAP7_75t_R FILLER_38_90 ();
 DECAPx10_ASAP7_75t_R FILLER_38_112 ();
 DECAPx10_ASAP7_75t_R FILLER_38_134 ();
 DECAPx10_ASAP7_75t_R FILLER_38_156 ();
 DECAPx10_ASAP7_75t_R FILLER_38_178 ();
 DECAPx10_ASAP7_75t_R FILLER_38_200 ();
 DECAPx10_ASAP7_75t_R FILLER_38_222 ();
 DECAPx10_ASAP7_75t_R FILLER_38_244 ();
 DECAPx10_ASAP7_75t_R FILLER_38_266 ();
 DECAPx10_ASAP7_75t_R FILLER_38_288 ();
 DECAPx10_ASAP7_75t_R FILLER_38_310 ();
 DECAPx10_ASAP7_75t_R FILLER_38_332 ();
 DECAPx10_ASAP7_75t_R FILLER_38_354 ();
 DECAPx10_ASAP7_75t_R FILLER_38_376 ();
 DECAPx10_ASAP7_75t_R FILLER_38_398 ();
 DECAPx10_ASAP7_75t_R FILLER_38_420 ();
 DECAPx6_ASAP7_75t_R FILLER_38_442 ();
 DECAPx2_ASAP7_75t_R FILLER_38_456 ();
 DECAPx10_ASAP7_75t_R FILLER_38_464 ();
 DECAPx10_ASAP7_75t_R FILLER_38_486 ();
 DECAPx6_ASAP7_75t_R FILLER_38_508 ();
 FILLER_ASAP7_75t_R FILLER_38_522 ();
 DECAPx2_ASAP7_75t_R FILLER_38_561 ();
 FILLER_ASAP7_75t_R FILLER_38_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_569 ();
 DECAPx2_ASAP7_75t_R FILLER_38_579 ();
 FILLER_ASAP7_75t_R FILLER_38_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_605 ();
 DECAPx4_ASAP7_75t_R FILLER_38_615 ();
 FILLER_ASAP7_75t_R FILLER_38_625 ();
 FILLER_ASAP7_75t_R FILLER_38_647 ();
 DECAPx4_ASAP7_75t_R FILLER_38_666 ();
 FILLER_ASAP7_75t_R FILLER_38_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_678 ();
 DECAPx1_ASAP7_75t_R FILLER_38_702 ();
 DECAPx1_ASAP7_75t_R FILLER_38_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_716 ();
 DECAPx6_ASAP7_75t_R FILLER_38_734 ();
 DECAPx4_ASAP7_75t_R FILLER_38_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_768 ();
 DECAPx2_ASAP7_75t_R FILLER_38_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_784 ();
 DECAPx6_ASAP7_75t_R FILLER_38_799 ();
 DECAPx1_ASAP7_75t_R FILLER_38_813 ();
 DECAPx4_ASAP7_75t_R FILLER_38_827 ();
 FILLER_ASAP7_75t_R FILLER_38_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_839 ();
 DECAPx1_ASAP7_75t_R FILLER_38_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_886 ();
 DECAPx1_ASAP7_75t_R FILLER_38_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_894 ();
 DECAPx2_ASAP7_75t_R FILLER_38_929 ();
 FILLER_ASAP7_75t_R FILLER_38_935 ();
 DECAPx4_ASAP7_75t_R FILLER_38_963 ();
 DECAPx1_ASAP7_75t_R FILLER_38_999 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1036 ();
 FILLER_ASAP7_75t_R FILLER_38_1042 ();
 DECAPx6_ASAP7_75t_R FILLER_38_1066 ();
 DECAPx6_ASAP7_75t_R FILLER_38_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1175 ();
 FILLER_ASAP7_75t_R FILLER_38_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1352 ();
 DECAPx4_ASAP7_75t_R FILLER_38_1374 ();
 FILLER_ASAP7_75t_R FILLER_38_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_39_2 ();
 DECAPx10_ASAP7_75t_R FILLER_39_24 ();
 DECAPx10_ASAP7_75t_R FILLER_39_46 ();
 DECAPx10_ASAP7_75t_R FILLER_39_68 ();
 DECAPx10_ASAP7_75t_R FILLER_39_90 ();
 DECAPx10_ASAP7_75t_R FILLER_39_112 ();
 DECAPx10_ASAP7_75t_R FILLER_39_134 ();
 DECAPx10_ASAP7_75t_R FILLER_39_156 ();
 DECAPx10_ASAP7_75t_R FILLER_39_178 ();
 DECAPx10_ASAP7_75t_R FILLER_39_200 ();
 DECAPx10_ASAP7_75t_R FILLER_39_222 ();
 DECAPx10_ASAP7_75t_R FILLER_39_244 ();
 DECAPx10_ASAP7_75t_R FILLER_39_266 ();
 DECAPx10_ASAP7_75t_R FILLER_39_288 ();
 DECAPx10_ASAP7_75t_R FILLER_39_310 ();
 DECAPx10_ASAP7_75t_R FILLER_39_332 ();
 DECAPx10_ASAP7_75t_R FILLER_39_354 ();
 DECAPx10_ASAP7_75t_R FILLER_39_376 ();
 DECAPx10_ASAP7_75t_R FILLER_39_398 ();
 DECAPx10_ASAP7_75t_R FILLER_39_420 ();
 DECAPx10_ASAP7_75t_R FILLER_39_442 ();
 DECAPx10_ASAP7_75t_R FILLER_39_464 ();
 DECAPx10_ASAP7_75t_R FILLER_39_486 ();
 DECAPx6_ASAP7_75t_R FILLER_39_508 ();
 DECAPx2_ASAP7_75t_R FILLER_39_522 ();
 DECAPx2_ASAP7_75t_R FILLER_39_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_563 ();
 DECAPx4_ASAP7_75t_R FILLER_39_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_597 ();
 DECAPx6_ASAP7_75t_R FILLER_39_604 ();
 DECAPx1_ASAP7_75t_R FILLER_39_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_622 ();
 FILLER_ASAP7_75t_R FILLER_39_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_654 ();
 DECAPx1_ASAP7_75t_R FILLER_39_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_673 ();
 DECAPx6_ASAP7_75t_R FILLER_39_688 ();
 DECAPx2_ASAP7_75t_R FILLER_39_702 ();
 DECAPx4_ASAP7_75t_R FILLER_39_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_732 ();
 DECAPx6_ASAP7_75t_R FILLER_39_742 ();
 DECAPx2_ASAP7_75t_R FILLER_39_756 ();
 DECAPx1_ASAP7_75t_R FILLER_39_768 ();
 DECAPx2_ASAP7_75t_R FILLER_39_780 ();
 FILLER_ASAP7_75t_R FILLER_39_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_788 ();
 DECAPx2_ASAP7_75t_R FILLER_39_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_801 ();
 DECAPx2_ASAP7_75t_R FILLER_39_828 ();
 FILLER_ASAP7_75t_R FILLER_39_834 ();
 FILLER_ASAP7_75t_R FILLER_39_862 ();
 DECAPx4_ASAP7_75t_R FILLER_39_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_894 ();
 DECAPx1_ASAP7_75t_R FILLER_39_905 ();
 DECAPx1_ASAP7_75t_R FILLER_39_912 ();
 DECAPx2_ASAP7_75t_R FILLER_39_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_940 ();
 FILLER_ASAP7_75t_R FILLER_39_967 ();
 DECAPx2_ASAP7_75t_R FILLER_39_979 ();
 FILLER_ASAP7_75t_R FILLER_39_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_987 ();
 DECAPx1_ASAP7_75t_R FILLER_39_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_995 ();
 DECAPx6_ASAP7_75t_R FILLER_39_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_39_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_39_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_39_1085 ();
 FILLER_ASAP7_75t_R FILLER_39_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1217 ();
 DECAPx6_ASAP7_75t_R FILLER_39_1227 ();
 FILLER_ASAP7_75t_R FILLER_39_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1349 ();
 DECAPx6_ASAP7_75t_R FILLER_39_1371 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1385 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_40_2 ();
 DECAPx10_ASAP7_75t_R FILLER_40_24 ();
 DECAPx10_ASAP7_75t_R FILLER_40_46 ();
 DECAPx10_ASAP7_75t_R FILLER_40_68 ();
 DECAPx10_ASAP7_75t_R FILLER_40_90 ();
 DECAPx10_ASAP7_75t_R FILLER_40_112 ();
 DECAPx10_ASAP7_75t_R FILLER_40_134 ();
 DECAPx10_ASAP7_75t_R FILLER_40_156 ();
 DECAPx10_ASAP7_75t_R FILLER_40_178 ();
 DECAPx10_ASAP7_75t_R FILLER_40_200 ();
 DECAPx10_ASAP7_75t_R FILLER_40_222 ();
 DECAPx10_ASAP7_75t_R FILLER_40_244 ();
 DECAPx10_ASAP7_75t_R FILLER_40_266 ();
 DECAPx10_ASAP7_75t_R FILLER_40_288 ();
 DECAPx10_ASAP7_75t_R FILLER_40_310 ();
 DECAPx10_ASAP7_75t_R FILLER_40_332 ();
 DECAPx10_ASAP7_75t_R FILLER_40_354 ();
 DECAPx10_ASAP7_75t_R FILLER_40_376 ();
 DECAPx10_ASAP7_75t_R FILLER_40_398 ();
 DECAPx10_ASAP7_75t_R FILLER_40_420 ();
 DECAPx6_ASAP7_75t_R FILLER_40_442 ();
 DECAPx2_ASAP7_75t_R FILLER_40_456 ();
 DECAPx10_ASAP7_75t_R FILLER_40_464 ();
 DECAPx10_ASAP7_75t_R FILLER_40_486 ();
 DECAPx6_ASAP7_75t_R FILLER_40_508 ();
 DECAPx1_ASAP7_75t_R FILLER_40_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_526 ();
 DECAPx4_ASAP7_75t_R FILLER_40_556 ();
 FILLER_ASAP7_75t_R FILLER_40_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_568 ();
 DECAPx10_ASAP7_75t_R FILLER_40_578 ();
 DECAPx2_ASAP7_75t_R FILLER_40_600 ();
 FILLER_ASAP7_75t_R FILLER_40_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_608 ();
 DECAPx1_ASAP7_75t_R FILLER_40_619 ();
 DECAPx2_ASAP7_75t_R FILLER_40_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_649 ();
 DECAPx2_ASAP7_75t_R FILLER_40_653 ();
 FILLER_ASAP7_75t_R FILLER_40_659 ();
 FILLER_ASAP7_75t_R FILLER_40_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_666 ();
 DECAPx4_ASAP7_75t_R FILLER_40_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_694 ();
 DECAPx1_ASAP7_75t_R FILLER_40_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_702 ();
 DECAPx2_ASAP7_75t_R FILLER_40_706 ();
 DECAPx2_ASAP7_75t_R FILLER_40_721 ();
 FILLER_ASAP7_75t_R FILLER_40_727 ();
 DECAPx1_ASAP7_75t_R FILLER_40_738 ();
 DECAPx2_ASAP7_75t_R FILLER_40_749 ();
 FILLER_ASAP7_75t_R FILLER_40_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_757 ();
 DECAPx2_ASAP7_75t_R FILLER_40_770 ();
 FILLER_ASAP7_75t_R FILLER_40_776 ();
 DECAPx2_ASAP7_75t_R FILLER_40_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_791 ();
 DECAPx1_ASAP7_75t_R FILLER_40_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_805 ();
 DECAPx1_ASAP7_75t_R FILLER_40_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_834 ();
 FILLER_ASAP7_75t_R FILLER_40_848 ();
 DECAPx6_ASAP7_75t_R FILLER_40_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_867 ();
 DECAPx6_ASAP7_75t_R FILLER_40_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_893 ();
 FILLER_ASAP7_75t_R FILLER_40_902 ();
 DECAPx2_ASAP7_75t_R FILLER_40_912 ();
 DECAPx1_ASAP7_75t_R FILLER_40_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_938 ();
 DECAPx2_ASAP7_75t_R FILLER_40_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_955 ();
 DECAPx2_ASAP7_75t_R FILLER_40_959 ();
 FILLER_ASAP7_75t_R FILLER_40_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_986 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1023 ();
 FILLER_ASAP7_75t_R FILLER_40_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1068 ();
 FILLER_ASAP7_75t_R FILLER_40_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_40_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1146 ();
 FILLER_ASAP7_75t_R FILLER_40_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1170 ();
 DECAPx4_ASAP7_75t_R FILLER_40_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1187 ();
 DECAPx6_ASAP7_75t_R FILLER_40_1203 ();
 FILLER_ASAP7_75t_R FILLER_40_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1219 ();
 DECAPx6_ASAP7_75t_R FILLER_40_1226 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1350 ();
 DECAPx6_ASAP7_75t_R FILLER_40_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_41_2 ();
 DECAPx10_ASAP7_75t_R FILLER_41_24 ();
 DECAPx10_ASAP7_75t_R FILLER_41_46 ();
 DECAPx10_ASAP7_75t_R FILLER_41_68 ();
 DECAPx10_ASAP7_75t_R FILLER_41_90 ();
 DECAPx10_ASAP7_75t_R FILLER_41_112 ();
 DECAPx10_ASAP7_75t_R FILLER_41_134 ();
 DECAPx10_ASAP7_75t_R FILLER_41_156 ();
 DECAPx10_ASAP7_75t_R FILLER_41_178 ();
 DECAPx10_ASAP7_75t_R FILLER_41_200 ();
 DECAPx10_ASAP7_75t_R FILLER_41_222 ();
 DECAPx10_ASAP7_75t_R FILLER_41_244 ();
 DECAPx10_ASAP7_75t_R FILLER_41_266 ();
 DECAPx10_ASAP7_75t_R FILLER_41_288 ();
 DECAPx10_ASAP7_75t_R FILLER_41_310 ();
 DECAPx10_ASAP7_75t_R FILLER_41_332 ();
 DECAPx10_ASAP7_75t_R FILLER_41_354 ();
 DECAPx10_ASAP7_75t_R FILLER_41_376 ();
 DECAPx10_ASAP7_75t_R FILLER_41_398 ();
 DECAPx10_ASAP7_75t_R FILLER_41_420 ();
 DECAPx10_ASAP7_75t_R FILLER_41_442 ();
 DECAPx10_ASAP7_75t_R FILLER_41_464 ();
 DECAPx10_ASAP7_75t_R FILLER_41_486 ();
 DECAPx2_ASAP7_75t_R FILLER_41_508 ();
 FILLER_ASAP7_75t_R FILLER_41_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_549 ();
 DECAPx6_ASAP7_75t_R FILLER_41_561 ();
 DECAPx1_ASAP7_75t_R FILLER_41_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_579 ();
 DECAPx4_ASAP7_75t_R FILLER_41_594 ();
 FILLER_ASAP7_75t_R FILLER_41_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_621 ();
 DECAPx1_ASAP7_75t_R FILLER_41_636 ();
 FILLER_ASAP7_75t_R FILLER_41_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_645 ();
 DECAPx2_ASAP7_75t_R FILLER_41_660 ();
 FILLER_ASAP7_75t_R FILLER_41_666 ();
 DECAPx1_ASAP7_75t_R FILLER_41_697 ();
 FILLER_ASAP7_75t_R FILLER_41_710 ();
 DECAPx4_ASAP7_75t_R FILLER_41_718 ();
 FILLER_ASAP7_75t_R FILLER_41_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_742 ();
 DECAPx1_ASAP7_75t_R FILLER_41_754 ();
 DECAPx1_ASAP7_75t_R FILLER_41_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_778 ();
 FILLER_ASAP7_75t_R FILLER_41_785 ();
 DECAPx2_ASAP7_75t_R FILLER_41_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_826 ();
 DECAPx2_ASAP7_75t_R FILLER_41_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_841 ();
 DECAPx6_ASAP7_75t_R FILLER_41_850 ();
 DECAPx1_ASAP7_75t_R FILLER_41_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_868 ();
 DECAPx4_ASAP7_75t_R FILLER_41_877 ();
 FILLER_ASAP7_75t_R FILLER_41_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_906 ();
 DECAPx2_ASAP7_75t_R FILLER_41_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_923 ();
 DECAPx4_ASAP7_75t_R FILLER_41_934 ();
 FILLER_ASAP7_75t_R FILLER_41_944 ();
 DECAPx4_ASAP7_75t_R FILLER_41_956 ();
 FILLER_ASAP7_75t_R FILLER_41_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_974 ();
 FILLER_ASAP7_75t_R FILLER_41_979 ();
 DECAPx2_ASAP7_75t_R FILLER_41_987 ();
 FILLER_ASAP7_75t_R FILLER_41_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_995 ();
 FILLER_ASAP7_75t_R FILLER_41_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_41_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1112 ();
 FILLER_ASAP7_75t_R FILLER_41_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1120 ();
 DECAPx6_ASAP7_75t_R FILLER_41_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1159 ();
 FILLER_ASAP7_75t_R FILLER_41_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_41_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_41_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1386 ();
 DECAPx10_ASAP7_75t_R FILLER_42_2 ();
 DECAPx10_ASAP7_75t_R FILLER_42_24 ();
 DECAPx10_ASAP7_75t_R FILLER_42_46 ();
 DECAPx10_ASAP7_75t_R FILLER_42_68 ();
 DECAPx10_ASAP7_75t_R FILLER_42_90 ();
 DECAPx10_ASAP7_75t_R FILLER_42_112 ();
 DECAPx10_ASAP7_75t_R FILLER_42_134 ();
 DECAPx10_ASAP7_75t_R FILLER_42_156 ();
 DECAPx10_ASAP7_75t_R FILLER_42_178 ();
 DECAPx10_ASAP7_75t_R FILLER_42_200 ();
 DECAPx10_ASAP7_75t_R FILLER_42_222 ();
 DECAPx10_ASAP7_75t_R FILLER_42_244 ();
 DECAPx10_ASAP7_75t_R FILLER_42_266 ();
 DECAPx10_ASAP7_75t_R FILLER_42_288 ();
 DECAPx10_ASAP7_75t_R FILLER_42_310 ();
 DECAPx10_ASAP7_75t_R FILLER_42_332 ();
 DECAPx10_ASAP7_75t_R FILLER_42_354 ();
 DECAPx10_ASAP7_75t_R FILLER_42_376 ();
 DECAPx10_ASAP7_75t_R FILLER_42_398 ();
 DECAPx10_ASAP7_75t_R FILLER_42_420 ();
 DECAPx6_ASAP7_75t_R FILLER_42_442 ();
 DECAPx2_ASAP7_75t_R FILLER_42_456 ();
 DECAPx10_ASAP7_75t_R FILLER_42_464 ();
 DECAPx10_ASAP7_75t_R FILLER_42_486 ();
 DECAPx6_ASAP7_75t_R FILLER_42_508 ();
 FILLER_ASAP7_75t_R FILLER_42_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_524 ();
 DECAPx4_ASAP7_75t_R FILLER_42_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_545 ();
 DECAPx1_ASAP7_75t_R FILLER_42_594 ();
 FILLER_ASAP7_75t_R FILLER_42_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_635 ();
 DECAPx10_ASAP7_75t_R FILLER_42_639 ();
 DECAPx2_ASAP7_75t_R FILLER_42_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_667 ();
 DECAPx6_ASAP7_75t_R FILLER_42_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_692 ();
 FILLER_ASAP7_75t_R FILLER_42_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_729 ();
 FILLER_ASAP7_75t_R FILLER_42_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_757 ();
 DECAPx2_ASAP7_75t_R FILLER_42_769 ();
 FILLER_ASAP7_75t_R FILLER_42_775 ();
 DECAPx1_ASAP7_75t_R FILLER_42_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_795 ();
 FILLER_ASAP7_75t_R FILLER_42_799 ();
 FILLER_ASAP7_75t_R FILLER_42_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_813 ();
 DECAPx2_ASAP7_75t_R FILLER_42_817 ();
 DECAPx6_ASAP7_75t_R FILLER_42_831 ();
 DECAPx2_ASAP7_75t_R FILLER_42_858 ();
 FILLER_ASAP7_75t_R FILLER_42_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_866 ();
 DECAPx4_ASAP7_75t_R FILLER_42_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_885 ();
 DECAPx4_ASAP7_75t_R FILLER_42_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_904 ();
 DECAPx6_ASAP7_75t_R FILLER_42_911 ();
 FILLER_ASAP7_75t_R FILLER_42_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_927 ();
 DECAPx2_ASAP7_75t_R FILLER_42_935 ();
 FILLER_ASAP7_75t_R FILLER_42_941 ();
 DECAPx4_ASAP7_75t_R FILLER_42_949 ();
 FILLER_ASAP7_75t_R FILLER_42_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_961 ();
 DECAPx1_ASAP7_75t_R FILLER_42_974 ();
 DECAPx2_ASAP7_75t_R FILLER_42_989 ();
 FILLER_ASAP7_75t_R FILLER_42_995 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_42_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1046 ();
 DECAPx6_ASAP7_75t_R FILLER_42_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_42_1080 ();
 FILLER_ASAP7_75t_R FILLER_42_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_42_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_43_2 ();
 DECAPx10_ASAP7_75t_R FILLER_43_24 ();
 DECAPx10_ASAP7_75t_R FILLER_43_46 ();
 DECAPx10_ASAP7_75t_R FILLER_43_68 ();
 DECAPx10_ASAP7_75t_R FILLER_43_90 ();
 DECAPx10_ASAP7_75t_R FILLER_43_112 ();
 DECAPx10_ASAP7_75t_R FILLER_43_134 ();
 DECAPx10_ASAP7_75t_R FILLER_43_156 ();
 DECAPx10_ASAP7_75t_R FILLER_43_178 ();
 DECAPx10_ASAP7_75t_R FILLER_43_200 ();
 DECAPx10_ASAP7_75t_R FILLER_43_222 ();
 DECAPx10_ASAP7_75t_R FILLER_43_244 ();
 DECAPx10_ASAP7_75t_R FILLER_43_266 ();
 DECAPx10_ASAP7_75t_R FILLER_43_288 ();
 DECAPx10_ASAP7_75t_R FILLER_43_310 ();
 DECAPx10_ASAP7_75t_R FILLER_43_332 ();
 DECAPx10_ASAP7_75t_R FILLER_43_354 ();
 DECAPx10_ASAP7_75t_R FILLER_43_376 ();
 DECAPx10_ASAP7_75t_R FILLER_43_398 ();
 DECAPx10_ASAP7_75t_R FILLER_43_420 ();
 DECAPx10_ASAP7_75t_R FILLER_43_442 ();
 DECAPx10_ASAP7_75t_R FILLER_43_464 ();
 DECAPx10_ASAP7_75t_R FILLER_43_486 ();
 DECAPx6_ASAP7_75t_R FILLER_43_508 ();
 DECAPx2_ASAP7_75t_R FILLER_43_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_528 ();
 DECAPx4_ASAP7_75t_R FILLER_43_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_551 ();
 DECAPx6_ASAP7_75t_R FILLER_43_563 ();
 FILLER_ASAP7_75t_R FILLER_43_577 ();
 DECAPx1_ASAP7_75t_R FILLER_43_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_590 ();
 DECAPx2_ASAP7_75t_R FILLER_43_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_600 ();
 DECAPx4_ASAP7_75t_R FILLER_43_615 ();
 DECAPx2_ASAP7_75t_R FILLER_43_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_637 ();
 DECAPx6_ASAP7_75t_R FILLER_43_652 ();
 DECAPx2_ASAP7_75t_R FILLER_43_666 ();
 DECAPx10_ASAP7_75t_R FILLER_43_681 ();
 DECAPx1_ASAP7_75t_R FILLER_43_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_707 ();
 DECAPx2_ASAP7_75t_R FILLER_43_731 ();
 FILLER_ASAP7_75t_R FILLER_43_737 ();
 DECAPx10_ASAP7_75t_R FILLER_43_750 ();
 DECAPx4_ASAP7_75t_R FILLER_43_772 ();
 DECAPx4_ASAP7_75t_R FILLER_43_791 ();
 DECAPx2_ASAP7_75t_R FILLER_43_814 ();
 DECAPx6_ASAP7_75t_R FILLER_43_823 ();
 FILLER_ASAP7_75t_R FILLER_43_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_839 ();
 DECAPx1_ASAP7_75t_R FILLER_43_866 ();
 DECAPx4_ASAP7_75t_R FILLER_43_878 ();
 FILLER_ASAP7_75t_R FILLER_43_888 ();
 DECAPx1_ASAP7_75t_R FILLER_43_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_904 ();
 DECAPx2_ASAP7_75t_R FILLER_43_915 ();
 FILLER_ASAP7_75t_R FILLER_43_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_923 ();
 DECAPx4_ASAP7_75t_R FILLER_43_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_998 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_43_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_43_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_43_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1077 ();
 DECAPx6_ASAP7_75t_R FILLER_43_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_43_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_43_1112 ();
 FILLER_ASAP7_75t_R FILLER_43_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_43_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_43_1159 ();
 FILLER_ASAP7_75t_R FILLER_43_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_43_1177 ();
 FILLER_ASAP7_75t_R FILLER_43_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1355 ();
 FILLER_ASAP7_75t_R FILLER_43_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1379 ();
 DECAPx10_ASAP7_75t_R FILLER_44_2 ();
 DECAPx10_ASAP7_75t_R FILLER_44_24 ();
 DECAPx10_ASAP7_75t_R FILLER_44_46 ();
 DECAPx10_ASAP7_75t_R FILLER_44_68 ();
 DECAPx10_ASAP7_75t_R FILLER_44_90 ();
 DECAPx10_ASAP7_75t_R FILLER_44_112 ();
 DECAPx10_ASAP7_75t_R FILLER_44_134 ();
 DECAPx10_ASAP7_75t_R FILLER_44_156 ();
 DECAPx10_ASAP7_75t_R FILLER_44_178 ();
 DECAPx10_ASAP7_75t_R FILLER_44_200 ();
 DECAPx10_ASAP7_75t_R FILLER_44_222 ();
 DECAPx10_ASAP7_75t_R FILLER_44_244 ();
 DECAPx10_ASAP7_75t_R FILLER_44_266 ();
 DECAPx10_ASAP7_75t_R FILLER_44_288 ();
 DECAPx10_ASAP7_75t_R FILLER_44_310 ();
 DECAPx10_ASAP7_75t_R FILLER_44_332 ();
 DECAPx10_ASAP7_75t_R FILLER_44_354 ();
 DECAPx10_ASAP7_75t_R FILLER_44_376 ();
 DECAPx10_ASAP7_75t_R FILLER_44_398 ();
 DECAPx10_ASAP7_75t_R FILLER_44_420 ();
 DECAPx6_ASAP7_75t_R FILLER_44_442 ();
 DECAPx2_ASAP7_75t_R FILLER_44_456 ();
 DECAPx10_ASAP7_75t_R FILLER_44_464 ();
 DECAPx10_ASAP7_75t_R FILLER_44_486 ();
 DECAPx4_ASAP7_75t_R FILLER_44_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_518 ();
 DECAPx2_ASAP7_75t_R FILLER_44_533 ();
 FILLER_ASAP7_75t_R FILLER_44_548 ();
 FILLER_ASAP7_75t_R FILLER_44_564 ();
 DECAPx4_ASAP7_75t_R FILLER_44_577 ();
 FILLER_ASAP7_75t_R FILLER_44_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_589 ();
 DECAPx6_ASAP7_75t_R FILLER_44_593 ();
 FILLER_ASAP7_75t_R FILLER_44_607 ();
 DECAPx4_ASAP7_75t_R FILLER_44_619 ();
 FILLER_ASAP7_75t_R FILLER_44_629 ();
 DECAPx1_ASAP7_75t_R FILLER_44_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_641 ();
 DECAPx2_ASAP7_75t_R FILLER_44_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_665 ();
 FILLER_ASAP7_75t_R FILLER_44_676 ();
 DECAPx1_ASAP7_75t_R FILLER_44_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_694 ();
 DECAPx1_ASAP7_75t_R FILLER_44_705 ();
 DECAPx2_ASAP7_75t_R FILLER_44_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_738 ();
 FILLER_ASAP7_75t_R FILLER_44_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_750 ();
 FILLER_ASAP7_75t_R FILLER_44_757 ();
 DECAPx4_ASAP7_75t_R FILLER_44_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_781 ();
 FILLER_ASAP7_75t_R FILLER_44_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_836 ();
 DECAPx6_ASAP7_75t_R FILLER_44_858 ();
 DECAPx1_ASAP7_75t_R FILLER_44_872 ();
 DECAPx1_ASAP7_75t_R FILLER_44_892 ();
 DECAPx2_ASAP7_75t_R FILLER_44_912 ();
 FILLER_ASAP7_75t_R FILLER_44_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_920 ();
 DECAPx4_ASAP7_75t_R FILLER_44_949 ();
 DECAPx4_ASAP7_75t_R FILLER_44_965 ();
 FILLER_ASAP7_75t_R FILLER_44_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1012 ();
 FILLER_ASAP7_75t_R FILLER_44_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1038 ();
 DECAPx4_ASAP7_75t_R FILLER_44_1093 ();
 FILLER_ASAP7_75t_R FILLER_44_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1142 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1214 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1230 ();
 FILLER_ASAP7_75t_R FILLER_44_1236 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_45_2 ();
 DECAPx10_ASAP7_75t_R FILLER_45_24 ();
 DECAPx10_ASAP7_75t_R FILLER_45_46 ();
 DECAPx10_ASAP7_75t_R FILLER_45_68 ();
 DECAPx10_ASAP7_75t_R FILLER_45_90 ();
 DECAPx10_ASAP7_75t_R FILLER_45_112 ();
 DECAPx10_ASAP7_75t_R FILLER_45_134 ();
 DECAPx10_ASAP7_75t_R FILLER_45_156 ();
 DECAPx10_ASAP7_75t_R FILLER_45_178 ();
 DECAPx10_ASAP7_75t_R FILLER_45_200 ();
 DECAPx10_ASAP7_75t_R FILLER_45_222 ();
 DECAPx10_ASAP7_75t_R FILLER_45_244 ();
 DECAPx10_ASAP7_75t_R FILLER_45_266 ();
 DECAPx10_ASAP7_75t_R FILLER_45_288 ();
 DECAPx10_ASAP7_75t_R FILLER_45_310 ();
 DECAPx10_ASAP7_75t_R FILLER_45_332 ();
 DECAPx10_ASAP7_75t_R FILLER_45_354 ();
 DECAPx10_ASAP7_75t_R FILLER_45_376 ();
 DECAPx10_ASAP7_75t_R FILLER_45_398 ();
 DECAPx10_ASAP7_75t_R FILLER_45_420 ();
 DECAPx10_ASAP7_75t_R FILLER_45_442 ();
 DECAPx10_ASAP7_75t_R FILLER_45_464 ();
 DECAPx10_ASAP7_75t_R FILLER_45_486 ();
 DECAPx2_ASAP7_75t_R FILLER_45_508 ();
 FILLER_ASAP7_75t_R FILLER_45_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_516 ();
 DECAPx4_ASAP7_75t_R FILLER_45_549 ();
 FILLER_ASAP7_75t_R FILLER_45_559 ();
 DECAPx4_ASAP7_75t_R FILLER_45_572 ();
 FILLER_ASAP7_75t_R FILLER_45_582 ();
 DECAPx2_ASAP7_75t_R FILLER_45_619 ();
 FILLER_ASAP7_75t_R FILLER_45_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_627 ();
 DECAPx2_ASAP7_75t_R FILLER_45_642 ();
 FILLER_ASAP7_75t_R FILLER_45_648 ();
 DECAPx2_ASAP7_75t_R FILLER_45_653 ();
 FILLER_ASAP7_75t_R FILLER_45_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_689 ();
 DECAPx1_ASAP7_75t_R FILLER_45_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_708 ();
 DECAPx2_ASAP7_75t_R FILLER_45_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_718 ();
 DECAPx6_ASAP7_75t_R FILLER_45_722 ();
 DECAPx2_ASAP7_75t_R FILLER_45_736 ();
 DECAPx6_ASAP7_75t_R FILLER_45_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_776 ();
 DECAPx4_ASAP7_75t_R FILLER_45_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_796 ();
 DECAPx2_ASAP7_75t_R FILLER_45_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_862 ();
 DECAPx2_ASAP7_75t_R FILLER_45_889 ();
 FILLER_ASAP7_75t_R FILLER_45_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_897 ();
 DECAPx1_ASAP7_75t_R FILLER_45_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_930 ();
 FILLER_ASAP7_75t_R FILLER_45_937 ();
 FILLER_ASAP7_75t_R FILLER_45_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_957 ();
 DECAPx2_ASAP7_75t_R FILLER_45_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_978 ();
 DECAPx2_ASAP7_75t_R FILLER_45_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_994 ();
 FILLER_ASAP7_75t_R FILLER_45_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_45_1067 ();
 FILLER_ASAP7_75t_R FILLER_45_1081 ();
 FILLER_ASAP7_75t_R FILLER_45_1089 ();
 DECAPx4_ASAP7_75t_R FILLER_45_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1128 ();
 FILLER_ASAP7_75t_R FILLER_45_1150 ();
 DECAPx4_ASAP7_75t_R FILLER_45_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1170 ();
 DECAPx4_ASAP7_75t_R FILLER_45_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1350 ();
 DECAPx6_ASAP7_75t_R FILLER_45_1372 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1386 ();
 DECAPx10_ASAP7_75t_R FILLER_46_2 ();
 DECAPx10_ASAP7_75t_R FILLER_46_24 ();
 DECAPx10_ASAP7_75t_R FILLER_46_46 ();
 DECAPx10_ASAP7_75t_R FILLER_46_68 ();
 DECAPx10_ASAP7_75t_R FILLER_46_90 ();
 DECAPx10_ASAP7_75t_R FILLER_46_112 ();
 DECAPx10_ASAP7_75t_R FILLER_46_134 ();
 DECAPx10_ASAP7_75t_R FILLER_46_156 ();
 DECAPx6_ASAP7_75t_R FILLER_46_178 ();
 FILLER_ASAP7_75t_R FILLER_46_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_194 ();
 DECAPx10_ASAP7_75t_R FILLER_46_247 ();
 DECAPx4_ASAP7_75t_R FILLER_46_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_308 ();
 DECAPx10_ASAP7_75t_R FILLER_46_339 ();
 DECAPx10_ASAP7_75t_R FILLER_46_361 ();
 DECAPx10_ASAP7_75t_R FILLER_46_383 ();
 DECAPx6_ASAP7_75t_R FILLER_46_405 ();
 FILLER_ASAP7_75t_R FILLER_46_419 ();
 DECAPx10_ASAP7_75t_R FILLER_46_424 ();
 DECAPx6_ASAP7_75t_R FILLER_46_446 ();
 FILLER_ASAP7_75t_R FILLER_46_460 ();
 DECAPx10_ASAP7_75t_R FILLER_46_464 ();
 DECAPx10_ASAP7_75t_R FILLER_46_486 ();
 DECAPx2_ASAP7_75t_R FILLER_46_508 ();
 FILLER_ASAP7_75t_R FILLER_46_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_516 ();
 DECAPx6_ASAP7_75t_R FILLER_46_535 ();
 FILLER_ASAP7_75t_R FILLER_46_549 ();
 DECAPx6_ASAP7_75t_R FILLER_46_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_568 ();
 DECAPx4_ASAP7_75t_R FILLER_46_591 ();
 FILLER_ASAP7_75t_R FILLER_46_601 ();
 DECAPx1_ASAP7_75t_R FILLER_46_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_656 ();
 DECAPx6_ASAP7_75t_R FILLER_46_671 ();
 DECAPx1_ASAP7_75t_R FILLER_46_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_689 ();
 DECAPx2_ASAP7_75t_R FILLER_46_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_702 ();
 FILLER_ASAP7_75t_R FILLER_46_706 ();
 DECAPx2_ASAP7_75t_R FILLER_46_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_728 ();
 DECAPx10_ASAP7_75t_R FILLER_46_738 ();
 DECAPx2_ASAP7_75t_R FILLER_46_760 ();
 FILLER_ASAP7_75t_R FILLER_46_766 ();
 DECAPx2_ASAP7_75t_R FILLER_46_771 ();
 FILLER_ASAP7_75t_R FILLER_46_777 ();
 DECAPx1_ASAP7_75t_R FILLER_46_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_793 ();
 FILLER_ASAP7_75t_R FILLER_46_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_799 ();
 DECAPx2_ASAP7_75t_R FILLER_46_849 ();
 FILLER_ASAP7_75t_R FILLER_46_855 ();
 DECAPx2_ASAP7_75t_R FILLER_46_867 ();
 FILLER_ASAP7_75t_R FILLER_46_873 ();
 DECAPx6_ASAP7_75t_R FILLER_46_886 ();
 FILLER_ASAP7_75t_R FILLER_46_900 ();
 DECAPx1_ASAP7_75t_R FILLER_46_910 ();
 DECAPx2_ASAP7_75t_R FILLER_46_917 ();
 FILLER_ASAP7_75t_R FILLER_46_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_925 ();
 FILLER_ASAP7_75t_R FILLER_46_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_944 ();
 FILLER_ASAP7_75t_R FILLER_46_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_954 ();
 DECAPx4_ASAP7_75t_R FILLER_46_965 ();
 FILLER_ASAP7_75t_R FILLER_46_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_977 ();
 DECAPx10_ASAP7_75t_R FILLER_46_987 ();
 FILLER_ASAP7_75t_R FILLER_46_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1022 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1044 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1096 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1204 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1378 ();
 FILLER_ASAP7_75t_R FILLER_46_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_47_2 ();
 DECAPx10_ASAP7_75t_R FILLER_47_24 ();
 DECAPx10_ASAP7_75t_R FILLER_47_46 ();
 DECAPx10_ASAP7_75t_R FILLER_47_68 ();
 DECAPx10_ASAP7_75t_R FILLER_47_90 ();
 DECAPx10_ASAP7_75t_R FILLER_47_112 ();
 DECAPx10_ASAP7_75t_R FILLER_47_134 ();
 DECAPx10_ASAP7_75t_R FILLER_47_156 ();
 DECAPx10_ASAP7_75t_R FILLER_47_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_212 ();
 FILLER_ASAP7_75t_R FILLER_47_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_218 ();
 FILLER_ASAP7_75t_R FILLER_47_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_225 ();
 DECAPx2_ASAP7_75t_R FILLER_47_262 ();
 FILLER_ASAP7_75t_R FILLER_47_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_270 ();
 FILLER_ASAP7_75t_R FILLER_47_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_276 ();
 DECAPx2_ASAP7_75t_R FILLER_47_281 ();
 FILLER_ASAP7_75t_R FILLER_47_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_289 ();
 FILLER_ASAP7_75t_R FILLER_47_316 ();
 DECAPx6_ASAP7_75t_R FILLER_47_350 ();
 FILLER_ASAP7_75t_R FILLER_47_364 ();
 FILLER_ASAP7_75t_R FILLER_47_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_386 ();
 DECAPx1_ASAP7_75t_R FILLER_47_393 ();
 DECAPx2_ASAP7_75t_R FILLER_47_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_406 ();
 DECAPx10_ASAP7_75t_R FILLER_47_433 ();
 DECAPx10_ASAP7_75t_R FILLER_47_455 ();
 DECAPx1_ASAP7_75t_R FILLER_47_477 ();
 DECAPx10_ASAP7_75t_R FILLER_47_487 ();
 DECAPx6_ASAP7_75t_R FILLER_47_509 ();
 DECAPx4_ASAP7_75t_R FILLER_47_529 ();
 DECAPx4_ASAP7_75t_R FILLER_47_554 ();
 FILLER_ASAP7_75t_R FILLER_47_564 ();
 DECAPx1_ASAP7_75t_R FILLER_47_580 ();
 DECAPx4_ASAP7_75t_R FILLER_47_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_605 ();
 DECAPx6_ASAP7_75t_R FILLER_47_620 ();
 DECAPx6_ASAP7_75t_R FILLER_47_637 ();
 DECAPx1_ASAP7_75t_R FILLER_47_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_655 ();
 DECAPx6_ASAP7_75t_R FILLER_47_672 ();
 DECAPx1_ASAP7_75t_R FILLER_47_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_693 ();
 DECAPx1_ASAP7_75t_R FILLER_47_697 ();
 DECAPx2_ASAP7_75t_R FILLER_47_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_721 ();
 DECAPx6_ASAP7_75t_R FILLER_47_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_779 ();
 DECAPx1_ASAP7_75t_R FILLER_47_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_818 ();
 FILLER_ASAP7_75t_R FILLER_47_837 ();
 DECAPx1_ASAP7_75t_R FILLER_47_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_853 ();
 FILLER_ASAP7_75t_R FILLER_47_880 ();
 DECAPx2_ASAP7_75t_R FILLER_47_892 ();
 FILLER_ASAP7_75t_R FILLER_47_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_900 ();
 DECAPx4_ASAP7_75t_R FILLER_47_911 ();
 FILLER_ASAP7_75t_R FILLER_47_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_923 ();
 DECAPx1_ASAP7_75t_R FILLER_47_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_930 ();
 DECAPx1_ASAP7_75t_R FILLER_47_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_952 ();
 FILLER_ASAP7_75t_R FILLER_47_957 ();
 DECAPx4_ASAP7_75t_R FILLER_47_995 ();
 FILLER_ASAP7_75t_R FILLER_47_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1007 ();
 FILLER_ASAP7_75t_R FILLER_47_1011 ();
 DECAPx4_ASAP7_75t_R FILLER_47_1018 ();
 FILLER_ASAP7_75t_R FILLER_47_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1035 ();
 FILLER_ASAP7_75t_R FILLER_47_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_47_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1100 ();
 FILLER_ASAP7_75t_R FILLER_47_1106 ();
 FILLER_ASAP7_75t_R FILLER_47_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1223 ();
 FILLER_ASAP7_75t_R FILLER_47_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1352 ();
 DECAPx4_ASAP7_75t_R FILLER_47_1374 ();
 FILLER_ASAP7_75t_R FILLER_47_1384 ();
 DECAPx10_ASAP7_75t_R FILLER_48_2 ();
 DECAPx10_ASAP7_75t_R FILLER_48_24 ();
 DECAPx10_ASAP7_75t_R FILLER_48_46 ();
 DECAPx10_ASAP7_75t_R FILLER_48_68 ();
 DECAPx10_ASAP7_75t_R FILLER_48_90 ();
 DECAPx10_ASAP7_75t_R FILLER_48_112 ();
 DECAPx10_ASAP7_75t_R FILLER_48_134 ();
 DECAPx6_ASAP7_75t_R FILLER_48_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_170 ();
 DECAPx4_ASAP7_75t_R FILLER_48_197 ();
 FILLER_ASAP7_75t_R FILLER_48_207 ();
 FILLER_ASAP7_75t_R FILLER_48_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_217 ();
 DECAPx1_ASAP7_75t_R FILLER_48_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_225 ();
 FILLER_ASAP7_75t_R FILLER_48_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_234 ();
 DECAPx1_ASAP7_75t_R FILLER_48_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_248 ();
 DECAPx1_ASAP7_75t_R FILLER_48_282 ();
 DECAPx2_ASAP7_75t_R FILLER_48_308 ();
 FILLER_ASAP7_75t_R FILLER_48_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_323 ();
 FILLER_ASAP7_75t_R FILLER_48_340 ();
 DECAPx2_ASAP7_75t_R FILLER_48_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_352 ();
 DECAPx4_ASAP7_75t_R FILLER_48_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_381 ();
 FILLER_ASAP7_75t_R FILLER_48_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_450 ();
 DECAPx1_ASAP7_75t_R FILLER_48_458 ();
 FILLER_ASAP7_75t_R FILLER_48_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_466 ();
 DECAPx1_ASAP7_75t_R FILLER_48_473 ();
 DECAPx6_ASAP7_75t_R FILLER_48_506 ();
 FILLER_ASAP7_75t_R FILLER_48_520 ();
 DECAPx2_ASAP7_75t_R FILLER_48_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_537 ();
 FILLER_ASAP7_75t_R FILLER_48_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_568 ();
 DECAPx6_ASAP7_75t_R FILLER_48_583 ();
 FILLER_ASAP7_75t_R FILLER_48_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_599 ();
 DECAPx2_ASAP7_75t_R FILLER_48_620 ();
 FILLER_ASAP7_75t_R FILLER_48_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_628 ();
 DECAPx2_ASAP7_75t_R FILLER_48_639 ();
 DECAPx2_ASAP7_75t_R FILLER_48_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_665 ();
 FILLER_ASAP7_75t_R FILLER_48_672 ();
 DECAPx2_ASAP7_75t_R FILLER_48_702 ();
 FILLER_ASAP7_75t_R FILLER_48_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_710 ();
 DECAPx2_ASAP7_75t_R FILLER_48_719 ();
 DECAPx1_ASAP7_75t_R FILLER_48_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_735 ();
 DECAPx10_ASAP7_75t_R FILLER_48_762 ();
 DECAPx6_ASAP7_75t_R FILLER_48_784 ();
 DECAPx2_ASAP7_75t_R FILLER_48_812 ();
 FILLER_ASAP7_75t_R FILLER_48_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_820 ();
 FILLER_ASAP7_75t_R FILLER_48_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_868 ();
 DECAPx1_ASAP7_75t_R FILLER_48_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_876 ();
 FILLER_ASAP7_75t_R FILLER_48_929 ();
 DECAPx6_ASAP7_75t_R FILLER_48_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_955 ();
 DECAPx2_ASAP7_75t_R FILLER_48_976 ();
 FILLER_ASAP7_75t_R FILLER_48_982 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1020 ();
 FILLER_ASAP7_75t_R FILLER_48_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1028 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1036 ();
 FILLER_ASAP7_75t_R FILLER_48_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1051 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1078 ();
 FILLER_ASAP7_75t_R FILLER_48_1092 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1102 ();
 FILLER_ASAP7_75t_R FILLER_48_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1175 ();
 DECAPx4_ASAP7_75t_R FILLER_48_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1207 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1215 ();
 FILLER_ASAP7_75t_R FILLER_48_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1349 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_49_2 ();
 DECAPx10_ASAP7_75t_R FILLER_49_24 ();
 DECAPx10_ASAP7_75t_R FILLER_49_46 ();
 DECAPx10_ASAP7_75t_R FILLER_49_68 ();
 DECAPx10_ASAP7_75t_R FILLER_49_90 ();
 DECAPx10_ASAP7_75t_R FILLER_49_112 ();
 DECAPx10_ASAP7_75t_R FILLER_49_134 ();
 DECAPx4_ASAP7_75t_R FILLER_49_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_166 ();
 FILLER_ASAP7_75t_R FILLER_49_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_175 ();
 FILLER_ASAP7_75t_R FILLER_49_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_181 ();
 FILLER_ASAP7_75t_R FILLER_49_201 ();
 DECAPx1_ASAP7_75t_R FILLER_49_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_237 ();
 DECAPx6_ASAP7_75t_R FILLER_49_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_258 ();
 DECAPx6_ASAP7_75t_R FILLER_49_271 ();
 FILLER_ASAP7_75t_R FILLER_49_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_293 ();
 DECAPx10_ASAP7_75t_R FILLER_49_297 ();
 DECAPx2_ASAP7_75t_R FILLER_49_319 ();
 FILLER_ASAP7_75t_R FILLER_49_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_327 ();
 DECAPx2_ASAP7_75t_R FILLER_49_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_337 ();
 DECAPx6_ASAP7_75t_R FILLER_49_341 ();
 FILLER_ASAP7_75t_R FILLER_49_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_357 ();
 FILLER_ASAP7_75t_R FILLER_49_364 ();
 FILLER_ASAP7_75t_R FILLER_49_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_371 ();
 DECAPx1_ASAP7_75t_R FILLER_49_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_393 ();
 DECAPx4_ASAP7_75t_R FILLER_49_397 ();
 FILLER_ASAP7_75t_R FILLER_49_407 ();
 FILLER_ASAP7_75t_R FILLER_49_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_417 ();
 FILLER_ASAP7_75t_R FILLER_49_424 ();
 FILLER_ASAP7_75t_R FILLER_49_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_464 ();
 FILLER_ASAP7_75t_R FILLER_49_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_513 ();
 DECAPx6_ASAP7_75t_R FILLER_49_557 ();
 FILLER_ASAP7_75t_R FILLER_49_571 ();
 DECAPx1_ASAP7_75t_R FILLER_49_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_580 ();
 DECAPx6_ASAP7_75t_R FILLER_49_587 ();
 FILLER_ASAP7_75t_R FILLER_49_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_603 ();
 FILLER_ASAP7_75t_R FILLER_49_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_613 ();
 FILLER_ASAP7_75t_R FILLER_49_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_635 ();
 DECAPx1_ASAP7_75t_R FILLER_49_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_654 ();
 DECAPx1_ASAP7_75t_R FILLER_49_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_693 ();
 DECAPx2_ASAP7_75t_R FILLER_49_708 ();
 DECAPx6_ASAP7_75t_R FILLER_49_722 ();
 FILLER_ASAP7_75t_R FILLER_49_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_738 ();
 DECAPx1_ASAP7_75t_R FILLER_49_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_770 ();
 DECAPx1_ASAP7_75t_R FILLER_49_807 ();
 FILLER_ASAP7_75t_R FILLER_49_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_824 ();
 FILLER_ASAP7_75t_R FILLER_49_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_830 ();
 DECAPx6_ASAP7_75t_R FILLER_49_844 ();
 DECAPx2_ASAP7_75t_R FILLER_49_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_864 ();
 DECAPx1_ASAP7_75t_R FILLER_49_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_879 ();
 FILLER_ASAP7_75t_R FILLER_49_890 ();
 DECAPx2_ASAP7_75t_R FILLER_49_895 ();
 DECAPx1_ASAP7_75t_R FILLER_49_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_913 ();
 DECAPx2_ASAP7_75t_R FILLER_49_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_923 ();
 DECAPx2_ASAP7_75t_R FILLER_49_926 ();
 DECAPx1_ASAP7_75t_R FILLER_49_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_942 ();
 FILLER_ASAP7_75t_R FILLER_49_953 ();
 DECAPx10_ASAP7_75t_R FILLER_49_963 ();
 FILLER_ASAP7_75t_R FILLER_49_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_987 ();
 FILLER_ASAP7_75t_R FILLER_49_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1055 ();
 FILLER_ASAP7_75t_R FILLER_49_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1063 ();
 FILLER_ASAP7_75t_R FILLER_49_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1126 ();
 FILLER_ASAP7_75t_R FILLER_49_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1175 ();
 FILLER_ASAP7_75t_R FILLER_49_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1201 ();
 DECAPx4_ASAP7_75t_R FILLER_49_1214 ();
 DECAPx6_ASAP7_75t_R FILLER_49_1243 ();
 FILLER_ASAP7_75t_R FILLER_49_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1337 ();
 DECAPx6_ASAP7_75t_R FILLER_49_1359 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1373 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1379 ();
 DECAPx10_ASAP7_75t_R FILLER_50_2 ();
 DECAPx10_ASAP7_75t_R FILLER_50_24 ();
 DECAPx10_ASAP7_75t_R FILLER_50_46 ();
 DECAPx10_ASAP7_75t_R FILLER_50_68 ();
 DECAPx10_ASAP7_75t_R FILLER_50_90 ();
 DECAPx10_ASAP7_75t_R FILLER_50_112 ();
 DECAPx10_ASAP7_75t_R FILLER_50_134 ();
 DECAPx2_ASAP7_75t_R FILLER_50_156 ();
 DECAPx2_ASAP7_75t_R FILLER_50_192 ();
 FILLER_ASAP7_75t_R FILLER_50_198 ();
 DECAPx10_ASAP7_75t_R FILLER_50_212 ();
 DECAPx2_ASAP7_75t_R FILLER_50_234 ();
 DECAPx1_ASAP7_75t_R FILLER_50_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_286 ();
 FILLER_ASAP7_75t_R FILLER_50_293 ();
 DECAPx2_ASAP7_75t_R FILLER_50_299 ();
 FILLER_ASAP7_75t_R FILLER_50_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_307 ();
 FILLER_ASAP7_75t_R FILLER_50_323 ();
 FILLER_ASAP7_75t_R FILLER_50_329 ();
 FILLER_ASAP7_75t_R FILLER_50_349 ();
 FILLER_ASAP7_75t_R FILLER_50_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_379 ();
 DECAPx2_ASAP7_75t_R FILLER_50_410 ();
 FILLER_ASAP7_75t_R FILLER_50_416 ();
 DECAPx2_ASAP7_75t_R FILLER_50_424 ();
 FILLER_ASAP7_75t_R FILLER_50_430 ();
 DECAPx1_ASAP7_75t_R FILLER_50_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_439 ();
 DECAPx6_ASAP7_75t_R FILLER_50_446 ();
 FILLER_ASAP7_75t_R FILLER_50_460 ();
 DECAPx2_ASAP7_75t_R FILLER_50_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_521 ();
 DECAPx4_ASAP7_75t_R FILLER_50_528 ();
 FILLER_ASAP7_75t_R FILLER_50_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_540 ();
 DECAPx6_ASAP7_75t_R FILLER_50_544 ();
 FILLER_ASAP7_75t_R FILLER_50_558 ();
 FILLER_ASAP7_75t_R FILLER_50_571 ();
 DECAPx2_ASAP7_75t_R FILLER_50_576 ();
 FILLER_ASAP7_75t_R FILLER_50_582 ();
 DECAPx10_ASAP7_75t_R FILLER_50_598 ();
 FILLER_ASAP7_75t_R FILLER_50_620 ();
 DECAPx1_ASAP7_75t_R FILLER_50_639 ();
 DECAPx2_ASAP7_75t_R FILLER_50_657 ();
 DECAPx4_ASAP7_75t_R FILLER_50_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_685 ();
 DECAPx6_ASAP7_75t_R FILLER_50_700 ();
 DECAPx6_ASAP7_75t_R FILLER_50_722 ();
 DECAPx1_ASAP7_75t_R FILLER_50_736 ();
 DECAPx4_ASAP7_75t_R FILLER_50_746 ();
 DECAPx4_ASAP7_75t_R FILLER_50_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_772 ();
 DECAPx2_ASAP7_75t_R FILLER_50_780 ();
 DECAPx6_ASAP7_75t_R FILLER_50_789 ();
 DECAPx2_ASAP7_75t_R FILLER_50_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_809 ();
 DECAPx2_ASAP7_75t_R FILLER_50_836 ();
 FILLER_ASAP7_75t_R FILLER_50_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_844 ();
 DECAPx4_ASAP7_75t_R FILLER_50_871 ();
 FILLER_ASAP7_75t_R FILLER_50_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_883 ();
 DECAPx6_ASAP7_75t_R FILLER_50_892 ();
 DECAPx1_ASAP7_75t_R FILLER_50_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_910 ();
 FILLER_ASAP7_75t_R FILLER_50_937 ();
 DECAPx10_ASAP7_75t_R FILLER_50_949 ();
 DECAPx10_ASAP7_75t_R FILLER_50_971 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1041 ();
 FILLER_ASAP7_75t_R FILLER_50_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1124 ();
 FILLER_ASAP7_75t_R FILLER_50_1130 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1154 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1222 ();
 FILLER_ASAP7_75t_R FILLER_50_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1246 ();
 FILLER_ASAP7_75t_R FILLER_50_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_51_2 ();
 DECAPx10_ASAP7_75t_R FILLER_51_24 ();
 DECAPx10_ASAP7_75t_R FILLER_51_46 ();
 DECAPx10_ASAP7_75t_R FILLER_51_68 ();
 DECAPx10_ASAP7_75t_R FILLER_51_90 ();
 DECAPx10_ASAP7_75t_R FILLER_51_112 ();
 DECAPx10_ASAP7_75t_R FILLER_51_134 ();
 DECAPx2_ASAP7_75t_R FILLER_51_156 ();
 FILLER_ASAP7_75t_R FILLER_51_162 ();
 DECAPx2_ASAP7_75t_R FILLER_51_173 ();
 FILLER_ASAP7_75t_R FILLER_51_179 ();
 DECAPx2_ASAP7_75t_R FILLER_51_187 ();
 FILLER_ASAP7_75t_R FILLER_51_193 ();
 FILLER_ASAP7_75t_R FILLER_51_221 ();
 DECAPx2_ASAP7_75t_R FILLER_51_229 ();
 FILLER_ASAP7_75t_R FILLER_51_235 ();
 DECAPx4_ASAP7_75t_R FILLER_51_263 ();
 FILLER_ASAP7_75t_R FILLER_51_273 ();
 DECAPx1_ASAP7_75t_R FILLER_51_301 ();
 DECAPx4_ASAP7_75t_R FILLER_51_363 ();
 FILLER_ASAP7_75t_R FILLER_51_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_375 ();
 DECAPx2_ASAP7_75t_R FILLER_51_414 ();
 DECAPx6_ASAP7_75t_R FILLER_51_446 ();
 DECAPx1_ASAP7_75t_R FILLER_51_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_464 ();
 DECAPx10_ASAP7_75t_R FILLER_51_471 ();
 DECAPx2_ASAP7_75t_R FILLER_51_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_499 ();
 DECAPx4_ASAP7_75t_R FILLER_51_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_516 ();
 DECAPx4_ASAP7_75t_R FILLER_51_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_537 ();
 DECAPx2_ASAP7_75t_R FILLER_51_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_596 ();
 DECAPx2_ASAP7_75t_R FILLER_51_603 ();
 FILLER_ASAP7_75t_R FILLER_51_609 ();
 DECAPx1_ASAP7_75t_R FILLER_51_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_626 ();
 DECAPx1_ASAP7_75t_R FILLER_51_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_634 ();
 DECAPx4_ASAP7_75t_R FILLER_51_638 ();
 FILLER_ASAP7_75t_R FILLER_51_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_650 ();
 DECAPx10_ASAP7_75t_R FILLER_51_661 ();
 DECAPx2_ASAP7_75t_R FILLER_51_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_689 ();
 DECAPx4_ASAP7_75t_R FILLER_51_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_712 ();
 DECAPx1_ASAP7_75t_R FILLER_51_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_725 ();
 DECAPx2_ASAP7_75t_R FILLER_51_762 ();
 FILLER_ASAP7_75t_R FILLER_51_768 ();
 DECAPx6_ASAP7_75t_R FILLER_51_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_793 ();
 DECAPx6_ASAP7_75t_R FILLER_51_820 ();
 DECAPx2_ASAP7_75t_R FILLER_51_834 ();
 DECAPx2_ASAP7_75t_R FILLER_51_853 ();
 DECAPx10_ASAP7_75t_R FILLER_51_862 ();
 DECAPx10_ASAP7_75t_R FILLER_51_884 ();
 DECAPx2_ASAP7_75t_R FILLER_51_906 ();
 FILLER_ASAP7_75t_R FILLER_51_912 ();
 FILLER_ASAP7_75t_R FILLER_51_922 ();
 DECAPx6_ASAP7_75t_R FILLER_51_929 ();
 DECAPx2_ASAP7_75t_R FILLER_51_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_956 ();
 DECAPx6_ASAP7_75t_R FILLER_51_989 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1020 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1041 ();
 FILLER_ASAP7_75t_R FILLER_51_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1069 ();
 FILLER_ASAP7_75t_R FILLER_51_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1085 ();
 FILLER_ASAP7_75t_R FILLER_51_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1163 ();
 DECAPx4_ASAP7_75t_R FILLER_51_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1194 ();
 FILLER_ASAP7_75t_R FILLER_51_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1229 ();
 FILLER_ASAP7_75t_R FILLER_51_1235 ();
 DECAPx4_ASAP7_75t_R FILLER_51_1247 ();
 FILLER_ASAP7_75t_R FILLER_51_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1354 ();
 DECAPx4_ASAP7_75t_R FILLER_51_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_52_2 ();
 DECAPx10_ASAP7_75t_R FILLER_52_24 ();
 DECAPx10_ASAP7_75t_R FILLER_52_46 ();
 DECAPx10_ASAP7_75t_R FILLER_52_68 ();
 DECAPx10_ASAP7_75t_R FILLER_52_90 ();
 DECAPx10_ASAP7_75t_R FILLER_52_112 ();
 DECAPx6_ASAP7_75t_R FILLER_52_134 ();
 FILLER_ASAP7_75t_R FILLER_52_148 ();
 DECAPx4_ASAP7_75t_R FILLER_52_180 ();
 FILLER_ASAP7_75t_R FILLER_52_190 ();
 DECAPx1_ASAP7_75t_R FILLER_52_198 ();
 FILLER_ASAP7_75t_R FILLER_52_208 ();
 FILLER_ASAP7_75t_R FILLER_52_213 ();
 FILLER_ASAP7_75t_R FILLER_52_219 ();
 DECAPx1_ASAP7_75t_R FILLER_52_247 ();
 DECAPx4_ASAP7_75t_R FILLER_52_254 ();
 DECAPx1_ASAP7_75t_R FILLER_52_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_283 ();
 FILLER_ASAP7_75t_R FILLER_52_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_295 ();
 DECAPx4_ASAP7_75t_R FILLER_52_322 ();
 FILLER_ASAP7_75t_R FILLER_52_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_350 ();
 DECAPx2_ASAP7_75t_R FILLER_52_355 ();
 FILLER_ASAP7_75t_R FILLER_52_361 ();
 FILLER_ASAP7_75t_R FILLER_52_372 ();
 DECAPx10_ASAP7_75t_R FILLER_52_378 ();
 FILLER_ASAP7_75t_R FILLER_52_400 ();
 DECAPx2_ASAP7_75t_R FILLER_52_428 ();
 FILLER_ASAP7_75t_R FILLER_52_434 ();
 DECAPx4_ASAP7_75t_R FILLER_52_464 ();
 FILLER_ASAP7_75t_R FILLER_52_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_503 ();
 DECAPx4_ASAP7_75t_R FILLER_52_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_520 ();
 DECAPx4_ASAP7_75t_R FILLER_52_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_535 ();
 DECAPx2_ASAP7_75t_R FILLER_52_550 ();
 FILLER_ASAP7_75t_R FILLER_52_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_558 ();
 DECAPx6_ASAP7_75t_R FILLER_52_566 ();
 FILLER_ASAP7_75t_R FILLER_52_580 ();
 FILLER_ASAP7_75t_R FILLER_52_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_622 ();
 DECAPx6_ASAP7_75t_R FILLER_52_634 ();
 DECAPx1_ASAP7_75t_R FILLER_52_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_662 ();
 DECAPx6_ASAP7_75t_R FILLER_52_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_691 ();
 DECAPx2_ASAP7_75t_R FILLER_52_704 ();
 FILLER_ASAP7_75t_R FILLER_52_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_712 ();
 DECAPx2_ASAP7_75t_R FILLER_52_721 ();
 FILLER_ASAP7_75t_R FILLER_52_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_729 ();
 FILLER_ASAP7_75t_R FILLER_52_738 ();
 DECAPx4_ASAP7_75t_R FILLER_52_743 ();
 FILLER_ASAP7_75t_R FILLER_52_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_802 ();
 DECAPx4_ASAP7_75t_R FILLER_52_813 ();
 DECAPx10_ASAP7_75t_R FILLER_52_849 ();
 DECAPx1_ASAP7_75t_R FILLER_52_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_875 ();
 DECAPx2_ASAP7_75t_R FILLER_52_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_914 ();
 DECAPx1_ASAP7_75t_R FILLER_52_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_947 ();
 DECAPx1_ASAP7_75t_R FILLER_52_974 ();
 DECAPx2_ASAP7_75t_R FILLER_52_999 ();
 FILLER_ASAP7_75t_R FILLER_52_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1013 ();
 FILLER_ASAP7_75t_R FILLER_52_1027 ();
 FILLER_ASAP7_75t_R FILLER_52_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1063 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1070 ();
 FILLER_ASAP7_75t_R FILLER_52_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1086 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1115 ();
 FILLER_ASAP7_75t_R FILLER_52_1127 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1153 ();
 FILLER_ASAP7_75t_R FILLER_52_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1225 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1250 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1264 ();
 FILLER_ASAP7_75t_R FILLER_52_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1345 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1367 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_53_2 ();
 DECAPx10_ASAP7_75t_R FILLER_53_24 ();
 DECAPx10_ASAP7_75t_R FILLER_53_46 ();
 DECAPx10_ASAP7_75t_R FILLER_53_68 ();
 DECAPx10_ASAP7_75t_R FILLER_53_90 ();
 DECAPx10_ASAP7_75t_R FILLER_53_112 ();
 DECAPx10_ASAP7_75t_R FILLER_53_134 ();
 DECAPx2_ASAP7_75t_R FILLER_53_156 ();
 FILLER_ASAP7_75t_R FILLER_53_162 ();
 DECAPx2_ASAP7_75t_R FILLER_53_170 ();
 FILLER_ASAP7_75t_R FILLER_53_176 ();
 DECAPx6_ASAP7_75t_R FILLER_53_204 ();
 DECAPx2_ASAP7_75t_R FILLER_53_218 ();
 DECAPx2_ASAP7_75t_R FILLER_53_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_239 ();
 DECAPx10_ASAP7_75t_R FILLER_53_244 ();
 DECAPx10_ASAP7_75t_R FILLER_53_266 ();
 DECAPx2_ASAP7_75t_R FILLER_53_288 ();
 FILLER_ASAP7_75t_R FILLER_53_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_309 ();
 DECAPx10_ASAP7_75t_R FILLER_53_313 ();
 DECAPx6_ASAP7_75t_R FILLER_53_335 ();
 DECAPx1_ASAP7_75t_R FILLER_53_349 ();
 FILLER_ASAP7_75t_R FILLER_53_379 ();
 FILLER_ASAP7_75t_R FILLER_53_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_395 ();
 DECAPx1_ASAP7_75t_R FILLER_53_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_403 ();
 DECAPx1_ASAP7_75t_R FILLER_53_408 ();
 FILLER_ASAP7_75t_R FILLER_53_418 ();
 DECAPx1_ASAP7_75t_R FILLER_53_430 ();
 FILLER_ASAP7_75t_R FILLER_53_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_449 ();
 FILLER_ASAP7_75t_R FILLER_53_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_526 ();
 DECAPx2_ASAP7_75t_R FILLER_53_547 ();
 DECAPx4_ASAP7_75t_R FILLER_53_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_577 ();
 DECAPx10_ASAP7_75t_R FILLER_53_581 ();
 FILLER_ASAP7_75t_R FILLER_53_603 ();
 DECAPx2_ASAP7_75t_R FILLER_53_614 ();
 DECAPx2_ASAP7_75t_R FILLER_53_634 ();
 DECAPx2_ASAP7_75t_R FILLER_53_654 ();
 DECAPx1_ASAP7_75t_R FILLER_53_677 ();
 DECAPx6_ASAP7_75t_R FILLER_53_695 ();
 FILLER_ASAP7_75t_R FILLER_53_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_711 ();
 DECAPx6_ASAP7_75t_R FILLER_53_730 ();
 DECAPx1_ASAP7_75t_R FILLER_53_744 ();
 FILLER_ASAP7_75t_R FILLER_53_761 ();
 DECAPx2_ASAP7_75t_R FILLER_53_773 ();
 DECAPx4_ASAP7_75t_R FILLER_53_799 ();
 FILLER_ASAP7_75t_R FILLER_53_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_838 ();
 FILLER_ASAP7_75t_R FILLER_53_846 ();
 DECAPx2_ASAP7_75t_R FILLER_53_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_913 ();
 DECAPx2_ASAP7_75t_R FILLER_53_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_923 ();
 DECAPx10_ASAP7_75t_R FILLER_53_926 ();
 DECAPx4_ASAP7_75t_R FILLER_53_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_958 ();
 DECAPx6_ASAP7_75t_R FILLER_53_969 ();
 DECAPx1_ASAP7_75t_R FILLER_53_983 ();
 FILLER_ASAP7_75t_R FILLER_53_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_995 ();
 FILLER_ASAP7_75t_R FILLER_53_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_53_1042 ();
 FILLER_ASAP7_75t_R FILLER_53_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1058 ();
 FILLER_ASAP7_75t_R FILLER_53_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1081 ();
 DECAPx4_ASAP7_75t_R FILLER_53_1108 ();
 FILLER_ASAP7_75t_R FILLER_53_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1176 ();
 FILLER_ASAP7_75t_R FILLER_53_1182 ();
 DECAPx6_ASAP7_75t_R FILLER_53_1196 ();
 FILLER_ASAP7_75t_R FILLER_53_1210 ();
 DECAPx1_ASAP7_75t_R FILLER_53_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1345 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1367 ();
 FILLER_ASAP7_75t_R FILLER_53_1389 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_54_2 ();
 DECAPx10_ASAP7_75t_R FILLER_54_24 ();
 DECAPx10_ASAP7_75t_R FILLER_54_46 ();
 DECAPx10_ASAP7_75t_R FILLER_54_68 ();
 DECAPx10_ASAP7_75t_R FILLER_54_90 ();
 DECAPx10_ASAP7_75t_R FILLER_54_112 ();
 DECAPx6_ASAP7_75t_R FILLER_54_134 ();
 DECAPx2_ASAP7_75t_R FILLER_54_148 ();
 DECAPx4_ASAP7_75t_R FILLER_54_180 ();
 FILLER_ASAP7_75t_R FILLER_54_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_195 ();
 FILLER_ASAP7_75t_R FILLER_54_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_210 ();
 DECAPx6_ASAP7_75t_R FILLER_54_217 ();
 FILLER_ASAP7_75t_R FILLER_54_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_233 ();
 FILLER_ASAP7_75t_R FILLER_54_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_262 ();
 DECAPx6_ASAP7_75t_R FILLER_54_272 ();
 DECAPx6_ASAP7_75t_R FILLER_54_301 ();
 DECAPx1_ASAP7_75t_R FILLER_54_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_319 ();
 DECAPx6_ASAP7_75t_R FILLER_54_332 ();
 FILLER_ASAP7_75t_R FILLER_54_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_348 ();
 DECAPx2_ASAP7_75t_R FILLER_54_373 ();
 FILLER_ASAP7_75t_R FILLER_54_379 ();
 DECAPx2_ASAP7_75t_R FILLER_54_387 ();
 FILLER_ASAP7_75t_R FILLER_54_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_395 ();
 DECAPx6_ASAP7_75t_R FILLER_54_399 ();
 DECAPx1_ASAP7_75t_R FILLER_54_413 ();
 DECAPx4_ASAP7_75t_R FILLER_54_426 ();
 FILLER_ASAP7_75t_R FILLER_54_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_438 ();
 DECAPx4_ASAP7_75t_R FILLER_54_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_455 ();
 FILLER_ASAP7_75t_R FILLER_54_460 ();
 FILLER_ASAP7_75t_R FILLER_54_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_472 ();
 FILLER_ASAP7_75t_R FILLER_54_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_478 ();
 DECAPx4_ASAP7_75t_R FILLER_54_489 ();
 FILLER_ASAP7_75t_R FILLER_54_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_501 ();
 DECAPx2_ASAP7_75t_R FILLER_54_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_514 ();
 DECAPx6_ASAP7_75t_R FILLER_54_518 ();
 DECAPx2_ASAP7_75t_R FILLER_54_532 ();
 DECAPx1_ASAP7_75t_R FILLER_54_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_554 ();
 DECAPx2_ASAP7_75t_R FILLER_54_569 ();
 FILLER_ASAP7_75t_R FILLER_54_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_577 ();
 DECAPx6_ASAP7_75t_R FILLER_54_620 ();
 FILLER_ASAP7_75t_R FILLER_54_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_636 ();
 DECAPx2_ASAP7_75t_R FILLER_54_654 ();
 FILLER_ASAP7_75t_R FILLER_54_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_662 ();
 FILLER_ASAP7_75t_R FILLER_54_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_668 ();
 FILLER_ASAP7_75t_R FILLER_54_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_685 ();
 DECAPx1_ASAP7_75t_R FILLER_54_702 ();
 DECAPx1_ASAP7_75t_R FILLER_54_754 ();
 FILLER_ASAP7_75t_R FILLER_54_768 ();
 DECAPx4_ASAP7_75t_R FILLER_54_790 ();
 FILLER_ASAP7_75t_R FILLER_54_800 ();
 DECAPx1_ASAP7_75t_R FILLER_54_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_816 ();
 FILLER_ASAP7_75t_R FILLER_54_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_826 ();
 DECAPx2_ASAP7_75t_R FILLER_54_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_836 ();
 FILLER_ASAP7_75t_R FILLER_54_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_848 ();
 DECAPx6_ASAP7_75t_R FILLER_54_881 ();
 FILLER_ASAP7_75t_R FILLER_54_895 ();
 DECAPx4_ASAP7_75t_R FILLER_54_926 ();
 FILLER_ASAP7_75t_R FILLER_54_936 ();
 DECAPx2_ASAP7_75t_R FILLER_54_951 ();
 FILLER_ASAP7_75t_R FILLER_54_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_988 ();
 DECAPx4_ASAP7_75t_R FILLER_54_997 ();
 FILLER_ASAP7_75t_R FILLER_54_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_54_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1042 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1107 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1148 ();
 FILLER_ASAP7_75t_R FILLER_54_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1182 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1231 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1247 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_55_2 ();
 DECAPx10_ASAP7_75t_R FILLER_55_24 ();
 DECAPx10_ASAP7_75t_R FILLER_55_46 ();
 DECAPx10_ASAP7_75t_R FILLER_55_68 ();
 DECAPx10_ASAP7_75t_R FILLER_55_90 ();
 DECAPx10_ASAP7_75t_R FILLER_55_112 ();
 DECAPx6_ASAP7_75t_R FILLER_55_134 ();
 FILLER_ASAP7_75t_R FILLER_55_148 ();
 DECAPx2_ASAP7_75t_R FILLER_55_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_159 ();
 FILLER_ASAP7_75t_R FILLER_55_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_168 ();
 DECAPx6_ASAP7_75t_R FILLER_55_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_198 ();
 FILLER_ASAP7_75t_R FILLER_55_225 ();
 FILLER_ASAP7_75t_R FILLER_55_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_281 ();
 DECAPx1_ASAP7_75t_R FILLER_55_308 ();
 FILLER_ASAP7_75t_R FILLER_55_315 ();
 DECAPx6_ASAP7_75t_R FILLER_55_343 ();
 FILLER_ASAP7_75t_R FILLER_55_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_359 ();
 FILLER_ASAP7_75t_R FILLER_55_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_380 ();
 DECAPx2_ASAP7_75t_R FILLER_55_407 ();
 DECAPx6_ASAP7_75t_R FILLER_55_419 ();
 DECAPx2_ASAP7_75t_R FILLER_55_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_439 ();
 FILLER_ASAP7_75t_R FILLER_55_452 ();
 DECAPx10_ASAP7_75t_R FILLER_55_457 ();
 DECAPx1_ASAP7_75t_R FILLER_55_479 ();
 DECAPx1_ASAP7_75t_R FILLER_55_489 ();
 DECAPx2_ASAP7_75t_R FILLER_55_496 ();
 FILLER_ASAP7_75t_R FILLER_55_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_522 ();
 DECAPx1_ASAP7_75t_R FILLER_55_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_536 ();
 FILLER_ASAP7_75t_R FILLER_55_547 ();
 FILLER_ASAP7_75t_R FILLER_55_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_554 ();
 DECAPx1_ASAP7_75t_R FILLER_55_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_576 ();
 DECAPx10_ASAP7_75t_R FILLER_55_591 ();
 DECAPx6_ASAP7_75t_R FILLER_55_613 ();
 FILLER_ASAP7_75t_R FILLER_55_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_629 ();
 DECAPx6_ASAP7_75t_R FILLER_55_647 ();
 FILLER_ASAP7_75t_R FILLER_55_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_663 ();
 FILLER_ASAP7_75t_R FILLER_55_667 ();
 DECAPx4_ASAP7_75t_R FILLER_55_683 ();
 FILLER_ASAP7_75t_R FILLER_55_693 ();
 DECAPx1_ASAP7_75t_R FILLER_55_703 ();
 DECAPx6_ASAP7_75t_R FILLER_55_717 ();
 FILLER_ASAP7_75t_R FILLER_55_731 ();
 FILLER_ASAP7_75t_R FILLER_55_749 ();
 DECAPx10_ASAP7_75t_R FILLER_55_754 ();
 DECAPx10_ASAP7_75t_R FILLER_55_776 ();
 DECAPx2_ASAP7_75t_R FILLER_55_798 ();
 FILLER_ASAP7_75t_R FILLER_55_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_816 ();
 DECAPx10_ASAP7_75t_R FILLER_55_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_845 ();
 DECAPx2_ASAP7_75t_R FILLER_55_852 ();
 FILLER_ASAP7_75t_R FILLER_55_858 ();
 DECAPx2_ASAP7_75t_R FILLER_55_886 ();
 FILLER_ASAP7_75t_R FILLER_55_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_894 ();
 FILLER_ASAP7_75t_R FILLER_55_898 ();
 DECAPx4_ASAP7_75t_R FILLER_55_903 ();
 FILLER_ASAP7_75t_R FILLER_55_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_915 ();
 FILLER_ASAP7_75t_R FILLER_55_922 ();
 DECAPx2_ASAP7_75t_R FILLER_55_926 ();
 FILLER_ASAP7_75t_R FILLER_55_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_934 ();
 DECAPx2_ASAP7_75t_R FILLER_55_961 ();
 DECAPx6_ASAP7_75t_R FILLER_55_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1014 ();
 FILLER_ASAP7_75t_R FILLER_55_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1023 ();
 DECAPx6_ASAP7_75t_R FILLER_55_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_55_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_55_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1120 ();
 FILLER_ASAP7_75t_R FILLER_55_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1129 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1140 ();
 FILLER_ASAP7_75t_R FILLER_55_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1199 ();
 DECAPx6_ASAP7_75t_R FILLER_55_1221 ();
 FILLER_ASAP7_75t_R FILLER_55_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1244 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1350 ();
 DECAPx6_ASAP7_75t_R FILLER_55_1372 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1386 ();
 DECAPx10_ASAP7_75t_R FILLER_56_2 ();
 DECAPx10_ASAP7_75t_R FILLER_56_24 ();
 DECAPx10_ASAP7_75t_R FILLER_56_46 ();
 DECAPx10_ASAP7_75t_R FILLER_56_68 ();
 DECAPx10_ASAP7_75t_R FILLER_56_90 ();
 DECAPx10_ASAP7_75t_R FILLER_56_112 ();
 FILLER_ASAP7_75t_R FILLER_56_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_162 ();
 FILLER_ASAP7_75t_R FILLER_56_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_175 ();
 DECAPx4_ASAP7_75t_R FILLER_56_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_212 ();
 DECAPx6_ASAP7_75t_R FILLER_56_242 ();
 FILLER_ASAP7_75t_R FILLER_56_262 ();
 FILLER_ASAP7_75t_R FILLER_56_290 ();
 DECAPx2_ASAP7_75t_R FILLER_56_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_330 ();
 DECAPx6_ASAP7_75t_R FILLER_56_343 ();
 DECAPx1_ASAP7_75t_R FILLER_56_357 ();
 DECAPx6_ASAP7_75t_R FILLER_56_367 ();
 DECAPx10_ASAP7_75t_R FILLER_56_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_435 ();
 DECAPx2_ASAP7_75t_R FILLER_56_464 ();
 FILLER_ASAP7_75t_R FILLER_56_470 ();
 DECAPx6_ASAP7_75t_R FILLER_56_504 ();
 DECAPx1_ASAP7_75t_R FILLER_56_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_552 ();
 DECAPx1_ASAP7_75t_R FILLER_56_567 ();
 DECAPx2_ASAP7_75t_R FILLER_56_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_614 ();
 DECAPx1_ASAP7_75t_R FILLER_56_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_626 ();
 DECAPx1_ASAP7_75t_R FILLER_56_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_662 ();
 DECAPx6_ASAP7_75t_R FILLER_56_677 ();
 FILLER_ASAP7_75t_R FILLER_56_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_693 ();
 DECAPx1_ASAP7_75t_R FILLER_56_702 ();
 DECAPx4_ASAP7_75t_R FILLER_56_724 ();
 FILLER_ASAP7_75t_R FILLER_56_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_736 ();
 DECAPx1_ASAP7_75t_R FILLER_56_783 ();
 DECAPx2_ASAP7_75t_R FILLER_56_795 ();
 DECAPx2_ASAP7_75t_R FILLER_56_811 ();
 FILLER_ASAP7_75t_R FILLER_56_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_819 ();
 DECAPx1_ASAP7_75t_R FILLER_56_846 ();
 DECAPx2_ASAP7_75t_R FILLER_56_858 ();
 DECAPx4_ASAP7_75t_R FILLER_56_867 ();
 FILLER_ASAP7_75t_R FILLER_56_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_879 ();
 FILLER_ASAP7_75t_R FILLER_56_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_908 ();
 DECAPx1_ASAP7_75t_R FILLER_56_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_920 ();
 DECAPx2_ASAP7_75t_R FILLER_56_935 ();
 FILLER_ASAP7_75t_R FILLER_56_941 ();
 DECAPx4_ASAP7_75t_R FILLER_56_952 ();
 FILLER_ASAP7_75t_R FILLER_56_962 ();
 FILLER_ASAP7_75t_R FILLER_56_971 ();
 DECAPx1_ASAP7_75t_R FILLER_56_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_980 ();
 DECAPx1_ASAP7_75t_R FILLER_56_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_988 ();
 FILLER_ASAP7_75t_R FILLER_56_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_56_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_56_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1148 ();
 FILLER_ASAP7_75t_R FILLER_56_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1222 ();
 FILLER_ASAP7_75t_R FILLER_56_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1230 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1258 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1370 ();
 FILLER_ASAP7_75t_R FILLER_56_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_56_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_57_2 ();
 DECAPx10_ASAP7_75t_R FILLER_57_24 ();
 DECAPx10_ASAP7_75t_R FILLER_57_46 ();
 DECAPx10_ASAP7_75t_R FILLER_57_68 ();
 DECAPx10_ASAP7_75t_R FILLER_57_90 ();
 DECAPx10_ASAP7_75t_R FILLER_57_112 ();
 DECAPx10_ASAP7_75t_R FILLER_57_134 ();
 DECAPx1_ASAP7_75t_R FILLER_57_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_160 ();
 DECAPx6_ASAP7_75t_R FILLER_57_173 ();
 DECAPx6_ASAP7_75t_R FILLER_57_202 ();
 DECAPx2_ASAP7_75t_R FILLER_57_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_229 ();
 DECAPx10_ASAP7_75t_R FILLER_57_233 ();
 DECAPx2_ASAP7_75t_R FILLER_57_255 ();
 FILLER_ASAP7_75t_R FILLER_57_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_263 ();
 FILLER_ASAP7_75t_R FILLER_57_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_278 ();
 DECAPx2_ASAP7_75t_R FILLER_57_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_315 ();
 DECAPx1_ASAP7_75t_R FILLER_57_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_324 ();
 FILLER_ASAP7_75t_R FILLER_57_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_416 ();
 DECAPx6_ASAP7_75t_R FILLER_57_446 ();
 FILLER_ASAP7_75t_R FILLER_57_460 ();
 DECAPx2_ASAP7_75t_R FILLER_57_488 ();
 FILLER_ASAP7_75t_R FILLER_57_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_496 ();
 DECAPx1_ASAP7_75t_R FILLER_57_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_507 ();
 DECAPx2_ASAP7_75t_R FILLER_57_511 ();
 FILLER_ASAP7_75t_R FILLER_57_517 ();
 DECAPx4_ASAP7_75t_R FILLER_57_550 ();
 FILLER_ASAP7_75t_R FILLER_57_560 ();
 DECAPx6_ASAP7_75t_R FILLER_57_565 ();
 FILLER_ASAP7_75t_R FILLER_57_579 ();
 DECAPx4_ASAP7_75t_R FILLER_57_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_626 ();
 DECAPx6_ASAP7_75t_R FILLER_57_630 ();
 FILLER_ASAP7_75t_R FILLER_57_644 ();
 DECAPx1_ASAP7_75t_R FILLER_57_660 ();
 DECAPx4_ASAP7_75t_R FILLER_57_667 ();
 DECAPx6_ASAP7_75t_R FILLER_57_694 ();
 DECAPx2_ASAP7_75t_R FILLER_57_708 ();
 DECAPx6_ASAP7_75t_R FILLER_57_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_736 ();
 DECAPx10_ASAP7_75t_R FILLER_57_744 ();
 DECAPx2_ASAP7_75t_R FILLER_57_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_772 ();
 FILLER_ASAP7_75t_R FILLER_57_783 ();
 DECAPx4_ASAP7_75t_R FILLER_57_811 ();
 FILLER_ASAP7_75t_R FILLER_57_821 ();
 DECAPx1_ASAP7_75t_R FILLER_57_831 ();
 DECAPx1_ASAP7_75t_R FILLER_57_838 ();
 FILLER_ASAP7_75t_R FILLER_57_848 ();
 FILLER_ASAP7_75t_R FILLER_57_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_860 ();
 FILLER_ASAP7_75t_R FILLER_57_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_869 ();
 DECAPx2_ASAP7_75t_R FILLER_57_873 ();
 FILLER_ASAP7_75t_R FILLER_57_901 ();
 DECAPx1_ASAP7_75t_R FILLER_57_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_940 ();
 DECAPx6_ASAP7_75t_R FILLER_57_967 ();
 FILLER_ASAP7_75t_R FILLER_57_981 ();
 DECAPx2_ASAP7_75t_R FILLER_57_989 ();
 FILLER_ASAP7_75t_R FILLER_57_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1000 ();
 DECAPx4_ASAP7_75t_R FILLER_57_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1025 ();
 FILLER_ASAP7_75t_R FILLER_57_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1036 ();
 FILLER_ASAP7_75t_R FILLER_57_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1056 ();
 DECAPx4_ASAP7_75t_R FILLER_57_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1095 ();
 FILLER_ASAP7_75t_R FILLER_57_1101 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1106 ();
 FILLER_ASAP7_75t_R FILLER_57_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1164 ();
 DECAPx4_ASAP7_75t_R FILLER_57_1171 ();
 FILLER_ASAP7_75t_R FILLER_57_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1203 ();
 FILLER_ASAP7_75t_R FILLER_57_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1356 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_58_2 ();
 DECAPx10_ASAP7_75t_R FILLER_58_24 ();
 DECAPx10_ASAP7_75t_R FILLER_58_46 ();
 DECAPx10_ASAP7_75t_R FILLER_58_68 ();
 DECAPx10_ASAP7_75t_R FILLER_58_90 ();
 DECAPx10_ASAP7_75t_R FILLER_58_112 ();
 DECAPx6_ASAP7_75t_R FILLER_58_134 ();
 DECAPx2_ASAP7_75t_R FILLER_58_148 ();
 DECAPx10_ASAP7_75t_R FILLER_58_184 ();
 DECAPx2_ASAP7_75t_R FILLER_58_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_224 ();
 DECAPx2_ASAP7_75t_R FILLER_58_228 ();
 FILLER_ASAP7_75t_R FILLER_58_266 ();
 FILLER_ASAP7_75t_R FILLER_58_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_300 ();
 DECAPx10_ASAP7_75t_R FILLER_58_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_329 ();
 DECAPx6_ASAP7_75t_R FILLER_58_336 ();
 DECAPx2_ASAP7_75t_R FILLER_58_350 ();
 DECAPx1_ASAP7_75t_R FILLER_58_362 ();
 FILLER_ASAP7_75t_R FILLER_58_401 ();
 DECAPx1_ASAP7_75t_R FILLER_58_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_432 ();
 DECAPx6_ASAP7_75t_R FILLER_58_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_493 ();
 FILLER_ASAP7_75t_R FILLER_58_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_522 ();
 DECAPx4_ASAP7_75t_R FILLER_58_529 ();
 FILLER_ASAP7_75t_R FILLER_58_549 ();
 DECAPx10_ASAP7_75t_R FILLER_58_568 ();
 DECAPx2_ASAP7_75t_R FILLER_58_590 ();
 FILLER_ASAP7_75t_R FILLER_58_596 ();
 FILLER_ASAP7_75t_R FILLER_58_612 ();
 DECAPx6_ASAP7_75t_R FILLER_58_628 ();
 FILLER_ASAP7_75t_R FILLER_58_642 ();
 DECAPx6_ASAP7_75t_R FILLER_58_661 ();
 DECAPx2_ASAP7_75t_R FILLER_58_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_712 ();
 DECAPx2_ASAP7_75t_R FILLER_58_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_729 ();
 FILLER_ASAP7_75t_R FILLER_58_740 ();
 DECAPx2_ASAP7_75t_R FILLER_58_745 ();
 DECAPx1_ASAP7_75t_R FILLER_58_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_799 ();
 DECAPx2_ASAP7_75t_R FILLER_58_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_823 ();
 DECAPx1_ASAP7_75t_R FILLER_58_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_882 ();
 DECAPx1_ASAP7_75t_R FILLER_58_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_893 ();
 DECAPx6_ASAP7_75t_R FILLER_58_900 ();
 FILLER_ASAP7_75t_R FILLER_58_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_916 ();
 DECAPx2_ASAP7_75t_R FILLER_58_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_957 ();
 DECAPx2_ASAP7_75t_R FILLER_58_965 ();
 FILLER_ASAP7_75t_R FILLER_58_997 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1007 ();
 FILLER_ASAP7_75t_R FILLER_58_1029 ();
 FILLER_ASAP7_75t_R FILLER_58_1037 ();
 DECAPx4_ASAP7_75t_R FILLER_58_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1081 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1097 ();
 FILLER_ASAP7_75t_R FILLER_58_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1136 ();
 FILLER_ASAP7_75t_R FILLER_58_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1180 ();
 FILLER_ASAP7_75t_R FILLER_58_1186 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1254 ();
 FILLER_ASAP7_75t_R FILLER_58_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1378 ();
 FILLER_ASAP7_75t_R FILLER_58_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_59_2 ();
 DECAPx10_ASAP7_75t_R FILLER_59_24 ();
 DECAPx10_ASAP7_75t_R FILLER_59_46 ();
 DECAPx10_ASAP7_75t_R FILLER_59_68 ();
 DECAPx10_ASAP7_75t_R FILLER_59_90 ();
 DECAPx4_ASAP7_75t_R FILLER_59_112 ();
 FILLER_ASAP7_75t_R FILLER_59_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_124 ();
 DECAPx4_ASAP7_75t_R FILLER_59_157 ();
 FILLER_ASAP7_75t_R FILLER_59_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_172 ();
 DECAPx1_ASAP7_75t_R FILLER_59_199 ();
 FILLER_ASAP7_75t_R FILLER_59_209 ();
 FILLER_ASAP7_75t_R FILLER_59_237 ();
 FILLER_ASAP7_75t_R FILLER_59_251 ();
 DECAPx1_ASAP7_75t_R FILLER_59_283 ();
 DECAPx1_ASAP7_75t_R FILLER_59_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_297 ();
 DECAPx6_ASAP7_75t_R FILLER_59_324 ();
 DECAPx1_ASAP7_75t_R FILLER_59_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_342 ();
 DECAPx1_ASAP7_75t_R FILLER_59_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_353 ();
 DECAPx6_ASAP7_75t_R FILLER_59_360 ();
 FILLER_ASAP7_75t_R FILLER_59_374 ();
 FILLER_ASAP7_75t_R FILLER_59_412 ();
 DECAPx1_ASAP7_75t_R FILLER_59_426 ();
 FILLER_ASAP7_75t_R FILLER_59_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_438 ();
 FILLER_ASAP7_75t_R FILLER_59_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_453 ();
 DECAPx10_ASAP7_75t_R FILLER_59_457 ();
 FILLER_ASAP7_75t_R FILLER_59_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_481 ();
 DECAPx2_ASAP7_75t_R FILLER_59_488 ();
 FILLER_ASAP7_75t_R FILLER_59_494 ();
 DECAPx6_ASAP7_75t_R FILLER_59_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_516 ();
 DECAPx4_ASAP7_75t_R FILLER_59_521 ();
 DECAPx1_ASAP7_75t_R FILLER_59_534 ();
 DECAPx6_ASAP7_75t_R FILLER_59_544 ();
 DECAPx1_ASAP7_75t_R FILLER_59_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_582 ();
 DECAPx4_ASAP7_75t_R FILLER_59_586 ();
 FILLER_ASAP7_75t_R FILLER_59_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_598 ();
 DECAPx4_ASAP7_75t_R FILLER_59_602 ();
 FILLER_ASAP7_75t_R FILLER_59_629 ();
 DECAPx2_ASAP7_75t_R FILLER_59_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_640 ();
 DECAPx1_ASAP7_75t_R FILLER_59_658 ();
 DECAPx2_ASAP7_75t_R FILLER_59_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_685 ();
 DECAPx2_ASAP7_75t_R FILLER_59_697 ();
 FILLER_ASAP7_75t_R FILLER_59_703 ();
 DECAPx6_ASAP7_75t_R FILLER_59_713 ();
 DECAPx2_ASAP7_75t_R FILLER_59_753 ();
 DECAPx6_ASAP7_75t_R FILLER_59_765 ();
 DECAPx1_ASAP7_75t_R FILLER_59_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_783 ();
 DECAPx4_ASAP7_75t_R FILLER_59_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_808 ();
 DECAPx10_ASAP7_75t_R FILLER_59_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_839 ();
 DECAPx6_ASAP7_75t_R FILLER_59_862 ();
 DECAPx1_ASAP7_75t_R FILLER_59_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_880 ();
 DECAPx2_ASAP7_75t_R FILLER_59_887 ();
 FILLER_ASAP7_75t_R FILLER_59_893 ();
 DECAPx2_ASAP7_75t_R FILLER_59_903 ();
 FILLER_ASAP7_75t_R FILLER_59_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_911 ();
 DECAPx6_ASAP7_75t_R FILLER_59_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_948 ();
 FILLER_ASAP7_75t_R FILLER_59_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_961 ();
 FILLER_ASAP7_75t_R FILLER_59_982 ();
 FILLER_ASAP7_75t_R FILLER_59_993 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1011 ();
 DECAPx6_ASAP7_75t_R FILLER_59_1023 ();
 DECAPx6_ASAP7_75t_R FILLER_59_1055 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1081 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1106 ();
 FILLER_ASAP7_75t_R FILLER_59_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1140 ();
 FILLER_ASAP7_75t_R FILLER_59_1147 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1186 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1193 ();
 DECAPx6_ASAP7_75t_R FILLER_59_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1223 ();
 FILLER_ASAP7_75t_R FILLER_59_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1231 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1235 ();
 FILLER_ASAP7_75t_R FILLER_59_1241 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1340 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1384 ();
 FILLER_ASAP7_75t_R FILLER_59_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_60_2 ();
 DECAPx10_ASAP7_75t_R FILLER_60_24 ();
 DECAPx10_ASAP7_75t_R FILLER_60_46 ();
 DECAPx10_ASAP7_75t_R FILLER_60_68 ();
 DECAPx10_ASAP7_75t_R FILLER_60_90 ();
 DECAPx6_ASAP7_75t_R FILLER_60_112 ();
 FILLER_ASAP7_75t_R FILLER_60_126 ();
 FILLER_ASAP7_75t_R FILLER_60_164 ();
 DECAPx4_ASAP7_75t_R FILLER_60_172 ();
 FILLER_ASAP7_75t_R FILLER_60_182 ();
 DECAPx10_ASAP7_75t_R FILLER_60_225 ();
 FILLER_ASAP7_75t_R FILLER_60_247 ();
 DECAPx4_ASAP7_75t_R FILLER_60_252 ();
 FILLER_ASAP7_75t_R FILLER_60_262 ();
 FILLER_ASAP7_75t_R FILLER_60_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_296 ();
 FILLER_ASAP7_75t_R FILLER_60_310 ();
 FILLER_ASAP7_75t_R FILLER_60_372 ();
 DECAPx1_ASAP7_75t_R FILLER_60_380 ();
 FILLER_ASAP7_75t_R FILLER_60_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_426 ();
 DECAPx2_ASAP7_75t_R FILLER_60_453 ();
 FILLER_ASAP7_75t_R FILLER_60_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_461 ();
 DECAPx2_ASAP7_75t_R FILLER_60_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_476 ();
 DECAPx2_ASAP7_75t_R FILLER_60_506 ();
 DECAPx10_ASAP7_75t_R FILLER_60_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_540 ();
 DECAPx1_ASAP7_75t_R FILLER_60_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_554 ();
 FILLER_ASAP7_75t_R FILLER_60_584 ();
 DECAPx1_ASAP7_75t_R FILLER_60_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_622 ();
 FILLER_ASAP7_75t_R FILLER_60_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_653 ();
 FILLER_ASAP7_75t_R FILLER_60_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_684 ();
 DECAPx2_ASAP7_75t_R FILLER_60_696 ();
 FILLER_ASAP7_75t_R FILLER_60_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_704 ();
 DECAPx4_ASAP7_75t_R FILLER_60_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_723 ();
 DECAPx6_ASAP7_75t_R FILLER_60_732 ();
 DECAPx1_ASAP7_75t_R FILLER_60_746 ();
 FILLER_ASAP7_75t_R FILLER_60_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_758 ();
 DECAPx4_ASAP7_75t_R FILLER_60_771 ();
 FILLER_ASAP7_75t_R FILLER_60_781 ();
 DECAPx1_ASAP7_75t_R FILLER_60_790 ();
 DECAPx1_ASAP7_75t_R FILLER_60_810 ();
 DECAPx1_ASAP7_75t_R FILLER_60_822 ();
 DECAPx10_ASAP7_75t_R FILLER_60_834 ();
 DECAPx6_ASAP7_75t_R FILLER_60_856 ();
 FILLER_ASAP7_75t_R FILLER_60_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_872 ();
 DECAPx2_ASAP7_75t_R FILLER_60_879 ();
 FILLER_ASAP7_75t_R FILLER_60_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_887 ();
 DECAPx2_ASAP7_75t_R FILLER_60_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_925 ();
 DECAPx6_ASAP7_75t_R FILLER_60_932 ();
 FILLER_ASAP7_75t_R FILLER_60_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_948 ();
 DECAPx10_ASAP7_75t_R FILLER_60_975 ();
 DECAPx1_ASAP7_75t_R FILLER_60_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1028 ();
 DECAPx4_ASAP7_75t_R FILLER_60_1053 ();
 FILLER_ASAP7_75t_R FILLER_60_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1100 ();
 FILLER_ASAP7_75t_R FILLER_60_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_60_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_60_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_60_1171 ();
 FILLER_ASAP7_75t_R FILLER_60_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1185 ();
 FILLER_ASAP7_75t_R FILLER_60_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1216 ();
 DECAPx2_ASAP7_75t_R FILLER_60_1251 ();
 FILLER_ASAP7_75t_R FILLER_60_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1370 ();
 FILLER_ASAP7_75t_R FILLER_60_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_61_2 ();
 DECAPx10_ASAP7_75t_R FILLER_61_24 ();
 DECAPx10_ASAP7_75t_R FILLER_61_46 ();
 DECAPx10_ASAP7_75t_R FILLER_61_68 ();
 DECAPx10_ASAP7_75t_R FILLER_61_90 ();
 DECAPx4_ASAP7_75t_R FILLER_61_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_141 ();
 DECAPx1_ASAP7_75t_R FILLER_61_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_160 ();
 DECAPx6_ASAP7_75t_R FILLER_61_190 ();
 DECAPx1_ASAP7_75t_R FILLER_61_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_208 ();
 DECAPx2_ASAP7_75t_R FILLER_61_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_224 ();
 DECAPx2_ASAP7_75t_R FILLER_61_235 ();
 FILLER_ASAP7_75t_R FILLER_61_241 ();
 DECAPx6_ASAP7_75t_R FILLER_61_253 ();
 DECAPx1_ASAP7_75t_R FILLER_61_267 ();
 DECAPx1_ASAP7_75t_R FILLER_61_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_278 ();
 DECAPx6_ASAP7_75t_R FILLER_61_283 ();
 FILLER_ASAP7_75t_R FILLER_61_297 ();
 DECAPx2_ASAP7_75t_R FILLER_61_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_311 ();
 DECAPx2_ASAP7_75t_R FILLER_61_315 ();
 FILLER_ASAP7_75t_R FILLER_61_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_330 ();
 DECAPx4_ASAP7_75t_R FILLER_61_344 ();
 FILLER_ASAP7_75t_R FILLER_61_354 ();
 DECAPx10_ASAP7_75t_R FILLER_61_359 ();
 FILLER_ASAP7_75t_R FILLER_61_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_383 ();
 DECAPx2_ASAP7_75t_R FILLER_61_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_396 ();
 DECAPx6_ASAP7_75t_R FILLER_61_400 ();
 FILLER_ASAP7_75t_R FILLER_61_414 ();
 DECAPx6_ASAP7_75t_R FILLER_61_446 ();
 FILLER_ASAP7_75t_R FILLER_61_460 ();
 DECAPx1_ASAP7_75t_R FILLER_61_497 ();
 DECAPx2_ASAP7_75t_R FILLER_61_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_533 ();
 DECAPx1_ASAP7_75t_R FILLER_61_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_552 ();
 DECAPx4_ASAP7_75t_R FILLER_61_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_566 ();
 DECAPx2_ASAP7_75t_R FILLER_61_573 ();
 FILLER_ASAP7_75t_R FILLER_61_579 ();
 FILLER_ASAP7_75t_R FILLER_61_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_600 ();
 DECAPx6_ASAP7_75t_R FILLER_61_629 ();
 FILLER_ASAP7_75t_R FILLER_61_643 ();
 DECAPx1_ASAP7_75t_R FILLER_61_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_652 ();
 DECAPx2_ASAP7_75t_R FILLER_61_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_665 ();
 DECAPx10_ASAP7_75t_R FILLER_61_675 ();
 DECAPx10_ASAP7_75t_R FILLER_61_697 ();
 DECAPx4_ASAP7_75t_R FILLER_61_719 ();
 FILLER_ASAP7_75t_R FILLER_61_729 ();
 FILLER_ASAP7_75t_R FILLER_61_745 ();
 DECAPx2_ASAP7_75t_R FILLER_61_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_761 ();
 DECAPx2_ASAP7_75t_R FILLER_61_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_780 ();
 DECAPx1_ASAP7_75t_R FILLER_61_807 ();
 DECAPx2_ASAP7_75t_R FILLER_61_819 ();
 FILLER_ASAP7_75t_R FILLER_61_851 ();
 DECAPx2_ASAP7_75t_R FILLER_61_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_873 ();
 DECAPx4_ASAP7_75t_R FILLER_61_900 ();
 FILLER_ASAP7_75t_R FILLER_61_910 ();
 DECAPx10_ASAP7_75t_R FILLER_61_933 ();
 DECAPx1_ASAP7_75t_R FILLER_61_955 ();
 DECAPx1_ASAP7_75t_R FILLER_61_966 ();
 DECAPx10_ASAP7_75t_R FILLER_61_976 ();
 FILLER_ASAP7_75t_R FILLER_61_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1008 ();
 FILLER_ASAP7_75t_R FILLER_61_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_61_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1069 ();
 FILLER_ASAP7_75t_R FILLER_61_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1127 ();
 FILLER_ASAP7_75t_R FILLER_61_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1156 ();
 DECAPx6_ASAP7_75t_R FILLER_61_1168 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1186 ();
 FILLER_ASAP7_75t_R FILLER_61_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1208 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1246 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_62_2 ();
 DECAPx10_ASAP7_75t_R FILLER_62_24 ();
 DECAPx10_ASAP7_75t_R FILLER_62_46 ();
 DECAPx10_ASAP7_75t_R FILLER_62_68 ();
 DECAPx10_ASAP7_75t_R FILLER_62_90 ();
 DECAPx10_ASAP7_75t_R FILLER_62_112 ();
 DECAPx1_ASAP7_75t_R FILLER_62_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_138 ();
 DECAPx4_ASAP7_75t_R FILLER_62_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_152 ();
 DECAPx4_ASAP7_75t_R FILLER_62_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_169 ();
 FILLER_ASAP7_75t_R FILLER_62_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_181 ();
 DECAPx1_ASAP7_75t_R FILLER_62_186 ();
 DECAPx1_ASAP7_75t_R FILLER_62_196 ();
 DECAPx4_ASAP7_75t_R FILLER_62_210 ();
 DECAPx2_ASAP7_75t_R FILLER_62_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_262 ();
 DECAPx6_ASAP7_75t_R FILLER_62_266 ();
 DECAPx1_ASAP7_75t_R FILLER_62_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_284 ();
 DECAPx10_ASAP7_75t_R FILLER_62_288 ();
 DECAPx4_ASAP7_75t_R FILLER_62_310 ();
 FILLER_ASAP7_75t_R FILLER_62_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_322 ();
 DECAPx2_ASAP7_75t_R FILLER_62_329 ();
 FILLER_ASAP7_75t_R FILLER_62_335 ();
 FILLER_ASAP7_75t_R FILLER_62_350 ();
 DECAPx6_ASAP7_75t_R FILLER_62_370 ();
 DECAPx6_ASAP7_75t_R FILLER_62_390 ();
 FILLER_ASAP7_75t_R FILLER_62_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_406 ();
 FILLER_ASAP7_75t_R FILLER_62_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_418 ();
 FILLER_ASAP7_75t_R FILLER_62_445 ();
 DECAPx2_ASAP7_75t_R FILLER_62_453 ();
 DECAPx10_ASAP7_75t_R FILLER_62_473 ();
 DECAPx2_ASAP7_75t_R FILLER_62_495 ();
 FILLER_ASAP7_75t_R FILLER_62_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_503 ();
 DECAPx1_ASAP7_75t_R FILLER_62_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_514 ();
 DECAPx4_ASAP7_75t_R FILLER_62_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_528 ();
 DECAPx2_ASAP7_75t_R FILLER_62_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_551 ();
 DECAPx2_ASAP7_75t_R FILLER_62_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_561 ();
 DECAPx6_ASAP7_75t_R FILLER_62_576 ();
 DECAPx1_ASAP7_75t_R FILLER_62_590 ();
 DECAPx6_ASAP7_75t_R FILLER_62_597 ();
 DECAPx1_ASAP7_75t_R FILLER_62_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_615 ();
 FILLER_ASAP7_75t_R FILLER_62_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_624 ();
 DECAPx10_ASAP7_75t_R FILLER_62_642 ();
 DECAPx10_ASAP7_75t_R FILLER_62_664 ();
 DECAPx2_ASAP7_75t_R FILLER_62_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_719 ();
 FILLER_ASAP7_75t_R FILLER_62_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_732 ();
 DECAPx2_ASAP7_75t_R FILLER_62_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_749 ();
 FILLER_ASAP7_75t_R FILLER_62_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_799 ();
 DECAPx1_ASAP7_75t_R FILLER_62_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_807 ();
 DECAPx6_ASAP7_75t_R FILLER_62_814 ();
 FILLER_ASAP7_75t_R FILLER_62_835 ();
 DECAPx2_ASAP7_75t_R FILLER_62_846 ();
 FILLER_ASAP7_75t_R FILLER_62_852 ();
 FILLER_ASAP7_75t_R FILLER_62_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_869 ();
 DECAPx2_ASAP7_75t_R FILLER_62_891 ();
 DECAPx2_ASAP7_75t_R FILLER_62_911 ();
 FILLER_ASAP7_75t_R FILLER_62_917 ();
 FILLER_ASAP7_75t_R FILLER_62_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_933 ();
 DECAPx6_ASAP7_75t_R FILLER_62_960 ();
 DECAPx1_ASAP7_75t_R FILLER_62_974 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1028 ();
 FILLER_ASAP7_75t_R FILLER_62_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1118 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1132 ();
 FILLER_ASAP7_75t_R FILLER_62_1142 ();
 FILLER_ASAP7_75t_R FILLER_62_1150 ();
 FILLER_ASAP7_75t_R FILLER_62_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1198 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1210 ();
 FILLER_ASAP7_75t_R FILLER_62_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1218 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1246 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1350 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_63_2 ();
 DECAPx10_ASAP7_75t_R FILLER_63_24 ();
 DECAPx10_ASAP7_75t_R FILLER_63_46 ();
 DECAPx10_ASAP7_75t_R FILLER_63_68 ();
 DECAPx10_ASAP7_75t_R FILLER_63_90 ();
 DECAPx4_ASAP7_75t_R FILLER_63_112 ();
 FILLER_ASAP7_75t_R FILLER_63_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_124 ();
 DECAPx6_ASAP7_75t_R FILLER_63_135 ();
 DECAPx1_ASAP7_75t_R FILLER_63_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_160 ();
 DECAPx6_ASAP7_75t_R FILLER_63_167 ();
 DECAPx1_ASAP7_75t_R FILLER_63_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_212 ();
 FILLER_ASAP7_75t_R FILLER_63_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_221 ();
 DECAPx2_ASAP7_75t_R FILLER_63_225 ();
 FILLER_ASAP7_75t_R FILLER_63_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_241 ();
 DECAPx1_ASAP7_75t_R FILLER_63_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_308 ();
 DECAPx6_ASAP7_75t_R FILLER_63_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_378 ();
 FILLER_ASAP7_75t_R FILLER_63_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_387 ();
 DECAPx1_ASAP7_75t_R FILLER_63_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_395 ();
 DECAPx6_ASAP7_75t_R FILLER_63_406 ();
 FILLER_ASAP7_75t_R FILLER_63_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_429 ();
 FILLER_ASAP7_75t_R FILLER_63_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_444 ();
 DECAPx1_ASAP7_75t_R FILLER_63_477 ();
 DECAPx2_ASAP7_75t_R FILLER_63_491 ();
 FILLER_ASAP7_75t_R FILLER_63_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_499 ();
 DECAPx2_ASAP7_75t_R FILLER_63_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_532 ();
 DECAPx1_ASAP7_75t_R FILLER_63_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_551 ();
 DECAPx10_ASAP7_75t_R FILLER_63_555 ();
 FILLER_ASAP7_75t_R FILLER_63_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_579 ();
 DECAPx4_ASAP7_75t_R FILLER_63_594 ();
 FILLER_ASAP7_75t_R FILLER_63_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_606 ();
 DECAPx4_ASAP7_75t_R FILLER_63_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_637 ();
 DECAPx1_ASAP7_75t_R FILLER_63_641 ();
 DECAPx6_ASAP7_75t_R FILLER_63_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_700 ();
 DECAPx4_ASAP7_75t_R FILLER_63_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_747 ();
 DECAPx2_ASAP7_75t_R FILLER_63_756 ();
 FILLER_ASAP7_75t_R FILLER_63_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_764 ();
 FILLER_ASAP7_75t_R FILLER_63_780 ();
 DECAPx10_ASAP7_75t_R FILLER_63_791 ();
 DECAPx2_ASAP7_75t_R FILLER_63_813 ();
 DECAPx2_ASAP7_75t_R FILLER_63_835 ();
 FILLER_ASAP7_75t_R FILLER_63_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_853 ();
 DECAPx2_ASAP7_75t_R FILLER_63_868 ();
 FILLER_ASAP7_75t_R FILLER_63_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_876 ();
 FILLER_ASAP7_75t_R FILLER_63_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_893 ();
 DECAPx2_ASAP7_75t_R FILLER_63_907 ();
 FILLER_ASAP7_75t_R FILLER_63_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_915 ();
 DECAPx1_ASAP7_75t_R FILLER_63_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_936 ();
 DECAPx6_ASAP7_75t_R FILLER_63_943 ();
 FILLER_ASAP7_75t_R FILLER_63_957 ();
 FILLER_ASAP7_75t_R FILLER_63_965 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1053 ();
 DECAPx4_ASAP7_75t_R FILLER_63_1075 ();
 FILLER_ASAP7_75t_R FILLER_63_1085 ();
 FILLER_ASAP7_75t_R FILLER_63_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1116 ();
 FILLER_ASAP7_75t_R FILLER_63_1123 ();
 DECAPx4_ASAP7_75t_R FILLER_63_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1158 ();
 FILLER_ASAP7_75t_R FILLER_63_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1173 ();
 FILLER_ASAP7_75t_R FILLER_63_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1182 ();
 FILLER_ASAP7_75t_R FILLER_63_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1348 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1370 ();
 DECAPx10_ASAP7_75t_R FILLER_64_2 ();
 DECAPx10_ASAP7_75t_R FILLER_64_24 ();
 DECAPx10_ASAP7_75t_R FILLER_64_46 ();
 DECAPx10_ASAP7_75t_R FILLER_64_68 ();
 DECAPx6_ASAP7_75t_R FILLER_64_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_115 ();
 DECAPx2_ASAP7_75t_R FILLER_64_119 ();
 DECAPx1_ASAP7_75t_R FILLER_64_139 ();
 FILLER_ASAP7_75t_R FILLER_64_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_158 ();
 DECAPx4_ASAP7_75t_R FILLER_64_185 ();
 FILLER_ASAP7_75t_R FILLER_64_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_206 ();
 DECAPx2_ASAP7_75t_R FILLER_64_233 ();
 DECAPx2_ASAP7_75t_R FILLER_64_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_258 ();
 DECAPx2_ASAP7_75t_R FILLER_64_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_271 ();
 FILLER_ASAP7_75t_R FILLER_64_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_326 ();
 DECAPx10_ASAP7_75t_R FILLER_64_330 ();
 FILLER_ASAP7_75t_R FILLER_64_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_354 ();
 FILLER_ASAP7_75t_R FILLER_64_370 ();
 DECAPx10_ASAP7_75t_R FILLER_64_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_446 ();
 DECAPx2_ASAP7_75t_R FILLER_64_453 ();
 FILLER_ASAP7_75t_R FILLER_64_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_461 ();
 FILLER_ASAP7_75t_R FILLER_64_496 ();
 DECAPx1_ASAP7_75t_R FILLER_64_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_534 ();
 FILLER_ASAP7_75t_R FILLER_64_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_557 ();
 DECAPx4_ASAP7_75t_R FILLER_64_595 ();
 FILLER_ASAP7_75t_R FILLER_64_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_627 ();
 DECAPx2_ASAP7_75t_R FILLER_64_631 ();
 DECAPx6_ASAP7_75t_R FILLER_64_651 ();
 DECAPx2_ASAP7_75t_R FILLER_64_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_679 ();
 DECAPx1_ASAP7_75t_R FILLER_64_690 ();
 DECAPx2_ASAP7_75t_R FILLER_64_700 ();
 FILLER_ASAP7_75t_R FILLER_64_706 ();
 DECAPx1_ASAP7_75t_R FILLER_64_711 ();
 DECAPx4_ASAP7_75t_R FILLER_64_718 ();
 DECAPx1_ASAP7_75t_R FILLER_64_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_750 ();
 DECAPx10_ASAP7_75t_R FILLER_64_757 ();
 DECAPx4_ASAP7_75t_R FILLER_64_779 ();
 DECAPx2_ASAP7_75t_R FILLER_64_795 ();
 FILLER_ASAP7_75t_R FILLER_64_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_817 ();
 DECAPx10_ASAP7_75t_R FILLER_64_824 ();
 DECAPx2_ASAP7_75t_R FILLER_64_852 ();
 FILLER_ASAP7_75t_R FILLER_64_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_860 ();
 DECAPx10_ASAP7_75t_R FILLER_64_865 ();
 DECAPx2_ASAP7_75t_R FILLER_64_887 ();
 DECAPx10_ASAP7_75t_R FILLER_64_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_938 ();
 FILLER_ASAP7_75t_R FILLER_64_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_953 ();
 DECAPx1_ASAP7_75t_R FILLER_64_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1096 ();
 DECAPx4_ASAP7_75t_R FILLER_64_1105 ();
 FILLER_ASAP7_75t_R FILLER_64_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1133 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1149 ();
 FILLER_ASAP7_75t_R FILLER_64_1169 ();
 FILLER_ASAP7_75t_R FILLER_64_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1205 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1218 ();
 FILLER_ASAP7_75t_R FILLER_64_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1227 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1234 ();
 DECAPx1_ASAP7_75t_R FILLER_64_1248 ();
 DECAPx4_ASAP7_75t_R FILLER_64_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1354 ();
 DECAPx4_ASAP7_75t_R FILLER_64_1376 ();
 DECAPx1_ASAP7_75t_R FILLER_64_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_65_2 ();
 DECAPx10_ASAP7_75t_R FILLER_65_24 ();
 DECAPx10_ASAP7_75t_R FILLER_65_46 ();
 DECAPx10_ASAP7_75t_R FILLER_65_68 ();
 DECAPx4_ASAP7_75t_R FILLER_65_90 ();
 FILLER_ASAP7_75t_R FILLER_65_100 ();
 DECAPx1_ASAP7_75t_R FILLER_65_179 ();
 DECAPx1_ASAP7_75t_R FILLER_65_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_191 ();
 DECAPx4_ASAP7_75t_R FILLER_65_198 ();
 FILLER_ASAP7_75t_R FILLER_65_208 ();
 DECAPx2_ASAP7_75t_R FILLER_65_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_223 ();
 DECAPx1_ASAP7_75t_R FILLER_65_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_235 ();
 DECAPx10_ASAP7_75t_R FILLER_65_239 ();
 DECAPx6_ASAP7_75t_R FILLER_65_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_275 ();
 DECAPx1_ASAP7_75t_R FILLER_65_308 ();
 FILLER_ASAP7_75t_R FILLER_65_319 ();
 DECAPx10_ASAP7_75t_R FILLER_65_347 ();
 DECAPx2_ASAP7_75t_R FILLER_65_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_375 ();
 DECAPx6_ASAP7_75t_R FILLER_65_382 ();
 DECAPx1_ASAP7_75t_R FILLER_65_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_407 ();
 DECAPx4_ASAP7_75t_R FILLER_65_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_447 ();
 DECAPx4_ASAP7_75t_R FILLER_65_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_484 ();
 FILLER_ASAP7_75t_R FILLER_65_488 ();
 FILLER_ASAP7_75t_R FILLER_65_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_518 ();
 DECAPx10_ASAP7_75t_R FILLER_65_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_553 ();
 DECAPx1_ASAP7_75t_R FILLER_65_577 ();
 DECAPx4_ASAP7_75t_R FILLER_65_584 ();
 FILLER_ASAP7_75t_R FILLER_65_594 ();
 DECAPx2_ASAP7_75t_R FILLER_65_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_625 ();
 DECAPx1_ASAP7_75t_R FILLER_65_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_648 ();
 DECAPx1_ASAP7_75t_R FILLER_65_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_662 ();
 DECAPx10_ASAP7_75t_R FILLER_65_670 ();
 DECAPx1_ASAP7_75t_R FILLER_65_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_696 ();
 FILLER_ASAP7_75t_R FILLER_65_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_705 ();
 DECAPx1_ASAP7_75t_R FILLER_65_712 ();
 DECAPx1_ASAP7_75t_R FILLER_65_723 ();
 DECAPx2_ASAP7_75t_R FILLER_65_741 ();
 DECAPx2_ASAP7_75t_R FILLER_65_759 ();
 FILLER_ASAP7_75t_R FILLER_65_765 ();
 FILLER_ASAP7_75t_R FILLER_65_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_775 ();
 FILLER_ASAP7_75t_R FILLER_65_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_784 ();
 DECAPx1_ASAP7_75t_R FILLER_65_801 ();
 DECAPx1_ASAP7_75t_R FILLER_65_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_816 ();
 DECAPx1_ASAP7_75t_R FILLER_65_827 ();
 DECAPx4_ASAP7_75t_R FILLER_65_841 ();
 DECAPx1_ASAP7_75t_R FILLER_65_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_868 ();
 FILLER_ASAP7_75t_R FILLER_65_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_877 ();
 FILLER_ASAP7_75t_R FILLER_65_901 ();
 FILLER_ASAP7_75t_R FILLER_65_915 ();
 DECAPx1_ASAP7_75t_R FILLER_65_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_940 ();
 FILLER_ASAP7_75t_R FILLER_65_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_963 ();
 DECAPx10_ASAP7_75t_R FILLER_65_976 ();
 DECAPx2_ASAP7_75t_R FILLER_65_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1073 ();
 FILLER_ASAP7_75t_R FILLER_65_1084 ();
 FILLER_ASAP7_75t_R FILLER_65_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1103 ();
 FILLER_ASAP7_75t_R FILLER_65_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1157 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1188 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1247 ();
 FILLER_ASAP7_75t_R FILLER_65_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1349 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_66_2 ();
 DECAPx10_ASAP7_75t_R FILLER_66_24 ();
 DECAPx10_ASAP7_75t_R FILLER_66_46 ();
 DECAPx10_ASAP7_75t_R FILLER_66_68 ();
 DECAPx4_ASAP7_75t_R FILLER_66_90 ();
 FILLER_ASAP7_75t_R FILLER_66_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_102 ();
 DECAPx10_ASAP7_75t_R FILLER_66_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_137 ();
 DECAPx6_ASAP7_75t_R FILLER_66_166 ();
 FILLER_ASAP7_75t_R FILLER_66_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_188 ();
 DECAPx2_ASAP7_75t_R FILLER_66_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_221 ();
 FILLER_ASAP7_75t_R FILLER_66_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_250 ();
 DECAPx1_ASAP7_75t_R FILLER_66_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_281 ();
 FILLER_ASAP7_75t_R FILLER_66_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_290 ();
 DECAPx10_ASAP7_75t_R FILLER_66_294 ();
 DECAPx2_ASAP7_75t_R FILLER_66_316 ();
 DECAPx2_ASAP7_75t_R FILLER_66_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_335 ();
 DECAPx4_ASAP7_75t_R FILLER_66_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_375 ();
 DECAPx10_ASAP7_75t_R FILLER_66_392 ();
 DECAPx6_ASAP7_75t_R FILLER_66_414 ();
 FILLER_ASAP7_75t_R FILLER_66_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_430 ();
 DECAPx1_ASAP7_75t_R FILLER_66_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_461 ();
 FILLER_ASAP7_75t_R FILLER_66_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_472 ();
 DECAPx2_ASAP7_75t_R FILLER_66_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_485 ();
 DECAPx1_ASAP7_75t_R FILLER_66_489 ();
 FILLER_ASAP7_75t_R FILLER_66_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_505 ();
 DECAPx4_ASAP7_75t_R FILLER_66_512 ();
 FILLER_ASAP7_75t_R FILLER_66_522 ();
 FILLER_ASAP7_75t_R FILLER_66_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_529 ();
 DECAPx2_ASAP7_75t_R FILLER_66_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_551 ();
 DECAPx4_ASAP7_75t_R FILLER_66_566 ();
 FILLER_ASAP7_75t_R FILLER_66_576 ();
 DECAPx2_ASAP7_75t_R FILLER_66_598 ();
 FILLER_ASAP7_75t_R FILLER_66_604 ();
 DECAPx2_ASAP7_75t_R FILLER_66_623 ();
 FILLER_ASAP7_75t_R FILLER_66_629 ();
 DECAPx4_ASAP7_75t_R FILLER_66_634 ();
 FILLER_ASAP7_75t_R FILLER_66_644 ();
 FILLER_ASAP7_75t_R FILLER_66_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_657 ();
 DECAPx6_ASAP7_75t_R FILLER_66_676 ();
 FILLER_ASAP7_75t_R FILLER_66_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_692 ();
 FILLER_ASAP7_75t_R FILLER_66_703 ();
 FILLER_ASAP7_75t_R FILLER_66_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_714 ();
 FILLER_ASAP7_75t_R FILLER_66_721 ();
 DECAPx2_ASAP7_75t_R FILLER_66_736 ();
 FILLER_ASAP7_75t_R FILLER_66_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_744 ();
 FILLER_ASAP7_75t_R FILLER_66_752 ();
 DECAPx1_ASAP7_75t_R FILLER_66_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_773 ();
 FILLER_ASAP7_75t_R FILLER_66_783 ();
 FILLER_ASAP7_75t_R FILLER_66_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_804 ();
 FILLER_ASAP7_75t_R FILLER_66_811 ();
 FILLER_ASAP7_75t_R FILLER_66_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_822 ();
 FILLER_ASAP7_75t_R FILLER_66_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_832 ();
 FILLER_ASAP7_75t_R FILLER_66_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_863 ();
 DECAPx1_ASAP7_75t_R FILLER_66_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_884 ();
 DECAPx6_ASAP7_75t_R FILLER_66_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_914 ();
 DECAPx6_ASAP7_75t_R FILLER_66_918 ();
 DECAPx2_ASAP7_75t_R FILLER_66_932 ();
 FILLER_ASAP7_75t_R FILLER_66_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_952 ();
 DECAPx2_ASAP7_75t_R FILLER_66_959 ();
 FILLER_ASAP7_75t_R FILLER_66_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_979 ();
 DECAPx1_ASAP7_75t_R FILLER_66_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_66_1066 ();
 FILLER_ASAP7_75t_R FILLER_66_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1094 ();
 FILLER_ASAP7_75t_R FILLER_66_1116 ();
 FILLER_ASAP7_75t_R FILLER_66_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1133 ();
 FILLER_ASAP7_75t_R FILLER_66_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1223 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1254 ();
 FILLER_ASAP7_75t_R FILLER_66_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1349 ();
 DECAPx6_ASAP7_75t_R FILLER_66_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_67_2 ();
 DECAPx10_ASAP7_75t_R FILLER_67_24 ();
 DECAPx10_ASAP7_75t_R FILLER_67_46 ();
 DECAPx10_ASAP7_75t_R FILLER_67_68 ();
 FILLER_ASAP7_75t_R FILLER_67_90 ();
 DECAPx4_ASAP7_75t_R FILLER_67_118 ();
 FILLER_ASAP7_75t_R FILLER_67_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_130 ();
 DECAPx1_ASAP7_75t_R FILLER_67_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_194 ();
 FILLER_ASAP7_75t_R FILLER_67_201 ();
 DECAPx2_ASAP7_75t_R FILLER_67_206 ();
 DECAPx4_ASAP7_75t_R FILLER_67_216 ();
 FILLER_ASAP7_75t_R FILLER_67_226 ();
 DECAPx6_ASAP7_75t_R FILLER_67_234 ();
 FILLER_ASAP7_75t_R FILLER_67_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_273 ();
 DECAPx2_ASAP7_75t_R FILLER_67_300 ();
 FILLER_ASAP7_75t_R FILLER_67_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_308 ();
 DECAPx1_ASAP7_75t_R FILLER_67_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_339 ();
 DECAPx1_ASAP7_75t_R FILLER_67_347 ();
 DECAPx2_ASAP7_75t_R FILLER_67_403 ();
 FILLER_ASAP7_75t_R FILLER_67_409 ();
 FILLER_ASAP7_75t_R FILLER_67_423 ();
 FILLER_ASAP7_75t_R FILLER_67_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_430 ();
 DECAPx6_ASAP7_75t_R FILLER_67_455 ();
 FILLER_ASAP7_75t_R FILLER_67_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_471 ();
 DECAPx2_ASAP7_75t_R FILLER_67_498 ();
 DECAPx1_ASAP7_75t_R FILLER_67_536 ();
 DECAPx4_ASAP7_75t_R FILLER_67_554 ();
 FILLER_ASAP7_75t_R FILLER_67_564 ();
 DECAPx1_ASAP7_75t_R FILLER_67_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_612 ();
 DECAPx1_ASAP7_75t_R FILLER_67_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_657 ();
 DECAPx1_ASAP7_75t_R FILLER_67_685 ();
 FILLER_ASAP7_75t_R FILLER_67_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_726 ();
 DECAPx4_ASAP7_75t_R FILLER_67_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_745 ();
 DECAPx4_ASAP7_75t_R FILLER_67_763 ();
 FILLER_ASAP7_75t_R FILLER_67_773 ();
 DECAPx1_ASAP7_75t_R FILLER_67_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_786 ();
 DECAPx1_ASAP7_75t_R FILLER_67_794 ();
 DECAPx2_ASAP7_75t_R FILLER_67_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_836 ();
 DECAPx4_ASAP7_75t_R FILLER_67_843 ();
 FILLER_ASAP7_75t_R FILLER_67_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_855 ();
 DECAPx1_ASAP7_75t_R FILLER_67_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_866 ();
 FILLER_ASAP7_75t_R FILLER_67_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_879 ();
 DECAPx2_ASAP7_75t_R FILLER_67_899 ();
 FILLER_ASAP7_75t_R FILLER_67_905 ();
 DECAPx2_ASAP7_75t_R FILLER_67_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_923 ();
 DECAPx1_ASAP7_75t_R FILLER_67_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_946 ();
 DECAPx1_ASAP7_75t_R FILLER_67_954 ();
 DECAPx4_ASAP7_75t_R FILLER_67_971 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1036 ();
 DECAPx4_ASAP7_75t_R FILLER_67_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1061 ();
 FILLER_ASAP7_75t_R FILLER_67_1083 ();
 FILLER_ASAP7_75t_R FILLER_67_1095 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1113 ();
 DECAPx4_ASAP7_75t_R FILLER_67_1134 ();
 FILLER_ASAP7_75t_R FILLER_67_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1160 ();
 DECAPx4_ASAP7_75t_R FILLER_67_1176 ();
 FILLER_ASAP7_75t_R FILLER_67_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1203 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1236 ();
 FILLER_ASAP7_75t_R FILLER_67_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1385 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_68_2 ();
 DECAPx10_ASAP7_75t_R FILLER_68_24 ();
 DECAPx10_ASAP7_75t_R FILLER_68_46 ();
 DECAPx4_ASAP7_75t_R FILLER_68_68 ();
 FILLER_ASAP7_75t_R FILLER_68_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_83 ();
 DECAPx1_ASAP7_75t_R FILLER_68_90 ();
 DECAPx2_ASAP7_75t_R FILLER_68_100 ();
 DECAPx2_ASAP7_75t_R FILLER_68_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_115 ();
 DECAPx1_ASAP7_75t_R FILLER_68_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_124 ();
 FILLER_ASAP7_75t_R FILLER_68_132 ();
 FILLER_ASAP7_75t_R FILLER_68_181 ();
 DECAPx6_ASAP7_75t_R FILLER_68_186 ();
 DECAPx2_ASAP7_75t_R FILLER_68_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_206 ();
 DECAPx1_ASAP7_75t_R FILLER_68_233 ();
 FILLER_ASAP7_75t_R FILLER_68_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_245 ();
 DECAPx2_ASAP7_75t_R FILLER_68_272 ();
 FILLER_ASAP7_75t_R FILLER_68_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_280 ();
 DECAPx6_ASAP7_75t_R FILLER_68_329 ();
 DECAPx1_ASAP7_75t_R FILLER_68_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_357 ();
 DECAPx2_ASAP7_75t_R FILLER_68_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_380 ();
 DECAPx1_ASAP7_75t_R FILLER_68_413 ();
 DECAPx2_ASAP7_75t_R FILLER_68_423 ();
 FILLER_ASAP7_75t_R FILLER_68_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_431 ();
 DECAPx2_ASAP7_75t_R FILLER_68_436 ();
 FILLER_ASAP7_75t_R FILLER_68_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_444 ();
 FILLER_ASAP7_75t_R FILLER_68_448 ();
 DECAPx2_ASAP7_75t_R FILLER_68_454 ();
 FILLER_ASAP7_75t_R FILLER_68_460 ();
 DECAPx1_ASAP7_75t_R FILLER_68_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_468 ();
 DECAPx1_ASAP7_75t_R FILLER_68_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_479 ();
 DECAPx1_ASAP7_75t_R FILLER_68_486 ();
 DECAPx4_ASAP7_75t_R FILLER_68_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_504 ();
 DECAPx4_ASAP7_75t_R FILLER_68_523 ();
 FILLER_ASAP7_75t_R FILLER_68_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_535 ();
 DECAPx6_ASAP7_75t_R FILLER_68_548 ();
 FILLER_ASAP7_75t_R FILLER_68_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_578 ();
 DECAPx10_ASAP7_75t_R FILLER_68_585 ();
 DECAPx1_ASAP7_75t_R FILLER_68_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_611 ();
 DECAPx2_ASAP7_75t_R FILLER_68_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_650 ();
 DECAPx6_ASAP7_75t_R FILLER_68_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_703 ();
 FILLER_ASAP7_75t_R FILLER_68_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_709 ();
 DECAPx4_ASAP7_75t_R FILLER_68_717 ();
 FILLER_ASAP7_75t_R FILLER_68_727 ();
 DECAPx2_ASAP7_75t_R FILLER_68_742 ();
 FILLER_ASAP7_75t_R FILLER_68_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_754 ();
 DECAPx10_ASAP7_75t_R FILLER_68_761 ();
 DECAPx2_ASAP7_75t_R FILLER_68_783 ();
 FILLER_ASAP7_75t_R FILLER_68_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_791 ();
 DECAPx6_ASAP7_75t_R FILLER_68_814 ();
 FILLER_ASAP7_75t_R FILLER_68_828 ();
 DECAPx10_ASAP7_75t_R FILLER_68_836 ();
 FILLER_ASAP7_75t_R FILLER_68_858 ();
 DECAPx2_ASAP7_75t_R FILLER_68_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_878 ();
 DECAPx2_ASAP7_75t_R FILLER_68_889 ();
 DECAPx2_ASAP7_75t_R FILLER_68_902 ();
 DECAPx2_ASAP7_75t_R FILLER_68_916 ();
 DECAPx2_ASAP7_75t_R FILLER_68_929 ();
 DECAPx1_ASAP7_75t_R FILLER_68_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_959 ();
 DECAPx1_ASAP7_75t_R FILLER_68_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_971 ();
 DECAPx1_ASAP7_75t_R FILLER_68_979 ();
 DECAPx2_ASAP7_75t_R FILLER_68_989 ();
 DECAPx6_ASAP7_75t_R FILLER_68_998 ();
 FILLER_ASAP7_75t_R FILLER_68_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_68_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_68_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1109 ();
 FILLER_ASAP7_75t_R FILLER_68_1115 ();
 DECAPx6_ASAP7_75t_R FILLER_68_1129 ();
 FILLER_ASAP7_75t_R FILLER_68_1157 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1167 ();
 FILLER_ASAP7_75t_R FILLER_68_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1175 ();
 FILLER_ASAP7_75t_R FILLER_68_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1234 ();
 FILLER_ASAP7_75t_R FILLER_68_1253 ();
 FILLER_ASAP7_75t_R FILLER_68_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_68_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_68_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_69_2 ();
 DECAPx10_ASAP7_75t_R FILLER_69_24 ();
 DECAPx6_ASAP7_75t_R FILLER_69_46 ();
 DECAPx1_ASAP7_75t_R FILLER_69_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_64 ();
 FILLER_ASAP7_75t_R FILLER_69_95 ();
 DECAPx1_ASAP7_75t_R FILLER_69_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_107 ();
 DECAPx2_ASAP7_75t_R FILLER_69_144 ();
 DECAPx2_ASAP7_75t_R FILLER_69_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_163 ();
 DECAPx6_ASAP7_75t_R FILLER_69_167 ();
 DECAPx1_ASAP7_75t_R FILLER_69_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_185 ();
 DECAPx4_ASAP7_75t_R FILLER_69_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_223 ();
 DECAPx2_ASAP7_75t_R FILLER_69_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_256 ();
 DECAPx4_ASAP7_75t_R FILLER_69_266 ();
 FILLER_ASAP7_75t_R FILLER_69_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_278 ();
 FILLER_ASAP7_75t_R FILLER_69_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_291 ();
 DECAPx1_ASAP7_75t_R FILLER_69_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_312 ();
 DECAPx6_ASAP7_75t_R FILLER_69_319 ();
 DECAPx1_ASAP7_75t_R FILLER_69_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_337 ();
 DECAPx10_ASAP7_75t_R FILLER_69_364 ();
 FILLER_ASAP7_75t_R FILLER_69_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_400 ();
 FILLER_ASAP7_75t_R FILLER_69_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_406 ();
 DECAPx2_ASAP7_75t_R FILLER_69_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_471 ();
 DECAPx1_ASAP7_75t_R FILLER_69_478 ();
 DECAPx6_ASAP7_75t_R FILLER_69_485 ();
 FILLER_ASAP7_75t_R FILLER_69_499 ();
 DECAPx6_ASAP7_75t_R FILLER_69_519 ();
 DECAPx10_ASAP7_75t_R FILLER_69_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_561 ();
 DECAPx6_ASAP7_75t_R FILLER_69_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_596 ();
 DECAPx4_ASAP7_75t_R FILLER_69_600 ();
 FILLER_ASAP7_75t_R FILLER_69_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_618 ();
 DECAPx6_ASAP7_75t_R FILLER_69_625 ();
 FILLER_ASAP7_75t_R FILLER_69_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_641 ();
 DECAPx2_ASAP7_75t_R FILLER_69_656 ();
 FILLER_ASAP7_75t_R FILLER_69_662 ();
 DECAPx2_ASAP7_75t_R FILLER_69_671 ();
 DECAPx10_ASAP7_75t_R FILLER_69_689 ();
 DECAPx2_ASAP7_75t_R FILLER_69_711 ();
 FILLER_ASAP7_75t_R FILLER_69_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_727 ();
 FILLER_ASAP7_75t_R FILLER_69_735 ();
 DECAPx6_ASAP7_75t_R FILLER_69_743 ();
 DECAPx2_ASAP7_75t_R FILLER_69_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_763 ();
 DECAPx1_ASAP7_75t_R FILLER_69_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_786 ();
 DECAPx1_ASAP7_75t_R FILLER_69_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_804 ();
 DECAPx2_ASAP7_75t_R FILLER_69_819 ();
 FILLER_ASAP7_75t_R FILLER_69_835 ();
 DECAPx1_ASAP7_75t_R FILLER_69_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_849 ();
 DECAPx6_ASAP7_75t_R FILLER_69_856 ();
 DECAPx1_ASAP7_75t_R FILLER_69_870 ();
 DECAPx6_ASAP7_75t_R FILLER_69_880 ();
 FILLER_ASAP7_75t_R FILLER_69_894 ();
 DECAPx1_ASAP7_75t_R FILLER_69_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_907 ();
 DECAPx4_ASAP7_75t_R FILLER_69_914 ();
 DECAPx2_ASAP7_75t_R FILLER_69_933 ();
 DECAPx1_ASAP7_75t_R FILLER_69_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_956 ();
 DECAPx2_ASAP7_75t_R FILLER_69_963 ();
 FILLER_ASAP7_75t_R FILLER_69_969 ();
 FILLER_ASAP7_75t_R FILLER_69_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_989 ();
 DECAPx1_ASAP7_75t_R FILLER_69_997 ();
 DECAPx1_ASAP7_75t_R FILLER_69_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1047 ();
 FILLER_ASAP7_75t_R FILLER_69_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_69_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1089 ();
 DECAPx6_ASAP7_75t_R FILLER_69_1113 ();
 FILLER_ASAP7_75t_R FILLER_69_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1129 ();
 FILLER_ASAP7_75t_R FILLER_69_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1152 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1174 ();
 FILLER_ASAP7_75t_R FILLER_69_1184 ();
 DECAPx1_ASAP7_75t_R FILLER_69_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1350 ();
 DECAPx6_ASAP7_75t_R FILLER_69_1372 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1386 ();
 DECAPx10_ASAP7_75t_R FILLER_70_2 ();
 DECAPx10_ASAP7_75t_R FILLER_70_24 ();
 DECAPx10_ASAP7_75t_R FILLER_70_46 ();
 DECAPx4_ASAP7_75t_R FILLER_70_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_78 ();
 FILLER_ASAP7_75t_R FILLER_70_85 ();
 DECAPx4_ASAP7_75t_R FILLER_70_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_127 ();
 DECAPx1_ASAP7_75t_R FILLER_70_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_138 ();
 DECAPx2_ASAP7_75t_R FILLER_70_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_178 ();
 DECAPx6_ASAP7_75t_R FILLER_70_205 ();
 FILLER_ASAP7_75t_R FILLER_70_219 ();
 DECAPx2_ASAP7_75t_R FILLER_70_224 ();
 FILLER_ASAP7_75t_R FILLER_70_237 ();
 DECAPx2_ASAP7_75t_R FILLER_70_242 ();
 DECAPx10_ASAP7_75t_R FILLER_70_255 ();
 DECAPx10_ASAP7_75t_R FILLER_70_277 ();
 DECAPx6_ASAP7_75t_R FILLER_70_299 ();
 DECAPx1_ASAP7_75t_R FILLER_70_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_333 ();
 FILLER_ASAP7_75t_R FILLER_70_354 ();
 DECAPx2_ASAP7_75t_R FILLER_70_362 ();
 FILLER_ASAP7_75t_R FILLER_70_368 ();
 DECAPx2_ASAP7_75t_R FILLER_70_377 ();
 FILLER_ASAP7_75t_R FILLER_70_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_385 ();
 FILLER_ASAP7_75t_R FILLER_70_389 ();
 DECAPx6_ASAP7_75t_R FILLER_70_394 ();
 FILLER_ASAP7_75t_R FILLER_70_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_410 ();
 DECAPx1_ASAP7_75t_R FILLER_70_417 ();
 DECAPx1_ASAP7_75t_R FILLER_70_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_461 ();
 DECAPx1_ASAP7_75t_R FILLER_70_464 ();
 DECAPx6_ASAP7_75t_R FILLER_70_494 ();
 DECAPx4_ASAP7_75t_R FILLER_70_560 ();
 FILLER_ASAP7_75t_R FILLER_70_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_582 ();
 DECAPx2_ASAP7_75t_R FILLER_70_586 ();
 FILLER_ASAP7_75t_R FILLER_70_592 ();
 DECAPx6_ASAP7_75t_R FILLER_70_611 ();
 DECAPx2_ASAP7_75t_R FILLER_70_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_631 ();
 DECAPx6_ASAP7_75t_R FILLER_70_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_681 ();
 DECAPx1_ASAP7_75t_R FILLER_70_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_692 ();
 FILLER_ASAP7_75t_R FILLER_70_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_767 ();
 DECAPx1_ASAP7_75t_R FILLER_70_781 ();
 FILLER_ASAP7_75t_R FILLER_70_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_804 ();
 DECAPx6_ASAP7_75t_R FILLER_70_815 ();
 FILLER_ASAP7_75t_R FILLER_70_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_838 ();
 DECAPx4_ASAP7_75t_R FILLER_70_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_871 ();
 DECAPx2_ASAP7_75t_R FILLER_70_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_888 ();
 DECAPx2_ASAP7_75t_R FILLER_70_913 ();
 DECAPx4_ASAP7_75t_R FILLER_70_933 ();
 FILLER_ASAP7_75t_R FILLER_70_943 ();
 FILLER_ASAP7_75t_R FILLER_70_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_964 ();
 FILLER_ASAP7_75t_R FILLER_70_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_987 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1014 ();
 FILLER_ASAP7_75t_R FILLER_70_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1025 ();
 FILLER_ASAP7_75t_R FILLER_70_1031 ();
 DECAPx4_ASAP7_75t_R FILLER_70_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1052 ();
 FILLER_ASAP7_75t_R FILLER_70_1071 ();
 FILLER_ASAP7_75t_R FILLER_70_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1089 ();
 FILLER_ASAP7_75t_R FILLER_70_1095 ();
 FILLER_ASAP7_75t_R FILLER_70_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_70_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1123 ();
 FILLER_ASAP7_75t_R FILLER_70_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1132 ();
 DECAPx4_ASAP7_75t_R FILLER_70_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1160 ();
 FILLER_ASAP7_75t_R FILLER_70_1166 ();
 FILLER_ASAP7_75t_R FILLER_70_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1192 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1220 ();
 FILLER_ASAP7_75t_R FILLER_70_1226 ();
 DECAPx4_ASAP7_75t_R FILLER_70_1231 ();
 FILLER_ASAP7_75t_R FILLER_70_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1351 ();
 DECAPx4_ASAP7_75t_R FILLER_70_1373 ();
 FILLER_ASAP7_75t_R FILLER_70_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_71_2 ();
 DECAPx6_ASAP7_75t_R FILLER_71_24 ();
 FILLER_ASAP7_75t_R FILLER_71_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_40 ();
 DECAPx6_ASAP7_75t_R FILLER_71_67 ();
 DECAPx2_ASAP7_75t_R FILLER_71_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_87 ();
 FILLER_ASAP7_75t_R FILLER_71_100 ();
 DECAPx6_ASAP7_75t_R FILLER_71_105 ();
 DECAPx1_ASAP7_75t_R FILLER_71_119 ();
 DECAPx1_ASAP7_75t_R FILLER_71_129 ();
 DECAPx10_ASAP7_75t_R FILLER_71_136 ();
 FILLER_ASAP7_75t_R FILLER_71_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_160 ();
 FILLER_ASAP7_75t_R FILLER_71_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_178 ();
 DECAPx2_ASAP7_75t_R FILLER_71_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_220 ();
 DECAPx1_ASAP7_75t_R FILLER_71_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_231 ();
 FILLER_ASAP7_75t_R FILLER_71_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_243 ();
 DECAPx1_ASAP7_75t_R FILLER_71_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_274 ();
 DECAPx1_ASAP7_75t_R FILLER_71_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_292 ();
 DECAPx2_ASAP7_75t_R FILLER_71_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_302 ();
 DECAPx2_ASAP7_75t_R FILLER_71_335 ();
 DECAPx1_ASAP7_75t_R FILLER_71_367 ();
 DECAPx10_ASAP7_75t_R FILLER_71_397 ();
 DECAPx6_ASAP7_75t_R FILLER_71_419 ();
 FILLER_ASAP7_75t_R FILLER_71_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_435 ();
 DECAPx1_ASAP7_75t_R FILLER_71_455 ();
 DECAPx2_ASAP7_75t_R FILLER_71_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_468 ();
 DECAPx2_ASAP7_75t_R FILLER_71_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_481 ();
 FILLER_ASAP7_75t_R FILLER_71_485 ();
 DECAPx6_ASAP7_75t_R FILLER_71_491 ();
 FILLER_ASAP7_75t_R FILLER_71_505 ();
 DECAPx1_ASAP7_75t_R FILLER_71_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_523 ();
 FILLER_ASAP7_75t_R FILLER_71_527 ();
 DECAPx2_ASAP7_75t_R FILLER_71_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_551 ();
 DECAPx4_ASAP7_75t_R FILLER_71_560 ();
 FILLER_ASAP7_75t_R FILLER_71_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_603 ();
 FILLER_ASAP7_75t_R FILLER_71_618 ();
 DECAPx4_ASAP7_75t_R FILLER_71_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_639 ();
 DECAPx10_ASAP7_75t_R FILLER_71_653 ();
 DECAPx6_ASAP7_75t_R FILLER_71_675 ();
 DECAPx1_ASAP7_75t_R FILLER_71_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_707 ();
 DECAPx4_ASAP7_75t_R FILLER_71_711 ();
 DECAPx4_ASAP7_75t_R FILLER_71_734 ();
 DECAPx4_ASAP7_75t_R FILLER_71_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_768 ();
 DECAPx2_ASAP7_75t_R FILLER_71_782 ();
 FILLER_ASAP7_75t_R FILLER_71_788 ();
 DECAPx2_ASAP7_75t_R FILLER_71_797 ();
 DECAPx4_ASAP7_75t_R FILLER_71_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_819 ();
 FILLER_ASAP7_75t_R FILLER_71_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_846 ();
 FILLER_ASAP7_75t_R FILLER_71_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_855 ();
 FILLER_ASAP7_75t_R FILLER_71_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_874 ();
 FILLER_ASAP7_75t_R FILLER_71_879 ();
 DECAPx2_ASAP7_75t_R FILLER_71_887 ();
 FILLER_ASAP7_75t_R FILLER_71_893 ();
 FILLER_ASAP7_75t_R FILLER_71_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_923 ();
 DECAPx1_ASAP7_75t_R FILLER_71_926 ();
 DECAPx4_ASAP7_75t_R FILLER_71_933 ();
 FILLER_ASAP7_75t_R FILLER_71_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_945 ();
 DECAPx2_ASAP7_75t_R FILLER_71_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_965 ();
 FILLER_ASAP7_75t_R FILLER_71_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_980 ();
 DECAPx6_ASAP7_75t_R FILLER_71_988 ();
 FILLER_ASAP7_75t_R FILLER_71_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1015 ();
 FILLER_ASAP7_75t_R FILLER_71_1025 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_71_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_71_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1108 ();
 FILLER_ASAP7_75t_R FILLER_71_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1121 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1166 ();
 FILLER_ASAP7_75t_R FILLER_71_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1187 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1213 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1223 ();
 FILLER_ASAP7_75t_R FILLER_71_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1343 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1365 ();
 DECAPx1_ASAP7_75t_R FILLER_71_1387 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_72_2 ();
 DECAPx10_ASAP7_75t_R FILLER_72_24 ();
 DECAPx6_ASAP7_75t_R FILLER_72_46 ();
 FILLER_ASAP7_75t_R FILLER_72_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_88 ();
 DECAPx6_ASAP7_75t_R FILLER_72_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_117 ();
 DECAPx6_ASAP7_75t_R FILLER_72_144 ();
 FILLER_ASAP7_75t_R FILLER_72_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_186 ();
 DECAPx2_ASAP7_75t_R FILLER_72_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_206 ();
 DECAPx1_ASAP7_75t_R FILLER_72_213 ();
 DECAPx2_ASAP7_75t_R FILLER_72_243 ();
 FILLER_ASAP7_75t_R FILLER_72_249 ();
 DECAPx4_ASAP7_75t_R FILLER_72_329 ();
 FILLER_ASAP7_75t_R FILLER_72_352 ();
 DECAPx2_ASAP7_75t_R FILLER_72_357 ();
 FILLER_ASAP7_75t_R FILLER_72_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_365 ();
 DECAPx1_ASAP7_75t_R FILLER_72_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_386 ();
 FILLER_ASAP7_75t_R FILLER_72_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_393 ();
 DECAPx1_ASAP7_75t_R FILLER_72_420 ();
 DECAPx10_ASAP7_75t_R FILLER_72_427 ();
 DECAPx4_ASAP7_75t_R FILLER_72_449 ();
 FILLER_ASAP7_75t_R FILLER_72_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_461 ();
 FILLER_ASAP7_75t_R FILLER_72_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_493 ();
 DECAPx4_ASAP7_75t_R FILLER_72_520 ();
 DECAPx2_ASAP7_75t_R FILLER_72_562 ();
 DECAPx2_ASAP7_75t_R FILLER_72_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_584 ();
 DECAPx1_ASAP7_75t_R FILLER_72_608 ();
 DECAPx4_ASAP7_75t_R FILLER_72_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_631 ();
 DECAPx1_ASAP7_75t_R FILLER_72_653 ();
 DECAPx1_ASAP7_75t_R FILLER_72_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_679 ();
 FILLER_ASAP7_75t_R FILLER_72_688 ();
 DECAPx10_ASAP7_75t_R FILLER_72_697 ();
 DECAPx1_ASAP7_75t_R FILLER_72_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_723 ();
 DECAPx6_ASAP7_75t_R FILLER_72_730 ();
 FILLER_ASAP7_75t_R FILLER_72_744 ();
 DECAPx6_ASAP7_75t_R FILLER_72_749 ();
 DECAPx1_ASAP7_75t_R FILLER_72_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_767 ();
 DECAPx2_ASAP7_75t_R FILLER_72_781 ();
 FILLER_ASAP7_75t_R FILLER_72_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_789 ();
 DECAPx4_ASAP7_75t_R FILLER_72_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_816 ();
 DECAPx6_ASAP7_75t_R FILLER_72_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_847 ();
 FILLER_ASAP7_75t_R FILLER_72_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_856 ();
 DECAPx2_ASAP7_75t_R FILLER_72_862 ();
 DECAPx1_ASAP7_75t_R FILLER_72_876 ();
 DECAPx1_ASAP7_75t_R FILLER_72_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_890 ();
 DECAPx2_ASAP7_75t_R FILLER_72_908 ();
 FILLER_ASAP7_75t_R FILLER_72_914 ();
 FILLER_ASAP7_75t_R FILLER_72_942 ();
 DECAPx6_ASAP7_75t_R FILLER_72_980 ();
 DECAPx1_ASAP7_75t_R FILLER_72_994 ();
 FILLER_ASAP7_75t_R FILLER_72_1011 ();
 FILLER_ASAP7_75t_R FILLER_72_1016 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1063 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1081 ();
 FILLER_ASAP7_75t_R FILLER_72_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_72_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1134 ();
 FILLER_ASAP7_75t_R FILLER_72_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1150 ();
 FILLER_ASAP7_75t_R FILLER_72_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1238 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_73_2 ();
 DECAPx4_ASAP7_75t_R FILLER_73_24 ();
 DECAPx4_ASAP7_75t_R FILLER_73_161 ();
 FILLER_ASAP7_75t_R FILLER_73_171 ();
 DECAPx1_ASAP7_75t_R FILLER_73_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_207 ();
 DECAPx4_ASAP7_75t_R FILLER_73_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_221 ();
 DECAPx10_ASAP7_75t_R FILLER_73_228 ();
 DECAPx1_ASAP7_75t_R FILLER_73_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_268 ();
 DECAPx4_ASAP7_75t_R FILLER_73_272 ();
 DECAPx6_ASAP7_75t_R FILLER_73_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_302 ();
 DECAPx2_ASAP7_75t_R FILLER_73_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_316 ();
 DECAPx4_ASAP7_75t_R FILLER_73_320 ();
 FILLER_ASAP7_75t_R FILLER_73_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_332 ();
 DECAPx1_ASAP7_75t_R FILLER_73_365 ();
 FILLER_ASAP7_75t_R FILLER_73_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_397 ();
 FILLER_ASAP7_75t_R FILLER_73_404 ();
 FILLER_ASAP7_75t_R FILLER_73_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_450 ();
 DECAPx6_ASAP7_75t_R FILLER_73_454 ();
 DECAPx6_ASAP7_75t_R FILLER_73_474 ();
 DECAPx2_ASAP7_75t_R FILLER_73_488 ();
 DECAPx2_ASAP7_75t_R FILLER_73_500 ();
 FILLER_ASAP7_75t_R FILLER_73_506 ();
 DECAPx2_ASAP7_75t_R FILLER_73_511 ();
 DECAPx6_ASAP7_75t_R FILLER_73_521 ();
 DECAPx1_ASAP7_75t_R FILLER_73_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_550 ();
 DECAPx10_ASAP7_75t_R FILLER_73_554 ();
 DECAPx10_ASAP7_75t_R FILLER_73_576 ();
 FILLER_ASAP7_75t_R FILLER_73_598 ();
 DECAPx2_ASAP7_75t_R FILLER_73_609 ();
 FILLER_ASAP7_75t_R FILLER_73_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_617 ();
 DECAPx4_ASAP7_75t_R FILLER_73_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_649 ();
 DECAPx4_ASAP7_75t_R FILLER_73_671 ();
 FILLER_ASAP7_75t_R FILLER_73_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_696 ();
 DECAPx2_ASAP7_75t_R FILLER_73_704 ();
 FILLER_ASAP7_75t_R FILLER_73_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_712 ();
 DECAPx2_ASAP7_75t_R FILLER_73_716 ();
 FILLER_ASAP7_75t_R FILLER_73_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_734 ();
 DECAPx1_ASAP7_75t_R FILLER_73_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_746 ();
 DECAPx4_ASAP7_75t_R FILLER_73_761 ();
 FILLER_ASAP7_75t_R FILLER_73_771 ();
 DECAPx1_ASAP7_75t_R FILLER_73_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_784 ();
 DECAPx6_ASAP7_75t_R FILLER_73_808 ();
 DECAPx6_ASAP7_75t_R FILLER_73_828 ();
 DECAPx2_ASAP7_75t_R FILLER_73_852 ();
 FILLER_ASAP7_75t_R FILLER_73_858 ();
 DECAPx1_ASAP7_75t_R FILLER_73_878 ();
 DECAPx4_ASAP7_75t_R FILLER_73_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_911 ();
 DECAPx6_ASAP7_75t_R FILLER_73_926 ();
 DECAPx1_ASAP7_75t_R FILLER_73_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_944 ();
 FILLER_ASAP7_75t_R FILLER_73_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_961 ();
 DECAPx6_ASAP7_75t_R FILLER_73_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_998 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1025 ();
 FILLER_ASAP7_75t_R FILLER_73_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1059 ();
 FILLER_ASAP7_75t_R FILLER_73_1065 ();
 FILLER_ASAP7_75t_R FILLER_73_1091 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1103 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_73_1139 ();
 FILLER_ASAP7_75t_R FILLER_73_1161 ();
 DECAPx6_ASAP7_75t_R FILLER_73_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1219 ();
 DECAPx6_ASAP7_75t_R FILLER_73_1241 ();
 FILLER_ASAP7_75t_R FILLER_73_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1257 ();
 FILLER_ASAP7_75t_R FILLER_73_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1345 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1367 ();
 FILLER_ASAP7_75t_R FILLER_73_1389 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_74_2 ();
 DECAPx6_ASAP7_75t_R FILLER_74_24 ();
 DECAPx1_ASAP7_75t_R FILLER_74_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_58 ();
 DECAPx1_ASAP7_75t_R FILLER_74_63 ();
 FILLER_ASAP7_75t_R FILLER_74_73 ();
 DECAPx6_ASAP7_75t_R FILLER_74_87 ();
 FILLER_ASAP7_75t_R FILLER_74_101 ();
 DECAPx10_ASAP7_75t_R FILLER_74_109 ();
 DECAPx1_ASAP7_75t_R FILLER_74_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_135 ();
 DECAPx6_ASAP7_75t_R FILLER_74_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_160 ();
 DECAPx6_ASAP7_75t_R FILLER_74_164 ();
 DECAPx1_ASAP7_75t_R FILLER_74_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_182 ();
 DECAPx2_ASAP7_75t_R FILLER_74_189 ();
 DECAPx1_ASAP7_75t_R FILLER_74_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_202 ();
 DECAPx2_ASAP7_75t_R FILLER_74_210 ();
 FILLER_ASAP7_75t_R FILLER_74_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_244 ();
 DECAPx1_ASAP7_75t_R FILLER_74_255 ();
 DECAPx4_ASAP7_75t_R FILLER_74_262 ();
 FILLER_ASAP7_75t_R FILLER_74_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_274 ();
 DECAPx10_ASAP7_75t_R FILLER_74_282 ();
 DECAPx1_ASAP7_75t_R FILLER_74_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_308 ();
 DECAPx1_ASAP7_75t_R FILLER_74_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_320 ();
 DECAPx2_ASAP7_75t_R FILLER_74_324 ();
 FILLER_ASAP7_75t_R FILLER_74_330 ();
 DECAPx1_ASAP7_75t_R FILLER_74_338 ();
 DECAPx10_ASAP7_75t_R FILLER_74_348 ();
 FILLER_ASAP7_75t_R FILLER_74_370 ();
 DECAPx6_ASAP7_75t_R FILLER_74_378 ();
 DECAPx1_ASAP7_75t_R FILLER_74_392 ();
 DECAPx2_ASAP7_75t_R FILLER_74_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_408 ();
 DECAPx6_ASAP7_75t_R FILLER_74_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_435 ();
 DECAPx1_ASAP7_75t_R FILLER_74_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_483 ();
 DECAPx2_ASAP7_75t_R FILLER_74_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_500 ();
 DECAPx2_ASAP7_75t_R FILLER_74_527 ();
 DECAPx6_ASAP7_75t_R FILLER_74_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_550 ();
 DECAPx4_ASAP7_75t_R FILLER_74_569 ();
 FILLER_ASAP7_75t_R FILLER_74_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_581 ();
 DECAPx10_ASAP7_75t_R FILLER_74_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_622 ();
 DECAPx4_ASAP7_75t_R FILLER_74_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_643 ();
 FILLER_ASAP7_75t_R FILLER_74_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_652 ();
 DECAPx2_ASAP7_75t_R FILLER_74_671 ();
 FILLER_ASAP7_75t_R FILLER_74_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_679 ();
 FILLER_ASAP7_75t_R FILLER_74_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_690 ();
 FILLER_ASAP7_75t_R FILLER_74_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_726 ();
 DECAPx2_ASAP7_75t_R FILLER_74_769 ();
 FILLER_ASAP7_75t_R FILLER_74_775 ();
 DECAPx4_ASAP7_75t_R FILLER_74_783 ();
 DECAPx2_ASAP7_75t_R FILLER_74_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_809 ();
 FILLER_ASAP7_75t_R FILLER_74_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_836 ();
 FILLER_ASAP7_75t_R FILLER_74_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_859 ();
 DECAPx1_ASAP7_75t_R FILLER_74_885 ();
 DECAPx2_ASAP7_75t_R FILLER_74_897 ();
 FILLER_ASAP7_75t_R FILLER_74_903 ();
 DECAPx2_ASAP7_75t_R FILLER_74_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_917 ();
 FILLER_ASAP7_75t_R FILLER_74_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_957 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1051 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1102 ();
 FILLER_ASAP7_75t_R FILLER_74_1112 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1156 ();
 FILLER_ASAP7_75t_R FILLER_74_1162 ();
 FILLER_ASAP7_75t_R FILLER_74_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1196 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1203 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1239 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1251 ();
 FILLER_ASAP7_75t_R FILLER_74_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1388 ();
 FILLER_ASAP7_75t_R FILLER_75_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_4 ();
 DECAPx4_ASAP7_75t_R FILLER_75_34 ();
 FILLER_ASAP7_75t_R FILLER_75_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_46 ();
 DECAPx6_ASAP7_75t_R FILLER_75_59 ();
 DECAPx1_ASAP7_75t_R FILLER_75_73 ();
 DECAPx1_ASAP7_75t_R FILLER_75_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_96 ();
 DECAPx2_ASAP7_75t_R FILLER_75_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_106 ();
 DECAPx6_ASAP7_75t_R FILLER_75_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_125 ();
 DECAPx4_ASAP7_75t_R FILLER_75_136 ();
 DECAPx4_ASAP7_75t_R FILLER_75_172 ();
 FILLER_ASAP7_75t_R FILLER_75_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_184 ();
 FILLER_ASAP7_75t_R FILLER_75_195 ();
 DECAPx2_ASAP7_75t_R FILLER_75_223 ();
 DECAPx2_ASAP7_75t_R FILLER_75_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_244 ();
 FILLER_ASAP7_75t_R FILLER_75_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_254 ();
 FILLER_ASAP7_75t_R FILLER_75_333 ();
 DECAPx1_ASAP7_75t_R FILLER_75_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_372 ();
 DECAPx2_ASAP7_75t_R FILLER_75_399 ();
 FILLER_ASAP7_75t_R FILLER_75_405 ();
 DECAPx2_ASAP7_75t_R FILLER_75_410 ();
 DECAPx4_ASAP7_75t_R FILLER_75_422 ();
 FILLER_ASAP7_75t_R FILLER_75_442 ();
 DECAPx2_ASAP7_75t_R FILLER_75_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_556 ();
 FILLER_ASAP7_75t_R FILLER_75_560 ();
 DECAPx10_ASAP7_75t_R FILLER_75_588 ();
 DECAPx6_ASAP7_75t_R FILLER_75_610 ();
 DECAPx10_ASAP7_75t_R FILLER_75_634 ();
 DECAPx2_ASAP7_75t_R FILLER_75_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_662 ();
 DECAPx1_ASAP7_75t_R FILLER_75_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_698 ();
 DECAPx2_ASAP7_75t_R FILLER_75_705 ();
 FILLER_ASAP7_75t_R FILLER_75_711 ();
 DECAPx1_ASAP7_75t_R FILLER_75_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_732 ();
 DECAPx1_ASAP7_75t_R FILLER_75_743 ();
 DECAPx1_ASAP7_75t_R FILLER_75_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_754 ();
 DECAPx2_ASAP7_75t_R FILLER_75_765 ();
 FILLER_ASAP7_75t_R FILLER_75_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_773 ();
 DECAPx2_ASAP7_75t_R FILLER_75_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_798 ();
 FILLER_ASAP7_75t_R FILLER_75_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_807 ();
 FILLER_ASAP7_75t_R FILLER_75_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_822 ();
 DECAPx2_ASAP7_75t_R FILLER_75_850 ();
 DECAPx2_ASAP7_75t_R FILLER_75_874 ();
 DECAPx4_ASAP7_75t_R FILLER_75_892 ();
 FILLER_ASAP7_75t_R FILLER_75_902 ();
 DECAPx2_ASAP7_75t_R FILLER_75_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_923 ();
 DECAPx2_ASAP7_75t_R FILLER_75_926 ();
 DECAPx4_ASAP7_75t_R FILLER_75_935 ();
 DECAPx6_ASAP7_75t_R FILLER_75_951 ();
 FILLER_ASAP7_75t_R FILLER_75_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_979 ();
 DECAPx10_ASAP7_75t_R FILLER_75_987 ();
 DECAPx4_ASAP7_75t_R FILLER_75_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_75_1045 ();
 FILLER_ASAP7_75t_R FILLER_75_1055 ();
 DECAPx4_ASAP7_75t_R FILLER_75_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1090 ();
 FILLER_ASAP7_75t_R FILLER_75_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1110 ();
 FILLER_ASAP7_75t_R FILLER_75_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1129 ();
 DECAPx4_ASAP7_75t_R FILLER_75_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1185 ();
 FILLER_ASAP7_75t_R FILLER_75_1191 ();
 FILLER_ASAP7_75t_R FILLER_75_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1231 ();
 FILLER_ASAP7_75t_R FILLER_75_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_75_1362 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_76_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_8 ();
 DECAPx10_ASAP7_75t_R FILLER_76_45 ();
 FILLER_ASAP7_75t_R FILLER_76_67 ();
 DECAPx1_ASAP7_75t_R FILLER_76_75 ();
 FILLER_ASAP7_75t_R FILLER_76_131 ();
 FILLER_ASAP7_75t_R FILLER_76_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_142 ();
 FILLER_ASAP7_75t_R FILLER_76_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_148 ();
 FILLER_ASAP7_75t_R FILLER_76_182 ();
 DECAPx2_ASAP7_75t_R FILLER_76_202 ();
 FILLER_ASAP7_75t_R FILLER_76_208 ();
 DECAPx10_ASAP7_75t_R FILLER_76_219 ();
 DECAPx1_ASAP7_75t_R FILLER_76_241 ();
 FILLER_ASAP7_75t_R FILLER_76_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_277 ();
 DECAPx1_ASAP7_75t_R FILLER_76_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_296 ();
 DECAPx1_ASAP7_75t_R FILLER_76_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_310 ();
 DECAPx1_ASAP7_75t_R FILLER_76_373 ();
 FILLER_ASAP7_75t_R FILLER_76_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_385 ();
 DECAPx2_ASAP7_75t_R FILLER_76_441 ();
 FILLER_ASAP7_75t_R FILLER_76_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_449 ();
 DECAPx2_ASAP7_75t_R FILLER_76_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_464 ();
 FILLER_ASAP7_75t_R FILLER_76_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_471 ();
 DECAPx10_ASAP7_75t_R FILLER_76_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_500 ();
 DECAPx2_ASAP7_75t_R FILLER_76_507 ();
 FILLER_ASAP7_75t_R FILLER_76_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_518 ();
 DECAPx2_ASAP7_75t_R FILLER_76_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_531 ();
 FILLER_ASAP7_75t_R FILLER_76_575 ();
 FILLER_ASAP7_75t_R FILLER_76_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_582 ();
 DECAPx2_ASAP7_75t_R FILLER_76_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_630 ();
 DECAPx1_ASAP7_75t_R FILLER_76_638 ();
 DECAPx10_ASAP7_75t_R FILLER_76_652 ();
 DECAPx2_ASAP7_75t_R FILLER_76_674 ();
 FILLER_ASAP7_75t_R FILLER_76_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_690 ();
 DECAPx4_ASAP7_75t_R FILLER_76_703 ();
 DECAPx1_ASAP7_75t_R FILLER_76_756 ();
 FILLER_ASAP7_75t_R FILLER_76_794 ();
 DECAPx2_ASAP7_75t_R FILLER_76_802 ();
 FILLER_ASAP7_75t_R FILLER_76_808 ();
 FILLER_ASAP7_75t_R FILLER_76_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_820 ();
 DECAPx4_ASAP7_75t_R FILLER_76_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_839 ();
 DECAPx6_ASAP7_75t_R FILLER_76_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_860 ();
 DECAPx10_ASAP7_75t_R FILLER_76_869 ();
 DECAPx2_ASAP7_75t_R FILLER_76_891 ();
 DECAPx6_ASAP7_75t_R FILLER_76_945 ();
 DECAPx2_ASAP7_75t_R FILLER_76_959 ();
 FILLER_ASAP7_75t_R FILLER_76_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_978 ();
 DECAPx1_ASAP7_75t_R FILLER_76_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_990 ();
 DECAPx1_ASAP7_75t_R FILLER_76_998 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1008 ();
 FILLER_ASAP7_75t_R FILLER_76_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1062 ();
 FILLER_ASAP7_75t_R FILLER_76_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1088 ();
 FILLER_ASAP7_75t_R FILLER_76_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_76_1120 ();
 FILLER_ASAP7_75t_R FILLER_76_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1145 ();
 FILLER_ASAP7_75t_R FILLER_76_1151 ();
 FILLER_ASAP7_75t_R FILLER_76_1163 ();
 DECAPx4_ASAP7_75t_R FILLER_76_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1190 ();
 FILLER_ASAP7_75t_R FILLER_76_1197 ();
 FILLER_ASAP7_75t_R FILLER_76_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_77_2 ();
 DECAPx1_ASAP7_75t_R FILLER_77_26 ();
 DECAPx1_ASAP7_75t_R FILLER_77_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_64 ();
 DECAPx6_ASAP7_75t_R FILLER_77_91 ();
 DECAPx1_ASAP7_75t_R FILLER_77_124 ();
 DECAPx1_ASAP7_75t_R FILLER_77_154 ();
 DECAPx10_ASAP7_75t_R FILLER_77_174 ();
 DECAPx6_ASAP7_75t_R FILLER_77_196 ();
 DECAPx1_ASAP7_75t_R FILLER_77_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_214 ();
 DECAPx1_ASAP7_75t_R FILLER_77_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_245 ();
 DECAPx2_ASAP7_75t_R FILLER_77_252 ();
 FILLER_ASAP7_75t_R FILLER_77_258 ();
 FILLER_ASAP7_75t_R FILLER_77_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_265 ();
 DECAPx4_ASAP7_75t_R FILLER_77_279 ();
 DECAPx6_ASAP7_75t_R FILLER_77_302 ();
 DECAPx2_ASAP7_75t_R FILLER_77_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_355 ();
 DECAPx6_ASAP7_75t_R FILLER_77_362 ();
 DECAPx2_ASAP7_75t_R FILLER_77_382 ();
 FILLER_ASAP7_75t_R FILLER_77_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_390 ();
 DECAPx4_ASAP7_75t_R FILLER_77_403 ();
 FILLER_ASAP7_75t_R FILLER_77_413 ();
 FILLER_ASAP7_75t_R FILLER_77_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_449 ();
 DECAPx6_ASAP7_75t_R FILLER_77_456 ();
 FILLER_ASAP7_75t_R FILLER_77_470 ();
 DECAPx10_ASAP7_75t_R FILLER_77_498 ();
 FILLER_ASAP7_75t_R FILLER_77_520 ();
 DECAPx2_ASAP7_75t_R FILLER_77_532 ();
 FILLER_ASAP7_75t_R FILLER_77_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_540 ();
 DECAPx6_ASAP7_75t_R FILLER_77_547 ();
 DECAPx2_ASAP7_75t_R FILLER_77_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_567 ();
 DECAPx2_ASAP7_75t_R FILLER_77_574 ();
 FILLER_ASAP7_75t_R FILLER_77_645 ();
 DECAPx1_ASAP7_75t_R FILLER_77_661 ();
 DECAPx1_ASAP7_75t_R FILLER_77_677 ();
 DECAPx4_ASAP7_75t_R FILLER_77_701 ();
 FILLER_ASAP7_75t_R FILLER_77_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_720 ();
 FILLER_ASAP7_75t_R FILLER_77_757 ();
 DECAPx6_ASAP7_75t_R FILLER_77_775 ();
 FILLER_ASAP7_75t_R FILLER_77_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_791 ();
 DECAPx4_ASAP7_75t_R FILLER_77_798 ();
 FILLER_ASAP7_75t_R FILLER_77_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_810 ();
 DECAPx2_ASAP7_75t_R FILLER_77_818 ();
 FILLER_ASAP7_75t_R FILLER_77_830 ();
 DECAPx2_ASAP7_75t_R FILLER_77_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_858 ();
 DECAPx2_ASAP7_75t_R FILLER_77_869 ();
 FILLER_ASAP7_75t_R FILLER_77_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_877 ();
 DECAPx2_ASAP7_75t_R FILLER_77_892 ();
 FILLER_ASAP7_75t_R FILLER_77_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_900 ();
 DECAPx2_ASAP7_75t_R FILLER_77_915 ();
 DECAPx6_ASAP7_75t_R FILLER_77_926 ();
 FILLER_ASAP7_75t_R FILLER_77_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_958 ();
 DECAPx6_ASAP7_75t_R FILLER_77_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_989 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1028 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1032 ();
 FILLER_ASAP7_75t_R FILLER_77_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1062 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1079 ();
 FILLER_ASAP7_75t_R FILLER_77_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1088 ();
 FILLER_ASAP7_75t_R FILLER_77_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1122 ();
 DECAPx4_ASAP7_75t_R FILLER_77_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1154 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1168 ();
 DECAPx4_ASAP7_75t_R FILLER_77_1180 ();
 FILLER_ASAP7_75t_R FILLER_77_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1192 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1215 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1233 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1238 ();
 DECAPx4_ASAP7_75t_R FILLER_77_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1338 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1360 ();
 DECAPx2_ASAP7_75t_R FILLER_78_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_8 ();
 DECAPx1_ASAP7_75t_R FILLER_78_15 ();
 DECAPx10_ASAP7_75t_R FILLER_78_22 ();
 DECAPx1_ASAP7_75t_R FILLER_78_70 ();
 DECAPx1_ASAP7_75t_R FILLER_78_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_87 ();
 DECAPx6_ASAP7_75t_R FILLER_78_92 ();
 DECAPx1_ASAP7_75t_R FILLER_78_106 ();
 DECAPx10_ASAP7_75t_R FILLER_78_116 ();
 DECAPx6_ASAP7_75t_R FILLER_78_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_158 ();
 DECAPx6_ASAP7_75t_R FILLER_78_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_206 ();
 DECAPx4_ASAP7_75t_R FILLER_78_213 ();
 DECAPx2_ASAP7_75t_R FILLER_78_311 ();
 FILLER_ASAP7_75t_R FILLER_78_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_319 ();
 DECAPx1_ASAP7_75t_R FILLER_78_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_340 ();
 DECAPx6_ASAP7_75t_R FILLER_78_348 ();
 DECAPx2_ASAP7_75t_R FILLER_78_362 ();
 DECAPx2_ASAP7_75t_R FILLER_78_394 ();
 FILLER_ASAP7_75t_R FILLER_78_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_402 ();
 DECAPx6_ASAP7_75t_R FILLER_78_406 ();
 DECAPx1_ASAP7_75t_R FILLER_78_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_424 ();
 FILLER_ASAP7_75t_R FILLER_78_431 ();
 DECAPx2_ASAP7_75t_R FILLER_78_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_486 ();
 DECAPx1_ASAP7_75t_R FILLER_78_490 ();
 DECAPx2_ASAP7_75t_R FILLER_78_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_507 ();
 FILLER_ASAP7_75t_R FILLER_78_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_513 ();
 DECAPx2_ASAP7_75t_R FILLER_78_520 ();
 FILLER_ASAP7_75t_R FILLER_78_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_528 ();
 DECAPx1_ASAP7_75t_R FILLER_78_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_577 ();
 DECAPx2_ASAP7_75t_R FILLER_78_581 ();
 FILLER_ASAP7_75t_R FILLER_78_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_589 ();
 DECAPx2_ASAP7_75t_R FILLER_78_597 ();
 DECAPx6_ASAP7_75t_R FILLER_78_609 ();
 FILLER_ASAP7_75t_R FILLER_78_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_635 ();
 DECAPx2_ASAP7_75t_R FILLER_78_643 ();
 DECAPx10_ASAP7_75t_R FILLER_78_667 ();
 FILLER_ASAP7_75t_R FILLER_78_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_691 ();
 DECAPx2_ASAP7_75t_R FILLER_78_718 ();
 FILLER_ASAP7_75t_R FILLER_78_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_726 ();
 FILLER_ASAP7_75t_R FILLER_78_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_753 ();
 DECAPx6_ASAP7_75t_R FILLER_78_765 ();
 FILLER_ASAP7_75t_R FILLER_78_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_781 ();
 DECAPx4_ASAP7_75t_R FILLER_78_799 ();
 DECAPx6_ASAP7_75t_R FILLER_78_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_829 ();
 DECAPx4_ASAP7_75t_R FILLER_78_850 ();
 FILLER_ASAP7_75t_R FILLER_78_860 ();
 DECAPx2_ASAP7_75t_R FILLER_78_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_874 ();
 DECAPx10_ASAP7_75t_R FILLER_78_881 ();
 DECAPx10_ASAP7_75t_R FILLER_78_909 ();
 DECAPx1_ASAP7_75t_R FILLER_78_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_935 ();
 DECAPx2_ASAP7_75t_R FILLER_78_968 ();
 FILLER_ASAP7_75t_R FILLER_78_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_982 ();
 DECAPx4_ASAP7_75t_R FILLER_78_990 ();
 FILLER_ASAP7_75t_R FILLER_78_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1002 ();
 FILLER_ASAP7_75t_R FILLER_78_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_78_1077 ();
 FILLER_ASAP7_75t_R FILLER_78_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1113 ();
 FILLER_ASAP7_75t_R FILLER_78_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_78_1136 ();
 FILLER_ASAP7_75t_R FILLER_78_1146 ();
 DECAPx4_ASAP7_75t_R FILLER_78_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_78_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1236 ();
 FILLER_ASAP7_75t_R FILLER_78_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1338 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1360 ();
 FILLER_ASAP7_75t_R FILLER_78_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_78_1388 ();
 FILLER_ASAP7_75t_R FILLER_79_2 ();
 DECAPx1_ASAP7_75t_R FILLER_79_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_52 ();
 FILLER_ASAP7_75t_R FILLER_79_56 ();
 FILLER_ASAP7_75t_R FILLER_79_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_67 ();
 DECAPx6_ASAP7_75t_R FILLER_79_72 ();
 DECAPx1_ASAP7_75t_R FILLER_79_86 ();
 DECAPx4_ASAP7_75t_R FILLER_79_116 ();
 FILLER_ASAP7_75t_R FILLER_79_126 ();
 DECAPx2_ASAP7_75t_R FILLER_79_138 ();
 FILLER_ASAP7_75t_R FILLER_79_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_149 ();
 DECAPx1_ASAP7_75t_R FILLER_79_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_161 ();
 DECAPx2_ASAP7_75t_R FILLER_79_165 ();
 FILLER_ASAP7_75t_R FILLER_79_196 ();
 FILLER_ASAP7_75t_R FILLER_79_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_226 ();
 DECAPx2_ASAP7_75t_R FILLER_79_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_239 ();
 DECAPx10_ASAP7_75t_R FILLER_79_256 ();
 DECAPx6_ASAP7_75t_R FILLER_79_281 ();
 DECAPx1_ASAP7_75t_R FILLER_79_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_299 ();
 FILLER_ASAP7_75t_R FILLER_79_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_313 ();
 DECAPx6_ASAP7_75t_R FILLER_79_320 ();
 DECAPx2_ASAP7_75t_R FILLER_79_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_340 ();
 FILLER_ASAP7_75t_R FILLER_79_367 ();
 DECAPx4_ASAP7_75t_R FILLER_79_375 ();
 FILLER_ASAP7_75t_R FILLER_79_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_387 ();
 DECAPx4_ASAP7_75t_R FILLER_79_414 ();
 FILLER_ASAP7_75t_R FILLER_79_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_435 ();
 DECAPx1_ASAP7_75t_R FILLER_79_451 ();
 DECAPx4_ASAP7_75t_R FILLER_79_481 ();
 FILLER_ASAP7_75t_R FILLER_79_491 ();
 DECAPx2_ASAP7_75t_R FILLER_79_522 ();
 FILLER_ASAP7_75t_R FILLER_79_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_530 ();
 DECAPx2_ASAP7_75t_R FILLER_79_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_563 ();
 FILLER_ASAP7_75t_R FILLER_79_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_592 ();
 DECAPx10_ASAP7_75t_R FILLER_79_600 ();
 DECAPx1_ASAP7_75t_R FILLER_79_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_626 ();
 DECAPx10_ASAP7_75t_R FILLER_79_634 ();
 DECAPx1_ASAP7_75t_R FILLER_79_656 ();
 FILLER_ASAP7_75t_R FILLER_79_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_688 ();
 DECAPx4_ASAP7_75t_R FILLER_79_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_705 ();
 DECAPx2_ASAP7_75t_R FILLER_79_709 ();
 DECAPx2_ASAP7_75t_R FILLER_79_725 ();
 DECAPx4_ASAP7_75t_R FILLER_79_744 ();
 FILLER_ASAP7_75t_R FILLER_79_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_756 ();
 DECAPx6_ASAP7_75t_R FILLER_79_767 ();
 DECAPx1_ASAP7_75t_R FILLER_79_781 ();
 DECAPx2_ASAP7_75t_R FILLER_79_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_798 ();
 DECAPx4_ASAP7_75t_R FILLER_79_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_840 ();
 FILLER_ASAP7_75t_R FILLER_79_847 ();
 DECAPx10_ASAP7_75t_R FILLER_79_855 ();
 DECAPx2_ASAP7_75t_R FILLER_79_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_883 ();
 DECAPx1_ASAP7_75t_R FILLER_79_890 ();
 DECAPx1_ASAP7_75t_R FILLER_79_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_905 ();
 DECAPx1_ASAP7_75t_R FILLER_79_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_917 ();
 DECAPx10_ASAP7_75t_R FILLER_79_939 ();
 DECAPx6_ASAP7_75t_R FILLER_79_961 ();
 FILLER_ASAP7_75t_R FILLER_79_975 ();
 DECAPx6_ASAP7_75t_R FILLER_79_991 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1018 ();
 FILLER_ASAP7_75t_R FILLER_79_1024 ();
 DECAPx6_ASAP7_75t_R FILLER_79_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1085 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1107 ();
 FILLER_ASAP7_75t_R FILLER_79_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1145 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1182 ();
 FILLER_ASAP7_75t_R FILLER_79_1188 ();
 DECAPx6_ASAP7_75t_R FILLER_79_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1223 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1336 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1358 ();
 DECAPx4_ASAP7_75t_R FILLER_80_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_12 ();
 DECAPx2_ASAP7_75t_R FILLER_80_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_28 ();
 DECAPx2_ASAP7_75t_R FILLER_80_33 ();
 FILLER_ASAP7_75t_R FILLER_80_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_41 ();
 DECAPx4_ASAP7_75t_R FILLER_80_48 ();
 FILLER_ASAP7_75t_R FILLER_80_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_72 ();
 DECAPx2_ASAP7_75t_R FILLER_80_76 ();
 FILLER_ASAP7_75t_R FILLER_80_86 ();
 DECAPx1_ASAP7_75t_R FILLER_80_100 ();
 DECAPx2_ASAP7_75t_R FILLER_80_107 ();
 FILLER_ASAP7_75t_R FILLER_80_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_119 ();
 FILLER_ASAP7_75t_R FILLER_80_146 ();
 DECAPx6_ASAP7_75t_R FILLER_80_174 ();
 FILLER_ASAP7_75t_R FILLER_80_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_190 ();
 DECAPx1_ASAP7_75t_R FILLER_80_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_211 ();
 DECAPx10_ASAP7_75t_R FILLER_80_215 ();
 DECAPx2_ASAP7_75t_R FILLER_80_263 ();
 DECAPx4_ASAP7_75t_R FILLER_80_275 ();
 DECAPx1_ASAP7_75t_R FILLER_80_292 ();
 DECAPx1_ASAP7_75t_R FILLER_80_299 ();
 DECAPx2_ASAP7_75t_R FILLER_80_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_343 ();
 DECAPx1_ASAP7_75t_R FILLER_80_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_354 ();
 FILLER_ASAP7_75t_R FILLER_80_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_360 ();
 DECAPx1_ASAP7_75t_R FILLER_80_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_382 ();
 FILLER_ASAP7_75t_R FILLER_80_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_429 ();
 DECAPx6_ASAP7_75t_R FILLER_80_433 ();
 DECAPx1_ASAP7_75t_R FILLER_80_447 ();
 FILLER_ASAP7_75t_R FILLER_80_460 ();
 DECAPx1_ASAP7_75t_R FILLER_80_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_468 ();
 FILLER_ASAP7_75t_R FILLER_80_472 ();
 DECAPx4_ASAP7_75t_R FILLER_80_477 ();
 DECAPx2_ASAP7_75t_R FILLER_80_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_503 ();
 FILLER_ASAP7_75t_R FILLER_80_530 ();
 FILLER_ASAP7_75t_R FILLER_80_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_560 ();
 DECAPx2_ASAP7_75t_R FILLER_80_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_594 ();
 DECAPx1_ASAP7_75t_R FILLER_80_621 ();
 DECAPx4_ASAP7_75t_R FILLER_80_638 ();
 DECAPx1_ASAP7_75t_R FILLER_80_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_657 ();
 FILLER_ASAP7_75t_R FILLER_80_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_670 ();
 DECAPx1_ASAP7_75t_R FILLER_80_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_686 ();
 DECAPx2_ASAP7_75t_R FILLER_80_695 ();
 DECAPx10_ASAP7_75t_R FILLER_80_704 ();
 DECAPx2_ASAP7_75t_R FILLER_80_726 ();
 FILLER_ASAP7_75t_R FILLER_80_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_734 ();
 DECAPx2_ASAP7_75t_R FILLER_80_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_777 ();
 DECAPx6_ASAP7_75t_R FILLER_80_788 ();
 DECAPx2_ASAP7_75t_R FILLER_80_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_808 ();
 DECAPx6_ASAP7_75t_R FILLER_80_823 ();
 DECAPx1_ASAP7_75t_R FILLER_80_837 ();
 DECAPx4_ASAP7_75t_R FILLER_80_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_885 ();
 FILLER_ASAP7_75t_R FILLER_80_932 ();
 DECAPx2_ASAP7_75t_R FILLER_80_942 ();
 FILLER_ASAP7_75t_R FILLER_80_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_983 ();
 DECAPx1_ASAP7_75t_R FILLER_80_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1012 ();
 FILLER_ASAP7_75t_R FILLER_80_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1097 ();
 FILLER_ASAP7_75t_R FILLER_80_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1150 ();
 FILLER_ASAP7_75t_R FILLER_80_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1163 ();
 DECAPx4_ASAP7_75t_R FILLER_80_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1190 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1214 ();
 DECAPx4_ASAP7_75t_R FILLER_80_1225 ();
 FILLER_ASAP7_75t_R FILLER_80_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1335 ();
 DECAPx4_ASAP7_75t_R FILLER_80_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1367 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_81_2 ();
 DECAPx1_ASAP7_75t_R FILLER_81_16 ();
 DECAPx4_ASAP7_75t_R FILLER_81_46 ();
 FILLER_ASAP7_75t_R FILLER_81_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_58 ();
 DECAPx1_ASAP7_75t_R FILLER_81_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_95 ();
 DECAPx2_ASAP7_75t_R FILLER_81_99 ();
 DECAPx2_ASAP7_75t_R FILLER_81_111 ();
 FILLER_ASAP7_75t_R FILLER_81_117 ();
 FILLER_ASAP7_75t_R FILLER_81_122 ();
 DECAPx6_ASAP7_75t_R FILLER_81_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_153 ();
 DECAPx1_ASAP7_75t_R FILLER_81_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_164 ();
 FILLER_ASAP7_75t_R FILLER_81_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_179 ();
 DECAPx1_ASAP7_75t_R FILLER_81_186 ();
 DECAPx6_ASAP7_75t_R FILLER_81_196 ();
 DECAPx2_ASAP7_75t_R FILLER_81_210 ();
 DECAPx6_ASAP7_75t_R FILLER_81_224 ();
 FILLER_ASAP7_75t_R FILLER_81_238 ();
 DECAPx1_ASAP7_75t_R FILLER_81_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_255 ();
 DECAPx4_ASAP7_75t_R FILLER_81_308 ();
 DECAPx4_ASAP7_75t_R FILLER_81_321 ();
 FILLER_ASAP7_75t_R FILLER_81_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_359 ();
 DECAPx1_ASAP7_75t_R FILLER_81_386 ();
 FILLER_ASAP7_75t_R FILLER_81_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_414 ();
 DECAPx6_ASAP7_75t_R FILLER_81_441 ();
 DECAPx6_ASAP7_75t_R FILLER_81_461 ();
 DECAPx2_ASAP7_75t_R FILLER_81_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_481 ();
 FILLER_ASAP7_75t_R FILLER_81_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_502 ();
 DECAPx1_ASAP7_75t_R FILLER_81_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_514 ();
 DECAPx4_ASAP7_75t_R FILLER_81_521 ();
 FILLER_ASAP7_75t_R FILLER_81_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_540 ();
 FILLER_ASAP7_75t_R FILLER_81_550 ();
 DECAPx1_ASAP7_75t_R FILLER_81_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_588 ();
 DECAPx2_ASAP7_75t_R FILLER_81_615 ();
 FILLER_ASAP7_75t_R FILLER_81_621 ();
 DECAPx6_ASAP7_75t_R FILLER_81_653 ();
 DECAPx2_ASAP7_75t_R FILLER_81_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_673 ();
 DECAPx2_ASAP7_75t_R FILLER_81_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_713 ();
 DECAPx4_ASAP7_75t_R FILLER_81_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_748 ();
 DECAPx2_ASAP7_75t_R FILLER_81_755 ();
 FILLER_ASAP7_75t_R FILLER_81_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_776 ();
 DECAPx6_ASAP7_75t_R FILLER_81_787 ();
 DECAPx2_ASAP7_75t_R FILLER_81_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_807 ();
 DECAPx1_ASAP7_75t_R FILLER_81_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_836 ();
 DECAPx4_ASAP7_75t_R FILLER_81_845 ();
 DECAPx1_ASAP7_75t_R FILLER_81_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_869 ();
 FILLER_ASAP7_75t_R FILLER_81_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_899 ();
 FILLER_ASAP7_75t_R FILLER_81_916 ();
 DECAPx2_ASAP7_75t_R FILLER_81_960 ();
 DECAPx1_ASAP7_75t_R FILLER_81_972 ();
 FILLER_ASAP7_75t_R FILLER_81_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_984 ();
 FILLER_ASAP7_75t_R FILLER_81_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1035 ();
 FILLER_ASAP7_75t_R FILLER_81_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1048 ();
 FILLER_ASAP7_75t_R FILLER_81_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1078 ();
 FILLER_ASAP7_75t_R FILLER_81_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1119 ();
 FILLER_ASAP7_75t_R FILLER_81_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1185 ();
 FILLER_ASAP7_75t_R FILLER_81_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1213 ();
 FILLER_ASAP7_75t_R FILLER_81_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1244 ();
 DECAPx4_ASAP7_75t_R FILLER_81_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1296 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1302 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1346 ();
 DECAPx4_ASAP7_75t_R FILLER_81_1358 ();
 FILLER_ASAP7_75t_R FILLER_82_34 ();
 DECAPx4_ASAP7_75t_R FILLER_82_66 ();
 FILLER_ASAP7_75t_R FILLER_82_76 ();
 DECAPx4_ASAP7_75t_R FILLER_82_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_140 ();
 FILLER_ASAP7_75t_R FILLER_82_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_150 ();
 DECAPx2_ASAP7_75t_R FILLER_82_154 ();
 FILLER_ASAP7_75t_R FILLER_82_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_179 ();
 FILLER_ASAP7_75t_R FILLER_82_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_212 ();
 DECAPx2_ASAP7_75t_R FILLER_82_233 ();
 FILLER_ASAP7_75t_R FILLER_82_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_241 ();
 DECAPx4_ASAP7_75t_R FILLER_82_248 ();
 FILLER_ASAP7_75t_R FILLER_82_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_260 ();
 DECAPx2_ASAP7_75t_R FILLER_82_268 ();
 DECAPx2_ASAP7_75t_R FILLER_82_277 ();
 FILLER_ASAP7_75t_R FILLER_82_283 ();
 DECAPx4_ASAP7_75t_R FILLER_82_291 ();
 FILLER_ASAP7_75t_R FILLER_82_301 ();
 DECAPx4_ASAP7_75t_R FILLER_82_329 ();
 FILLER_ASAP7_75t_R FILLER_82_339 ();
 DECAPx4_ASAP7_75t_R FILLER_82_350 ();
 FILLER_ASAP7_75t_R FILLER_82_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_362 ();
 DECAPx6_ASAP7_75t_R FILLER_82_369 ();
 FILLER_ASAP7_75t_R FILLER_82_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_385 ();
 DECAPx1_ASAP7_75t_R FILLER_82_392 ();
 DECAPx6_ASAP7_75t_R FILLER_82_399 ();
 FILLER_ASAP7_75t_R FILLER_82_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_415 ();
 FILLER_ASAP7_75t_R FILLER_82_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_425 ();
 DECAPx4_ASAP7_75t_R FILLER_82_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_442 ();
 DECAPx2_ASAP7_75t_R FILLER_82_450 ();
 FILLER_ASAP7_75t_R FILLER_82_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_461 ();
 DECAPx10_ASAP7_75t_R FILLER_82_464 ();
 DECAPx2_ASAP7_75t_R FILLER_82_486 ();
 DECAPx10_ASAP7_75t_R FILLER_82_518 ();
 DECAPx2_ASAP7_75t_R FILLER_82_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_546 ();
 DECAPx4_ASAP7_75t_R FILLER_82_550 ();
 FILLER_ASAP7_75t_R FILLER_82_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_562 ();
 FILLER_ASAP7_75t_R FILLER_82_570 ();
 DECAPx4_ASAP7_75t_R FILLER_82_575 ();
 FILLER_ASAP7_75t_R FILLER_82_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_587 ();
 DECAPx1_ASAP7_75t_R FILLER_82_600 ();
 FILLER_ASAP7_75t_R FILLER_82_607 ();
 DECAPx4_ASAP7_75t_R FILLER_82_612 ();
 FILLER_ASAP7_75t_R FILLER_82_622 ();
 DECAPx6_ASAP7_75t_R FILLER_82_638 ();
 FILLER_ASAP7_75t_R FILLER_82_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_654 ();
 DECAPx4_ASAP7_75t_R FILLER_82_670 ();
 DECAPx2_ASAP7_75t_R FILLER_82_697 ();
 DECAPx10_ASAP7_75t_R FILLER_82_715 ();
 DECAPx2_ASAP7_75t_R FILLER_82_737 ();
 FILLER_ASAP7_75t_R FILLER_82_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_745 ();
 DECAPx2_ASAP7_75t_R FILLER_82_766 ();
 FILLER_ASAP7_75t_R FILLER_82_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_794 ();
 FILLER_ASAP7_75t_R FILLER_82_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_813 ();
 DECAPx2_ASAP7_75t_R FILLER_82_827 ();
 FILLER_ASAP7_75t_R FILLER_82_833 ();
 DECAPx4_ASAP7_75t_R FILLER_82_848 ();
 FILLER_ASAP7_75t_R FILLER_82_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_881 ();
 DECAPx1_ASAP7_75t_R FILLER_82_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_893 ();
 DECAPx6_ASAP7_75t_R FILLER_82_897 ();
 DECAPx1_ASAP7_75t_R FILLER_82_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_915 ();
 FILLER_ASAP7_75t_R FILLER_82_934 ();
 FILLER_ASAP7_75t_R FILLER_82_944 ();
 DECAPx2_ASAP7_75t_R FILLER_82_981 ();
 FILLER_ASAP7_75t_R FILLER_82_987 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1019 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1081 ();
 FILLER_ASAP7_75t_R FILLER_82_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_82_1155 ();
 FILLER_ASAP7_75t_R FILLER_82_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1194 ();
 FILLER_ASAP7_75t_R FILLER_82_1208 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1263 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1277 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1281 ();
 FILLER_ASAP7_75t_R FILLER_82_1289 ();
 FILLER_ASAP7_75t_R FILLER_82_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1349 ();
 FILLER_ASAP7_75t_R FILLER_82_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1388 ();
 FILLER_ASAP7_75t_R FILLER_83_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_26 ();
 FILLER_ASAP7_75t_R FILLER_83_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_37 ();
 DECAPx1_ASAP7_75t_R FILLER_83_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_54 ();
 DECAPx2_ASAP7_75t_R FILLER_83_58 ();
 DECAPx6_ASAP7_75t_R FILLER_83_68 ();
 DECAPx2_ASAP7_75t_R FILLER_83_100 ();
 FILLER_ASAP7_75t_R FILLER_83_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_108 ();
 DECAPx6_ASAP7_75t_R FILLER_83_115 ();
 DECAPx2_ASAP7_75t_R FILLER_83_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_135 ();
 FILLER_ASAP7_75t_R FILLER_83_162 ();
 DECAPx2_ASAP7_75t_R FILLER_83_170 ();
 DECAPx1_ASAP7_75t_R FILLER_83_182 ();
 DECAPx2_ASAP7_75t_R FILLER_83_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_204 ();
 DECAPx2_ASAP7_75t_R FILLER_83_239 ();
 DECAPx1_ASAP7_75t_R FILLER_83_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_255 ();
 DECAPx1_ASAP7_75t_R FILLER_83_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_266 ();
 DECAPx10_ASAP7_75t_R FILLER_83_275 ();
 DECAPx2_ASAP7_75t_R FILLER_83_297 ();
 FILLER_ASAP7_75t_R FILLER_83_303 ();
 DECAPx4_ASAP7_75t_R FILLER_83_321 ();
 DECAPx6_ASAP7_75t_R FILLER_83_337 ();
 DECAPx2_ASAP7_75t_R FILLER_83_351 ();
 DECAPx6_ASAP7_75t_R FILLER_83_363 ();
 DECAPx1_ASAP7_75t_R FILLER_83_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_381 ();
 DECAPx1_ASAP7_75t_R FILLER_83_411 ();
 DECAPx2_ASAP7_75t_R FILLER_83_473 ();
 FILLER_ASAP7_75t_R FILLER_83_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_484 ();
 FILLER_ASAP7_75t_R FILLER_83_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_491 ();
 FILLER_ASAP7_75t_R FILLER_83_499 ();
 FILLER_ASAP7_75t_R FILLER_83_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_543 ();
 DECAPx6_ASAP7_75t_R FILLER_83_547 ();
 DECAPx1_ASAP7_75t_R FILLER_83_561 ();
 DECAPx10_ASAP7_75t_R FILLER_83_591 ();
 DECAPx2_ASAP7_75t_R FILLER_83_613 ();
 DECAPx1_ASAP7_75t_R FILLER_83_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_629 ();
 DECAPx2_ASAP7_75t_R FILLER_83_640 ();
 FILLER_ASAP7_75t_R FILLER_83_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_683 ();
 DECAPx1_ASAP7_75t_R FILLER_83_710 ();
 DECAPx6_ASAP7_75t_R FILLER_83_748 ();
 FILLER_ASAP7_75t_R FILLER_83_762 ();
 FILLER_ASAP7_75t_R FILLER_83_774 ();
 DECAPx2_ASAP7_75t_R FILLER_83_786 ();
 DECAPx6_ASAP7_75t_R FILLER_83_812 ();
 DECAPx1_ASAP7_75t_R FILLER_83_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_841 ();
 FILLER_ASAP7_75t_R FILLER_83_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_857 ();
 DECAPx2_ASAP7_75t_R FILLER_83_865 ();
 FILLER_ASAP7_75t_R FILLER_83_871 ();
 DECAPx1_ASAP7_75t_R FILLER_83_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_883 ();
 DECAPx2_ASAP7_75t_R FILLER_83_892 ();
 FILLER_ASAP7_75t_R FILLER_83_898 ();
 DECAPx2_ASAP7_75t_R FILLER_83_910 ();
 FILLER_ASAP7_75t_R FILLER_83_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_934 ();
 DECAPx6_ASAP7_75t_R FILLER_83_942 ();
 DECAPx2_ASAP7_75t_R FILLER_83_964 ();
 DECAPx4_ASAP7_75t_R FILLER_83_973 ();
 FILLER_ASAP7_75t_R FILLER_83_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_985 ();
 DECAPx2_ASAP7_75t_R FILLER_83_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1002 ();
 DECAPx4_ASAP7_75t_R FILLER_83_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_83_1023 ();
 FILLER_ASAP7_75t_R FILLER_83_1043 ();
 DECAPx4_ASAP7_75t_R FILLER_83_1061 ();
 FILLER_ASAP7_75t_R FILLER_83_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1073 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1080 ();
 FILLER_ASAP7_75t_R FILLER_83_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1144 ();
 FILLER_ASAP7_75t_R FILLER_83_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1180 ();
 FILLER_ASAP7_75t_R FILLER_83_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1206 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1239 ();
 FILLER_ASAP7_75t_R FILLER_83_1245 ();
 FILLER_ASAP7_75t_R FILLER_83_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1281 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1307 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1323 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1329 ();
 DECAPx1_ASAP7_75t_R FILLER_83_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1350 ();
 FILLER_ASAP7_75t_R FILLER_83_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1373 ();
 DECAPx4_ASAP7_75t_R FILLER_84_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_12 ();
 DECAPx10_ASAP7_75t_R FILLER_84_19 ();
 DECAPx10_ASAP7_75t_R FILLER_84_41 ();
 DECAPx6_ASAP7_75t_R FILLER_84_63 ();
 FILLER_ASAP7_75t_R FILLER_84_103 ();
 FILLER_ASAP7_75t_R FILLER_84_117 ();
 DECAPx2_ASAP7_75t_R FILLER_84_122 ();
 FILLER_ASAP7_75t_R FILLER_84_128 ();
 DECAPx2_ASAP7_75t_R FILLER_84_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_145 ();
 DECAPx4_ASAP7_75t_R FILLER_84_152 ();
 FILLER_ASAP7_75t_R FILLER_84_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_179 ();
 DECAPx2_ASAP7_75t_R FILLER_84_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_192 ();
 DECAPx1_ASAP7_75t_R FILLER_84_201 ();
 DECAPx1_ASAP7_75t_R FILLER_84_211 ();
 DECAPx2_ASAP7_75t_R FILLER_84_221 ();
 FILLER_ASAP7_75t_R FILLER_84_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_258 ();
 DECAPx4_ASAP7_75t_R FILLER_84_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_295 ();
 DECAPx10_ASAP7_75t_R FILLER_84_302 ();
 FILLER_ASAP7_75t_R FILLER_84_324 ();
 DECAPx1_ASAP7_75t_R FILLER_84_346 ();
 DECAPx4_ASAP7_75t_R FILLER_84_370 ();
 FILLER_ASAP7_75t_R FILLER_84_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_382 ();
 FILLER_ASAP7_75t_R FILLER_84_389 ();
 DECAPx6_ASAP7_75t_R FILLER_84_397 ();
 DECAPx2_ASAP7_75t_R FILLER_84_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_417 ();
 DECAPx2_ASAP7_75t_R FILLER_84_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_430 ();
 DECAPx1_ASAP7_75t_R FILLER_84_442 ();
 DECAPx1_ASAP7_75t_R FILLER_84_452 ();
 FILLER_ASAP7_75t_R FILLER_84_464 ();
 FILLER_ASAP7_75t_R FILLER_84_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_494 ();
 FILLER_ASAP7_75t_R FILLER_84_514 ();
 DECAPx1_ASAP7_75t_R FILLER_84_519 ();
 DECAPx2_ASAP7_75t_R FILLER_84_556 ();
 FILLER_ASAP7_75t_R FILLER_84_562 ();
 DECAPx2_ASAP7_75t_R FILLER_84_570 ();
 FILLER_ASAP7_75t_R FILLER_84_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_578 ();
 DECAPx10_ASAP7_75t_R FILLER_84_588 ();
 DECAPx1_ASAP7_75t_R FILLER_84_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_614 ();
 DECAPx6_ASAP7_75t_R FILLER_84_631 ();
 FILLER_ASAP7_75t_R FILLER_84_645 ();
 FILLER_ASAP7_75t_R FILLER_84_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_659 ();
 DECAPx2_ASAP7_75t_R FILLER_84_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_678 ();
 DECAPx2_ASAP7_75t_R FILLER_84_693 ();
 DECAPx1_ASAP7_75t_R FILLER_84_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_706 ();
 DECAPx10_ASAP7_75t_R FILLER_84_713 ();
 FILLER_ASAP7_75t_R FILLER_84_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_771 ();
 DECAPx2_ASAP7_75t_R FILLER_84_782 ();
 FILLER_ASAP7_75t_R FILLER_84_788 ();
 FILLER_ASAP7_75t_R FILLER_84_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_812 ();
 DECAPx1_ASAP7_75t_R FILLER_84_819 ();
 DECAPx1_ASAP7_75t_R FILLER_84_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_839 ();
 DECAPx2_ASAP7_75t_R FILLER_84_873 ();
 FILLER_ASAP7_75t_R FILLER_84_879 ();
 FILLER_ASAP7_75t_R FILLER_84_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_893 ();
 DECAPx6_ASAP7_75t_R FILLER_84_905 ();
 DECAPx1_ASAP7_75t_R FILLER_84_919 ();
 DECAPx10_ASAP7_75t_R FILLER_84_929 ();
 DECAPx2_ASAP7_75t_R FILLER_84_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_957 ();
 DECAPx6_ASAP7_75t_R FILLER_84_964 ();
 FILLER_ASAP7_75t_R FILLER_84_984 ();
 DECAPx10_ASAP7_75t_R FILLER_84_996 ();
 DECAPx6_ASAP7_75t_R FILLER_84_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1058 ();
 FILLER_ASAP7_75t_R FILLER_84_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1091 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1122 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1143 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1163 ();
 FILLER_ASAP7_75t_R FILLER_84_1173 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1182 ();
 DECAPx6_ASAP7_75t_R FILLER_84_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1227 ();
 DECAPx6_ASAP7_75t_R FILLER_84_1231 ();
 FILLER_ASAP7_75t_R FILLER_84_1245 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1254 ();
 FILLER_ASAP7_75t_R FILLER_84_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1262 ();
 DECAPx6_ASAP7_75t_R FILLER_84_1275 ();
 FILLER_ASAP7_75t_R FILLER_84_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1294 ();
 DECAPx6_ASAP7_75t_R FILLER_84_1301 ();
 FILLER_ASAP7_75t_R FILLER_84_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1328 ();
 FILLER_ASAP7_75t_R FILLER_84_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1336 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1367 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1388 ();
 FILLER_ASAP7_75t_R FILLER_85_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_4 ();
 DECAPx1_ASAP7_75t_R FILLER_85_35 ();
 DECAPx2_ASAP7_75t_R FILLER_85_45 ();
 FILLER_ASAP7_75t_R FILLER_85_51 ();
 DECAPx2_ASAP7_75t_R FILLER_85_83 ();
 FILLER_ASAP7_75t_R FILLER_85_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_91 ();
 DECAPx2_ASAP7_75t_R FILLER_85_95 ();
 DECAPx4_ASAP7_75t_R FILLER_85_153 ();
 FILLER_ASAP7_75t_R FILLER_85_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_165 ();
 DECAPx10_ASAP7_75t_R FILLER_85_174 ();
 DECAPx4_ASAP7_75t_R FILLER_85_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_220 ();
 DECAPx1_ASAP7_75t_R FILLER_85_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_289 ();
 DECAPx2_ASAP7_75t_R FILLER_85_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_312 ();
 FILLER_ASAP7_75t_R FILLER_85_349 ();
 DECAPx1_ASAP7_75t_R FILLER_85_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_376 ();
 DECAPx2_ASAP7_75t_R FILLER_85_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_390 ();
 DECAPx4_ASAP7_75t_R FILLER_85_399 ();
 DECAPx4_ASAP7_75t_R FILLER_85_415 ();
 FILLER_ASAP7_75t_R FILLER_85_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_427 ();
 DECAPx4_ASAP7_75t_R FILLER_85_442 ();
 FILLER_ASAP7_75t_R FILLER_85_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_466 ();
 FILLER_ASAP7_75t_R FILLER_85_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_501 ();
 DECAPx4_ASAP7_75t_R FILLER_85_512 ();
 DECAPx2_ASAP7_75t_R FILLER_85_554 ();
 FILLER_ASAP7_75t_R FILLER_85_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_565 ();
 FILLER_ASAP7_75t_R FILLER_85_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_612 ();
 DECAPx6_ASAP7_75t_R FILLER_85_644 ();
 FILLER_ASAP7_75t_R FILLER_85_658 ();
 DECAPx10_ASAP7_75t_R FILLER_85_670 ();
 DECAPx10_ASAP7_75t_R FILLER_85_692 ();
 DECAPx10_ASAP7_75t_R FILLER_85_714 ();
 DECAPx10_ASAP7_75t_R FILLER_85_736 ();
 DECAPx4_ASAP7_75t_R FILLER_85_758 ();
 FILLER_ASAP7_75t_R FILLER_85_768 ();
 DECAPx6_ASAP7_75t_R FILLER_85_787 ();
 DECAPx4_ASAP7_75t_R FILLER_85_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_859 ();
 DECAPx4_ASAP7_75t_R FILLER_85_870 ();
 DECAPx1_ASAP7_75t_R FILLER_85_887 ();
 DECAPx6_ASAP7_75t_R FILLER_85_907 ();
 FILLER_ASAP7_75t_R FILLER_85_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_923 ();
 DECAPx2_ASAP7_75t_R FILLER_85_926 ();
 FILLER_ASAP7_75t_R FILLER_85_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_934 ();
 DECAPx2_ASAP7_75t_R FILLER_85_942 ();
 FILLER_ASAP7_75t_R FILLER_85_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_974 ();
 DECAPx1_ASAP7_75t_R FILLER_85_980 ();
 FILLER_ASAP7_75t_R FILLER_85_993 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1037 ();
 FILLER_ASAP7_75t_R FILLER_85_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1058 ();
 FILLER_ASAP7_75t_R FILLER_85_1064 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1084 ();
 FILLER_ASAP7_75t_R FILLER_85_1094 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1114 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1141 ();
 FILLER_ASAP7_75t_R FILLER_85_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1149 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1174 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1181 ();
 FILLER_ASAP7_75t_R FILLER_85_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1208 ();
 FILLER_ASAP7_75t_R FILLER_85_1230 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1258 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1272 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1284 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1310 ();
 FILLER_ASAP7_75t_R FILLER_85_1317 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1322 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1338 ();
 FILLER_ASAP7_75t_R FILLER_85_1348 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1350 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_86_2 ();
 FILLER_ASAP7_75t_R FILLER_86_8 ();
 DECAPx1_ASAP7_75t_R FILLER_86_16 ();
 DECAPx2_ASAP7_75t_R FILLER_86_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_55 ();
 FILLER_ASAP7_75t_R FILLER_86_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_64 ();
 DECAPx1_ASAP7_75t_R FILLER_86_74 ();
 DECAPx10_ASAP7_75t_R FILLER_86_81 ();
 DECAPx2_ASAP7_75t_R FILLER_86_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_109 ();
 DECAPx2_ASAP7_75t_R FILLER_86_122 ();
 DECAPx6_ASAP7_75t_R FILLER_86_134 ();
 DECAPx2_ASAP7_75t_R FILLER_86_151 ();
 FILLER_ASAP7_75t_R FILLER_86_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_159 ();
 DECAPx1_ASAP7_75t_R FILLER_86_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_205 ();
 DECAPx4_ASAP7_75t_R FILLER_86_230 ();
 FILLER_ASAP7_75t_R FILLER_86_240 ();
 DECAPx2_ASAP7_75t_R FILLER_86_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_262 ();
 DECAPx4_ASAP7_75t_R FILLER_86_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_302 ();
 DECAPx2_ASAP7_75t_R FILLER_86_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_329 ();
 FILLER_ASAP7_75t_R FILLER_86_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_344 ();
 FILLER_ASAP7_75t_R FILLER_86_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_367 ();
 DECAPx2_ASAP7_75t_R FILLER_86_376 ();
 FILLER_ASAP7_75t_R FILLER_86_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_384 ();
 DECAPx1_ASAP7_75t_R FILLER_86_399 ();
 DECAPx4_ASAP7_75t_R FILLER_86_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_427 ();
 DECAPx1_ASAP7_75t_R FILLER_86_470 ();
 DECAPx2_ASAP7_75t_R FILLER_86_480 ();
 FILLER_ASAP7_75t_R FILLER_86_486 ();
 DECAPx4_ASAP7_75t_R FILLER_86_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_501 ();
 DECAPx6_ASAP7_75t_R FILLER_86_509 ();
 DECAPx2_ASAP7_75t_R FILLER_86_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_536 ();
 FILLER_ASAP7_75t_R FILLER_86_540 ();
 DECAPx1_ASAP7_75t_R FILLER_86_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_578 ();
 DECAPx10_ASAP7_75t_R FILLER_86_615 ();
 FILLER_ASAP7_75t_R FILLER_86_637 ();
 DECAPx4_ASAP7_75t_R FILLER_86_645 ();
 DECAPx4_ASAP7_75t_R FILLER_86_661 ();
 FILLER_ASAP7_75t_R FILLER_86_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_673 ();
 DECAPx2_ASAP7_75t_R FILLER_86_677 ();
 DECAPx2_ASAP7_75t_R FILLER_86_686 ();
 DECAPx10_ASAP7_75t_R FILLER_86_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_740 ();
 DECAPx4_ASAP7_75t_R FILLER_86_767 ();
 DECAPx10_ASAP7_75t_R FILLER_86_784 ();
 DECAPx10_ASAP7_75t_R FILLER_86_806 ();
 DECAPx10_ASAP7_75t_R FILLER_86_828 ();
 DECAPx10_ASAP7_75t_R FILLER_86_850 ();
 DECAPx4_ASAP7_75t_R FILLER_86_872 ();
 FILLER_ASAP7_75t_R FILLER_86_882 ();
 DECAPx1_ASAP7_75t_R FILLER_86_897 ();
 FILLER_ASAP7_75t_R FILLER_86_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_924 ();
 FILLER_ASAP7_75t_R FILLER_86_933 ();
 DECAPx1_ASAP7_75t_R FILLER_86_945 ();
 DECAPx1_ASAP7_75t_R FILLER_86_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_959 ();
 FILLER_ASAP7_75t_R FILLER_86_996 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1024 ();
 FILLER_ASAP7_75t_R FILLER_86_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1096 ();
 FILLER_ASAP7_75t_R FILLER_86_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1117 ();
 FILLER_ASAP7_75t_R FILLER_86_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1143 ();
 FILLER_ASAP7_75t_R FILLER_86_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1151 ();
 DECAPx4_ASAP7_75t_R FILLER_86_1162 ();
 FILLER_ASAP7_75t_R FILLER_86_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1174 ();
 DECAPx4_ASAP7_75t_R FILLER_86_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1206 ();
 DECAPx4_ASAP7_75t_R FILLER_86_1233 ();
 FILLER_ASAP7_75t_R FILLER_86_1249 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1257 ();
 FILLER_ASAP7_75t_R FILLER_86_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1271 ();
 FILLER_ASAP7_75t_R FILLER_86_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1330 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1344 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1361 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_87_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_8 ();
 DECAPx6_ASAP7_75t_R FILLER_87_21 ();
 FILLER_ASAP7_75t_R FILLER_87_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_43 ();
 DECAPx1_ASAP7_75t_R FILLER_87_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_62 ();
 FILLER_ASAP7_75t_R FILLER_87_93 ();
 FILLER_ASAP7_75t_R FILLER_87_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_107 ();
 DECAPx10_ASAP7_75t_R FILLER_87_174 ();
 DECAPx6_ASAP7_75t_R FILLER_87_196 ();
 FILLER_ASAP7_75t_R FILLER_87_210 ();
 DECAPx6_ASAP7_75t_R FILLER_87_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_240 ();
 FILLER_ASAP7_75t_R FILLER_87_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_249 ();
 DECAPx2_ASAP7_75t_R FILLER_87_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_262 ();
 DECAPx2_ASAP7_75t_R FILLER_87_269 ();
 FILLER_ASAP7_75t_R FILLER_87_275 ();
 DECAPx6_ASAP7_75t_R FILLER_87_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_304 ();
 DECAPx4_ASAP7_75t_R FILLER_87_313 ();
 FILLER_ASAP7_75t_R FILLER_87_323 ();
 DECAPx6_ASAP7_75t_R FILLER_87_331 ();
 DECAPx1_ASAP7_75t_R FILLER_87_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_349 ();
 DECAPx1_ASAP7_75t_R FILLER_87_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_362 ();
 FILLER_ASAP7_75t_R FILLER_87_383 ();
 DECAPx1_ASAP7_75t_R FILLER_87_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_409 ();
 DECAPx4_ASAP7_75t_R FILLER_87_418 ();
 DECAPx1_ASAP7_75t_R FILLER_87_442 ();
 DECAPx1_ASAP7_75t_R FILLER_87_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_458 ();
 DECAPx10_ASAP7_75t_R FILLER_87_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_489 ();
 DECAPx6_ASAP7_75t_R FILLER_87_496 ();
 DECAPx1_ASAP7_75t_R FILLER_87_510 ();
 DECAPx2_ASAP7_75t_R FILLER_87_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_526 ();
 DECAPx6_ASAP7_75t_R FILLER_87_530 ();
 FILLER_ASAP7_75t_R FILLER_87_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_546 ();
 DECAPx4_ASAP7_75t_R FILLER_87_557 ();
 DECAPx2_ASAP7_75t_R FILLER_87_571 ();
 DECAPx4_ASAP7_75t_R FILLER_87_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_605 ();
 DECAPx4_ASAP7_75t_R FILLER_87_610 ();
 FILLER_ASAP7_75t_R FILLER_87_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_622 ();
 DECAPx2_ASAP7_75t_R FILLER_87_629 ();
 FILLER_ASAP7_75t_R FILLER_87_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_637 ();
 FILLER_ASAP7_75t_R FILLER_87_651 ();
 DECAPx1_ASAP7_75t_R FILLER_87_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_707 ();
 FILLER_ASAP7_75t_R FILLER_87_759 ();
 DECAPx2_ASAP7_75t_R FILLER_87_768 ();
 DECAPx10_ASAP7_75t_R FILLER_87_806 ();
 FILLER_ASAP7_75t_R FILLER_87_828 ();
 DECAPx1_ASAP7_75t_R FILLER_87_837 ();
 DECAPx1_ASAP7_75t_R FILLER_87_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_852 ();
 FILLER_ASAP7_75t_R FILLER_87_859 ();
 FILLER_ASAP7_75t_R FILLER_87_864 ();
 DECAPx2_ASAP7_75t_R FILLER_87_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_926 ();
 DECAPx6_ASAP7_75t_R FILLER_87_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_957 ();
 FILLER_ASAP7_75t_R FILLER_87_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_973 ();
 DECAPx6_ASAP7_75t_R FILLER_87_977 ();
 DECAPx2_ASAP7_75t_R FILLER_87_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_997 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1030 ();
 FILLER_ASAP7_75t_R FILLER_87_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1039 ();
 DECAPx6_ASAP7_75t_R FILLER_87_1060 ();
 FILLER_ASAP7_75t_R FILLER_87_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1102 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1129 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1137 ();
 FILLER_ASAP7_75t_R FILLER_87_1147 ();
 FILLER_ASAP7_75t_R FILLER_87_1171 ();
 FILLER_ASAP7_75t_R FILLER_87_1203 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1221 ();
 FILLER_ASAP7_75t_R FILLER_87_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1227 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1290 ();
 FILLER_ASAP7_75t_R FILLER_87_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1300 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1304 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1317 ();
 FILLER_ASAP7_75t_R FILLER_87_1323 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1325 ();
 FILLER_ASAP7_75t_R FILLER_87_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_32 ();
 FILLER_ASAP7_75t_R FILLER_88_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_61 ();
 DECAPx2_ASAP7_75t_R FILLER_88_118 ();
 DECAPx6_ASAP7_75t_R FILLER_88_127 ();
 FILLER_ASAP7_75t_R FILLER_88_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_143 ();
 DECAPx6_ASAP7_75t_R FILLER_88_156 ();
 DECAPx1_ASAP7_75t_R FILLER_88_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_174 ();
 FILLER_ASAP7_75t_R FILLER_88_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_183 ();
 DECAPx6_ASAP7_75t_R FILLER_88_190 ();
 DECAPx1_ASAP7_75t_R FILLER_88_204 ();
 DECAPx2_ASAP7_75t_R FILLER_88_224 ();
 DECAPx6_ASAP7_75t_R FILLER_88_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_250 ();
 DECAPx4_ASAP7_75t_R FILLER_88_257 ();
 FILLER_ASAP7_75t_R FILLER_88_273 ();
 DECAPx4_ASAP7_75t_R FILLER_88_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_293 ();
 DECAPx2_ASAP7_75t_R FILLER_88_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_306 ();
 DECAPx4_ASAP7_75t_R FILLER_88_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_343 ();
 DECAPx1_ASAP7_75t_R FILLER_88_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_399 ();
 DECAPx1_ASAP7_75t_R FILLER_88_406 ();
 DECAPx2_ASAP7_75t_R FILLER_88_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_455 ();
 DECAPx2_ASAP7_75t_R FILLER_88_464 ();
 FILLER_ASAP7_75t_R FILLER_88_470 ();
 DECAPx2_ASAP7_75t_R FILLER_88_478 ();
 FILLER_ASAP7_75t_R FILLER_88_484 ();
 DECAPx10_ASAP7_75t_R FILLER_88_538 ();
 DECAPx10_ASAP7_75t_R FILLER_88_560 ();
 DECAPx6_ASAP7_75t_R FILLER_88_582 ();
 DECAPx1_ASAP7_75t_R FILLER_88_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_600 ();
 DECAPx2_ASAP7_75t_R FILLER_88_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_613 ();
 DECAPx2_ASAP7_75t_R FILLER_88_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_641 ();
 FILLER_ASAP7_75t_R FILLER_88_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_682 ();
 DECAPx4_ASAP7_75t_R FILLER_88_695 ();
 DECAPx1_ASAP7_75t_R FILLER_88_720 ();
 FILLER_ASAP7_75t_R FILLER_88_740 ();
 DECAPx4_ASAP7_75t_R FILLER_88_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_759 ();
 DECAPx2_ASAP7_75t_R FILLER_88_789 ();
 DECAPx1_ASAP7_75t_R FILLER_88_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_833 ();
 DECAPx2_ASAP7_75t_R FILLER_88_866 ();
 FILLER_ASAP7_75t_R FILLER_88_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_874 ();
 DECAPx10_ASAP7_75t_R FILLER_88_894 ();
 DECAPx1_ASAP7_75t_R FILLER_88_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_920 ();
 DECAPx1_ASAP7_75t_R FILLER_88_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_935 ();
 DECAPx2_ASAP7_75t_R FILLER_88_949 ();
 DECAPx10_ASAP7_75t_R FILLER_88_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_985 ();
 FILLER_ASAP7_75t_R FILLER_88_996 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1005 ();
 FILLER_ASAP7_75t_R FILLER_88_1011 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1026 ();
 FILLER_ASAP7_75t_R FILLER_88_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1069 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1077 ();
 FILLER_ASAP7_75t_R FILLER_88_1087 ();
 FILLER_ASAP7_75t_R FILLER_88_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1121 ();
 FILLER_ASAP7_75t_R FILLER_88_1145 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1175 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1201 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1225 ();
 FILLER_ASAP7_75t_R FILLER_88_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1237 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1277 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1299 ();
 FILLER_ASAP7_75t_R FILLER_88_1309 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1343 ();
 FILLER_ASAP7_75t_R FILLER_88_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1357 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_89_2 ();
 FILLER_ASAP7_75t_R FILLER_89_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_10 ();
 DECAPx6_ASAP7_75t_R FILLER_89_20 ();
 FILLER_ASAP7_75t_R FILLER_89_46 ();
 DECAPx1_ASAP7_75t_R FILLER_89_51 ();
 FILLER_ASAP7_75t_R FILLER_89_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_67 ();
 DECAPx1_ASAP7_75t_R FILLER_89_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_81 ();
 DECAPx1_ASAP7_75t_R FILLER_89_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_90 ();
 DECAPx10_ASAP7_75t_R FILLER_89_97 ();
 DECAPx6_ASAP7_75t_R FILLER_89_119 ();
 DECAPx2_ASAP7_75t_R FILLER_89_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_139 ();
 DECAPx4_ASAP7_75t_R FILLER_89_156 ();
 FILLER_ASAP7_75t_R FILLER_89_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_168 ();
 DECAPx2_ASAP7_75t_R FILLER_89_205 ();
 FILLER_ASAP7_75t_R FILLER_89_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_213 ();
 DECAPx10_ASAP7_75t_R FILLER_89_222 ();
 DECAPx1_ASAP7_75t_R FILLER_89_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_248 ();
 DECAPx6_ASAP7_75t_R FILLER_89_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_271 ();
 DECAPx2_ASAP7_75t_R FILLER_89_306 ();
 FILLER_ASAP7_75t_R FILLER_89_312 ();
 FILLER_ASAP7_75t_R FILLER_89_328 ();
 DECAPx1_ASAP7_75t_R FILLER_89_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_348 ();
 DECAPx6_ASAP7_75t_R FILLER_89_355 ();
 FILLER_ASAP7_75t_R FILLER_89_369 ();
 DECAPx2_ASAP7_75t_R FILLER_89_377 ();
 FILLER_ASAP7_75t_R FILLER_89_383 ();
 DECAPx6_ASAP7_75t_R FILLER_89_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_405 ();
 DECAPx10_ASAP7_75t_R FILLER_89_420 ();
 DECAPx1_ASAP7_75t_R FILLER_89_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_446 ();
 DECAPx6_ASAP7_75t_R FILLER_89_455 ();
 FILLER_ASAP7_75t_R FILLER_89_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_471 ();
 DECAPx1_ASAP7_75t_R FILLER_89_501 ();
 DECAPx1_ASAP7_75t_R FILLER_89_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_579 ();
 FILLER_ASAP7_75t_R FILLER_89_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_588 ();
 DECAPx1_ASAP7_75t_R FILLER_89_595 ();
 FILLER_ASAP7_75t_R FILLER_89_625 ();
 DECAPx2_ASAP7_75t_R FILLER_89_651 ();
 FILLER_ASAP7_75t_R FILLER_89_657 ();
 DECAPx6_ASAP7_75t_R FILLER_89_663 ();
 DECAPx1_ASAP7_75t_R FILLER_89_677 ();
 DECAPx4_ASAP7_75t_R FILLER_89_687 ();
 FILLER_ASAP7_75t_R FILLER_89_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_699 ();
 DECAPx1_ASAP7_75t_R FILLER_89_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_711 ();
 FILLER_ASAP7_75t_R FILLER_89_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_717 ();
 DECAPx4_ASAP7_75t_R FILLER_89_724 ();
 FILLER_ASAP7_75t_R FILLER_89_750 ();
 DECAPx2_ASAP7_75t_R FILLER_89_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_776 ();
 FILLER_ASAP7_75t_R FILLER_89_789 ();
 DECAPx2_ASAP7_75t_R FILLER_89_794 ();
 DECAPx2_ASAP7_75t_R FILLER_89_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_822 ();
 DECAPx2_ASAP7_75t_R FILLER_89_838 ();
 FILLER_ASAP7_75t_R FILLER_89_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_853 ();
 DECAPx4_ASAP7_75t_R FILLER_89_867 ();
 FILLER_ASAP7_75t_R FILLER_89_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_879 ();
 DECAPx2_ASAP7_75t_R FILLER_89_887 ();
 FILLER_ASAP7_75t_R FILLER_89_893 ();
 DECAPx4_ASAP7_75t_R FILLER_89_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_917 ();
 FILLER_ASAP7_75t_R FILLER_89_952 ();
 DECAPx1_ASAP7_75t_R FILLER_89_980 ();
 FILLER_ASAP7_75t_R FILLER_89_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1083 ();
 FILLER_ASAP7_75t_R FILLER_89_1089 ();
 FILLER_ASAP7_75t_R FILLER_89_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_89_1109 ();
 DECAPx4_ASAP7_75t_R FILLER_89_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1147 ();
 FILLER_ASAP7_75t_R FILLER_89_1161 ();
 FILLER_ASAP7_75t_R FILLER_89_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1214 ();
 FILLER_ASAP7_75t_R FILLER_89_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1222 ();
 DECAPx4_ASAP7_75t_R FILLER_89_1249 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1272 ();
 FILLER_ASAP7_75t_R FILLER_89_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1286 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1308 ();
 FILLER_ASAP7_75t_R FILLER_89_1314 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1316 ();
 DECAPx4_ASAP7_75t_R FILLER_89_1335 ();
 FILLER_ASAP7_75t_R FILLER_89_1345 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1347 ();
 FILLER_ASAP7_75t_R FILLER_89_1358 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1379 ();
 DECAPx2_ASAP7_75t_R FILLER_90_28 ();
 DECAPx6_ASAP7_75t_R FILLER_90_43 ();
 DECAPx1_ASAP7_75t_R FILLER_90_83 ();
 FILLER_ASAP7_75t_R FILLER_90_93 ();
 DECAPx2_ASAP7_75t_R FILLER_90_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_131 ();
 DECAPx2_ASAP7_75t_R FILLER_90_158 ();
 FILLER_ASAP7_75t_R FILLER_90_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_194 ();
 DECAPx2_ASAP7_75t_R FILLER_90_215 ();
 FILLER_ASAP7_75t_R FILLER_90_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_223 ();
 FILLER_ASAP7_75t_R FILLER_90_258 ();
 DECAPx2_ASAP7_75t_R FILLER_90_266 ();
 DECAPx2_ASAP7_75t_R FILLER_90_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_299 ();
 DECAPx6_ASAP7_75t_R FILLER_90_312 ();
 FILLER_ASAP7_75t_R FILLER_90_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_336 ();
 DECAPx10_ASAP7_75t_R FILLER_90_343 ();
 DECAPx6_ASAP7_75t_R FILLER_90_365 ();
 DECAPx2_ASAP7_75t_R FILLER_90_379 ();
 DECAPx4_ASAP7_75t_R FILLER_90_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_409 ();
 DECAPx10_ASAP7_75t_R FILLER_90_422 ();
 DECAPx1_ASAP7_75t_R FILLER_90_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_448 ();
 DECAPx2_ASAP7_75t_R FILLER_90_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_461 ();
 FILLER_ASAP7_75t_R FILLER_90_464 ();
 DECAPx2_ASAP7_75t_R FILLER_90_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_484 ();
 DECAPx4_ASAP7_75t_R FILLER_90_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_504 ();
 DECAPx6_ASAP7_75t_R FILLER_90_511 ();
 FILLER_ASAP7_75t_R FILLER_90_525 ();
 DECAPx2_ASAP7_75t_R FILLER_90_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_539 ();
 DECAPx2_ASAP7_75t_R FILLER_90_543 ();
 FILLER_ASAP7_75t_R FILLER_90_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_557 ();
 FILLER_ASAP7_75t_R FILLER_90_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_586 ();
 DECAPx6_ASAP7_75t_R FILLER_90_613 ();
 DECAPx6_ASAP7_75t_R FILLER_90_633 ();
 DECAPx2_ASAP7_75t_R FILLER_90_665 ();
 DECAPx6_ASAP7_75t_R FILLER_90_723 ();
 DECAPx2_ASAP7_75t_R FILLER_90_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_743 ();
 FILLER_ASAP7_75t_R FILLER_90_754 ();
 DECAPx10_ASAP7_75t_R FILLER_90_766 ();
 DECAPx4_ASAP7_75t_R FILLER_90_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_798 ();
 FILLER_ASAP7_75t_R FILLER_90_805 ();
 DECAPx6_ASAP7_75t_R FILLER_90_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_827 ();
 DECAPx2_ASAP7_75t_R FILLER_90_848 ();
 FILLER_ASAP7_75t_R FILLER_90_854 ();
 DECAPx6_ASAP7_75t_R FILLER_90_863 ();
 DECAPx1_ASAP7_75t_R FILLER_90_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_881 ();
 DECAPx2_ASAP7_75t_R FILLER_90_890 ();
 FILLER_ASAP7_75t_R FILLER_90_896 ();
 FILLER_ASAP7_75t_R FILLER_90_906 ();
 DECAPx2_ASAP7_75t_R FILLER_90_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_939 ();
 DECAPx6_ASAP7_75t_R FILLER_90_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_957 ();
 DECAPx2_ASAP7_75t_R FILLER_90_961 ();
 FILLER_ASAP7_75t_R FILLER_90_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_972 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1059 ();
 FILLER_ASAP7_75t_R FILLER_90_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1105 ();
 DECAPx6_ASAP7_75t_R FILLER_90_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1141 ();
 FILLER_ASAP7_75t_R FILLER_90_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1164 ();
 FILLER_ASAP7_75t_R FILLER_90_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1223 ();
 FILLER_ASAP7_75t_R FILLER_90_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1247 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1269 ();
 FILLER_ASAP7_75t_R FILLER_90_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1277 ();
 DECAPx6_ASAP7_75t_R FILLER_90_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1308 ();
 FILLER_ASAP7_75t_R FILLER_90_1330 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1332 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1339 ();
 FILLER_ASAP7_75t_R FILLER_90_1345 ();
 FILLER_ASAP7_75t_R FILLER_90_1357 ();
 FILLER_ASAP7_75t_R FILLER_90_1378 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_91_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_12 ();
 FILLER_ASAP7_75t_R FILLER_91_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_24 ();
 FILLER_ASAP7_75t_R FILLER_91_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_57 ();
 DECAPx4_ASAP7_75t_R FILLER_91_64 ();
 FILLER_ASAP7_75t_R FILLER_91_74 ();
 FILLER_ASAP7_75t_R FILLER_91_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_104 ();
 FILLER_ASAP7_75t_R FILLER_91_111 ();
 FILLER_ASAP7_75t_R FILLER_91_116 ();
 FILLER_ASAP7_75t_R FILLER_91_144 ();
 DECAPx4_ASAP7_75t_R FILLER_91_155 ();
 DECAPx6_ASAP7_75t_R FILLER_91_179 ();
 DECAPx2_ASAP7_75t_R FILLER_91_215 ();
 FILLER_ASAP7_75t_R FILLER_91_239 ();
 FILLER_ASAP7_75t_R FILLER_91_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_263 ();
 DECAPx2_ASAP7_75t_R FILLER_91_278 ();
 FILLER_ASAP7_75t_R FILLER_91_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_286 ();
 DECAPx4_ASAP7_75t_R FILLER_91_315 ();
 DECAPx1_ASAP7_75t_R FILLER_91_347 ();
 DECAPx1_ASAP7_75t_R FILLER_91_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_363 ();
 DECAPx2_ASAP7_75t_R FILLER_91_370 ();
 FILLER_ASAP7_75t_R FILLER_91_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_398 ();
 DECAPx6_ASAP7_75t_R FILLER_91_405 ();
 FILLER_ASAP7_75t_R FILLER_91_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_427 ();
 DECAPx4_ASAP7_75t_R FILLER_91_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_444 ();
 DECAPx4_ASAP7_75t_R FILLER_91_453 ();
 FILLER_ASAP7_75t_R FILLER_91_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_465 ();
 DECAPx4_ASAP7_75t_R FILLER_91_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_495 ();
 DECAPx6_ASAP7_75t_R FILLER_91_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_528 ();
 DECAPx1_ASAP7_75t_R FILLER_91_547 ();
 DECAPx2_ASAP7_75t_R FILLER_91_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_563 ();
 DECAPx1_ASAP7_75t_R FILLER_91_567 ();
 DECAPx1_ASAP7_75t_R FILLER_91_584 ();
 DECAPx1_ASAP7_75t_R FILLER_91_594 ();
 FILLER_ASAP7_75t_R FILLER_91_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_609 ();
 FILLER_ASAP7_75t_R FILLER_91_622 ();
 DECAPx10_ASAP7_75t_R FILLER_91_631 ();
 DECAPx1_ASAP7_75t_R FILLER_91_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_657 ();
 DECAPx4_ASAP7_75t_R FILLER_91_664 ();
 FILLER_ASAP7_75t_R FILLER_91_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_690 ();
 DECAPx1_ASAP7_75t_R FILLER_91_694 ();
 DECAPx4_ASAP7_75t_R FILLER_91_704 ();
 FILLER_ASAP7_75t_R FILLER_91_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_716 ();
 DECAPx2_ASAP7_75t_R FILLER_91_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_733 ();
 DECAPx6_ASAP7_75t_R FILLER_91_741 ();
 FILLER_ASAP7_75t_R FILLER_91_755 ();
 FILLER_ASAP7_75t_R FILLER_91_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_772 ();
 DECAPx6_ASAP7_75t_R FILLER_91_799 ();
 FILLER_ASAP7_75t_R FILLER_91_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_825 ();
 DECAPx6_ASAP7_75t_R FILLER_91_833 ();
 FILLER_ASAP7_75t_R FILLER_91_847 ();
 DECAPx4_ASAP7_75t_R FILLER_91_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_875 ();
 DECAPx4_ASAP7_75t_R FILLER_91_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_896 ();
 FILLER_ASAP7_75t_R FILLER_91_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_917 ();
 DECAPx1_ASAP7_75t_R FILLER_91_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_930 ();
 DECAPx2_ASAP7_75t_R FILLER_91_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_970 ();
 DECAPx2_ASAP7_75t_R FILLER_91_983 ();
 FILLER_ASAP7_75t_R FILLER_91_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_991 ();
 DECAPx4_ASAP7_75t_R FILLER_91_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1028 ();
 FILLER_ASAP7_75t_R FILLER_91_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_91_1087 ();
 FILLER_ASAP7_75t_R FILLER_91_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1099 ();
 DECAPx4_ASAP7_75t_R FILLER_91_1108 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1130 ();
 DECAPx4_ASAP7_75t_R FILLER_91_1141 ();
 FILLER_ASAP7_75t_R FILLER_91_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1180 ();
 DECAPx4_ASAP7_75t_R FILLER_91_1202 ();
 FILLER_ASAP7_75t_R FILLER_91_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1261 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1330 ();
 DECAPx4_ASAP7_75t_R FILLER_91_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_92_2 ();
 DECAPx2_ASAP7_75t_R FILLER_92_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_22 ();
 DECAPx1_ASAP7_75t_R FILLER_92_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_31 ();
 DECAPx6_ASAP7_75t_R FILLER_92_38 ();
 DECAPx1_ASAP7_75t_R FILLER_92_52 ();
 DECAPx2_ASAP7_75t_R FILLER_92_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_68 ();
 DECAPx2_ASAP7_75t_R FILLER_92_72 ();
 FILLER_ASAP7_75t_R FILLER_92_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_80 ();
 FILLER_ASAP7_75t_R FILLER_92_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_89 ();
 DECAPx1_ASAP7_75t_R FILLER_92_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_97 ();
 DECAPx2_ASAP7_75t_R FILLER_92_110 ();
 FILLER_ASAP7_75t_R FILLER_92_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_131 ();
 DECAPx4_ASAP7_75t_R FILLER_92_135 ();
 FILLER_ASAP7_75t_R FILLER_92_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_147 ();
 FILLER_ASAP7_75t_R FILLER_92_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_183 ();
 DECAPx4_ASAP7_75t_R FILLER_92_190 ();
 FILLER_ASAP7_75t_R FILLER_92_200 ();
 DECAPx1_ASAP7_75t_R FILLER_92_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_212 ();
 DECAPx1_ASAP7_75t_R FILLER_92_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_223 ();
 DECAPx2_ASAP7_75t_R FILLER_92_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_246 ();
 DECAPx1_ASAP7_75t_R FILLER_92_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_271 ();
 DECAPx10_ASAP7_75t_R FILLER_92_292 ();
 DECAPx6_ASAP7_75t_R FILLER_92_314 ();
 DECAPx1_ASAP7_75t_R FILLER_92_328 ();
 DECAPx6_ASAP7_75t_R FILLER_92_338 ();
 FILLER_ASAP7_75t_R FILLER_92_352 ();
 FILLER_ASAP7_75t_R FILLER_92_368 ();
 DECAPx4_ASAP7_75t_R FILLER_92_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_386 ();
 FILLER_ASAP7_75t_R FILLER_92_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_438 ();
 FILLER_ASAP7_75t_R FILLER_92_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_464 ();
 DECAPx1_ASAP7_75t_R FILLER_92_473 ();
 DECAPx2_ASAP7_75t_R FILLER_92_492 ();
 FILLER_ASAP7_75t_R FILLER_92_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_500 ();
 DECAPx10_ASAP7_75t_R FILLER_92_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_539 ();
 FILLER_ASAP7_75t_R FILLER_92_546 ();
 DECAPx10_ASAP7_75t_R FILLER_92_554 ();
 FILLER_ASAP7_75t_R FILLER_92_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_578 ();
 DECAPx6_ASAP7_75t_R FILLER_92_591 ();
 DECAPx1_ASAP7_75t_R FILLER_92_605 ();
 DECAPx4_ASAP7_75t_R FILLER_92_625 ();
 FILLER_ASAP7_75t_R FILLER_92_635 ();
 DECAPx2_ASAP7_75t_R FILLER_92_645 ();
 FILLER_ASAP7_75t_R FILLER_92_651 ();
 DECAPx4_ASAP7_75t_R FILLER_92_663 ();
 FILLER_ASAP7_75t_R FILLER_92_673 ();
 DECAPx2_ASAP7_75t_R FILLER_92_690 ();
 FILLER_ASAP7_75t_R FILLER_92_696 ();
 DECAPx2_ASAP7_75t_R FILLER_92_705 ();
 FILLER_ASAP7_75t_R FILLER_92_714 ();
 DECAPx2_ASAP7_75t_R FILLER_92_748 ();
 FILLER_ASAP7_75t_R FILLER_92_754 ();
 FILLER_ASAP7_75t_R FILLER_92_782 ();
 FILLER_ASAP7_75t_R FILLER_92_803 ();
 DECAPx2_ASAP7_75t_R FILLER_92_843 ();
 DECAPx2_ASAP7_75t_R FILLER_92_895 ();
 DECAPx4_ASAP7_75t_R FILLER_92_909 ();
 DECAPx10_ASAP7_75t_R FILLER_92_925 ();
 DECAPx1_ASAP7_75t_R FILLER_92_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_951 ();
 DECAPx2_ASAP7_75t_R FILLER_92_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_961 ();
 DECAPx10_ASAP7_75t_R FILLER_92_980 ();
 FILLER_ASAP7_75t_R FILLER_92_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1043 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1062 ();
 FILLER_ASAP7_75t_R FILLER_92_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1100 ();
 FILLER_ASAP7_75t_R FILLER_92_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1163 ();
 FILLER_ASAP7_75t_R FILLER_92_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1185 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1224 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1269 ();
 FILLER_ASAP7_75t_R FILLER_92_1289 ();
 FILLER_ASAP7_75t_R FILLER_92_1303 ();
 FILLER_ASAP7_75t_R FILLER_92_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1379 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_93_28 ();
 FILLER_ASAP7_75t_R FILLER_93_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_40 ();
 FILLER_ASAP7_75t_R FILLER_93_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_84 ();
 DECAPx6_ASAP7_75t_R FILLER_93_88 ();
 DECAPx2_ASAP7_75t_R FILLER_93_128 ();
 FILLER_ASAP7_75t_R FILLER_93_134 ();
 DECAPx1_ASAP7_75t_R FILLER_93_162 ();
 DECAPx10_ASAP7_75t_R FILLER_93_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_202 ();
 FILLER_ASAP7_75t_R FILLER_93_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_219 ();
 FILLER_ASAP7_75t_R FILLER_93_226 ();
 DECAPx10_ASAP7_75t_R FILLER_93_244 ();
 DECAPx2_ASAP7_75t_R FILLER_93_266 ();
 FILLER_ASAP7_75t_R FILLER_93_272 ();
 DECAPx10_ASAP7_75t_R FILLER_93_280 ();
 DECAPx1_ASAP7_75t_R FILLER_93_302 ();
 DECAPx2_ASAP7_75t_R FILLER_93_319 ();
 FILLER_ASAP7_75t_R FILLER_93_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_338 ();
 FILLER_ASAP7_75t_R FILLER_93_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_353 ();
 DECAPx1_ASAP7_75t_R FILLER_93_368 ();
 DECAPx4_ASAP7_75t_R FILLER_93_380 ();
 FILLER_ASAP7_75t_R FILLER_93_390 ();
 DECAPx1_ASAP7_75t_R FILLER_93_404 ();
 DECAPx4_ASAP7_75t_R FILLER_93_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_440 ();
 DECAPx1_ASAP7_75t_R FILLER_93_447 ();
 DECAPx2_ASAP7_75t_R FILLER_93_457 ();
 FILLER_ASAP7_75t_R FILLER_93_463 ();
 DECAPx2_ASAP7_75t_R FILLER_93_477 ();
 FILLER_ASAP7_75t_R FILLER_93_483 ();
 DECAPx1_ASAP7_75t_R FILLER_93_500 ();
 FILLER_ASAP7_75t_R FILLER_93_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_522 ();
 DECAPx2_ASAP7_75t_R FILLER_93_529 ();
 FILLER_ASAP7_75t_R FILLER_93_535 ();
 DECAPx1_ASAP7_75t_R FILLER_93_559 ();
 FILLER_ASAP7_75t_R FILLER_93_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_577 ();
 FILLER_ASAP7_75t_R FILLER_93_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_612 ();
 FILLER_ASAP7_75t_R FILLER_93_631 ();
 FILLER_ASAP7_75t_R FILLER_93_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_677 ();
 DECAPx4_ASAP7_75t_R FILLER_93_684 ();
 FILLER_ASAP7_75t_R FILLER_93_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_696 ();
 DECAPx2_ASAP7_75t_R FILLER_93_723 ();
 DECAPx4_ASAP7_75t_R FILLER_93_750 ();
 DECAPx1_ASAP7_75t_R FILLER_93_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_770 ();
 FILLER_ASAP7_75t_R FILLER_93_774 ();
 FILLER_ASAP7_75t_R FILLER_93_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_784 ();
 FILLER_ASAP7_75t_R FILLER_93_791 ();
 DECAPx6_ASAP7_75t_R FILLER_93_799 ();
 DECAPx2_ASAP7_75t_R FILLER_93_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_823 ();
 DECAPx2_ASAP7_75t_R FILLER_93_836 ();
 FILLER_ASAP7_75t_R FILLER_93_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_844 ();
 DECAPx2_ASAP7_75t_R FILLER_93_865 ();
 FILLER_ASAP7_75t_R FILLER_93_871 ();
 FILLER_ASAP7_75t_R FILLER_93_882 ();
 DECAPx1_ASAP7_75t_R FILLER_93_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_901 ();
 FILLER_ASAP7_75t_R FILLER_93_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_916 ();
 DECAPx6_ASAP7_75t_R FILLER_93_952 ();
 FILLER_ASAP7_75t_R FILLER_93_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_995 ();
 DECAPx4_ASAP7_75t_R FILLER_93_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1023 ();
 FILLER_ASAP7_75t_R FILLER_93_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1055 ();
 FILLER_ASAP7_75t_R FILLER_93_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1063 ();
 DECAPx4_ASAP7_75t_R FILLER_93_1072 ();
 FILLER_ASAP7_75t_R FILLER_93_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1129 ();
 FILLER_ASAP7_75t_R FILLER_93_1135 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1147 ();
 FILLER_ASAP7_75t_R FILLER_93_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1166 ();
 DECAPx4_ASAP7_75t_R FILLER_93_1188 ();
 FILLER_ASAP7_75t_R FILLER_93_1198 ();
 FILLER_ASAP7_75t_R FILLER_93_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1226 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1280 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1302 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1308 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1321 ();
 FILLER_ASAP7_75t_R FILLER_93_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1329 ();
 FILLER_ASAP7_75t_R FILLER_93_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_94_2 ();
 DECAPx2_ASAP7_75t_R FILLER_94_99 ();
 FILLER_ASAP7_75t_R FILLER_94_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_107 ();
 FILLER_ASAP7_75t_R FILLER_94_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_116 ();
 DECAPx2_ASAP7_75t_R FILLER_94_120 ();
 FILLER_ASAP7_75t_R FILLER_94_126 ();
 DECAPx6_ASAP7_75t_R FILLER_94_134 ();
 FILLER_ASAP7_75t_R FILLER_94_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_150 ();
 FILLER_ASAP7_75t_R FILLER_94_154 ();
 DECAPx2_ASAP7_75t_R FILLER_94_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_168 ();
 DECAPx6_ASAP7_75t_R FILLER_94_175 ();
 DECAPx2_ASAP7_75t_R FILLER_94_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_195 ();
 DECAPx2_ASAP7_75t_R FILLER_94_222 ();
 DECAPx10_ASAP7_75t_R FILLER_94_234 ();
 DECAPx4_ASAP7_75t_R FILLER_94_256 ();
 FILLER_ASAP7_75t_R FILLER_94_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_268 ();
 DECAPx2_ASAP7_75t_R FILLER_94_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_294 ();
 DECAPx2_ASAP7_75t_R FILLER_94_305 ();
 FILLER_ASAP7_75t_R FILLER_94_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_313 ();
 DECAPx1_ASAP7_75t_R FILLER_94_324 ();
 DECAPx1_ASAP7_75t_R FILLER_94_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_362 ();
 DECAPx2_ASAP7_75t_R FILLER_94_389 ();
 FILLER_ASAP7_75t_R FILLER_94_395 ();
 DECAPx6_ASAP7_75t_R FILLER_94_403 ();
 DECAPx2_ASAP7_75t_R FILLER_94_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_423 ();
 DECAPx1_ASAP7_75t_R FILLER_94_432 ();
 DECAPx2_ASAP7_75t_R FILLER_94_442 ();
 DECAPx2_ASAP7_75t_R FILLER_94_454 ();
 FILLER_ASAP7_75t_R FILLER_94_460 ();
 DECAPx1_ASAP7_75t_R FILLER_94_464 ();
 DECAPx6_ASAP7_75t_R FILLER_94_474 ();
 DECAPx4_ASAP7_75t_R FILLER_94_495 ();
 DECAPx2_ASAP7_75t_R FILLER_94_515 ();
 FILLER_ASAP7_75t_R FILLER_94_521 ();
 DECAPx4_ASAP7_75t_R FILLER_94_529 ();
 DECAPx6_ASAP7_75t_R FILLER_94_549 ();
 FILLER_ASAP7_75t_R FILLER_94_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_577 ();
 DECAPx4_ASAP7_75t_R FILLER_94_604 ();
 FILLER_ASAP7_75t_R FILLER_94_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_629 ();
 DECAPx6_ASAP7_75t_R FILLER_94_642 ();
 DECAPx2_ASAP7_75t_R FILLER_94_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_662 ();
 DECAPx2_ASAP7_75t_R FILLER_94_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_672 ();
 DECAPx2_ASAP7_75t_R FILLER_94_683 ();
 FILLER_ASAP7_75t_R FILLER_94_702 ();
 DECAPx1_ASAP7_75t_R FILLER_94_707 ();
 DECAPx1_ASAP7_75t_R FILLER_94_714 ();
 DECAPx4_ASAP7_75t_R FILLER_94_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_734 ();
 FILLER_ASAP7_75t_R FILLER_94_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_743 ();
 DECAPx1_ASAP7_75t_R FILLER_94_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_752 ();
 DECAPx10_ASAP7_75t_R FILLER_94_763 ();
 DECAPx6_ASAP7_75t_R FILLER_94_785 ();
 DECAPx2_ASAP7_75t_R FILLER_94_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_805 ();
 DECAPx4_ASAP7_75t_R FILLER_94_812 ();
 FILLER_ASAP7_75t_R FILLER_94_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_830 ();
 DECAPx6_ASAP7_75t_R FILLER_94_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_851 ();
 DECAPx6_ASAP7_75t_R FILLER_94_855 ();
 DECAPx1_ASAP7_75t_R FILLER_94_869 ();
 FILLER_ASAP7_75t_R FILLER_94_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_881 ();
 DECAPx2_ASAP7_75t_R FILLER_94_888 ();
 FILLER_ASAP7_75t_R FILLER_94_894 ();
 FILLER_ASAP7_75t_R FILLER_94_903 ();
 FILLER_ASAP7_75t_R FILLER_94_937 ();
 FILLER_ASAP7_75t_R FILLER_94_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_944 ();
 DECAPx4_ASAP7_75t_R FILLER_94_948 ();
 FILLER_ASAP7_75t_R FILLER_94_958 ();
 DECAPx1_ASAP7_75t_R FILLER_94_978 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1008 ();
 FILLER_ASAP7_75t_R FILLER_94_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1016 ();
 FILLER_ASAP7_75t_R FILLER_94_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1032 ();
 FILLER_ASAP7_75t_R FILLER_94_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1083 ();
 FILLER_ASAP7_75t_R FILLER_94_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1091 ();
 FILLER_ASAP7_75t_R FILLER_94_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1104 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1108 ();
 FILLER_ASAP7_75t_R FILLER_94_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1126 ();
 FILLER_ASAP7_75t_R FILLER_94_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1152 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1171 ();
 FILLER_ASAP7_75t_R FILLER_94_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1183 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1194 ();
 FILLER_ASAP7_75t_R FILLER_94_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1223 ();
 FILLER_ASAP7_75t_R FILLER_94_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1237 ();
 FILLER_ASAP7_75t_R FILLER_94_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1255 ();
 FILLER_ASAP7_75t_R FILLER_94_1277 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1279 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1297 ();
 DECAPx6_ASAP7_75t_R FILLER_94_1311 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1325 ();
 DECAPx6_ASAP7_75t_R FILLER_94_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1349 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1360 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1364 ();
 FILLER_ASAP7_75t_R FILLER_94_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1388 ();
 DECAPx1_ASAP7_75t_R FILLER_95_2 ();
 FILLER_ASAP7_75t_R FILLER_95_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_33 ();
 DECAPx1_ASAP7_75t_R FILLER_95_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_48 ();
 DECAPx6_ASAP7_75t_R FILLER_95_52 ();
 DECAPx1_ASAP7_75t_R FILLER_95_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_70 ();
 DECAPx6_ASAP7_75t_R FILLER_95_77 ();
 DECAPx1_ASAP7_75t_R FILLER_95_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_95 ();
 FILLER_ASAP7_75t_R FILLER_95_102 ();
 DECAPx6_ASAP7_75t_R FILLER_95_107 ();
 FILLER_ASAP7_75t_R FILLER_95_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_123 ();
 DECAPx6_ASAP7_75t_R FILLER_95_150 ();
 DECAPx1_ASAP7_75t_R FILLER_95_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_168 ();
 DECAPx1_ASAP7_75t_R FILLER_95_177 ();
 DECAPx1_ASAP7_75t_R FILLER_95_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_193 ();
 DECAPx6_ASAP7_75t_R FILLER_95_208 ();
 FILLER_ASAP7_75t_R FILLER_95_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_224 ();
 DECAPx4_ASAP7_75t_R FILLER_95_231 ();
 FILLER_ASAP7_75t_R FILLER_95_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_243 ();
 DECAPx6_ASAP7_75t_R FILLER_95_250 ();
 DECAPx2_ASAP7_75t_R FILLER_95_264 ();
 DECAPx1_ASAP7_75t_R FILLER_95_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_288 ();
 DECAPx1_ASAP7_75t_R FILLER_95_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_307 ();
 DECAPx2_ASAP7_75t_R FILLER_95_322 ();
 FILLER_ASAP7_75t_R FILLER_95_328 ();
 DECAPx2_ASAP7_75t_R FILLER_95_356 ();
 FILLER_ASAP7_75t_R FILLER_95_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_364 ();
 DECAPx4_ASAP7_75t_R FILLER_95_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_387 ();
 DECAPx1_ASAP7_75t_R FILLER_95_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_406 ();
 FILLER_ASAP7_75t_R FILLER_95_427 ();
 DECAPx2_ASAP7_75t_R FILLER_95_435 ();
 FILLER_ASAP7_75t_R FILLER_95_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_443 ();
 FILLER_ASAP7_75t_R FILLER_95_450 ();
 DECAPx1_ASAP7_75t_R FILLER_95_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_463 ();
 DECAPx10_ASAP7_75t_R FILLER_95_478 ();
 DECAPx2_ASAP7_75t_R FILLER_95_500 ();
 FILLER_ASAP7_75t_R FILLER_95_506 ();
 DECAPx1_ASAP7_75t_R FILLER_95_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_520 ();
 DECAPx1_ASAP7_75t_R FILLER_95_544 ();
 FILLER_ASAP7_75t_R FILLER_95_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_562 ();
 DECAPx2_ASAP7_75t_R FILLER_95_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_579 ();
 FILLER_ASAP7_75t_R FILLER_95_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_597 ();
 DECAPx4_ASAP7_75t_R FILLER_95_601 ();
 FILLER_ASAP7_75t_R FILLER_95_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_613 ();
 DECAPx2_ASAP7_75t_R FILLER_95_620 ();
 FILLER_ASAP7_75t_R FILLER_95_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_628 ();
 DECAPx2_ASAP7_75t_R FILLER_95_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_641 ();
 DECAPx6_ASAP7_75t_R FILLER_95_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_662 ();
 DECAPx2_ASAP7_75t_R FILLER_95_666 ();
 DECAPx1_ASAP7_75t_R FILLER_95_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_689 ();
 DECAPx2_ASAP7_75t_R FILLER_95_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_722 ();
 DECAPx10_ASAP7_75t_R FILLER_95_729 ();
 DECAPx2_ASAP7_75t_R FILLER_95_751 ();
 FILLER_ASAP7_75t_R FILLER_95_757 ();
 DECAPx2_ASAP7_75t_R FILLER_95_766 ();
 FILLER_ASAP7_75t_R FILLER_95_775 ();
 DECAPx6_ASAP7_75t_R FILLER_95_815 ();
 DECAPx6_ASAP7_75t_R FILLER_95_835 ();
 DECAPx4_ASAP7_75t_R FILLER_95_862 ();
 FILLER_ASAP7_75t_R FILLER_95_872 ();
 DECAPx2_ASAP7_75t_R FILLER_95_890 ();
 FILLER_ASAP7_75t_R FILLER_95_896 ();
 DECAPx2_ASAP7_75t_R FILLER_95_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_923 ();
 DECAPx10_ASAP7_75t_R FILLER_95_926 ();
 DECAPx4_ASAP7_75t_R FILLER_95_948 ();
 FILLER_ASAP7_75t_R FILLER_95_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_960 ();
 DECAPx2_ASAP7_75t_R FILLER_95_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_985 ();
 DECAPx6_ASAP7_75t_R FILLER_95_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1040 ();
 FILLER_ASAP7_75t_R FILLER_95_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1048 ();
 FILLER_ASAP7_75t_R FILLER_95_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1128 ();
 FILLER_ASAP7_75t_R FILLER_95_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_95_1173 ();
 FILLER_ASAP7_75t_R FILLER_95_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1271 ();
 FILLER_ASAP7_75t_R FILLER_95_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1339 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1367 ();
 DECAPx1_ASAP7_75t_R FILLER_96_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_6 ();
 FILLER_ASAP7_75t_R FILLER_96_13 ();
 DECAPx4_ASAP7_75t_R FILLER_96_18 ();
 DECAPx10_ASAP7_75t_R FILLER_96_34 ();
 FILLER_ASAP7_75t_R FILLER_96_56 ();
 DECAPx1_ASAP7_75t_R FILLER_96_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_68 ();
 DECAPx6_ASAP7_75t_R FILLER_96_72 ();
 FILLER_ASAP7_75t_R FILLER_96_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_88 ();
 DECAPx2_ASAP7_75t_R FILLER_96_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_124 ();
 DECAPx2_ASAP7_75t_R FILLER_96_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_137 ();
 DECAPx2_ASAP7_75t_R FILLER_96_141 ();
 FILLER_ASAP7_75t_R FILLER_96_147 ();
 FILLER_ASAP7_75t_R FILLER_96_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_161 ();
 DECAPx1_ASAP7_75t_R FILLER_96_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_180 ();
 DECAPx1_ASAP7_75t_R FILLER_96_189 ();
 DECAPx1_ASAP7_75t_R FILLER_96_209 ();
 DECAPx1_ASAP7_75t_R FILLER_96_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_252 ();
 DECAPx2_ASAP7_75t_R FILLER_96_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_265 ();
 DECAPx1_ASAP7_75t_R FILLER_96_274 ();
 FILLER_ASAP7_75t_R FILLER_96_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_288 ();
 FILLER_ASAP7_75t_R FILLER_96_303 ();
 DECAPx6_ASAP7_75t_R FILLER_96_325 ();
 DECAPx1_ASAP7_75t_R FILLER_96_339 ();
 FILLER_ASAP7_75t_R FILLER_96_357 ();
 DECAPx2_ASAP7_75t_R FILLER_96_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_395 ();
 FILLER_ASAP7_75t_R FILLER_96_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_406 ();
 DECAPx10_ASAP7_75t_R FILLER_96_421 ();
 DECAPx1_ASAP7_75t_R FILLER_96_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_461 ();
 DECAPx2_ASAP7_75t_R FILLER_96_486 ();
 FILLER_ASAP7_75t_R FILLER_96_492 ();
 DECAPx2_ASAP7_75t_R FILLER_96_502 ();
 DECAPx6_ASAP7_75t_R FILLER_96_521 ();
 FILLER_ASAP7_75t_R FILLER_96_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_537 ();
 DECAPx2_ASAP7_75t_R FILLER_96_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_580 ();
 DECAPx6_ASAP7_75t_R FILLER_96_588 ();
 DECAPx2_ASAP7_75t_R FILLER_96_602 ();
 FILLER_ASAP7_75t_R FILLER_96_614 ();
 DECAPx6_ASAP7_75t_R FILLER_96_622 ();
 FILLER_ASAP7_75t_R FILLER_96_636 ();
 FILLER_ASAP7_75t_R FILLER_96_674 ();
 DECAPx1_ASAP7_75t_R FILLER_96_688 ();
 FILLER_ASAP7_75t_R FILLER_96_698 ();
 DECAPx1_ASAP7_75t_R FILLER_96_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_710 ();
 DECAPx2_ASAP7_75t_R FILLER_96_749 ();
 FILLER_ASAP7_75t_R FILLER_96_755 ();
 DECAPx2_ASAP7_75t_R FILLER_96_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_789 ();
 DECAPx4_ASAP7_75t_R FILLER_96_809 ();
 FILLER_ASAP7_75t_R FILLER_96_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_825 ();
 DECAPx1_ASAP7_75t_R FILLER_96_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_837 ();
 FILLER_ASAP7_75t_R FILLER_96_864 ();
 DECAPx4_ASAP7_75t_R FILLER_96_876 ();
 DECAPx6_ASAP7_75t_R FILLER_96_892 ();
 DECAPx4_ASAP7_75t_R FILLER_96_912 ();
 FILLER_ASAP7_75t_R FILLER_96_931 ();
 DECAPx10_ASAP7_75t_R FILLER_96_939 ();
 DECAPx10_ASAP7_75t_R FILLER_96_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_983 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1010 ();
 FILLER_ASAP7_75t_R FILLER_96_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1037 ();
 DECAPx4_ASAP7_75t_R FILLER_96_1056 ();
 DECAPx4_ASAP7_75t_R FILLER_96_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1097 ();
 FILLER_ASAP7_75t_R FILLER_96_1112 ();
 DECAPx1_ASAP7_75t_R FILLER_96_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1169 ();
 FILLER_ASAP7_75t_R FILLER_96_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1177 ();
 FILLER_ASAP7_75t_R FILLER_96_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1216 ();
 FILLER_ASAP7_75t_R FILLER_96_1243 ();
 DECAPx1_ASAP7_75t_R FILLER_96_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1293 ();
 FILLER_ASAP7_75t_R FILLER_96_1306 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1321 ();
 FILLER_ASAP7_75t_R FILLER_96_1327 ();
 DECAPx1_ASAP7_75t_R FILLER_96_1342 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1363 ();
 FILLER_ASAP7_75t_R FILLER_96_1369 ();
 FILLER_ASAP7_75t_R FILLER_96_1378 ();
 DECAPx1_ASAP7_75t_R FILLER_96_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_97_2 ();
 FILLER_ASAP7_75t_R FILLER_97_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_53 ();
 DECAPx1_ASAP7_75t_R FILLER_97_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_91 ();
 DECAPx2_ASAP7_75t_R FILLER_97_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_104 ();
 FILLER_ASAP7_75t_R FILLER_97_137 ();
 DECAPx1_ASAP7_75t_R FILLER_97_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_150 ();
 DECAPx6_ASAP7_75t_R FILLER_97_154 ();
 FILLER_ASAP7_75t_R FILLER_97_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_188 ();
 FILLER_ASAP7_75t_R FILLER_97_201 ();
 DECAPx2_ASAP7_75t_R FILLER_97_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_215 ();
 FILLER_ASAP7_75t_R FILLER_97_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_226 ();
 FILLER_ASAP7_75t_R FILLER_97_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_251 ();
 DECAPx2_ASAP7_75t_R FILLER_97_258 ();
 DECAPx6_ASAP7_75t_R FILLER_97_297 ();
 DECAPx1_ASAP7_75t_R FILLER_97_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_321 ();
 DECAPx4_ASAP7_75t_R FILLER_97_329 ();
 FILLER_ASAP7_75t_R FILLER_97_339 ();
 DECAPx6_ASAP7_75t_R FILLER_97_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_361 ();
 DECAPx1_ASAP7_75t_R FILLER_97_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_372 ();
 FILLER_ASAP7_75t_R FILLER_97_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_381 ();
 DECAPx6_ASAP7_75t_R FILLER_97_388 ();
 DECAPx1_ASAP7_75t_R FILLER_97_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_412 ();
 DECAPx2_ASAP7_75t_R FILLER_97_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_425 ();
 DECAPx2_ASAP7_75t_R FILLER_97_454 ();
 FILLER_ASAP7_75t_R FILLER_97_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_462 ();
 FILLER_ASAP7_75t_R FILLER_97_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_485 ();
 FILLER_ASAP7_75t_R FILLER_97_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_496 ();
 DECAPx4_ASAP7_75t_R FILLER_97_511 ();
 FILLER_ASAP7_75t_R FILLER_97_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_523 ();
 DECAPx1_ASAP7_75t_R FILLER_97_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_547 ();
 DECAPx6_ASAP7_75t_R FILLER_97_560 ();
 DECAPx2_ASAP7_75t_R FILLER_97_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_580 ();
 DECAPx4_ASAP7_75t_R FILLER_97_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_630 ();
 DECAPx2_ASAP7_75t_R FILLER_97_637 ();
 FILLER_ASAP7_75t_R FILLER_97_643 ();
 DECAPx4_ASAP7_75t_R FILLER_97_662 ();
 DECAPx6_ASAP7_75t_R FILLER_97_679 ();
 DECAPx1_ASAP7_75t_R FILLER_97_693 ();
 DECAPx4_ASAP7_75t_R FILLER_97_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_713 ();
 DECAPx1_ASAP7_75t_R FILLER_97_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_725 ();
 DECAPx1_ASAP7_75t_R FILLER_97_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_733 ();
 FILLER_ASAP7_75t_R FILLER_97_752 ();
 DECAPx1_ASAP7_75t_R FILLER_97_773 ();
 DECAPx4_ASAP7_75t_R FILLER_97_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_806 ();
 FILLER_ASAP7_75t_R FILLER_97_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_865 ();
 DECAPx4_ASAP7_75t_R FILLER_97_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_908 ();
 DECAPx2_ASAP7_75t_R FILLER_97_915 ();
 FILLER_ASAP7_75t_R FILLER_97_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_923 ();
 DECAPx1_ASAP7_75t_R FILLER_97_926 ();
 DECAPx2_ASAP7_75t_R FILLER_97_963 ();
 DECAPx4_ASAP7_75t_R FILLER_97_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_989 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1046 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1057 ();
 FILLER_ASAP7_75t_R FILLER_97_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1076 ();
 FILLER_ASAP7_75t_R FILLER_97_1083 ();
 FILLER_ASAP7_75t_R FILLER_97_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1111 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1128 ();
 FILLER_ASAP7_75t_R FILLER_97_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1151 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1161 ();
 FILLER_ASAP7_75t_R FILLER_97_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1220 ();
 FILLER_ASAP7_75t_R FILLER_97_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1236 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1271 ();
 FILLER_ASAP7_75t_R FILLER_97_1277 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1285 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1324 ();
 FILLER_ASAP7_75t_R FILLER_97_1345 ();
 FILLER_ASAP7_75t_R FILLER_97_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1369 ();
 DECAPx1_ASAP7_75t_R FILLER_98_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_56 ();
 DECAPx1_ASAP7_75t_R FILLER_98_63 ();
 DECAPx4_ASAP7_75t_R FILLER_98_103 ();
 DECAPx2_ASAP7_75t_R FILLER_98_119 ();
 DECAPx2_ASAP7_75t_R FILLER_98_128 ();
 FILLER_ASAP7_75t_R FILLER_98_134 ();
 DECAPx1_ASAP7_75t_R FILLER_98_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_166 ();
 FILLER_ASAP7_75t_R FILLER_98_181 ();
 DECAPx10_ASAP7_75t_R FILLER_98_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_211 ();
 DECAPx4_ASAP7_75t_R FILLER_98_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_240 ();
 DECAPx4_ASAP7_75t_R FILLER_98_255 ();
 DECAPx4_ASAP7_75t_R FILLER_98_277 ();
 FILLER_ASAP7_75t_R FILLER_98_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_289 ();
 DECAPx4_ASAP7_75t_R FILLER_98_297 ();
 FILLER_ASAP7_75t_R FILLER_98_307 ();
 FILLER_ASAP7_75t_R FILLER_98_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_323 ();
 FILLER_ASAP7_75t_R FILLER_98_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_340 ();
 DECAPx4_ASAP7_75t_R FILLER_98_349 ();
 FILLER_ASAP7_75t_R FILLER_98_359 ();
 DECAPx10_ASAP7_75t_R FILLER_98_367 ();
 FILLER_ASAP7_75t_R FILLER_98_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_391 ();
 DECAPx4_ASAP7_75t_R FILLER_98_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_420 ();
 DECAPx1_ASAP7_75t_R FILLER_98_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_437 ();
 FILLER_ASAP7_75t_R FILLER_98_460 ();
 DECAPx2_ASAP7_75t_R FILLER_98_464 ();
 FILLER_ASAP7_75t_R FILLER_98_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_472 ();
 DECAPx4_ASAP7_75t_R FILLER_98_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_489 ();
 FILLER_ASAP7_75t_R FILLER_98_497 ();
 FILLER_ASAP7_75t_R FILLER_98_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_507 ();
 DECAPx1_ASAP7_75t_R FILLER_98_515 ();
 DECAPx4_ASAP7_75t_R FILLER_98_534 ();
 DECAPx6_ASAP7_75t_R FILLER_98_551 ();
 DECAPx1_ASAP7_75t_R FILLER_98_565 ();
 FILLER_ASAP7_75t_R FILLER_98_581 ();
 DECAPx2_ASAP7_75t_R FILLER_98_589 ();
 DECAPx4_ASAP7_75t_R FILLER_98_598 ();
 DECAPx1_ASAP7_75t_R FILLER_98_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_630 ();
 DECAPx1_ASAP7_75t_R FILLER_98_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_641 ();
 DECAPx1_ASAP7_75t_R FILLER_98_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_687 ();
 FILLER_ASAP7_75t_R FILLER_98_701 ();
 DECAPx4_ASAP7_75t_R FILLER_98_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_731 ();
 DECAPx2_ASAP7_75t_R FILLER_98_751 ();
 DECAPx4_ASAP7_75t_R FILLER_98_763 ();
 FILLER_ASAP7_75t_R FILLER_98_773 ();
 FILLER_ASAP7_75t_R FILLER_98_781 ();
 DECAPx1_ASAP7_75t_R FILLER_98_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_799 ();
 DECAPx6_ASAP7_75t_R FILLER_98_810 ();
 FILLER_ASAP7_75t_R FILLER_98_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_826 ();
 DECAPx2_ASAP7_75t_R FILLER_98_839 ();
 FILLER_ASAP7_75t_R FILLER_98_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_847 ();
 FILLER_ASAP7_75t_R FILLER_98_854 ();
 FILLER_ASAP7_75t_R FILLER_98_868 ();
 DECAPx4_ASAP7_75t_R FILLER_98_877 ();
 DECAPx1_ASAP7_75t_R FILLER_98_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_907 ();
 DECAPx1_ASAP7_75t_R FILLER_98_916 ();
 DECAPx1_ASAP7_75t_R FILLER_98_962 ();
 DECAPx1_ASAP7_75t_R FILLER_98_992 ();
 DECAPx4_ASAP7_75t_R FILLER_98_1002 ();
 DECAPx6_ASAP7_75t_R FILLER_98_1022 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1040 ();
 DECAPx4_ASAP7_75t_R FILLER_98_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1067 ();
 FILLER_ASAP7_75t_R FILLER_98_1087 ();
 DECAPx4_ASAP7_75t_R FILLER_98_1107 ();
 FILLER_ASAP7_75t_R FILLER_98_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1129 ();
 FILLER_ASAP7_75t_R FILLER_98_1135 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1149 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1215 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1254 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1276 ();
 FILLER_ASAP7_75t_R FILLER_98_1302 ();
 DECAPx4_ASAP7_75t_R FILLER_98_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1327 ();
 DECAPx4_ASAP7_75t_R FILLER_98_1340 ();
 FILLER_ASAP7_75t_R FILLER_98_1350 ();
 FILLER_ASAP7_75t_R FILLER_98_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1367 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_99_2 ();
 FILLER_ASAP7_75t_R FILLER_99_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_14 ();
 DECAPx1_ASAP7_75t_R FILLER_99_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_22 ();
 DECAPx1_ASAP7_75t_R FILLER_99_27 ();
 DECAPx6_ASAP7_75t_R FILLER_99_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_82 ();
 DECAPx1_ASAP7_75t_R FILLER_99_115 ();
 DECAPx2_ASAP7_75t_R FILLER_99_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_128 ();
 DECAPx4_ASAP7_75t_R FILLER_99_135 ();
 DECAPx4_ASAP7_75t_R FILLER_99_151 ();
 FILLER_ASAP7_75t_R FILLER_99_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_163 ();
 DECAPx4_ASAP7_75t_R FILLER_99_184 ();
 FILLER_ASAP7_75t_R FILLER_99_200 ();
 DECAPx4_ASAP7_75t_R FILLER_99_214 ();
 FILLER_ASAP7_75t_R FILLER_99_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_226 ();
 DECAPx2_ASAP7_75t_R FILLER_99_233 ();
 DECAPx2_ASAP7_75t_R FILLER_99_253 ();
 DECAPx1_ASAP7_75t_R FILLER_99_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_269 ();
 DECAPx6_ASAP7_75t_R FILLER_99_276 ();
 FILLER_ASAP7_75t_R FILLER_99_290 ();
 DECAPx2_ASAP7_75t_R FILLER_99_300 ();
 FILLER_ASAP7_75t_R FILLER_99_314 ();
 FILLER_ASAP7_75t_R FILLER_99_324 ();
 DECAPx2_ASAP7_75t_R FILLER_99_348 ();
 FILLER_ASAP7_75t_R FILLER_99_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_356 ();
 DECAPx10_ASAP7_75t_R FILLER_99_369 ();
 DECAPx2_ASAP7_75t_R FILLER_99_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_423 ();
 DECAPx4_ASAP7_75t_R FILLER_99_432 ();
 FILLER_ASAP7_75t_R FILLER_99_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_450 ();
 DECAPx2_ASAP7_75t_R FILLER_99_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_463 ();
 FILLER_ASAP7_75t_R FILLER_99_476 ();
 FILLER_ASAP7_75t_R FILLER_99_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_511 ();
 FILLER_ASAP7_75t_R FILLER_99_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_522 ();
 DECAPx10_ASAP7_75t_R FILLER_99_529 ();
 DECAPx1_ASAP7_75t_R FILLER_99_551 ();
 DECAPx6_ASAP7_75t_R FILLER_99_584 ();
 DECAPx1_ASAP7_75t_R FILLER_99_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_602 ();
 DECAPx1_ASAP7_75t_R FILLER_99_613 ();
 DECAPx1_ASAP7_75t_R FILLER_99_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_636 ();
 DECAPx6_ASAP7_75t_R FILLER_99_643 ();
 DECAPx1_ASAP7_75t_R FILLER_99_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_689 ();
 DECAPx4_ASAP7_75t_R FILLER_99_697 ();
 FILLER_ASAP7_75t_R FILLER_99_707 ();
 DECAPx4_ASAP7_75t_R FILLER_99_728 ();
 DECAPx1_ASAP7_75t_R FILLER_99_751 ();
 DECAPx1_ASAP7_75t_R FILLER_99_799 ();
 DECAPx2_ASAP7_75t_R FILLER_99_821 ();
 DECAPx10_ASAP7_75t_R FILLER_99_839 ();
 FILLER_ASAP7_75t_R FILLER_99_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_863 ();
 DECAPx10_ASAP7_75t_R FILLER_99_871 ();
 DECAPx1_ASAP7_75t_R FILLER_99_908 ();
 FILLER_ASAP7_75t_R FILLER_99_922 ();
 FILLER_ASAP7_75t_R FILLER_99_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_928 ();
 DECAPx4_ASAP7_75t_R FILLER_99_935 ();
 FILLER_ASAP7_75t_R FILLER_99_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_947 ();
 DECAPx4_ASAP7_75t_R FILLER_99_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_980 ();
 FILLER_ASAP7_75t_R FILLER_99_984 ();
 DECAPx2_ASAP7_75t_R FILLER_99_992 ();
 FILLER_ASAP7_75t_R FILLER_99_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1000 ();
 FILLER_ASAP7_75t_R FILLER_99_1011 ();
 FILLER_ASAP7_75t_R FILLER_99_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1073 ();
 DECAPx4_ASAP7_75t_R FILLER_99_1088 ();
 FILLER_ASAP7_75t_R FILLER_99_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1209 ();
 DECAPx6_ASAP7_75t_R FILLER_99_1225 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1243 ();
 DECAPx4_ASAP7_75t_R FILLER_99_1262 ();
 FILLER_ASAP7_75t_R FILLER_99_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1280 ();
 DECAPx4_ASAP7_75t_R FILLER_99_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1330 ();
 DECAPx6_ASAP7_75t_R FILLER_99_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1378 ();
 FILLER_ASAP7_75t_R FILLER_99_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_100_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_6 ();
 DECAPx10_ASAP7_75t_R FILLER_100_13 ();
 FILLER_ASAP7_75t_R FILLER_100_35 ();
 DECAPx2_ASAP7_75t_R FILLER_100_43 ();
 DECAPx2_ASAP7_75t_R FILLER_100_75 ();
 FILLER_ASAP7_75t_R FILLER_100_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_83 ();
 DECAPx4_ASAP7_75t_R FILLER_100_90 ();
 DECAPx4_ASAP7_75t_R FILLER_100_152 ();
 FILLER_ASAP7_75t_R FILLER_100_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_192 ();
 DECAPx1_ASAP7_75t_R FILLER_100_207 ();
 DECAPx4_ASAP7_75t_R FILLER_100_217 ();
 FILLER_ASAP7_75t_R FILLER_100_227 ();
 DECAPx4_ASAP7_75t_R FILLER_100_235 ();
 FILLER_ASAP7_75t_R FILLER_100_245 ();
 DECAPx1_ASAP7_75t_R FILLER_100_253 ();
 DECAPx1_ASAP7_75t_R FILLER_100_263 ();
 DECAPx1_ASAP7_75t_R FILLER_100_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_277 ();
 FILLER_ASAP7_75t_R FILLER_100_285 ();
 DECAPx2_ASAP7_75t_R FILLER_100_302 ();
 DECAPx2_ASAP7_75t_R FILLER_100_331 ();
 FILLER_ASAP7_75t_R FILLER_100_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_339 ();
 DECAPx1_ASAP7_75t_R FILLER_100_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_350 ();
 DECAPx1_ASAP7_75t_R FILLER_100_377 ();
 DECAPx4_ASAP7_75t_R FILLER_100_389 ();
 FILLER_ASAP7_75t_R FILLER_100_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_401 ();
 FILLER_ASAP7_75t_R FILLER_100_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_426 ();
 DECAPx1_ASAP7_75t_R FILLER_100_435 ();
 DECAPx2_ASAP7_75t_R FILLER_100_453 ();
 FILLER_ASAP7_75t_R FILLER_100_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_461 ();
 DECAPx1_ASAP7_75t_R FILLER_100_464 ();
 DECAPx4_ASAP7_75t_R FILLER_100_476 ();
 FILLER_ASAP7_75t_R FILLER_100_486 ();
 DECAPx6_ASAP7_75t_R FILLER_100_496 ();
 FILLER_ASAP7_75t_R FILLER_100_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_512 ();
 DECAPx6_ASAP7_75t_R FILLER_100_521 ();
 DECAPx1_ASAP7_75t_R FILLER_100_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_539 ();
 FILLER_ASAP7_75t_R FILLER_100_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_557 ();
 DECAPx1_ASAP7_75t_R FILLER_100_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_570 ();
 DECAPx4_ASAP7_75t_R FILLER_100_585 ();
 DECAPx1_ASAP7_75t_R FILLER_100_601 ();
 DECAPx2_ASAP7_75t_R FILLER_100_608 ();
 DECAPx4_ASAP7_75t_R FILLER_100_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_650 ();
 DECAPx6_ASAP7_75t_R FILLER_100_665 ();
 FILLER_ASAP7_75t_R FILLER_100_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_681 ();
 DECAPx4_ASAP7_75t_R FILLER_100_694 ();
 DECAPx2_ASAP7_75t_R FILLER_100_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_713 ();
 FILLER_ASAP7_75t_R FILLER_100_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_719 ();
 FILLER_ASAP7_75t_R FILLER_100_728 ();
 FILLER_ASAP7_75t_R FILLER_100_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_754 ();
 DECAPx2_ASAP7_75t_R FILLER_100_762 ();
 FILLER_ASAP7_75t_R FILLER_100_768 ();
 FILLER_ASAP7_75t_R FILLER_100_773 ();
 DECAPx1_ASAP7_75t_R FILLER_100_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_782 ();
 DECAPx4_ASAP7_75t_R FILLER_100_803 ();
 FILLER_ASAP7_75t_R FILLER_100_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_815 ();
 DECAPx1_ASAP7_75t_R FILLER_100_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_827 ();
 FILLER_ASAP7_75t_R FILLER_100_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_840 ();
 FILLER_ASAP7_75t_R FILLER_100_847 ();
 FILLER_ASAP7_75t_R FILLER_100_855 ();
 DECAPx2_ASAP7_75t_R FILLER_100_870 ();
 FILLER_ASAP7_75t_R FILLER_100_876 ();
 FILLER_ASAP7_75t_R FILLER_100_890 ();
 DECAPx6_ASAP7_75t_R FILLER_100_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_924 ();
 DECAPx10_ASAP7_75t_R FILLER_100_931 ();
 DECAPx6_ASAP7_75t_R FILLER_100_953 ();
 DECAPx1_ASAP7_75t_R FILLER_100_967 ();
 DECAPx4_ASAP7_75t_R FILLER_100_977 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1017 ();
 FILLER_ASAP7_75t_R FILLER_100_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1026 ();
 DECAPx4_ASAP7_75t_R FILLER_100_1030 ();
 FILLER_ASAP7_75t_R FILLER_100_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1067 ();
 FILLER_ASAP7_75t_R FILLER_100_1081 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1103 ();
 FILLER_ASAP7_75t_R FILLER_100_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1121 ();
 FILLER_ASAP7_75t_R FILLER_100_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1129 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1167 ();
 FILLER_ASAP7_75t_R FILLER_100_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1237 ();
 FILLER_ASAP7_75t_R FILLER_100_1243 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1294 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1316 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1320 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1357 ();
 DECAPx4_ASAP7_75t_R FILLER_100_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1377 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_101_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_62 ();
 FILLER_ASAP7_75t_R FILLER_101_72 ();
 DECAPx2_ASAP7_75t_R FILLER_101_78 ();
 FILLER_ASAP7_75t_R FILLER_101_84 ();
 DECAPx1_ASAP7_75t_R FILLER_101_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_96 ();
 DECAPx1_ASAP7_75t_R FILLER_101_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_104 ();
 DECAPx6_ASAP7_75t_R FILLER_101_111 ();
 FILLER_ASAP7_75t_R FILLER_101_125 ();
 FILLER_ASAP7_75t_R FILLER_101_133 ();
 DECAPx1_ASAP7_75t_R FILLER_101_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_168 ();
 FILLER_ASAP7_75t_R FILLER_101_175 ();
 DECAPx4_ASAP7_75t_R FILLER_101_183 ();
 FILLER_ASAP7_75t_R FILLER_101_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_195 ();
 DECAPx2_ASAP7_75t_R FILLER_101_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_208 ();
 FILLER_ASAP7_75t_R FILLER_101_241 ();
 DECAPx1_ASAP7_75t_R FILLER_101_269 ();
 DECAPx6_ASAP7_75t_R FILLER_101_279 ();
 FILLER_ASAP7_75t_R FILLER_101_293 ();
 DECAPx6_ASAP7_75t_R FILLER_101_318 ();
 DECAPx1_ASAP7_75t_R FILLER_101_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_336 ();
 FILLER_ASAP7_75t_R FILLER_101_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_358 ();
 DECAPx6_ASAP7_75t_R FILLER_101_373 ();
 DECAPx2_ASAP7_75t_R FILLER_101_387 ();
 DECAPx2_ASAP7_75t_R FILLER_101_411 ();
 FILLER_ASAP7_75t_R FILLER_101_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_419 ();
 DECAPx1_ASAP7_75t_R FILLER_101_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_438 ();
 FILLER_ASAP7_75t_R FILLER_101_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_455 ();
 DECAPx1_ASAP7_75t_R FILLER_101_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_490 ();
 DECAPx2_ASAP7_75t_R FILLER_101_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_550 ();
 DECAPx4_ASAP7_75t_R FILLER_101_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_577 ();
 FILLER_ASAP7_75t_R FILLER_101_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_590 ();
 DECAPx1_ASAP7_75t_R FILLER_101_617 ();
 FILLER_ASAP7_75t_R FILLER_101_638 ();
 FILLER_ASAP7_75t_R FILLER_101_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_660 ();
 DECAPx6_ASAP7_75t_R FILLER_101_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_691 ();
 DECAPx2_ASAP7_75t_R FILLER_101_699 ();
 DECAPx2_ASAP7_75t_R FILLER_101_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_714 ();
 DECAPx4_ASAP7_75t_R FILLER_101_718 ();
 FILLER_ASAP7_75t_R FILLER_101_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_730 ();
 DECAPx2_ASAP7_75t_R FILLER_101_749 ();
 DECAPx2_ASAP7_75t_R FILLER_101_761 ();
 FILLER_ASAP7_75t_R FILLER_101_767 ();
 DECAPx4_ASAP7_75t_R FILLER_101_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_811 ();
 DECAPx1_ASAP7_75t_R FILLER_101_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_868 ();
 DECAPx4_ASAP7_75t_R FILLER_101_887 ();
 FILLER_ASAP7_75t_R FILLER_101_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_899 ();
 DECAPx6_ASAP7_75t_R FILLER_101_908 ();
 FILLER_ASAP7_75t_R FILLER_101_922 ();
 FILLER_ASAP7_75t_R FILLER_101_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_928 ();
 DECAPx2_ASAP7_75t_R FILLER_101_936 ();
 DECAPx1_ASAP7_75t_R FILLER_101_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_955 ();
 DECAPx6_ASAP7_75t_R FILLER_101_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_989 ();
 DECAPx1_ASAP7_75t_R FILLER_101_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1004 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1026 ();
 FILLER_ASAP7_75t_R FILLER_101_1040 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1086 ();
 FILLER_ASAP7_75t_R FILLER_101_1097 ();
 FILLER_ASAP7_75t_R FILLER_101_1119 ();
 FILLER_ASAP7_75t_R FILLER_101_1131 ();
 FILLER_ASAP7_75t_R FILLER_101_1147 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1169 ();
 FILLER_ASAP7_75t_R FILLER_101_1179 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1211 ();
 FILLER_ASAP7_75t_R FILLER_101_1221 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1231 ();
 FILLER_ASAP7_75t_R FILLER_101_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1243 ();
 FILLER_ASAP7_75t_R FILLER_101_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1290 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1318 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1340 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1384 ();
 FILLER_ASAP7_75t_R FILLER_101_1390 ();
 DECAPx2_ASAP7_75t_R FILLER_102_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_8 ();
 DECAPx6_ASAP7_75t_R FILLER_102_45 ();
 DECAPx1_ASAP7_75t_R FILLER_102_59 ();
 DECAPx4_ASAP7_75t_R FILLER_102_93 ();
 FILLER_ASAP7_75t_R FILLER_102_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_110 ();
 DECAPx1_ASAP7_75t_R FILLER_102_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_121 ();
 DECAPx6_ASAP7_75t_R FILLER_102_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_152 ();
 DECAPx1_ASAP7_75t_R FILLER_102_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_160 ();
 DECAPx6_ASAP7_75t_R FILLER_102_165 ();
 DECAPx4_ASAP7_75t_R FILLER_102_185 ();
 DECAPx4_ASAP7_75t_R FILLER_102_201 ();
 FILLER_ASAP7_75t_R FILLER_102_211 ();
 DECAPx2_ASAP7_75t_R FILLER_102_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_227 ();
 DECAPx4_ASAP7_75t_R FILLER_102_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_257 ();
 DECAPx2_ASAP7_75t_R FILLER_102_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_292 ();
 DECAPx10_ASAP7_75t_R FILLER_102_305 ();
 DECAPx6_ASAP7_75t_R FILLER_102_327 ();
 DECAPx1_ASAP7_75t_R FILLER_102_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_351 ();
 DECAPx1_ASAP7_75t_R FILLER_102_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_368 ();
 DECAPx2_ASAP7_75t_R FILLER_102_383 ();
 DECAPx2_ASAP7_75t_R FILLER_102_431 ();
 FILLER_ASAP7_75t_R FILLER_102_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_439 ();
 DECAPx4_ASAP7_75t_R FILLER_102_450 ();
 FILLER_ASAP7_75t_R FILLER_102_460 ();
 DECAPx4_ASAP7_75t_R FILLER_102_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_491 ();
 DECAPx2_ASAP7_75t_R FILLER_102_506 ();
 DECAPx10_ASAP7_75t_R FILLER_102_542 ();
 FILLER_ASAP7_75t_R FILLER_102_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_566 ();
 DECAPx4_ASAP7_75t_R FILLER_102_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_583 ();
 DECAPx1_ASAP7_75t_R FILLER_102_590 ();
 DECAPx2_ASAP7_75t_R FILLER_102_600 ();
 FILLER_ASAP7_75t_R FILLER_102_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_608 ();
 DECAPx6_ASAP7_75t_R FILLER_102_621 ();
 DECAPx1_ASAP7_75t_R FILLER_102_635 ();
 DECAPx6_ASAP7_75t_R FILLER_102_659 ();
 DECAPx1_ASAP7_75t_R FILLER_102_697 ();
 DECAPx4_ASAP7_75t_R FILLER_102_713 ();
 DECAPx10_ASAP7_75t_R FILLER_102_729 ();
 DECAPx10_ASAP7_75t_R FILLER_102_751 ();
 DECAPx4_ASAP7_75t_R FILLER_102_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_783 ();
 DECAPx4_ASAP7_75t_R FILLER_102_791 ();
 DECAPx4_ASAP7_75t_R FILLER_102_817 ();
 FILLER_ASAP7_75t_R FILLER_102_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_829 ();
 DECAPx6_ASAP7_75t_R FILLER_102_836 ();
 FILLER_ASAP7_75t_R FILLER_102_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_852 ();
 DECAPx4_ASAP7_75t_R FILLER_102_859 ();
 FILLER_ASAP7_75t_R FILLER_102_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_871 ();
 DECAPx1_ASAP7_75t_R FILLER_102_890 ();
 DECAPx6_ASAP7_75t_R FILLER_102_900 ();
 FILLER_ASAP7_75t_R FILLER_102_914 ();
 FILLER_ASAP7_75t_R FILLER_102_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_930 ();
 FILLER_ASAP7_75t_R FILLER_102_966 ();
 DECAPx6_ASAP7_75t_R FILLER_102_985 ();
 DECAPx1_ASAP7_75t_R FILLER_102_999 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1013 ();
 FILLER_ASAP7_75t_R FILLER_102_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1021 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1063 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1077 ();
 FILLER_ASAP7_75t_R FILLER_102_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1114 ();
 FILLER_ASAP7_75t_R FILLER_102_1125 ();
 FILLER_ASAP7_75t_R FILLER_102_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1135 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1167 ();
 FILLER_ASAP7_75t_R FILLER_102_1193 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1265 ();
 FILLER_ASAP7_75t_R FILLER_102_1279 ();
 FILLER_ASAP7_75t_R FILLER_102_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1289 ();
 FILLER_ASAP7_75t_R FILLER_102_1296 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1298 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1307 ();
 FILLER_ASAP7_75t_R FILLER_102_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1323 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1340 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1344 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1377 ();
 FILLER_ASAP7_75t_R FILLER_102_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_103_2 ();
 FILLER_ASAP7_75t_R FILLER_103_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_19 ();
 DECAPx2_ASAP7_75t_R FILLER_103_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_46 ();
 DECAPx6_ASAP7_75t_R FILLER_103_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_64 ();
 DECAPx2_ASAP7_75t_R FILLER_103_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_80 ();
 DECAPx4_ASAP7_75t_R FILLER_103_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_147 ();
 DECAPx4_ASAP7_75t_R FILLER_103_160 ();
 FILLER_ASAP7_75t_R FILLER_103_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_172 ();
 FILLER_ASAP7_75t_R FILLER_103_187 ();
 DECAPx4_ASAP7_75t_R FILLER_103_203 ();
 DECAPx4_ASAP7_75t_R FILLER_103_219 ();
 FILLER_ASAP7_75t_R FILLER_103_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_261 ();
 DECAPx2_ASAP7_75t_R FILLER_103_268 ();
 DECAPx2_ASAP7_75t_R FILLER_103_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_288 ();
 DECAPx2_ASAP7_75t_R FILLER_103_307 ();
 DECAPx2_ASAP7_75t_R FILLER_103_325 ();
 FILLER_ASAP7_75t_R FILLER_103_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_333 ();
 DECAPx10_ASAP7_75t_R FILLER_103_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_376 ();
 DECAPx10_ASAP7_75t_R FILLER_103_385 ();
 DECAPx4_ASAP7_75t_R FILLER_103_407 ();
 DECAPx6_ASAP7_75t_R FILLER_103_430 ();
 DECAPx1_ASAP7_75t_R FILLER_103_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_448 ();
 DECAPx4_ASAP7_75t_R FILLER_103_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_465 ();
 DECAPx2_ASAP7_75t_R FILLER_103_472 ();
 FILLER_ASAP7_75t_R FILLER_103_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_500 ();
 FILLER_ASAP7_75t_R FILLER_103_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_511 ();
 FILLER_ASAP7_75t_R FILLER_103_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_536 ();
 DECAPx6_ASAP7_75t_R FILLER_103_543 ();
 DECAPx2_ASAP7_75t_R FILLER_103_557 ();
 DECAPx2_ASAP7_75t_R FILLER_103_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_579 ();
 DECAPx6_ASAP7_75t_R FILLER_103_606 ();
 DECAPx1_ASAP7_75t_R FILLER_103_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_636 ();
 DECAPx6_ASAP7_75t_R FILLER_103_643 ();
 DECAPx2_ASAP7_75t_R FILLER_103_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_663 ();
 DECAPx6_ASAP7_75t_R FILLER_103_671 ();
 DECAPx1_ASAP7_75t_R FILLER_103_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_706 ();
 FILLER_ASAP7_75t_R FILLER_103_713 ();
 DECAPx4_ASAP7_75t_R FILLER_103_731 ();
 FILLER_ASAP7_75t_R FILLER_103_741 ();
 FILLER_ASAP7_75t_R FILLER_103_754 ();
 DECAPx6_ASAP7_75t_R FILLER_103_762 ();
 DECAPx10_ASAP7_75t_R FILLER_103_786 ();
 DECAPx6_ASAP7_75t_R FILLER_103_808 ();
 FILLER_ASAP7_75t_R FILLER_103_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_824 ();
 DECAPx10_ASAP7_75t_R FILLER_103_831 ();
 DECAPx1_ASAP7_75t_R FILLER_103_853 ();
 DECAPx6_ASAP7_75t_R FILLER_103_864 ();
 FILLER_ASAP7_75t_R FILLER_103_884 ();
 FILLER_ASAP7_75t_R FILLER_103_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_912 ();
 DECAPx1_ASAP7_75t_R FILLER_103_932 ();
 FILLER_ASAP7_75t_R FILLER_103_972 ();
 FILLER_ASAP7_75t_R FILLER_103_994 ();
 FILLER_ASAP7_75t_R FILLER_103_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1004 ();
 FILLER_ASAP7_75t_R FILLER_103_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1044 ();
 FILLER_ASAP7_75t_R FILLER_103_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1062 ();
 DECAPx1_ASAP7_75t_R FILLER_103_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1096 ();
 FILLER_ASAP7_75t_R FILLER_103_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1126 ();
 FILLER_ASAP7_75t_R FILLER_103_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1163 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1185 ();
 FILLER_ASAP7_75t_R FILLER_103_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_103_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1231 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1245 ();
 FILLER_ASAP7_75t_R FILLER_103_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1253 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1267 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1291 ();
 FILLER_ASAP7_75t_R FILLER_103_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1299 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1306 ();
 FILLER_ASAP7_75t_R FILLER_103_1312 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1314 ();
 DECAPx1_ASAP7_75t_R FILLER_103_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1333 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1355 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1368 ();
 FILLER_ASAP7_75t_R FILLER_103_1390 ();
 FILLER_ASAP7_75t_R FILLER_104_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_4 ();
 DECAPx6_ASAP7_75t_R FILLER_104_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_31 ();
 DECAPx1_ASAP7_75t_R FILLER_104_62 ();
 DECAPx2_ASAP7_75t_R FILLER_104_72 ();
 FILLER_ASAP7_75t_R FILLER_104_78 ();
 DECAPx2_ASAP7_75t_R FILLER_104_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_98 ();
 FILLER_ASAP7_75t_R FILLER_104_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_104 ();
 DECAPx4_ASAP7_75t_R FILLER_104_115 ();
 FILLER_ASAP7_75t_R FILLER_104_125 ();
 DECAPx1_ASAP7_75t_R FILLER_104_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_143 ();
 DECAPx1_ASAP7_75t_R FILLER_104_170 ();
 FILLER_ASAP7_75t_R FILLER_104_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_184 ();
 FILLER_ASAP7_75t_R FILLER_104_191 ();
 DECAPx4_ASAP7_75t_R FILLER_104_201 ();
 DECAPx1_ASAP7_75t_R FILLER_104_225 ();
 DECAPx1_ASAP7_75t_R FILLER_104_235 ();
 DECAPx10_ASAP7_75t_R FILLER_104_251 ();
 DECAPx1_ASAP7_75t_R FILLER_104_273 ();
 FILLER_ASAP7_75t_R FILLER_104_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_285 ();
 DECAPx4_ASAP7_75t_R FILLER_104_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_312 ();
 FILLER_ASAP7_75t_R FILLER_104_335 ();
 FILLER_ASAP7_75t_R FILLER_104_345 ();
 DECAPx4_ASAP7_75t_R FILLER_104_353 ();
 FILLER_ASAP7_75t_R FILLER_104_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_365 ();
 FILLER_ASAP7_75t_R FILLER_104_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_382 ();
 DECAPx6_ASAP7_75t_R FILLER_104_401 ();
 DECAPx4_ASAP7_75t_R FILLER_104_429 ();
 FILLER_ASAP7_75t_R FILLER_104_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_441 ();
 DECAPx1_ASAP7_75t_R FILLER_104_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_474 ();
 DECAPx1_ASAP7_75t_R FILLER_104_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_495 ();
 DECAPx4_ASAP7_75t_R FILLER_104_510 ();
 DECAPx2_ASAP7_75t_R FILLER_104_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_579 ();
 DECAPx2_ASAP7_75t_R FILLER_104_587 ();
 FILLER_ASAP7_75t_R FILLER_104_593 ();
 DECAPx10_ASAP7_75t_R FILLER_104_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_620 ();
 DECAPx4_ASAP7_75t_R FILLER_104_631 ();
 FILLER_ASAP7_75t_R FILLER_104_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_650 ();
 DECAPx1_ASAP7_75t_R FILLER_104_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_661 ();
 DECAPx2_ASAP7_75t_R FILLER_104_668 ();
 FILLER_ASAP7_75t_R FILLER_104_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_676 ();
 DECAPx2_ASAP7_75t_R FILLER_104_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_690 ();
 DECAPx2_ASAP7_75t_R FILLER_104_698 ();
 FILLER_ASAP7_75t_R FILLER_104_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_706 ();
 DECAPx6_ASAP7_75t_R FILLER_104_713 ();
 FILLER_ASAP7_75t_R FILLER_104_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_735 ();
 FILLER_ASAP7_75t_R FILLER_104_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_744 ();
 DECAPx2_ASAP7_75t_R FILLER_104_765 ();
 DECAPx2_ASAP7_75t_R FILLER_104_783 ();
 FILLER_ASAP7_75t_R FILLER_104_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_791 ();
 DECAPx6_ASAP7_75t_R FILLER_104_802 ();
 DECAPx2_ASAP7_75t_R FILLER_104_816 ();
 FILLER_ASAP7_75t_R FILLER_104_834 ();
 DECAPx2_ASAP7_75t_R FILLER_104_848 ();
 FILLER_ASAP7_75t_R FILLER_104_854 ();
 FILLER_ASAP7_75t_R FILLER_104_863 ();
 DECAPx6_ASAP7_75t_R FILLER_104_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_893 ();
 DECAPx2_ASAP7_75t_R FILLER_104_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_913 ();
 FILLER_ASAP7_75t_R FILLER_104_917 ();
 FILLER_ASAP7_75t_R FILLER_104_925 ();
 DECAPx2_ASAP7_75t_R FILLER_104_984 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1042 ();
 FILLER_ASAP7_75t_R FILLER_104_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1059 ();
 FILLER_ASAP7_75t_R FILLER_104_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1067 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1100 ();
 FILLER_ASAP7_75t_R FILLER_104_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1161 ();
 FILLER_ASAP7_75t_R FILLER_104_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1186 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1212 ();
 FILLER_ASAP7_75t_R FILLER_104_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1233 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1280 ();
 DECAPx4_ASAP7_75t_R FILLER_104_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1315 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1352 ();
 FILLER_ASAP7_75t_R FILLER_104_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1363 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1388 ();
 DECAPx1_ASAP7_75t_R FILLER_105_32 ();
 DECAPx2_ASAP7_75t_R FILLER_105_42 ();
 FILLER_ASAP7_75t_R FILLER_105_48 ();
 FILLER_ASAP7_75t_R FILLER_105_56 ();
 DECAPx6_ASAP7_75t_R FILLER_105_90 ();
 DECAPx1_ASAP7_75t_R FILLER_105_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_108 ();
 DECAPx4_ASAP7_75t_R FILLER_105_115 ();
 FILLER_ASAP7_75t_R FILLER_105_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_158 ();
 DECAPx1_ASAP7_75t_R FILLER_105_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_171 ();
 DECAPx2_ASAP7_75t_R FILLER_105_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_192 ();
 DECAPx1_ASAP7_75t_R FILLER_105_207 ();
 DECAPx4_ASAP7_75t_R FILLER_105_217 ();
 FILLER_ASAP7_75t_R FILLER_105_227 ();
 DECAPx1_ASAP7_75t_R FILLER_105_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_239 ();
 DECAPx6_ASAP7_75t_R FILLER_105_254 ();
 DECAPx4_ASAP7_75t_R FILLER_105_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_292 ();
 DECAPx2_ASAP7_75t_R FILLER_105_299 ();
 FILLER_ASAP7_75t_R FILLER_105_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_307 ();
 DECAPx4_ASAP7_75t_R FILLER_105_342 ();
 FILLER_ASAP7_75t_R FILLER_105_352 ();
 DECAPx1_ASAP7_75t_R FILLER_105_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_366 ();
 DECAPx1_ASAP7_75t_R FILLER_105_375 ();
 DECAPx10_ASAP7_75t_R FILLER_105_403 ();
 FILLER_ASAP7_75t_R FILLER_105_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_427 ();
 DECAPx1_ASAP7_75t_R FILLER_105_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_439 ();
 DECAPx1_ASAP7_75t_R FILLER_105_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_460 ();
 DECAPx1_ASAP7_75t_R FILLER_105_475 ();
 DECAPx6_ASAP7_75t_R FILLER_105_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_520 ();
 DECAPx6_ASAP7_75t_R FILLER_105_527 ();
 FILLER_ASAP7_75t_R FILLER_105_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_543 ();
 DECAPx2_ASAP7_75t_R FILLER_105_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_562 ();
 DECAPx4_ASAP7_75t_R FILLER_105_569 ();
 FILLER_ASAP7_75t_R FILLER_105_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_587 ();
 DECAPx2_ASAP7_75t_R FILLER_105_594 ();
 FILLER_ASAP7_75t_R FILLER_105_626 ();
 DECAPx1_ASAP7_75t_R FILLER_105_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_665 ();
 DECAPx1_ASAP7_75t_R FILLER_105_673 ();
 DECAPx10_ASAP7_75t_R FILLER_105_688 ();
 DECAPx6_ASAP7_75t_R FILLER_105_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_724 ();
 DECAPx6_ASAP7_75t_R FILLER_105_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_765 ();
 DECAPx2_ASAP7_75t_R FILLER_105_778 ();
 FILLER_ASAP7_75t_R FILLER_105_784 ();
 DECAPx4_ASAP7_75t_R FILLER_105_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_801 ();
 FILLER_ASAP7_75t_R FILLER_105_827 ();
 DECAPx2_ASAP7_75t_R FILLER_105_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_865 ();
 DECAPx10_ASAP7_75t_R FILLER_105_879 ();
 DECAPx1_ASAP7_75t_R FILLER_105_901 ();
 FILLER_ASAP7_75t_R FILLER_105_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_914 ();
 FILLER_ASAP7_75t_R FILLER_105_922 ();
 DECAPx1_ASAP7_75t_R FILLER_105_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_930 ();
 FILLER_ASAP7_75t_R FILLER_105_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_946 ();
 FILLER_ASAP7_75t_R FILLER_105_954 ();
 DECAPx1_ASAP7_75t_R FILLER_105_962 ();
 DECAPx6_ASAP7_75t_R FILLER_105_972 ();
 DECAPx1_ASAP7_75t_R FILLER_105_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_998 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1017 ();
 FILLER_ASAP7_75t_R FILLER_105_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_105_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_105_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1084 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1101 ();
 FILLER_ASAP7_75t_R FILLER_105_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1116 ();
 FILLER_ASAP7_75t_R FILLER_105_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1128 ();
 DECAPx1_ASAP7_75t_R FILLER_105_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1149 ();
 FILLER_ASAP7_75t_R FILLER_105_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1162 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1197 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1220 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1237 ();
 DECAPx6_ASAP7_75t_R FILLER_105_1250 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1283 ();
 FILLER_ASAP7_75t_R FILLER_105_1290 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1326 ();
 FILLER_ASAP7_75t_R FILLER_105_1336 ();
 FILLER_ASAP7_75t_R FILLER_105_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1346 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1361 ();
 FILLER_ASAP7_75t_R FILLER_105_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1369 ();
 FILLER_ASAP7_75t_R FILLER_106_8 ();
 DECAPx2_ASAP7_75t_R FILLER_106_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_46 ();
 DECAPx1_ASAP7_75t_R FILLER_106_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_77 ();
 DECAPx2_ASAP7_75t_R FILLER_106_81 ();
 DECAPx4_ASAP7_75t_R FILLER_106_133 ();
 DECAPx10_ASAP7_75t_R FILLER_106_146 ();
 DECAPx2_ASAP7_75t_R FILLER_106_168 ();
 FILLER_ASAP7_75t_R FILLER_106_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_182 ();
 DECAPx4_ASAP7_75t_R FILLER_106_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_228 ();
 DECAPx2_ASAP7_75t_R FILLER_106_237 ();
 FILLER_ASAP7_75t_R FILLER_106_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_245 ();
 DECAPx2_ASAP7_75t_R FILLER_106_258 ();
 FILLER_ASAP7_75t_R FILLER_106_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_266 ();
 DECAPx6_ASAP7_75t_R FILLER_106_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_295 ();
 DECAPx4_ASAP7_75t_R FILLER_106_308 ();
 DECAPx6_ASAP7_75t_R FILLER_106_332 ();
 FILLER_ASAP7_75t_R FILLER_106_356 ();
 FILLER_ASAP7_75t_R FILLER_106_366 ();
 FILLER_ASAP7_75t_R FILLER_106_380 ();
 DECAPx2_ASAP7_75t_R FILLER_106_402 ();
 FILLER_ASAP7_75t_R FILLER_106_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_410 ();
 DECAPx4_ASAP7_75t_R FILLER_106_429 ();
 FILLER_ASAP7_75t_R FILLER_106_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_441 ();
 DECAPx1_ASAP7_75t_R FILLER_106_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_483 ();
 DECAPx4_ASAP7_75t_R FILLER_106_490 ();
 FILLER_ASAP7_75t_R FILLER_106_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_502 ();
 DECAPx1_ASAP7_75t_R FILLER_106_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_521 ();
 DECAPx6_ASAP7_75t_R FILLER_106_528 ();
 FILLER_ASAP7_75t_R FILLER_106_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_544 ();
 FILLER_ASAP7_75t_R FILLER_106_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_553 ();
 DECAPx6_ASAP7_75t_R FILLER_106_564 ();
 DECAPx1_ASAP7_75t_R FILLER_106_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_582 ();
 DECAPx2_ASAP7_75t_R FILLER_106_618 ();
 FILLER_ASAP7_75t_R FILLER_106_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_639 ();
 DECAPx4_ASAP7_75t_R FILLER_106_646 ();
 FILLER_ASAP7_75t_R FILLER_106_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_658 ();
 FILLER_ASAP7_75t_R FILLER_106_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_667 ();
 FILLER_ASAP7_75t_R FILLER_106_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_683 ();
 FILLER_ASAP7_75t_R FILLER_106_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_694 ();
 DECAPx1_ASAP7_75t_R FILLER_106_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_732 ();
 DECAPx4_ASAP7_75t_R FILLER_106_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_785 ();
 DECAPx1_ASAP7_75t_R FILLER_106_797 ();
 DECAPx1_ASAP7_75t_R FILLER_106_818 ();
 FILLER_ASAP7_75t_R FILLER_106_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_843 ();
 DECAPx2_ASAP7_75t_R FILLER_106_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_873 ();
 FILLER_ASAP7_75t_R FILLER_106_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_896 ();
 DECAPx2_ASAP7_75t_R FILLER_106_948 ();
 FILLER_ASAP7_75t_R FILLER_106_960 ();
 DECAPx10_ASAP7_75t_R FILLER_106_974 ();
 FILLER_ASAP7_75t_R FILLER_106_996 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1023 ();
 DECAPx6_ASAP7_75t_R FILLER_106_1030 ();
 FILLER_ASAP7_75t_R FILLER_106_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1148 ();
 DECAPx4_ASAP7_75t_R FILLER_106_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1258 ();
 DECAPx6_ASAP7_75t_R FILLER_106_1280 ();
 FILLER_ASAP7_75t_R FILLER_106_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1296 ();
 FILLER_ASAP7_75t_R FILLER_106_1317 ();
 FILLER_ASAP7_75t_R FILLER_106_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1337 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1348 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1354 ();
 FILLER_ASAP7_75t_R FILLER_106_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1388 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_14 ();
 DECAPx2_ASAP7_75t_R FILLER_107_33 ();
 FILLER_ASAP7_75t_R FILLER_107_39 ();
 DECAPx2_ASAP7_75t_R FILLER_107_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_60 ();
 DECAPx2_ASAP7_75t_R FILLER_107_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_70 ();
 DECAPx4_ASAP7_75t_R FILLER_107_75 ();
 FILLER_ASAP7_75t_R FILLER_107_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_87 ();
 DECAPx2_ASAP7_75t_R FILLER_107_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_103 ();
 DECAPx4_ASAP7_75t_R FILLER_107_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_179 ();
 DECAPx1_ASAP7_75t_R FILLER_107_188 ();
 DECAPx2_ASAP7_75t_R FILLER_107_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_204 ();
 DECAPx10_ASAP7_75t_R FILLER_107_225 ();
 FILLER_ASAP7_75t_R FILLER_107_255 ();
 DECAPx1_ASAP7_75t_R FILLER_107_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_287 ();
 DECAPx2_ASAP7_75t_R FILLER_107_312 ();
 DECAPx6_ASAP7_75t_R FILLER_107_326 ();
 DECAPx2_ASAP7_75t_R FILLER_107_340 ();
 DECAPx1_ASAP7_75t_R FILLER_107_352 ();
 DECAPx6_ASAP7_75t_R FILLER_107_375 ();
 DECAPx1_ASAP7_75t_R FILLER_107_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_393 ();
 DECAPx6_ASAP7_75t_R FILLER_107_400 ();
 FILLER_ASAP7_75t_R FILLER_107_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_416 ();
 FILLER_ASAP7_75t_R FILLER_107_441 ();
 DECAPx6_ASAP7_75t_R FILLER_107_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_477 ();
 DECAPx10_ASAP7_75t_R FILLER_107_484 ();
 DECAPx1_ASAP7_75t_R FILLER_107_506 ();
 DECAPx1_ASAP7_75t_R FILLER_107_518 ();
 DECAPx10_ASAP7_75t_R FILLER_107_538 ();
 FILLER_ASAP7_75t_R FILLER_107_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_562 ();
 DECAPx2_ASAP7_75t_R FILLER_107_570 ();
 FILLER_ASAP7_75t_R FILLER_107_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_578 ();
 DECAPx1_ASAP7_75t_R FILLER_107_582 ();
 DECAPx2_ASAP7_75t_R FILLER_107_592 ();
 FILLER_ASAP7_75t_R FILLER_107_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_603 ();
 DECAPx6_ASAP7_75t_R FILLER_107_610 ();
 DECAPx1_ASAP7_75t_R FILLER_107_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_628 ();
 DECAPx6_ASAP7_75t_R FILLER_107_635 ();
 DECAPx2_ASAP7_75t_R FILLER_107_656 ();
 FILLER_ASAP7_75t_R FILLER_107_662 ();
 FILLER_ASAP7_75t_R FILLER_107_676 ();
 DECAPx4_ASAP7_75t_R FILLER_107_684 ();
 FILLER_ASAP7_75t_R FILLER_107_694 ();
 FILLER_ASAP7_75t_R FILLER_107_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_711 ();
 DECAPx2_ASAP7_75t_R FILLER_107_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_730 ();
 DECAPx6_ASAP7_75t_R FILLER_107_737 ();
 DECAPx1_ASAP7_75t_R FILLER_107_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_755 ();
 FILLER_ASAP7_75t_R FILLER_107_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_787 ();
 DECAPx1_ASAP7_75t_R FILLER_107_813 ();
 DECAPx1_ASAP7_75t_R FILLER_107_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_827 ();
 DECAPx2_ASAP7_75t_R FILLER_107_834 ();
 FILLER_ASAP7_75t_R FILLER_107_849 ();
 DECAPx2_ASAP7_75t_R FILLER_107_861 ();
 FILLER_ASAP7_75t_R FILLER_107_867 ();
 DECAPx1_ASAP7_75t_R FILLER_107_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_894 ();
 FILLER_ASAP7_75t_R FILLER_107_910 ();
 FILLER_ASAP7_75t_R FILLER_107_926 ();
 FILLER_ASAP7_75t_R FILLER_107_962 ();
 DECAPx4_ASAP7_75t_R FILLER_107_981 ();
 FILLER_ASAP7_75t_R FILLER_107_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1038 ();
 FILLER_ASAP7_75t_R FILLER_107_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1062 ();
 FILLER_ASAP7_75t_R FILLER_107_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_107_1085 ();
 FILLER_ASAP7_75t_R FILLER_107_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_107_1116 ();
 FILLER_ASAP7_75t_R FILLER_107_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_107_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1148 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1155 ();
 FILLER_ASAP7_75t_R FILLER_107_1169 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_107_1191 ();
 FILLER_ASAP7_75t_R FILLER_107_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1234 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1260 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1280 ();
 FILLER_ASAP7_75t_R FILLER_107_1294 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1303 ();
 FILLER_ASAP7_75t_R FILLER_107_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1333 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1347 ();
 FILLER_ASAP7_75t_R FILLER_107_1353 ();
 DECAPx1_ASAP7_75t_R FILLER_107_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_8 ();
 FILLER_ASAP7_75t_R FILLER_108_21 ();
 FILLER_ASAP7_75t_R FILLER_108_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_29 ();
 DECAPx4_ASAP7_75t_R FILLER_108_60 ();
 DECAPx1_ASAP7_75t_R FILLER_108_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_84 ();
 FILLER_ASAP7_75t_R FILLER_108_115 ();
 DECAPx6_ASAP7_75t_R FILLER_108_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_177 ();
 FILLER_ASAP7_75t_R FILLER_108_192 ();
 FILLER_ASAP7_75t_R FILLER_108_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_210 ();
 DECAPx2_ASAP7_75t_R FILLER_108_225 ();
 FILLER_ASAP7_75t_R FILLER_108_231 ();
 DECAPx2_ASAP7_75t_R FILLER_108_241 ();
 FILLER_ASAP7_75t_R FILLER_108_247 ();
 FILLER_ASAP7_75t_R FILLER_108_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_265 ();
 DECAPx6_ASAP7_75t_R FILLER_108_278 ();
 FILLER_ASAP7_75t_R FILLER_108_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_294 ();
 DECAPx6_ASAP7_75t_R FILLER_108_315 ();
 DECAPx4_ASAP7_75t_R FILLER_108_345 ();
 FILLER_ASAP7_75t_R FILLER_108_355 ();
 DECAPx1_ASAP7_75t_R FILLER_108_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_367 ();
 DECAPx6_ASAP7_75t_R FILLER_108_374 ();
 FILLER_ASAP7_75t_R FILLER_108_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_427 ();
 DECAPx10_ASAP7_75t_R FILLER_108_438 ();
 FILLER_ASAP7_75t_R FILLER_108_460 ();
 DECAPx4_ASAP7_75t_R FILLER_108_464 ();
 FILLER_ASAP7_75t_R FILLER_108_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_476 ();
 DECAPx2_ASAP7_75t_R FILLER_108_485 ();
 DECAPx4_ASAP7_75t_R FILLER_108_507 ();
 DECAPx2_ASAP7_75t_R FILLER_108_531 ();
 FILLER_ASAP7_75t_R FILLER_108_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_564 ();
 DECAPx4_ASAP7_75t_R FILLER_108_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_601 ();
 DECAPx10_ASAP7_75t_R FILLER_108_608 ();
 FILLER_ASAP7_75t_R FILLER_108_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_642 ();
 FILLER_ASAP7_75t_R FILLER_108_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_655 ();
 FILLER_ASAP7_75t_R FILLER_108_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_670 ();
 DECAPx2_ASAP7_75t_R FILLER_108_687 ();
 FILLER_ASAP7_75t_R FILLER_108_693 ();
 FILLER_ASAP7_75t_R FILLER_108_709 ();
 DECAPx4_ASAP7_75t_R FILLER_108_719 ();
 FILLER_ASAP7_75t_R FILLER_108_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_731 ();
 FILLER_ASAP7_75t_R FILLER_108_739 ();
 DECAPx1_ASAP7_75t_R FILLER_108_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_757 ();
 DECAPx2_ASAP7_75t_R FILLER_108_764 ();
 FILLER_ASAP7_75t_R FILLER_108_770 ();
 DECAPx4_ASAP7_75t_R FILLER_108_782 ();
 FILLER_ASAP7_75t_R FILLER_108_792 ();
 DECAPx4_ASAP7_75t_R FILLER_108_804 ();
 DECAPx4_ASAP7_75t_R FILLER_108_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_851 ();
 DECAPx4_ASAP7_75t_R FILLER_108_865 ();
 FILLER_ASAP7_75t_R FILLER_108_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_877 ();
 FILLER_ASAP7_75t_R FILLER_108_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_940 ();
 DECAPx2_ASAP7_75t_R FILLER_108_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_970 ();
 DECAPx2_ASAP7_75t_R FILLER_108_982 ();
 FILLER_ASAP7_75t_R FILLER_108_988 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1141 ();
 FILLER_ASAP7_75t_R FILLER_108_1147 ();
 FILLER_ASAP7_75t_R FILLER_108_1157 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1169 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1185 ();
 FILLER_ASAP7_75t_R FILLER_108_1199 ();
 FILLER_ASAP7_75t_R FILLER_108_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1282 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1296 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1308 ();
 FILLER_ASAP7_75t_R FILLER_108_1318 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1326 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1332 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1388 ();
 DECAPx1_ASAP7_75t_R FILLER_109_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_12 ();
 DECAPx1_ASAP7_75t_R FILLER_109_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_35 ();
 FILLER_ASAP7_75t_R FILLER_109_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_44 ();
 DECAPx4_ASAP7_75t_R FILLER_109_48 ();
 FILLER_ASAP7_75t_R FILLER_109_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_97 ();
 DECAPx1_ASAP7_75t_R FILLER_109_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_128 ();
 DECAPx2_ASAP7_75t_R FILLER_109_135 ();
 FILLER_ASAP7_75t_R FILLER_109_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_143 ();
 DECAPx2_ASAP7_75t_R FILLER_109_147 ();
 FILLER_ASAP7_75t_R FILLER_109_153 ();
 DECAPx2_ASAP7_75t_R FILLER_109_168 ();
 FILLER_ASAP7_75t_R FILLER_109_174 ();
 DECAPx4_ASAP7_75t_R FILLER_109_182 ();
 FILLER_ASAP7_75t_R FILLER_109_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_217 ();
 FILLER_ASAP7_75t_R FILLER_109_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_226 ();
 FILLER_ASAP7_75t_R FILLER_109_247 ();
 FILLER_ASAP7_75t_R FILLER_109_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_265 ();
 DECAPx1_ASAP7_75t_R FILLER_109_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_289 ();
 DECAPx1_ASAP7_75t_R FILLER_109_298 ();
 DECAPx10_ASAP7_75t_R FILLER_109_308 ();
 FILLER_ASAP7_75t_R FILLER_109_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_332 ();
 DECAPx6_ASAP7_75t_R FILLER_109_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_361 ();
 DECAPx10_ASAP7_75t_R FILLER_109_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_390 ();
 DECAPx4_ASAP7_75t_R FILLER_109_409 ();
 FILLER_ASAP7_75t_R FILLER_109_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_451 ();
 DECAPx2_ASAP7_75t_R FILLER_109_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_465 ();
 DECAPx1_ASAP7_75t_R FILLER_109_484 ();
 DECAPx1_ASAP7_75t_R FILLER_109_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_499 ();
 DECAPx2_ASAP7_75t_R FILLER_109_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_522 ();
 FILLER_ASAP7_75t_R FILLER_109_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_553 ();
 DECAPx2_ASAP7_75t_R FILLER_109_573 ();
 FILLER_ASAP7_75t_R FILLER_109_579 ();
 DECAPx6_ASAP7_75t_R FILLER_109_655 ();
 FILLER_ASAP7_75t_R FILLER_109_669 ();
 DECAPx1_ASAP7_75t_R FILLER_109_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_709 ();
 DECAPx4_ASAP7_75t_R FILLER_109_713 ();
 DECAPx4_ASAP7_75t_R FILLER_109_752 ();
 FILLER_ASAP7_75t_R FILLER_109_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_764 ();
 DECAPx6_ASAP7_75t_R FILLER_109_777 ();
 DECAPx1_ASAP7_75t_R FILLER_109_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_795 ();
 DECAPx1_ASAP7_75t_R FILLER_109_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_812 ();
 DECAPx4_ASAP7_75t_R FILLER_109_821 ();
 FILLER_ASAP7_75t_R FILLER_109_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_833 ();
 FILLER_ASAP7_75t_R FILLER_109_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_850 ();
 DECAPx4_ASAP7_75t_R FILLER_109_863 ();
 DECAPx2_ASAP7_75t_R FILLER_109_888 ();
 FILLER_ASAP7_75t_R FILLER_109_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_896 ();
 DECAPx1_ASAP7_75t_R FILLER_109_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_908 ();
 FILLER_ASAP7_75t_R FILLER_109_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_932 ();
 DECAPx2_ASAP7_75t_R FILLER_109_940 ();
 FILLER_ASAP7_75t_R FILLER_109_946 ();
 DECAPx4_ASAP7_75t_R FILLER_109_954 ();
 DECAPx1_ASAP7_75t_R FILLER_109_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_974 ();
 DECAPx2_ASAP7_75t_R FILLER_109_989 ();
 FILLER_ASAP7_75t_R FILLER_109_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_997 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1144 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1215 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1237 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1317 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1335 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1360 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1372 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1386 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_28 ();
 DECAPx1_ASAP7_75t_R FILLER_110_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_39 ();
 DECAPx2_ASAP7_75t_R FILLER_110_44 ();
 FILLER_ASAP7_75t_R FILLER_110_50 ();
 DECAPx2_ASAP7_75t_R FILLER_110_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_67 ();
 DECAPx10_ASAP7_75t_R FILLER_110_74 ();
 DECAPx1_ASAP7_75t_R FILLER_110_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_100 ();
 FILLER_ASAP7_75t_R FILLER_110_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_118 ();
 DECAPx10_ASAP7_75t_R FILLER_110_145 ();
 DECAPx10_ASAP7_75t_R FILLER_110_167 ();
 FILLER_ASAP7_75t_R FILLER_110_189 ();
 DECAPx4_ASAP7_75t_R FILLER_110_197 ();
 FILLER_ASAP7_75t_R FILLER_110_213 ();
 DECAPx6_ASAP7_75t_R FILLER_110_221 ();
 FILLER_ASAP7_75t_R FILLER_110_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_250 ();
 DECAPx2_ASAP7_75t_R FILLER_110_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_272 ();
 DECAPx6_ASAP7_75t_R FILLER_110_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_301 ();
 DECAPx1_ASAP7_75t_R FILLER_110_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_314 ();
 DECAPx1_ASAP7_75t_R FILLER_110_327 ();
 DECAPx1_ASAP7_75t_R FILLER_110_345 ();
 FILLER_ASAP7_75t_R FILLER_110_355 ();
 DECAPx4_ASAP7_75t_R FILLER_110_371 ();
 DECAPx10_ASAP7_75t_R FILLER_110_388 ();
 DECAPx4_ASAP7_75t_R FILLER_110_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_427 ();
 DECAPx2_ASAP7_75t_R FILLER_110_435 ();
 DECAPx4_ASAP7_75t_R FILLER_110_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_464 ();
 FILLER_ASAP7_75t_R FILLER_110_483 ();
 DECAPx10_ASAP7_75t_R FILLER_110_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_533 ();
 DECAPx4_ASAP7_75t_R FILLER_110_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_558 ();
 DECAPx2_ASAP7_75t_R FILLER_110_620 ();
 FILLER_ASAP7_75t_R FILLER_110_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_628 ();
 FILLER_ASAP7_75t_R FILLER_110_636 ();
 DECAPx2_ASAP7_75t_R FILLER_110_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_647 ();
 FILLER_ASAP7_75t_R FILLER_110_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_656 ();
 DECAPx1_ASAP7_75t_R FILLER_110_669 ();
 DECAPx4_ASAP7_75t_R FILLER_110_691 ();
 FILLER_ASAP7_75t_R FILLER_110_701 ();
 DECAPx2_ASAP7_75t_R FILLER_110_709 ();
 DECAPx10_ASAP7_75t_R FILLER_110_729 ();
 DECAPx6_ASAP7_75t_R FILLER_110_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_765 ();
 DECAPx1_ASAP7_75t_R FILLER_110_773 ();
 DECAPx10_ASAP7_75t_R FILLER_110_783 ();
 DECAPx2_ASAP7_75t_R FILLER_110_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_811 ();
 DECAPx1_ASAP7_75t_R FILLER_110_835 ();
 DECAPx4_ASAP7_75t_R FILLER_110_862 ();
 FILLER_ASAP7_75t_R FILLER_110_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_882 ();
 DECAPx1_ASAP7_75t_R FILLER_110_923 ();
 FILLER_ASAP7_75t_R FILLER_110_941 ();
 FILLER_ASAP7_75t_R FILLER_110_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_957 ();
 DECAPx2_ASAP7_75t_R FILLER_110_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_974 ();
 FILLER_ASAP7_75t_R FILLER_110_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_993 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1034 ();
 FILLER_ASAP7_75t_R FILLER_110_1040 ();
 FILLER_ASAP7_75t_R FILLER_110_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1131 ();
 FILLER_ASAP7_75t_R FILLER_110_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1200 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1211 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1228 ();
 FILLER_ASAP7_75t_R FILLER_110_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1246 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1324 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1336 ();
 FILLER_ASAP7_75t_R FILLER_110_1346 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1348 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1355 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1376 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_111_99 ();
 DECAPx1_ASAP7_75t_R FILLER_111_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_129 ();
 DECAPx2_ASAP7_75t_R FILLER_111_139 ();
 FILLER_ASAP7_75t_R FILLER_111_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_174 ();
 DECAPx1_ASAP7_75t_R FILLER_111_178 ();
 DECAPx4_ASAP7_75t_R FILLER_111_198 ();
 FILLER_ASAP7_75t_R FILLER_111_208 ();
 DECAPx10_ASAP7_75t_R FILLER_111_230 ();
 FILLER_ASAP7_75t_R FILLER_111_252 ();
 DECAPx2_ASAP7_75t_R FILLER_111_264 ();
 FILLER_ASAP7_75t_R FILLER_111_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_272 ();
 FILLER_ASAP7_75t_R FILLER_111_287 ();
 DECAPx6_ASAP7_75t_R FILLER_111_297 ();
 DECAPx1_ASAP7_75t_R FILLER_111_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_324 ();
 DECAPx1_ASAP7_75t_R FILLER_111_333 ();
 DECAPx1_ASAP7_75t_R FILLER_111_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_361 ();
 FILLER_ASAP7_75t_R FILLER_111_376 ();
 DECAPx2_ASAP7_75t_R FILLER_111_386 ();
 DECAPx4_ASAP7_75t_R FILLER_111_398 ();
 FILLER_ASAP7_75t_R FILLER_111_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_428 ();
 DECAPx1_ASAP7_75t_R FILLER_111_435 ();
 DECAPx4_ASAP7_75t_R FILLER_111_449 ();
 FILLER_ASAP7_75t_R FILLER_111_459 ();
 DECAPx2_ASAP7_75t_R FILLER_111_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_479 ();
 DECAPx2_ASAP7_75t_R FILLER_111_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_493 ();
 DECAPx4_ASAP7_75t_R FILLER_111_512 ();
 FILLER_ASAP7_75t_R FILLER_111_522 ();
 DECAPx4_ASAP7_75t_R FILLER_111_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_541 ();
 DECAPx4_ASAP7_75t_R FILLER_111_548 ();
 FILLER_ASAP7_75t_R FILLER_111_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_560 ();
 DECAPx2_ASAP7_75t_R FILLER_111_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_573 ();
 DECAPx2_ASAP7_75t_R FILLER_111_577 ();
 FILLER_ASAP7_75t_R FILLER_111_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_585 ();
 DECAPx2_ASAP7_75t_R FILLER_111_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_598 ();
 DECAPx4_ASAP7_75t_R FILLER_111_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_612 ();
 DECAPx2_ASAP7_75t_R FILLER_111_635 ();
 FILLER_ASAP7_75t_R FILLER_111_641 ();
 DECAPx4_ASAP7_75t_R FILLER_111_650 ();
 DECAPx2_ASAP7_75t_R FILLER_111_667 ();
 FILLER_ASAP7_75t_R FILLER_111_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_678 ();
 DECAPx6_ASAP7_75t_R FILLER_111_686 ();
 FILLER_ASAP7_75t_R FILLER_111_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_708 ();
 DECAPx2_ASAP7_75t_R FILLER_111_736 ();
 FILLER_ASAP7_75t_R FILLER_111_742 ();
 FILLER_ASAP7_75t_R FILLER_111_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_759 ();
 DECAPx2_ASAP7_75t_R FILLER_111_768 ();
 FILLER_ASAP7_75t_R FILLER_111_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_776 ();
 DECAPx6_ASAP7_75t_R FILLER_111_794 ();
 DECAPx1_ASAP7_75t_R FILLER_111_808 ();
 DECAPx2_ASAP7_75t_R FILLER_111_819 ();
 FILLER_ASAP7_75t_R FILLER_111_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_827 ();
 FILLER_ASAP7_75t_R FILLER_111_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_847 ();
 DECAPx2_ASAP7_75t_R FILLER_111_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_889 ();
 DECAPx1_ASAP7_75t_R FILLER_111_906 ();
 FILLER_ASAP7_75t_R FILLER_111_916 ();
 FILLER_ASAP7_75t_R FILLER_111_941 ();
 DECAPx4_ASAP7_75t_R FILLER_111_962 ();
 DECAPx10_ASAP7_75t_R FILLER_111_980 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1054 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1095 ();
 FILLER_ASAP7_75t_R FILLER_111_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1131 ();
 FILLER_ASAP7_75t_R FILLER_111_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1154 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1171 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1189 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1208 ();
 FILLER_ASAP7_75t_R FILLER_111_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1246 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1278 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1304 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1312 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1319 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1335 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1369 ();
 DECAPx1_ASAP7_75t_R FILLER_112_8 ();
 DECAPx1_ASAP7_75t_R FILLER_112_18 ();
 DECAPx4_ASAP7_75t_R FILLER_112_37 ();
 FILLER_ASAP7_75t_R FILLER_112_47 ();
 DECAPx4_ASAP7_75t_R FILLER_112_55 ();
 DECAPx2_ASAP7_75t_R FILLER_112_75 ();
 FILLER_ASAP7_75t_R FILLER_112_81 ();
 DECAPx1_ASAP7_75t_R FILLER_112_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_90 ();
 DECAPx2_ASAP7_75t_R FILLER_112_97 ();
 FILLER_ASAP7_75t_R FILLER_112_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_105 ();
 DECAPx6_ASAP7_75t_R FILLER_112_116 ();
 FILLER_ASAP7_75t_R FILLER_112_130 ();
 FILLER_ASAP7_75t_R FILLER_112_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_160 ();
 DECAPx1_ASAP7_75t_R FILLER_112_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_198 ();
 DECAPx4_ASAP7_75t_R FILLER_112_207 ();
 FILLER_ASAP7_75t_R FILLER_112_217 ();
 DECAPx6_ASAP7_75t_R FILLER_112_227 ();
 FILLER_ASAP7_75t_R FILLER_112_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_243 ();
 DECAPx4_ASAP7_75t_R FILLER_112_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_274 ();
 FILLER_ASAP7_75t_R FILLER_112_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_285 ();
 DECAPx2_ASAP7_75t_R FILLER_112_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_306 ();
 FILLER_ASAP7_75t_R FILLER_112_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_323 ();
 DECAPx1_ASAP7_75t_R FILLER_112_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_342 ();
 DECAPx1_ASAP7_75t_R FILLER_112_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_377 ();
 DECAPx4_ASAP7_75t_R FILLER_112_397 ();
 FILLER_ASAP7_75t_R FILLER_112_407 ();
 DECAPx1_ASAP7_75t_R FILLER_112_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_431 ();
 DECAPx1_ASAP7_75t_R FILLER_112_440 ();
 FILLER_ASAP7_75t_R FILLER_112_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_466 ();
 DECAPx10_ASAP7_75t_R FILLER_112_477 ();
 DECAPx1_ASAP7_75t_R FILLER_112_502 ();
 FILLER_ASAP7_75t_R FILLER_112_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_529 ();
 DECAPx2_ASAP7_75t_R FILLER_112_538 ();
 FILLER_ASAP7_75t_R FILLER_112_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_546 ();
 DECAPx6_ASAP7_75t_R FILLER_112_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_567 ();
 DECAPx4_ASAP7_75t_R FILLER_112_575 ();
 FILLER_ASAP7_75t_R FILLER_112_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_613 ();
 DECAPx6_ASAP7_75t_R FILLER_112_624 ();
 DECAPx1_ASAP7_75t_R FILLER_112_638 ();
 DECAPx2_ASAP7_75t_R FILLER_112_648 ();
 FILLER_ASAP7_75t_R FILLER_112_654 ();
 DECAPx4_ASAP7_75t_R FILLER_112_668 ();
 DECAPx2_ASAP7_75t_R FILLER_112_685 ();
 FILLER_ASAP7_75t_R FILLER_112_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_693 ();
 DECAPx1_ASAP7_75t_R FILLER_112_713 ();
 FILLER_ASAP7_75t_R FILLER_112_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_749 ();
 FILLER_ASAP7_75t_R FILLER_112_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_776 ();
 DECAPx1_ASAP7_75t_R FILLER_112_832 ();
 FILLER_ASAP7_75t_R FILLER_112_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_858 ();
 DECAPx1_ASAP7_75t_R FILLER_112_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_886 ();
 FILLER_ASAP7_75t_R FILLER_112_896 ();
 DECAPx2_ASAP7_75t_R FILLER_112_904 ();
 DECAPx1_ASAP7_75t_R FILLER_112_917 ();
 DECAPx1_ASAP7_75t_R FILLER_112_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_950 ();
 FILLER_ASAP7_75t_R FILLER_112_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_960 ();
 DECAPx2_ASAP7_75t_R FILLER_112_971 ();
 FILLER_ASAP7_75t_R FILLER_112_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_989 ();
 DECAPx6_ASAP7_75t_R FILLER_112_997 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1037 ();
 FILLER_ASAP7_75t_R FILLER_112_1046 ();
 FILLER_ASAP7_75t_R FILLER_112_1055 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1077 ();
 FILLER_ASAP7_75t_R FILLER_112_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1102 ();
 FILLER_ASAP7_75t_R FILLER_112_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1176 ();
 FILLER_ASAP7_75t_R FILLER_112_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1184 ();
 FILLER_ASAP7_75t_R FILLER_112_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1214 ();
 FILLER_ASAP7_75t_R FILLER_112_1230 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1300 ();
 DECAPx4_ASAP7_75t_R FILLER_112_1307 ();
 FILLER_ASAP7_75t_R FILLER_112_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1319 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1347 ();
 FILLER_ASAP7_75t_R FILLER_112_1353 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1370 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_113_32 ();
 FILLER_ASAP7_75t_R FILLER_113_46 ();
 DECAPx1_ASAP7_75t_R FILLER_113_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_64 ();
 DECAPx2_ASAP7_75t_R FILLER_113_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_78 ();
 DECAPx2_ASAP7_75t_R FILLER_113_137 ();
 FILLER_ASAP7_75t_R FILLER_113_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_161 ();
 DECAPx2_ASAP7_75t_R FILLER_113_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_183 ();
 DECAPx1_ASAP7_75t_R FILLER_113_190 ();
 DECAPx1_ASAP7_75t_R FILLER_113_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_218 ();
 DECAPx10_ASAP7_75t_R FILLER_113_245 ();
 DECAPx4_ASAP7_75t_R FILLER_113_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_283 ();
 DECAPx4_ASAP7_75t_R FILLER_113_296 ();
 FILLER_ASAP7_75t_R FILLER_113_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_308 ();
 DECAPx1_ASAP7_75t_R FILLER_113_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_319 ();
 DECAPx2_ASAP7_75t_R FILLER_113_326 ();
 FILLER_ASAP7_75t_R FILLER_113_332 ();
 DECAPx2_ASAP7_75t_R FILLER_113_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_367 ();
 FILLER_ASAP7_75t_R FILLER_113_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_376 ();
 FILLER_ASAP7_75t_R FILLER_113_385 ();
 DECAPx1_ASAP7_75t_R FILLER_113_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_407 ();
 FILLER_ASAP7_75t_R FILLER_113_421 ();
 DECAPx1_ASAP7_75t_R FILLER_113_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_446 ();
 DECAPx1_ASAP7_75t_R FILLER_113_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_469 ();
 DECAPx1_ASAP7_75t_R FILLER_113_480 ();
 DECAPx6_ASAP7_75t_R FILLER_113_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_508 ();
 DECAPx1_ASAP7_75t_R FILLER_113_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_521 ();
 FILLER_ASAP7_75t_R FILLER_113_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_544 ();
 FILLER_ASAP7_75t_R FILLER_113_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_573 ();
 DECAPx2_ASAP7_75t_R FILLER_113_580 ();
 DECAPx2_ASAP7_75t_R FILLER_113_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_598 ();
 DECAPx10_ASAP7_75t_R FILLER_113_602 ();
 DECAPx2_ASAP7_75t_R FILLER_113_624 ();
 DECAPx2_ASAP7_75t_R FILLER_113_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_646 ();
 FILLER_ASAP7_75t_R FILLER_113_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_659 ();
 DECAPx2_ASAP7_75t_R FILLER_113_666 ();
 DECAPx4_ASAP7_75t_R FILLER_113_684 ();
 FILLER_ASAP7_75t_R FILLER_113_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_696 ();
 DECAPx2_ASAP7_75t_R FILLER_113_703 ();
 FILLER_ASAP7_75t_R FILLER_113_709 ();
 DECAPx6_ASAP7_75t_R FILLER_113_731 ();
 DECAPx6_ASAP7_75t_R FILLER_113_760 ();
 DECAPx6_ASAP7_75t_R FILLER_113_793 ();
 DECAPx1_ASAP7_75t_R FILLER_113_807 ();
 DECAPx2_ASAP7_75t_R FILLER_113_825 ();
 DECAPx2_ASAP7_75t_R FILLER_113_837 ();
 DECAPx6_ASAP7_75t_R FILLER_113_850 ();
 FILLER_ASAP7_75t_R FILLER_113_864 ();
 DECAPx2_ASAP7_75t_R FILLER_113_874 ();
 DECAPx2_ASAP7_75t_R FILLER_113_886 ();
 DECAPx1_ASAP7_75t_R FILLER_113_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_923 ();
 DECAPx10_ASAP7_75t_R FILLER_113_926 ();
 DECAPx4_ASAP7_75t_R FILLER_113_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_958 ();
 DECAPx1_ASAP7_75t_R FILLER_113_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_973 ();
 FILLER_ASAP7_75t_R FILLER_113_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_983 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1022 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1029 ();
 FILLER_ASAP7_75t_R FILLER_113_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1160 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1201 ();
 FILLER_ASAP7_75t_R FILLER_113_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1209 ();
 FILLER_ASAP7_75t_R FILLER_113_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1219 ();
 FILLER_ASAP7_75t_R FILLER_113_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1233 ();
 FILLER_ASAP7_75t_R FILLER_113_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1300 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1313 ();
 FILLER_ASAP7_75t_R FILLER_113_1327 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1341 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1371 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1380 ();
 FILLER_ASAP7_75t_R FILLER_113_1390 ();
 DECAPx1_ASAP7_75t_R FILLER_114_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_6 ();
 FILLER_ASAP7_75t_R FILLER_114_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_41 ();
 DECAPx1_ASAP7_75t_R FILLER_114_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_49 ();
 DECAPx1_ASAP7_75t_R FILLER_114_76 ();
 FILLER_ASAP7_75t_R FILLER_114_84 ();
 DECAPx2_ASAP7_75t_R FILLER_114_92 ();
 DECAPx1_ASAP7_75t_R FILLER_114_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_105 ();
 DECAPx2_ASAP7_75t_R FILLER_114_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_118 ();
 DECAPx2_ASAP7_75t_R FILLER_114_122 ();
 DECAPx10_ASAP7_75t_R FILLER_114_134 ();
 DECAPx6_ASAP7_75t_R FILLER_114_156 ();
 FILLER_ASAP7_75t_R FILLER_114_170 ();
 FILLER_ASAP7_75t_R FILLER_114_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_178 ();
 DECAPx4_ASAP7_75t_R FILLER_114_185 ();
 FILLER_ASAP7_75t_R FILLER_114_195 ();
 FILLER_ASAP7_75t_R FILLER_114_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_219 ();
 DECAPx10_ASAP7_75t_R FILLER_114_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_250 ();
 DECAPx2_ASAP7_75t_R FILLER_114_257 ();
 DECAPx10_ASAP7_75t_R FILLER_114_275 ();
 DECAPx1_ASAP7_75t_R FILLER_114_304 ();
 DECAPx2_ASAP7_75t_R FILLER_114_316 ();
 FILLER_ASAP7_75t_R FILLER_114_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_324 ();
 DECAPx10_ASAP7_75t_R FILLER_114_337 ();
 DECAPx2_ASAP7_75t_R FILLER_114_359 ();
 FILLER_ASAP7_75t_R FILLER_114_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_373 ();
 FILLER_ASAP7_75t_R FILLER_114_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_390 ();
 DECAPx4_ASAP7_75t_R FILLER_114_403 ();
 FILLER_ASAP7_75t_R FILLER_114_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_415 ();
 DECAPx4_ASAP7_75t_R FILLER_114_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_434 ();
 DECAPx6_ASAP7_75t_R FILLER_114_443 ();
 DECAPx1_ASAP7_75t_R FILLER_114_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_461 ();
 DECAPx2_ASAP7_75t_R FILLER_114_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_470 ();
 FILLER_ASAP7_75t_R FILLER_114_489 ();
 DECAPx2_ASAP7_75t_R FILLER_114_523 ();
 FILLER_ASAP7_75t_R FILLER_114_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_531 ();
 FILLER_ASAP7_75t_R FILLER_114_540 ();
 FILLER_ASAP7_75t_R FILLER_114_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_552 ();
 DECAPx1_ASAP7_75t_R FILLER_114_569 ();
 DECAPx10_ASAP7_75t_R FILLER_114_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_621 ();
 FILLER_ASAP7_75t_R FILLER_114_645 ();
 DECAPx4_ASAP7_75t_R FILLER_114_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_677 ();
 DECAPx2_ASAP7_75t_R FILLER_114_688 ();
 FILLER_ASAP7_75t_R FILLER_114_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_722 ();
 DECAPx6_ASAP7_75t_R FILLER_114_729 ();
 FILLER_ASAP7_75t_R FILLER_114_743 ();
 DECAPx6_ASAP7_75t_R FILLER_114_757 ();
 DECAPx1_ASAP7_75t_R FILLER_114_771 ();
 DECAPx2_ASAP7_75t_R FILLER_114_789 ();
 FILLER_ASAP7_75t_R FILLER_114_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_797 ();
 DECAPx2_ASAP7_75t_R FILLER_114_804 ();
 FILLER_ASAP7_75t_R FILLER_114_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_812 ();
 DECAPx1_ASAP7_75t_R FILLER_114_819 ();
 DECAPx10_ASAP7_75t_R FILLER_114_829 ();
 DECAPx6_ASAP7_75t_R FILLER_114_851 ();
 FILLER_ASAP7_75t_R FILLER_114_879 ();
 DECAPx1_ASAP7_75t_R FILLER_114_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_892 ();
 DECAPx4_ASAP7_75t_R FILLER_114_899 ();
 FILLER_ASAP7_75t_R FILLER_114_909 ();
 FILLER_ASAP7_75t_R FILLER_114_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_919 ();
 DECAPx6_ASAP7_75t_R FILLER_114_926 ();
 FILLER_ASAP7_75t_R FILLER_114_946 ();
 DECAPx10_ASAP7_75t_R FILLER_114_956 ();
 DECAPx6_ASAP7_75t_R FILLER_114_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1019 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1061 ();
 FILLER_ASAP7_75t_R FILLER_114_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1083 ();
 FILLER_ASAP7_75t_R FILLER_114_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1105 ();
 FILLER_ASAP7_75t_R FILLER_114_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1132 ();
 FILLER_ASAP7_75t_R FILLER_114_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1140 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1161 ();
 FILLER_ASAP7_75t_R FILLER_114_1167 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1178 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1210 ();
 FILLER_ASAP7_75t_R FILLER_114_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1235 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1288 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1318 ();
 FILLER_ASAP7_75t_R FILLER_114_1328 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1330 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1356 ();
 FILLER_ASAP7_75t_R FILLER_114_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1377 ();
 FILLER_ASAP7_75t_R FILLER_114_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1388 ();
 FILLER_ASAP7_75t_R FILLER_115_8 ();
 FILLER_ASAP7_75t_R FILLER_115_25 ();
 FILLER_ASAP7_75t_R FILLER_115_53 ();
 DECAPx4_ASAP7_75t_R FILLER_115_87 ();
 FILLER_ASAP7_75t_R FILLER_115_97 ();
 DECAPx4_ASAP7_75t_R FILLER_115_111 ();
 DECAPx2_ASAP7_75t_R FILLER_115_151 ();
 DECAPx4_ASAP7_75t_R FILLER_115_164 ();
 FILLER_ASAP7_75t_R FILLER_115_174 ();
 FILLER_ASAP7_75t_R FILLER_115_190 ();
 DECAPx4_ASAP7_75t_R FILLER_115_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_214 ();
 DECAPx6_ASAP7_75t_R FILLER_115_223 ();
 FILLER_ASAP7_75t_R FILLER_115_237 ();
 FILLER_ASAP7_75t_R FILLER_115_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_255 ();
 DECAPx2_ASAP7_75t_R FILLER_115_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_276 ();
 FILLER_ASAP7_75t_R FILLER_115_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_285 ();
 DECAPx1_ASAP7_75t_R FILLER_115_302 ();
 FILLER_ASAP7_75t_R FILLER_115_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_322 ();
 DECAPx2_ASAP7_75t_R FILLER_115_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_343 ();
 DECAPx4_ASAP7_75t_R FILLER_115_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_364 ();
 DECAPx10_ASAP7_75t_R FILLER_115_383 ();
 FILLER_ASAP7_75t_R FILLER_115_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_407 ();
 DECAPx10_ASAP7_75t_R FILLER_115_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_448 ();
 FILLER_ASAP7_75t_R FILLER_115_459 ();
 DECAPx6_ASAP7_75t_R FILLER_115_471 ();
 FILLER_ASAP7_75t_R FILLER_115_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_514 ();
 DECAPx2_ASAP7_75t_R FILLER_115_521 ();
 FILLER_ASAP7_75t_R FILLER_115_527 ();
 DECAPx4_ASAP7_75t_R FILLER_115_535 ();
 FILLER_ASAP7_75t_R FILLER_115_545 ();
 DECAPx6_ASAP7_75t_R FILLER_115_559 ();
 DECAPx1_ASAP7_75t_R FILLER_115_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_584 ();
 DECAPx2_ASAP7_75t_R FILLER_115_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_630 ();
 DECAPx10_ASAP7_75t_R FILLER_115_637 ();
 DECAPx2_ASAP7_75t_R FILLER_115_666 ();
 FILLER_ASAP7_75t_R FILLER_115_672 ();
 FILLER_ASAP7_75t_R FILLER_115_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_689 ();
 DECAPx1_ASAP7_75t_R FILLER_115_710 ();
 DECAPx2_ASAP7_75t_R FILLER_115_723 ();
 FILLER_ASAP7_75t_R FILLER_115_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_731 ();
 DECAPx2_ASAP7_75t_R FILLER_115_738 ();
 DECAPx1_ASAP7_75t_R FILLER_115_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_755 ();
 FILLER_ASAP7_75t_R FILLER_115_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_770 ();
 DECAPx4_ASAP7_75t_R FILLER_115_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_792 ();
 DECAPx2_ASAP7_75t_R FILLER_115_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_823 ();
 DECAPx2_ASAP7_75t_R FILLER_115_875 ();
 FILLER_ASAP7_75t_R FILLER_115_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_883 ();
 DECAPx1_ASAP7_75t_R FILLER_115_891 ();
 DECAPx1_ASAP7_75t_R FILLER_115_901 ();
 DECAPx4_ASAP7_75t_R FILLER_115_914 ();
 DECAPx1_ASAP7_75t_R FILLER_115_944 ();
 DECAPx1_ASAP7_75t_R FILLER_115_958 ();
 DECAPx10_ASAP7_75t_R FILLER_115_987 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1111 ();
 DECAPx6_ASAP7_75t_R FILLER_115_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1174 ();
 FILLER_ASAP7_75t_R FILLER_115_1182 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1206 ();
 FILLER_ASAP7_75t_R FILLER_115_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_115_1225 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1247 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1268 ();
 FILLER_ASAP7_75t_R FILLER_115_1274 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1276 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1299 ();
 FILLER_ASAP7_75t_R FILLER_115_1305 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1333 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1344 ();
 FILLER_ASAP7_75t_R FILLER_115_1350 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1352 ();
 DECAPx6_ASAP7_75t_R FILLER_115_1370 ();
 FILLER_ASAP7_75t_R FILLER_115_1384 ();
 FILLER_ASAP7_75t_R FILLER_116_8 ();
 DECAPx4_ASAP7_75t_R FILLER_116_38 ();
 FILLER_ASAP7_75t_R FILLER_116_48 ();
 DECAPx2_ASAP7_75t_R FILLER_116_60 ();
 FILLER_ASAP7_75t_R FILLER_116_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_68 ();
 DECAPx4_ASAP7_75t_R FILLER_116_72 ();
 DECAPx2_ASAP7_75t_R FILLER_116_88 ();
 FILLER_ASAP7_75t_R FILLER_116_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_123 ();
 DECAPx2_ASAP7_75t_R FILLER_116_130 ();
 FILLER_ASAP7_75t_R FILLER_116_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_190 ();
 DECAPx4_ASAP7_75t_R FILLER_116_203 ();
 FILLER_ASAP7_75t_R FILLER_116_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_259 ();
 DECAPx2_ASAP7_75t_R FILLER_116_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_274 ();
 DECAPx2_ASAP7_75t_R FILLER_116_302 ();
 FILLER_ASAP7_75t_R FILLER_116_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_310 ();
 DECAPx1_ASAP7_75t_R FILLER_116_317 ();
 DECAPx6_ASAP7_75t_R FILLER_116_329 ();
 DECAPx2_ASAP7_75t_R FILLER_116_343 ();
 DECAPx6_ASAP7_75t_R FILLER_116_369 ();
 DECAPx1_ASAP7_75t_R FILLER_116_383 ();
 FILLER_ASAP7_75t_R FILLER_116_400 ();
 DECAPx2_ASAP7_75t_R FILLER_116_405 ();
 DECAPx1_ASAP7_75t_R FILLER_116_443 ();
 DECAPx2_ASAP7_75t_R FILLER_116_453 ();
 FILLER_ASAP7_75t_R FILLER_116_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_461 ();
 FILLER_ASAP7_75t_R FILLER_116_464 ();
 DECAPx6_ASAP7_75t_R FILLER_116_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_507 ();
 FILLER_ASAP7_75t_R FILLER_116_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_542 ();
 DECAPx2_ASAP7_75t_R FILLER_116_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_555 ();
 DECAPx10_ASAP7_75t_R FILLER_116_565 ();
 DECAPx4_ASAP7_75t_R FILLER_116_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_609 ();
 DECAPx2_ASAP7_75t_R FILLER_116_622 ();
 FILLER_ASAP7_75t_R FILLER_116_628 ();
 DECAPx4_ASAP7_75t_R FILLER_116_640 ();
 FILLER_ASAP7_75t_R FILLER_116_650 ();
 DECAPx1_ASAP7_75t_R FILLER_116_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_668 ();
 DECAPx4_ASAP7_75t_R FILLER_116_688 ();
 FILLER_ASAP7_75t_R FILLER_116_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_700 ();
 FILLER_ASAP7_75t_R FILLER_116_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_709 ();
 DECAPx4_ASAP7_75t_R FILLER_116_716 ();
 FILLER_ASAP7_75t_R FILLER_116_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_745 ();
 FILLER_ASAP7_75t_R FILLER_116_777 ();
 DECAPx4_ASAP7_75t_R FILLER_116_783 ();
 FILLER_ASAP7_75t_R FILLER_116_796 ();
 FILLER_ASAP7_75t_R FILLER_116_801 ();
 DECAPx6_ASAP7_75t_R FILLER_116_813 ();
 FILLER_ASAP7_75t_R FILLER_116_833 ();
 DECAPx4_ASAP7_75t_R FILLER_116_847 ();
 DECAPx6_ASAP7_75t_R FILLER_116_873 ();
 DECAPx2_ASAP7_75t_R FILLER_116_900 ();
 DECAPx2_ASAP7_75t_R FILLER_116_912 ();
 FILLER_ASAP7_75t_R FILLER_116_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_920 ();
 FILLER_ASAP7_75t_R FILLER_116_943 ();
 DECAPx10_ASAP7_75t_R FILLER_116_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_980 ();
 DECAPx1_ASAP7_75t_R FILLER_116_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_992 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1063 ();
 FILLER_ASAP7_75t_R FILLER_116_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1171 ();
 FILLER_ASAP7_75t_R FILLER_116_1177 ();
 FILLER_ASAP7_75t_R FILLER_116_1182 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1195 ();
 FILLER_ASAP7_75t_R FILLER_116_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1228 ();
 FILLER_ASAP7_75t_R FILLER_116_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1239 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1257 ();
 FILLER_ASAP7_75t_R FILLER_116_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1277 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1289 ();
 FILLER_ASAP7_75t_R FILLER_116_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1306 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1348 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1391 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_18 ();
 DECAPx4_ASAP7_75t_R FILLER_117_31 ();
 FILLER_ASAP7_75t_R FILLER_117_41 ();
 DECAPx6_ASAP7_75t_R FILLER_117_57 ();
 FILLER_ASAP7_75t_R FILLER_117_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_100 ();
 DECAPx1_ASAP7_75t_R FILLER_117_107 ();
 DECAPx2_ASAP7_75t_R FILLER_117_114 ();
 FILLER_ASAP7_75t_R FILLER_117_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_122 ();
 DECAPx6_ASAP7_75t_R FILLER_117_126 ();
 DECAPx1_ASAP7_75t_R FILLER_117_166 ();
 DECAPx2_ASAP7_75t_R FILLER_117_173 ();
 DECAPx1_ASAP7_75t_R FILLER_117_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_197 ();
 DECAPx4_ASAP7_75t_R FILLER_117_204 ();
 DECAPx1_ASAP7_75t_R FILLER_117_221 ();
 FILLER_ASAP7_75t_R FILLER_117_251 ();
 DECAPx4_ASAP7_75t_R FILLER_117_265 ();
 FILLER_ASAP7_75t_R FILLER_117_275 ();
 DECAPx6_ASAP7_75t_R FILLER_117_283 ();
 FILLER_ASAP7_75t_R FILLER_117_312 ();
 DECAPx2_ASAP7_75t_R FILLER_117_326 ();
 FILLER_ASAP7_75t_R FILLER_117_332 ();
 DECAPx10_ASAP7_75t_R FILLER_117_344 ();
 FILLER_ASAP7_75t_R FILLER_117_366 ();
 DECAPx2_ASAP7_75t_R FILLER_117_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_381 ();
 FILLER_ASAP7_75t_R FILLER_117_385 ();
 DECAPx1_ASAP7_75t_R FILLER_117_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_417 ();
 FILLER_ASAP7_75t_R FILLER_117_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_439 ();
 FILLER_ASAP7_75t_R FILLER_117_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_456 ();
 FILLER_ASAP7_75t_R FILLER_117_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_465 ();
 DECAPx6_ASAP7_75t_R FILLER_117_495 ();
 DECAPx2_ASAP7_75t_R FILLER_117_509 ();
 DECAPx2_ASAP7_75t_R FILLER_117_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_528 ();
 FILLER_ASAP7_75t_R FILLER_117_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_534 ();
 DECAPx10_ASAP7_75t_R FILLER_117_568 ();
 DECAPx6_ASAP7_75t_R FILLER_117_590 ();
 DECAPx1_ASAP7_75t_R FILLER_117_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_608 ();
 DECAPx2_ASAP7_75t_R FILLER_117_615 ();
 FILLER_ASAP7_75t_R FILLER_117_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_649 ();
 DECAPx1_ASAP7_75t_R FILLER_117_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_673 ();
 FILLER_ASAP7_75t_R FILLER_117_686 ();
 DECAPx10_ASAP7_75t_R FILLER_117_692 ();
 DECAPx6_ASAP7_75t_R FILLER_117_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_728 ();
 FILLER_ASAP7_75t_R FILLER_117_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_746 ();
 DECAPx4_ASAP7_75t_R FILLER_117_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_778 ();
 DECAPx10_ASAP7_75t_R FILLER_117_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_823 ();
 FILLER_ASAP7_75t_R FILLER_117_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_829 ();
 FILLER_ASAP7_75t_R FILLER_117_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_841 ();
 DECAPx2_ASAP7_75t_R FILLER_117_849 ();
 DECAPx2_ASAP7_75t_R FILLER_117_874 ();
 DECAPx2_ASAP7_75t_R FILLER_117_888 ();
 FILLER_ASAP7_75t_R FILLER_117_894 ();
 FILLER_ASAP7_75t_R FILLER_117_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_940 ();
 DECAPx6_ASAP7_75t_R FILLER_117_960 ();
 FILLER_ASAP7_75t_R FILLER_117_974 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1008 ();
 FILLER_ASAP7_75t_R FILLER_117_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1034 ();
 FILLER_ASAP7_75t_R FILLER_117_1056 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1064 ();
 FILLER_ASAP7_75t_R FILLER_117_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1119 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1163 ();
 FILLER_ASAP7_75t_R FILLER_117_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1186 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1193 ();
 FILLER_ASAP7_75t_R FILLER_117_1203 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1240 ();
 FILLER_ASAP7_75t_R FILLER_117_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1290 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1301 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1342 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_118_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_18 ();
 FILLER_ASAP7_75t_R FILLER_118_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_47 ();
 FILLER_ASAP7_75t_R FILLER_118_64 ();
 DECAPx4_ASAP7_75t_R FILLER_118_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_79 ();
 FILLER_ASAP7_75t_R FILLER_118_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_88 ();
 FILLER_ASAP7_75t_R FILLER_118_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_94 ();
 DECAPx2_ASAP7_75t_R FILLER_118_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_141 ();
 FILLER_ASAP7_75t_R FILLER_118_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_154 ();
 DECAPx10_ASAP7_75t_R FILLER_118_158 ();
 DECAPx4_ASAP7_75t_R FILLER_118_180 ();
 FILLER_ASAP7_75t_R FILLER_118_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_200 ();
 DECAPx4_ASAP7_75t_R FILLER_118_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_224 ();
 DECAPx2_ASAP7_75t_R FILLER_118_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_250 ();
 DECAPx2_ASAP7_75t_R FILLER_118_265 ();
 DECAPx10_ASAP7_75t_R FILLER_118_277 ();
 DECAPx2_ASAP7_75t_R FILLER_118_307 ();
 DECAPx6_ASAP7_75t_R FILLER_118_321 ();
 DECAPx4_ASAP7_75t_R FILLER_118_345 ();
 FILLER_ASAP7_75t_R FILLER_118_365 ();
 DECAPx1_ASAP7_75t_R FILLER_118_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_397 ();
 DECAPx6_ASAP7_75t_R FILLER_118_408 ();
 DECAPx2_ASAP7_75t_R FILLER_118_422 ();
 FILLER_ASAP7_75t_R FILLER_118_446 ();
 FILLER_ASAP7_75t_R FILLER_118_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_466 ();
 FILLER_ASAP7_75t_R FILLER_118_493 ();
 DECAPx4_ASAP7_75t_R FILLER_118_501 ();
 FILLER_ASAP7_75t_R FILLER_118_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_513 ();
 DECAPx10_ASAP7_75t_R FILLER_118_520 ();
 DECAPx4_ASAP7_75t_R FILLER_118_542 ();
 FILLER_ASAP7_75t_R FILLER_118_552 ();
 DECAPx2_ASAP7_75t_R FILLER_118_592 ();
 FILLER_ASAP7_75t_R FILLER_118_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_603 ();
 DECAPx10_ASAP7_75t_R FILLER_118_607 ();
 DECAPx1_ASAP7_75t_R FILLER_118_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_633 ();
 DECAPx2_ASAP7_75t_R FILLER_118_642 ();
 FILLER_ASAP7_75t_R FILLER_118_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_650 ();
 DECAPx4_ASAP7_75t_R FILLER_118_663 ();
 FILLER_ASAP7_75t_R FILLER_118_673 ();
 DECAPx4_ASAP7_75t_R FILLER_118_681 ();
 FILLER_ASAP7_75t_R FILLER_118_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_693 ();
 FILLER_ASAP7_75t_R FILLER_118_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_704 ();
 FILLER_ASAP7_75t_R FILLER_118_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_722 ();
 DECAPx4_ASAP7_75t_R FILLER_118_732 ();
 DECAPx10_ASAP7_75t_R FILLER_118_748 ();
 DECAPx1_ASAP7_75t_R FILLER_118_770 ();
 DECAPx2_ASAP7_75t_R FILLER_118_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_816 ();
 FILLER_ASAP7_75t_R FILLER_118_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_829 ();
 FILLER_ASAP7_75t_R FILLER_118_868 ();
 DECAPx10_ASAP7_75t_R FILLER_118_882 ();
 DECAPx6_ASAP7_75t_R FILLER_118_904 ();
 DECAPx6_ASAP7_75t_R FILLER_118_943 ();
 DECAPx2_ASAP7_75t_R FILLER_118_957 ();
 FILLER_ASAP7_75t_R FILLER_118_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_987 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1014 ();
 FILLER_ASAP7_75t_R FILLER_118_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1022 ();
 FILLER_ASAP7_75t_R FILLER_118_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1114 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1252 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1259 ();
 FILLER_ASAP7_75t_R FILLER_118_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1274 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1307 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1329 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1339 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1349 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1361 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1388 ();
 DECAPx1_ASAP7_75t_R FILLER_119_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_32 ();
 DECAPx6_ASAP7_75t_R FILLER_119_36 ();
 FILLER_ASAP7_75t_R FILLER_119_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_82 ();
 DECAPx2_ASAP7_75t_R FILLER_119_93 ();
 FILLER_ASAP7_75t_R FILLER_119_99 ();
 DECAPx2_ASAP7_75t_R FILLER_119_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_113 ();
 FILLER_ASAP7_75t_R FILLER_119_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_119 ();
 DECAPx2_ASAP7_75t_R FILLER_119_153 ();
 FILLER_ASAP7_75t_R FILLER_119_159 ();
 FILLER_ASAP7_75t_R FILLER_119_164 ();
 DECAPx6_ASAP7_75t_R FILLER_119_173 ();
 DECAPx1_ASAP7_75t_R FILLER_119_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_191 ();
 DECAPx6_ASAP7_75t_R FILLER_119_198 ();
 FILLER_ASAP7_75t_R FILLER_119_212 ();
 DECAPx10_ASAP7_75t_R FILLER_119_220 ();
 DECAPx4_ASAP7_75t_R FILLER_119_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_252 ();
 DECAPx2_ASAP7_75t_R FILLER_119_289 ();
 FILLER_ASAP7_75t_R FILLER_119_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_297 ();
 DECAPx6_ASAP7_75t_R FILLER_119_331 ();
 FILLER_ASAP7_75t_R FILLER_119_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_347 ();
 DECAPx1_ASAP7_75t_R FILLER_119_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_370 ();
 DECAPx10_ASAP7_75t_R FILLER_119_377 ();
 DECAPx6_ASAP7_75t_R FILLER_119_399 ();
 DECAPx1_ASAP7_75t_R FILLER_119_413 ();
 DECAPx6_ASAP7_75t_R FILLER_119_424 ();
 DECAPx1_ASAP7_75t_R FILLER_119_438 ();
 DECAPx1_ASAP7_75t_R FILLER_119_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_460 ();
 DECAPx2_ASAP7_75t_R FILLER_119_473 ();
 FILLER_ASAP7_75t_R FILLER_119_485 ();
 DECAPx2_ASAP7_75t_R FILLER_119_501 ();
 FILLER_ASAP7_75t_R FILLER_119_507 ();
 FILLER_ASAP7_75t_R FILLER_119_517 ();
 DECAPx2_ASAP7_75t_R FILLER_119_527 ();
 DECAPx1_ASAP7_75t_R FILLER_119_549 ();
 DECAPx1_ASAP7_75t_R FILLER_119_567 ();
 DECAPx2_ASAP7_75t_R FILLER_119_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_633 ();
 DECAPx2_ASAP7_75t_R FILLER_119_642 ();
 FILLER_ASAP7_75t_R FILLER_119_648 ();
 DECAPx6_ASAP7_75t_R FILLER_119_670 ();
 DECAPx1_ASAP7_75t_R FILLER_119_684 ();
 DECAPx2_ASAP7_75t_R FILLER_119_713 ();
 FILLER_ASAP7_75t_R FILLER_119_719 ();
 DECAPx2_ASAP7_75t_R FILLER_119_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_748 ();
 DECAPx4_ASAP7_75t_R FILLER_119_758 ();
 DECAPx6_ASAP7_75t_R FILLER_119_782 ();
 FILLER_ASAP7_75t_R FILLER_119_796 ();
 DECAPx2_ASAP7_75t_R FILLER_119_806 ();
 FILLER_ASAP7_75t_R FILLER_119_812 ();
 DECAPx10_ASAP7_75t_R FILLER_119_824 ();
 FILLER_ASAP7_75t_R FILLER_119_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_848 ();
 DECAPx2_ASAP7_75t_R FILLER_119_855 ();
 DECAPx10_ASAP7_75t_R FILLER_119_864 ();
 DECAPx1_ASAP7_75t_R FILLER_119_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_905 ();
 DECAPx4_ASAP7_75t_R FILLER_119_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_923 ();
 FILLER_ASAP7_75t_R FILLER_119_926 ();
 DECAPx2_ASAP7_75t_R FILLER_119_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_972 ();
 DECAPx1_ASAP7_75t_R FILLER_119_998 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1070 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1084 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1101 ();
 FILLER_ASAP7_75t_R FILLER_119_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1123 ();
 FILLER_ASAP7_75t_R FILLER_119_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1156 ();
 FILLER_ASAP7_75t_R FILLER_119_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1173 ();
 FILLER_ASAP7_75t_R FILLER_119_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1229 ();
 DECAPx6_ASAP7_75t_R FILLER_119_1251 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1287 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1309 ();
 DECAPx6_ASAP7_75t_R FILLER_119_1322 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1368 ();
 FILLER_ASAP7_75t_R FILLER_119_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1385 ();
 DECAPx4_ASAP7_75t_R FILLER_120_27 ();
 FILLER_ASAP7_75t_R FILLER_120_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_39 ();
 DECAPx2_ASAP7_75t_R FILLER_120_49 ();
 FILLER_ASAP7_75t_R FILLER_120_55 ();
 DECAPx10_ASAP7_75t_R FILLER_120_63 ();
 FILLER_ASAP7_75t_R FILLER_120_85 ();
 DECAPx10_ASAP7_75t_R FILLER_120_91 ();
 DECAPx2_ASAP7_75t_R FILLER_120_113 ();
 FILLER_ASAP7_75t_R FILLER_120_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_133 ();
 DECAPx2_ASAP7_75t_R FILLER_120_137 ();
 FILLER_ASAP7_75t_R FILLER_120_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_172 ();
 DECAPx1_ASAP7_75t_R FILLER_120_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_183 ();
 DECAPx2_ASAP7_75t_R FILLER_120_206 ();
 DECAPx4_ASAP7_75t_R FILLER_120_226 ();
 FILLER_ASAP7_75t_R FILLER_120_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_238 ();
 DECAPx2_ASAP7_75t_R FILLER_120_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_251 ();
 DECAPx6_ASAP7_75t_R FILLER_120_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_272 ();
 DECAPx4_ASAP7_75t_R FILLER_120_289 ();
 DECAPx6_ASAP7_75t_R FILLER_120_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_320 ();
 FILLER_ASAP7_75t_R FILLER_120_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_335 ();
 DECAPx1_ASAP7_75t_R FILLER_120_346 ();
 DECAPx1_ASAP7_75t_R FILLER_120_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_439 ();
 DECAPx2_ASAP7_75t_R FILLER_120_454 ();
 FILLER_ASAP7_75t_R FILLER_120_460 ();
 FILLER_ASAP7_75t_R FILLER_120_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_466 ();
 DECAPx6_ASAP7_75t_R FILLER_120_473 ();
 FILLER_ASAP7_75t_R FILLER_120_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_509 ();
 FILLER_ASAP7_75t_R FILLER_120_524 ();
 FILLER_ASAP7_75t_R FILLER_120_545 ();
 FILLER_ASAP7_75t_R FILLER_120_550 ();
 DECAPx2_ASAP7_75t_R FILLER_120_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_577 ();
 DECAPx6_ASAP7_75t_R FILLER_120_610 ();
 DECAPx1_ASAP7_75t_R FILLER_120_624 ();
 DECAPx2_ASAP7_75t_R FILLER_120_631 ();
 DECAPx1_ASAP7_75t_R FILLER_120_645 ();
 DECAPx1_ASAP7_75t_R FILLER_120_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_667 ();
 DECAPx2_ASAP7_75t_R FILLER_120_684 ();
 FILLER_ASAP7_75t_R FILLER_120_690 ();
 DECAPx1_ASAP7_75t_R FILLER_120_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_704 ();
 DECAPx1_ASAP7_75t_R FILLER_120_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_718 ();
 DECAPx4_ASAP7_75t_R FILLER_120_731 ();
 FILLER_ASAP7_75t_R FILLER_120_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_743 ();
 FILLER_ASAP7_75t_R FILLER_120_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_767 ();
 FILLER_ASAP7_75t_R FILLER_120_784 ();
 DECAPx2_ASAP7_75t_R FILLER_120_802 ();
 FILLER_ASAP7_75t_R FILLER_120_808 ();
 DECAPx2_ASAP7_75t_R FILLER_120_813 ();
 FILLER_ASAP7_75t_R FILLER_120_819 ();
 DECAPx4_ASAP7_75t_R FILLER_120_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_843 ();
 DECAPx2_ASAP7_75t_R FILLER_120_861 ();
 FILLER_ASAP7_75t_R FILLER_120_867 ();
 DECAPx1_ASAP7_75t_R FILLER_120_875 ();
 FILLER_ASAP7_75t_R FILLER_120_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_895 ();
 FILLER_ASAP7_75t_R FILLER_120_905 ();
 FILLER_ASAP7_75t_R FILLER_120_919 ();
 DECAPx6_ASAP7_75t_R FILLER_120_961 ();
 DECAPx2_ASAP7_75t_R FILLER_120_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_981 ();
 DECAPx6_ASAP7_75t_R FILLER_120_994 ();
 FILLER_ASAP7_75t_R FILLER_120_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1086 ();
 DECAPx6_ASAP7_75t_R FILLER_120_1149 ();
 FILLER_ASAP7_75t_R FILLER_120_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1202 ();
 FILLER_ASAP7_75t_R FILLER_120_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1236 ();
 DECAPx6_ASAP7_75t_R FILLER_120_1256 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1270 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1294 ();
 FILLER_ASAP7_75t_R FILLER_120_1300 ();
 FILLER_ASAP7_75t_R FILLER_120_1312 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1314 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1323 ();
 FILLER_ASAP7_75t_R FILLER_120_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1331 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1342 ();
 FILLER_ASAP7_75t_R FILLER_120_1348 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_121_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_30 ();
 DECAPx1_ASAP7_75t_R FILLER_121_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_77 ();
 FILLER_ASAP7_75t_R FILLER_121_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_83 ();
 DECAPx10_ASAP7_75t_R FILLER_121_110 ();
 DECAPx6_ASAP7_75t_R FILLER_121_132 ();
 FILLER_ASAP7_75t_R FILLER_121_146 ();
 DECAPx2_ASAP7_75t_R FILLER_121_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_160 ();
 DECAPx4_ASAP7_75t_R FILLER_121_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_218 ();
 DECAPx2_ASAP7_75t_R FILLER_121_233 ();
 DECAPx2_ASAP7_75t_R FILLER_121_247 ();
 DECAPx2_ASAP7_75t_R FILLER_121_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_286 ();
 DECAPx1_ASAP7_75t_R FILLER_121_294 ();
 DECAPx10_ASAP7_75t_R FILLER_121_306 ();
 DECAPx10_ASAP7_75t_R FILLER_121_328 ();
 DECAPx10_ASAP7_75t_R FILLER_121_350 ();
 DECAPx4_ASAP7_75t_R FILLER_121_372 ();
 FILLER_ASAP7_75t_R FILLER_121_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_384 ();
 FILLER_ASAP7_75t_R FILLER_121_395 ();
 DECAPx1_ASAP7_75t_R FILLER_121_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_423 ();
 DECAPx4_ASAP7_75t_R FILLER_121_427 ();
 FILLER_ASAP7_75t_R FILLER_121_449 ();
 FILLER_ASAP7_75t_R FILLER_121_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_459 ();
 DECAPx6_ASAP7_75t_R FILLER_121_472 ();
 FILLER_ASAP7_75t_R FILLER_121_486 ();
 DECAPx1_ASAP7_75t_R FILLER_121_520 ();
 FILLER_ASAP7_75t_R FILLER_121_530 ();
 DECAPx2_ASAP7_75t_R FILLER_121_558 ();
 DECAPx1_ASAP7_75t_R FILLER_121_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_574 ();
 FILLER_ASAP7_75t_R FILLER_121_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_616 ();
 DECAPx4_ASAP7_75t_R FILLER_121_658 ();
 DECAPx1_ASAP7_75t_R FILLER_121_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_692 ();
 DECAPx6_ASAP7_75t_R FILLER_121_701 ();
 DECAPx1_ASAP7_75t_R FILLER_121_715 ();
 DECAPx6_ASAP7_75t_R FILLER_121_725 ();
 FILLER_ASAP7_75t_R FILLER_121_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_741 ();
 DECAPx2_ASAP7_75t_R FILLER_121_754 ();
 DECAPx1_ASAP7_75t_R FILLER_121_766 ();
 DECAPx4_ASAP7_75t_R FILLER_121_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_786 ();
 DECAPx4_ASAP7_75t_R FILLER_121_795 ();
 FILLER_ASAP7_75t_R FILLER_121_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_807 ();
 DECAPx1_ASAP7_75t_R FILLER_121_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_821 ();
 DECAPx2_ASAP7_75t_R FILLER_121_834 ();
 FILLER_ASAP7_75t_R FILLER_121_840 ();
 DECAPx2_ASAP7_75t_R FILLER_121_861 ();
 DECAPx1_ASAP7_75t_R FILLER_121_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_881 ();
 DECAPx1_ASAP7_75t_R FILLER_121_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_895 ();
 DECAPx1_ASAP7_75t_R FILLER_121_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_909 ();
 DECAPx1_ASAP7_75t_R FILLER_121_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_923 ();
 FILLER_ASAP7_75t_R FILLER_121_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_939 ();
 DECAPx10_ASAP7_75t_R FILLER_121_967 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1015 ();
 FILLER_ASAP7_75t_R FILLER_121_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1030 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1088 ();
 FILLER_ASAP7_75t_R FILLER_121_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1152 ();
 FILLER_ASAP7_75t_R FILLER_121_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1193 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1249 ();
 FILLER_ASAP7_75t_R FILLER_121_1277 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1279 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1339 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1346 ();
 FILLER_ASAP7_75t_R FILLER_121_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1358 ();
 FILLER_ASAP7_75t_R FILLER_121_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1369 ();
 FILLER_ASAP7_75t_R FILLER_122_8 ();
 DECAPx1_ASAP7_75t_R FILLER_122_25 ();
 FILLER_ASAP7_75t_R FILLER_122_33 ();
 FILLER_ASAP7_75t_R FILLER_122_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_96 ();
 DECAPx2_ASAP7_75t_R FILLER_122_127 ();
 FILLER_ASAP7_75t_R FILLER_122_133 ();
 DECAPx4_ASAP7_75t_R FILLER_122_165 ();
 DECAPx1_ASAP7_75t_R FILLER_122_178 ();
 DECAPx4_ASAP7_75t_R FILLER_122_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_226 ();
 DECAPx6_ASAP7_75t_R FILLER_122_253 ();
 DECAPx4_ASAP7_75t_R FILLER_122_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_285 ();
 FILLER_ASAP7_75t_R FILLER_122_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_308 ();
 FILLER_ASAP7_75t_R FILLER_122_315 ();
 DECAPx10_ASAP7_75t_R FILLER_122_324 ();
 FILLER_ASAP7_75t_R FILLER_122_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_367 ();
 DECAPx1_ASAP7_75t_R FILLER_122_386 ();
 DECAPx6_ASAP7_75t_R FILLER_122_400 ();
 DECAPx1_ASAP7_75t_R FILLER_122_414 ();
 DECAPx4_ASAP7_75t_R FILLER_122_428 ();
 FILLER_ASAP7_75t_R FILLER_122_438 ();
 FILLER_ASAP7_75t_R FILLER_122_448 ();
 DECAPx1_ASAP7_75t_R FILLER_122_458 ();
 DECAPx6_ASAP7_75t_R FILLER_122_490 ();
 DECAPx1_ASAP7_75t_R FILLER_122_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_508 ();
 DECAPx6_ASAP7_75t_R FILLER_122_518 ();
 FILLER_ASAP7_75t_R FILLER_122_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_534 ();
 DECAPx10_ASAP7_75t_R FILLER_122_538 ();
 FILLER_ASAP7_75t_R FILLER_122_560 ();
 DECAPx4_ASAP7_75t_R FILLER_122_606 ();
 FILLER_ASAP7_75t_R FILLER_122_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_618 ();
 DECAPx4_ASAP7_75t_R FILLER_122_631 ();
 FILLER_ASAP7_75t_R FILLER_122_641 ();
 DECAPx2_ASAP7_75t_R FILLER_122_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_700 ();
 DECAPx2_ASAP7_75t_R FILLER_122_707 ();
 FILLER_ASAP7_75t_R FILLER_122_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_715 ();
 DECAPx4_ASAP7_75t_R FILLER_122_725 ();
 DECAPx6_ASAP7_75t_R FILLER_122_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_769 ();
 DECAPx1_ASAP7_75t_R FILLER_122_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_780 ();
 DECAPx4_ASAP7_75t_R FILLER_122_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_807 ();
 DECAPx2_ASAP7_75t_R FILLER_122_839 ();
 FILLER_ASAP7_75t_R FILLER_122_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_847 ();
 DECAPx4_ASAP7_75t_R FILLER_122_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_890 ();
 FILLER_ASAP7_75t_R FILLER_122_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_899 ();
 DECAPx2_ASAP7_75t_R FILLER_122_915 ();
 DECAPx4_ASAP7_75t_R FILLER_122_933 ();
 FILLER_ASAP7_75t_R FILLER_122_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_945 ();
 FILLER_ASAP7_75t_R FILLER_122_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_957 ();
 DECAPx4_ASAP7_75t_R FILLER_122_965 ();
 FILLER_ASAP7_75t_R FILLER_122_993 ();
 FILLER_ASAP7_75t_R FILLER_122_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1003 ();
 FILLER_ASAP7_75t_R FILLER_122_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1123 ();
 FILLER_ASAP7_75t_R FILLER_122_1129 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1213 ();
 FILLER_ASAP7_75t_R FILLER_122_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1250 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1295 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1301 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1322 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1340 ();
 FILLER_ASAP7_75t_R FILLER_122_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1388 ();
 DECAPx1_ASAP7_75t_R FILLER_123_2 ();
 DECAPx2_ASAP7_75t_R FILLER_123_32 ();
 FILLER_ASAP7_75t_R FILLER_123_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_67 ();
 DECAPx4_ASAP7_75t_R FILLER_123_74 ();
 FILLER_ASAP7_75t_R FILLER_123_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_93 ();
 FILLER_ASAP7_75t_R FILLER_123_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_111 ();
 DECAPx1_ASAP7_75t_R FILLER_123_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_151 ();
 FILLER_ASAP7_75t_R FILLER_123_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_186 ();
 DECAPx6_ASAP7_75t_R FILLER_123_193 ();
 DECAPx2_ASAP7_75t_R FILLER_123_207 ();
 DECAPx6_ASAP7_75t_R FILLER_123_221 ();
 DECAPx2_ASAP7_75t_R FILLER_123_235 ();
 FILLER_ASAP7_75t_R FILLER_123_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_269 ();
 DECAPx2_ASAP7_75t_R FILLER_123_276 ();
 FILLER_ASAP7_75t_R FILLER_123_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_284 ();
 FILLER_ASAP7_75t_R FILLER_123_315 ();
 DECAPx2_ASAP7_75t_R FILLER_123_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_386 ();
 DECAPx10_ASAP7_75t_R FILLER_123_397 ();
 DECAPx2_ASAP7_75t_R FILLER_123_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_435 ();
 FILLER_ASAP7_75t_R FILLER_123_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_458 ();
 DECAPx1_ASAP7_75t_R FILLER_123_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_477 ();
 DECAPx2_ASAP7_75t_R FILLER_123_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_496 ();
 DECAPx2_ASAP7_75t_R FILLER_123_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_506 ();
 DECAPx1_ASAP7_75t_R FILLER_123_525 ();
 FILLER_ASAP7_75t_R FILLER_123_539 ();
 DECAPx2_ASAP7_75t_R FILLER_123_547 ();
 DECAPx2_ASAP7_75t_R FILLER_123_556 ();
 FILLER_ASAP7_75t_R FILLER_123_562 ();
 FILLER_ASAP7_75t_R FILLER_123_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_624 ();
 DECAPx10_ASAP7_75t_R FILLER_123_642 ();
 DECAPx10_ASAP7_75t_R FILLER_123_664 ();
 DECAPx2_ASAP7_75t_R FILLER_123_686 ();
 FILLER_ASAP7_75t_R FILLER_123_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_694 ();
 DECAPx2_ASAP7_75t_R FILLER_123_728 ();
 DECAPx1_ASAP7_75t_R FILLER_123_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_761 ();
 FILLER_ASAP7_75t_R FILLER_123_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_776 ();
 FILLER_ASAP7_75t_R FILLER_123_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_786 ();
 DECAPx1_ASAP7_75t_R FILLER_123_803 ();
 DECAPx6_ASAP7_75t_R FILLER_123_832 ();
 FILLER_ASAP7_75t_R FILLER_123_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_848 ();
 DECAPx4_ASAP7_75t_R FILLER_123_855 ();
 FILLER_ASAP7_75t_R FILLER_123_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_867 ();
 DECAPx2_ASAP7_75t_R FILLER_123_874 ();
 DECAPx6_ASAP7_75t_R FILLER_123_886 ();
 DECAPx4_ASAP7_75t_R FILLER_123_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_916 ();
 FILLER_ASAP7_75t_R FILLER_123_938 ();
 DECAPx4_ASAP7_75t_R FILLER_123_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_993 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1020 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_123_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1116 ();
 FILLER_ASAP7_75t_R FILLER_123_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1135 ();
 FILLER_ASAP7_75t_R FILLER_123_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_123_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1171 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1197 ();
 FILLER_ASAP7_75t_R FILLER_123_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1249 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1265 ();
 DECAPx4_ASAP7_75t_R FILLER_123_1277 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_123_1294 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1316 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1330 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1341 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1366 ();
 FILLER_ASAP7_75t_R FILLER_123_1372 ();
 DECAPx10_ASAP7_75t_R FILLER_124_32 ();
 DECAPx2_ASAP7_75t_R FILLER_124_54 ();
 FILLER_ASAP7_75t_R FILLER_124_60 ();
 DECAPx10_ASAP7_75t_R FILLER_124_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_127 ();
 FILLER_ASAP7_75t_R FILLER_124_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_152 ();
 FILLER_ASAP7_75t_R FILLER_124_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_171 ();
 DECAPx6_ASAP7_75t_R FILLER_124_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_212 ();
 DECAPx4_ASAP7_75t_R FILLER_124_231 ();
 FILLER_ASAP7_75t_R FILLER_124_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_257 ();
 DECAPx6_ASAP7_75t_R FILLER_124_270 ();
 DECAPx2_ASAP7_75t_R FILLER_124_284 ();
 DECAPx2_ASAP7_75t_R FILLER_124_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_304 ();
 FILLER_ASAP7_75t_R FILLER_124_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_313 ();
 DECAPx6_ASAP7_75t_R FILLER_124_352 ();
 FILLER_ASAP7_75t_R FILLER_124_366 ();
 DECAPx6_ASAP7_75t_R FILLER_124_386 ();
 DECAPx2_ASAP7_75t_R FILLER_124_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_406 ();
 FILLER_ASAP7_75t_R FILLER_124_443 ();
 DECAPx4_ASAP7_75t_R FILLER_124_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_461 ();
 DECAPx2_ASAP7_75t_R FILLER_124_470 ();
 FILLER_ASAP7_75t_R FILLER_124_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_478 ();
 FILLER_ASAP7_75t_R FILLER_124_505 ();
 DECAPx2_ASAP7_75t_R FILLER_124_571 ();
 DECAPx6_ASAP7_75t_R FILLER_124_616 ();
 DECAPx1_ASAP7_75t_R FILLER_124_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_634 ();
 DECAPx2_ASAP7_75t_R FILLER_124_643 ();
 DECAPx1_ASAP7_75t_R FILLER_124_656 ();
 DECAPx4_ASAP7_75t_R FILLER_124_672 ();
 DECAPx1_ASAP7_75t_R FILLER_124_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_696 ();
 DECAPx2_ASAP7_75t_R FILLER_124_705 ();
 FILLER_ASAP7_75t_R FILLER_124_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_713 ();
 DECAPx1_ASAP7_75t_R FILLER_124_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_741 ();
 DECAPx6_ASAP7_75t_R FILLER_124_771 ();
 FILLER_ASAP7_75t_R FILLER_124_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_804 ();
 DECAPx4_ASAP7_75t_R FILLER_124_813 ();
 FILLER_ASAP7_75t_R FILLER_124_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_834 ();
 DECAPx6_ASAP7_75t_R FILLER_124_853 ();
 DECAPx2_ASAP7_75t_R FILLER_124_876 ();
 FILLER_ASAP7_75t_R FILLER_124_882 ();
 DECAPx1_ASAP7_75t_R FILLER_124_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_897 ();
 DECAPx10_ASAP7_75t_R FILLER_124_907 ();
 DECAPx10_ASAP7_75t_R FILLER_124_929 ();
 DECAPx6_ASAP7_75t_R FILLER_124_951 ();
 FILLER_ASAP7_75t_R FILLER_124_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_977 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1138 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1181 ();
 FILLER_ASAP7_75t_R FILLER_124_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1206 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1234 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1262 ();
 DECAPx6_ASAP7_75t_R FILLER_124_1278 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_124_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1341 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1373 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_125_23 ();
 FILLER_ASAP7_75t_R FILLER_125_37 ();
 DECAPx2_ASAP7_75t_R FILLER_125_48 ();
 DECAPx2_ASAP7_75t_R FILLER_125_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_86 ();
 FILLER_ASAP7_75t_R FILLER_125_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_95 ();
 DECAPx1_ASAP7_75t_R FILLER_125_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_106 ();
 DECAPx10_ASAP7_75t_R FILLER_125_110 ();
 DECAPx10_ASAP7_75t_R FILLER_125_132 ();
 DECAPx6_ASAP7_75t_R FILLER_125_154 ();
 DECAPx1_ASAP7_75t_R FILLER_125_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_172 ();
 DECAPx2_ASAP7_75t_R FILLER_125_180 ();
 FILLER_ASAP7_75t_R FILLER_125_189 ();
 DECAPx2_ASAP7_75t_R FILLER_125_197 ();
 FILLER_ASAP7_75t_R FILLER_125_203 ();
 DECAPx2_ASAP7_75t_R FILLER_125_239 ();
 FILLER_ASAP7_75t_R FILLER_125_245 ();
 FILLER_ASAP7_75t_R FILLER_125_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_255 ();
 DECAPx2_ASAP7_75t_R FILLER_125_264 ();
 DECAPx6_ASAP7_75t_R FILLER_125_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_290 ();
 FILLER_ASAP7_75t_R FILLER_125_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_299 ();
 DECAPx6_ASAP7_75t_R FILLER_125_306 ();
 DECAPx2_ASAP7_75t_R FILLER_125_320 ();
 DECAPx1_ASAP7_75t_R FILLER_125_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_340 ();
 DECAPx10_ASAP7_75t_R FILLER_125_344 ();
 DECAPx4_ASAP7_75t_R FILLER_125_366 ();
 DECAPx10_ASAP7_75t_R FILLER_125_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_446 ();
 DECAPx2_ASAP7_75t_R FILLER_125_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_463 ();
 DECAPx2_ASAP7_75t_R FILLER_125_474 ();
 DECAPx6_ASAP7_75t_R FILLER_125_486 ();
 DECAPx6_ASAP7_75t_R FILLER_125_506 ();
 DECAPx1_ASAP7_75t_R FILLER_125_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_538 ();
 DECAPx1_ASAP7_75t_R FILLER_125_545 ();
 DECAPx4_ASAP7_75t_R FILLER_125_559 ();
 FILLER_ASAP7_75t_R FILLER_125_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_571 ();
 DECAPx1_ASAP7_75t_R FILLER_125_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_600 ();
 DECAPx10_ASAP7_75t_R FILLER_125_604 ();
 DECAPx2_ASAP7_75t_R FILLER_125_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_632 ();
 DECAPx2_ASAP7_75t_R FILLER_125_676 ();
 FILLER_ASAP7_75t_R FILLER_125_682 ();
 DECAPx2_ASAP7_75t_R FILLER_125_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_716 ();
 DECAPx10_ASAP7_75t_R FILLER_125_734 ();
 DECAPx2_ASAP7_75t_R FILLER_125_756 ();
 FILLER_ASAP7_75t_R FILLER_125_762 ();
 DECAPx6_ASAP7_75t_R FILLER_125_776 ();
 DECAPx1_ASAP7_75t_R FILLER_125_790 ();
 DECAPx6_ASAP7_75t_R FILLER_125_797 ();
 FILLER_ASAP7_75t_R FILLER_125_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_813 ();
 FILLER_ASAP7_75t_R FILLER_125_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_824 ();
 DECAPx2_ASAP7_75t_R FILLER_125_831 ();
 FILLER_ASAP7_75t_R FILLER_125_837 ();
 DECAPx2_ASAP7_75t_R FILLER_125_859 ();
 FILLER_ASAP7_75t_R FILLER_125_865 ();
 DECAPx1_ASAP7_75t_R FILLER_125_876 ();
 DECAPx2_ASAP7_75t_R FILLER_125_911 ();
 DECAPx6_ASAP7_75t_R FILLER_125_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_940 ();
 DECAPx2_ASAP7_75t_R FILLER_125_948 ();
 FILLER_ASAP7_75t_R FILLER_125_954 ();
 DECAPx6_ASAP7_75t_R FILLER_125_963 ();
 DECAPx10_ASAP7_75t_R FILLER_125_987 ();
 FILLER_ASAP7_75t_R FILLER_125_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1042 ();
 FILLER_ASAP7_75t_R FILLER_125_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1101 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1108 ();
 FILLER_ASAP7_75t_R FILLER_125_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1138 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1164 ();
 FILLER_ASAP7_75t_R FILLER_125_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1201 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1256 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1260 ();
 FILLER_ASAP7_75t_R FILLER_125_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1308 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_8 ();
 DECAPx2_ASAP7_75t_R FILLER_126_21 ();
 FILLER_ASAP7_75t_R FILLER_126_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_29 ();
 DECAPx4_ASAP7_75t_R FILLER_126_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_66 ();
 DECAPx2_ASAP7_75t_R FILLER_126_119 ();
 DECAPx2_ASAP7_75t_R FILLER_126_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_137 ();
 DECAPx2_ASAP7_75t_R FILLER_126_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_154 ();
 DECAPx10_ASAP7_75t_R FILLER_126_162 ();
 DECAPx1_ASAP7_75t_R FILLER_126_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_188 ();
 DECAPx2_ASAP7_75t_R FILLER_126_203 ();
 FILLER_ASAP7_75t_R FILLER_126_215 ();
 FILLER_ASAP7_75t_R FILLER_126_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_227 ();
 FILLER_ASAP7_75t_R FILLER_126_234 ();
 DECAPx2_ASAP7_75t_R FILLER_126_262 ();
 FILLER_ASAP7_75t_R FILLER_126_268 ();
 DECAPx4_ASAP7_75t_R FILLER_126_282 ();
 FILLER_ASAP7_75t_R FILLER_126_292 ();
 DECAPx10_ASAP7_75t_R FILLER_126_308 ();
 DECAPx1_ASAP7_75t_R FILLER_126_330 ();
 DECAPx6_ASAP7_75t_R FILLER_126_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_356 ();
 DECAPx2_ASAP7_75t_R FILLER_126_371 ();
 FILLER_ASAP7_75t_R FILLER_126_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_379 ();
 DECAPx2_ASAP7_75t_R FILLER_126_390 ();
 FILLER_ASAP7_75t_R FILLER_126_396 ();
 DECAPx2_ASAP7_75t_R FILLER_126_428 ();
 FILLER_ASAP7_75t_R FILLER_126_444 ();
 DECAPx2_ASAP7_75t_R FILLER_126_456 ();
 DECAPx2_ASAP7_75t_R FILLER_126_464 ();
 DECAPx2_ASAP7_75t_R FILLER_126_480 ();
 FILLER_ASAP7_75t_R FILLER_126_486 ();
 FILLER_ASAP7_75t_R FILLER_126_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_500 ();
 DECAPx6_ASAP7_75t_R FILLER_126_507 ();
 DECAPx1_ASAP7_75t_R FILLER_126_521 ();
 DECAPx1_ASAP7_75t_R FILLER_126_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_551 ();
 DECAPx6_ASAP7_75t_R FILLER_126_562 ();
 DECAPx1_ASAP7_75t_R FILLER_126_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_580 ();
 DECAPx2_ASAP7_75t_R FILLER_126_607 ();
 FILLER_ASAP7_75t_R FILLER_126_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_623 ();
 DECAPx1_ASAP7_75t_R FILLER_126_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_656 ();
 FILLER_ASAP7_75t_R FILLER_126_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_667 ();
 DECAPx10_ASAP7_75t_R FILLER_126_675 ();
 DECAPx1_ASAP7_75t_R FILLER_126_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_701 ();
 DECAPx6_ASAP7_75t_R FILLER_126_712 ();
 DECAPx10_ASAP7_75t_R FILLER_126_745 ();
 DECAPx1_ASAP7_75t_R FILLER_126_777 ();
 DECAPx2_ASAP7_75t_R FILLER_126_805 ();
 FILLER_ASAP7_75t_R FILLER_126_811 ();
 DECAPx4_ASAP7_75t_R FILLER_126_829 ();
 FILLER_ASAP7_75t_R FILLER_126_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_841 ();
 FILLER_ASAP7_75t_R FILLER_126_845 ();
 DECAPx4_ASAP7_75t_R FILLER_126_875 ();
 DECAPx4_ASAP7_75t_R FILLER_126_888 ();
 FILLER_ASAP7_75t_R FILLER_126_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_916 ();
 FILLER_ASAP7_75t_R FILLER_126_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_926 ();
 FILLER_ASAP7_75t_R FILLER_126_939 ();
 FILLER_ASAP7_75t_R FILLER_126_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_953 ();
 DECAPx10_ASAP7_75t_R FILLER_126_964 ();
 FILLER_ASAP7_75t_R FILLER_126_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1062 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1073 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1080 ();
 FILLER_ASAP7_75t_R FILLER_126_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1092 ();
 DECAPx6_ASAP7_75t_R FILLER_126_1113 ();
 FILLER_ASAP7_75t_R FILLER_126_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1132 ();
 DECAPx6_ASAP7_75t_R FILLER_126_1155 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1195 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1216 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1228 ();
 FILLER_ASAP7_75t_R FILLER_126_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1238 ();
 DECAPx2_ASAP7_75t_R FILLER_126_1255 ();
 FILLER_ASAP7_75t_R FILLER_126_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1263 ();
 FILLER_ASAP7_75t_R FILLER_126_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1283 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1335 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1344 ();
 FILLER_ASAP7_75t_R FILLER_126_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1388 ();
 DECAPx1_ASAP7_75t_R FILLER_127_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_6 ();
 FILLER_ASAP7_75t_R FILLER_127_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_41 ();
 FILLER_ASAP7_75t_R FILLER_127_48 ();
 FILLER_ASAP7_75t_R FILLER_127_62 ();
 DECAPx1_ASAP7_75t_R FILLER_127_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_72 ();
 FILLER_ASAP7_75t_R FILLER_127_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_133 ();
 DECAPx2_ASAP7_75t_R FILLER_127_137 ();
 DECAPx2_ASAP7_75t_R FILLER_127_146 ();
 FILLER_ASAP7_75t_R FILLER_127_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_180 ();
 FILLER_ASAP7_75t_R FILLER_127_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_197 ();
 DECAPx4_ASAP7_75t_R FILLER_127_206 ();
 FILLER_ASAP7_75t_R FILLER_127_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_218 ();
 DECAPx6_ASAP7_75t_R FILLER_127_227 ();
 DECAPx2_ASAP7_75t_R FILLER_127_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_247 ();
 DECAPx1_ASAP7_75t_R FILLER_127_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_260 ();
 FILLER_ASAP7_75t_R FILLER_127_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_269 ();
 FILLER_ASAP7_75t_R FILLER_127_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_280 ();
 DECAPx1_ASAP7_75t_R FILLER_127_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_291 ();
 DECAPx4_ASAP7_75t_R FILLER_127_315 ();
 FILLER_ASAP7_75t_R FILLER_127_325 ();
 DECAPx1_ASAP7_75t_R FILLER_127_354 ();
 DECAPx4_ASAP7_75t_R FILLER_127_374 ();
 DECAPx1_ASAP7_75t_R FILLER_127_390 ();
 FILLER_ASAP7_75t_R FILLER_127_400 ();
 DECAPx4_ASAP7_75t_R FILLER_127_408 ();
 FILLER_ASAP7_75t_R FILLER_127_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_420 ();
 FILLER_ASAP7_75t_R FILLER_127_431 ();
 DECAPx2_ASAP7_75t_R FILLER_127_443 ();
 FILLER_ASAP7_75t_R FILLER_127_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_461 ();
 DECAPx2_ASAP7_75t_R FILLER_127_470 ();
 FILLER_ASAP7_75t_R FILLER_127_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_478 ();
 DECAPx1_ASAP7_75t_R FILLER_127_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_523 ();
 DECAPx6_ASAP7_75t_R FILLER_127_530 ();
 DECAPx2_ASAP7_75t_R FILLER_127_544 ();
 DECAPx2_ASAP7_75t_R FILLER_127_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_584 ();
 DECAPx1_ASAP7_75t_R FILLER_127_591 ();
 DECAPx1_ASAP7_75t_R FILLER_127_627 ();
 DECAPx1_ASAP7_75t_R FILLER_127_641 ();
 DECAPx10_ASAP7_75t_R FILLER_127_658 ();
 DECAPx4_ASAP7_75t_R FILLER_127_680 ();
 DECAPx6_ASAP7_75t_R FILLER_127_716 ();
 FILLER_ASAP7_75t_R FILLER_127_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_735 ();
 FILLER_ASAP7_75t_R FILLER_127_754 ();
 DECAPx1_ASAP7_75t_R FILLER_127_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_769 ();
 FILLER_ASAP7_75t_R FILLER_127_776 ();
 DECAPx1_ASAP7_75t_R FILLER_127_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_788 ();
 DECAPx10_ASAP7_75t_R FILLER_127_801 ();
 DECAPx2_ASAP7_75t_R FILLER_127_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_829 ();
 DECAPx6_ASAP7_75t_R FILLER_127_845 ();
 DECAPx2_ASAP7_75t_R FILLER_127_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_865 ();
 DECAPx2_ASAP7_75t_R FILLER_127_873 ();
 DECAPx2_ASAP7_75t_R FILLER_127_891 ();
 FILLER_ASAP7_75t_R FILLER_127_903 ();
 DECAPx1_ASAP7_75t_R FILLER_127_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_917 ();
 DECAPx1_ASAP7_75t_R FILLER_127_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_930 ();
 DECAPx1_ASAP7_75t_R FILLER_127_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_982 ();
 DECAPx2_ASAP7_75t_R FILLER_127_995 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1068 ();
 FILLER_ASAP7_75t_R FILLER_127_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1082 ();
 FILLER_ASAP7_75t_R FILLER_127_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1097 ();
 DECAPx4_ASAP7_75t_R FILLER_127_1110 ();
 FILLER_ASAP7_75t_R FILLER_127_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1141 ();
 DECAPx4_ASAP7_75t_R FILLER_127_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1220 ();
 DECAPx6_ASAP7_75t_R FILLER_127_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1286 ();
 FILLER_ASAP7_75t_R FILLER_127_1298 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1307 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1313 ();
 DECAPx6_ASAP7_75t_R FILLER_127_1320 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1346 ();
 FILLER_ASAP7_75t_R FILLER_127_1358 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_128_8 ();
 DECAPx1_ASAP7_75t_R FILLER_128_18 ();
 DECAPx2_ASAP7_75t_R FILLER_128_25 ();
 FILLER_ASAP7_75t_R FILLER_128_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_37 ();
 DECAPx1_ASAP7_75t_R FILLER_128_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_145 ();
 FILLER_ASAP7_75t_R FILLER_128_152 ();
 DECAPx1_ASAP7_75t_R FILLER_128_157 ();
 DECAPx2_ASAP7_75t_R FILLER_128_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_176 ();
 DECAPx1_ASAP7_75t_R FILLER_128_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_195 ();
 DECAPx2_ASAP7_75t_R FILLER_128_210 ();
 FILLER_ASAP7_75t_R FILLER_128_216 ();
 FILLER_ASAP7_75t_R FILLER_128_224 ();
 DECAPx1_ASAP7_75t_R FILLER_128_232 ();
 DECAPx4_ASAP7_75t_R FILLER_128_242 ();
 DECAPx1_ASAP7_75t_R FILLER_128_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_274 ();
 DECAPx4_ASAP7_75t_R FILLER_128_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_321 ();
 DECAPx2_ASAP7_75t_R FILLER_128_329 ();
 DECAPx2_ASAP7_75t_R FILLER_128_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_355 ();
 DECAPx6_ASAP7_75t_R FILLER_128_370 ();
 FILLER_ASAP7_75t_R FILLER_128_392 ();
 DECAPx6_ASAP7_75t_R FILLER_128_408 ();
 DECAPx2_ASAP7_75t_R FILLER_128_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_428 ();
 DECAPx2_ASAP7_75t_R FILLER_128_447 ();
 FILLER_ASAP7_75t_R FILLER_128_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_455 ();
 DECAPx2_ASAP7_75t_R FILLER_128_472 ();
 FILLER_ASAP7_75t_R FILLER_128_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_480 ();
 FILLER_ASAP7_75t_R FILLER_128_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_516 ();
 DECAPx2_ASAP7_75t_R FILLER_128_532 ();
 FILLER_ASAP7_75t_R FILLER_128_538 ();
 DECAPx2_ASAP7_75t_R FILLER_128_547 ();
 FILLER_ASAP7_75t_R FILLER_128_553 ();
 DECAPx10_ASAP7_75t_R FILLER_128_561 ();
 DECAPx2_ASAP7_75t_R FILLER_128_590 ();
 FILLER_ASAP7_75t_R FILLER_128_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_601 ();
 DECAPx2_ASAP7_75t_R FILLER_128_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_614 ();
 FILLER_ASAP7_75t_R FILLER_128_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_620 ();
 DECAPx1_ASAP7_75t_R FILLER_128_628 ();
 DECAPx10_ASAP7_75t_R FILLER_128_656 ();
 DECAPx6_ASAP7_75t_R FILLER_128_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_701 ();
 DECAPx2_ASAP7_75t_R FILLER_128_728 ();
 DECAPx2_ASAP7_75t_R FILLER_128_767 ();
 FILLER_ASAP7_75t_R FILLER_128_773 ();
 DECAPx6_ASAP7_75t_R FILLER_128_782 ();
 FILLER_ASAP7_75t_R FILLER_128_796 ();
 FILLER_ASAP7_75t_R FILLER_128_807 ();
 DECAPx1_ASAP7_75t_R FILLER_128_816 ();
 FILLER_ASAP7_75t_R FILLER_128_847 ();
 DECAPx2_ASAP7_75t_R FILLER_128_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_882 ();
 DECAPx1_ASAP7_75t_R FILLER_128_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_903 ();
 DECAPx2_ASAP7_75t_R FILLER_128_916 ();
 DECAPx2_ASAP7_75t_R FILLER_128_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_934 ();
 DECAPx2_ASAP7_75t_R FILLER_128_942 ();
 DECAPx4_ASAP7_75t_R FILLER_128_958 ();
 FILLER_ASAP7_75t_R FILLER_128_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_970 ();
 FILLER_ASAP7_75t_R FILLER_128_985 ();
 DECAPx4_ASAP7_75t_R FILLER_128_993 ();
 FILLER_ASAP7_75t_R FILLER_128_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_128_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_128_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1086 ();
 DECAPx4_ASAP7_75t_R FILLER_128_1096 ();
 FILLER_ASAP7_75t_R FILLER_128_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1108 ();
 FILLER_ASAP7_75t_R FILLER_128_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1179 ();
 FILLER_ASAP7_75t_R FILLER_128_1206 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1226 ();
 FILLER_ASAP7_75t_R FILLER_128_1240 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1249 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1282 ();
 FILLER_ASAP7_75t_R FILLER_128_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_128_1297 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1329 ();
 DECAPx4_ASAP7_75t_R FILLER_128_1343 ();
 FILLER_ASAP7_75t_R FILLER_128_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1355 ();
 DECAPx4_ASAP7_75t_R FILLER_128_1362 ();
 FILLER_ASAP7_75t_R FILLER_128_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_129_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_79 ();
 DECAPx1_ASAP7_75t_R FILLER_129_89 ();
 DECAPx10_ASAP7_75t_R FILLER_129_96 ();
 DECAPx4_ASAP7_75t_R FILLER_129_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_128 ();
 DECAPx1_ASAP7_75t_R FILLER_129_135 ();
 DECAPx2_ASAP7_75t_R FILLER_129_165 ();
 FILLER_ASAP7_75t_R FILLER_129_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_173 ();
 DECAPx1_ASAP7_75t_R FILLER_129_194 ();
 DECAPx6_ASAP7_75t_R FILLER_129_204 ();
 DECAPx1_ASAP7_75t_R FILLER_129_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_222 ();
 FILLER_ASAP7_75t_R FILLER_129_231 ();
 DECAPx10_ASAP7_75t_R FILLER_129_265 ();
 DECAPx2_ASAP7_75t_R FILLER_129_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_293 ();
 DECAPx1_ASAP7_75t_R FILLER_129_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_318 ();
 DECAPx1_ASAP7_75t_R FILLER_129_327 ();
 DECAPx2_ASAP7_75t_R FILLER_129_337 ();
 FILLER_ASAP7_75t_R FILLER_129_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_345 ();
 FILLER_ASAP7_75t_R FILLER_129_352 ();
 DECAPx2_ASAP7_75t_R FILLER_129_366 ();
 FILLER_ASAP7_75t_R FILLER_129_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_398 ();
 DECAPx4_ASAP7_75t_R FILLER_129_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_417 ();
 DECAPx4_ASAP7_75t_R FILLER_129_428 ();
 FILLER_ASAP7_75t_R FILLER_129_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_446 ();
 DECAPx2_ASAP7_75t_R FILLER_129_481 ();
 DECAPx1_ASAP7_75t_R FILLER_129_494 ();
 DECAPx1_ASAP7_75t_R FILLER_129_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_509 ();
 DECAPx2_ASAP7_75t_R FILLER_129_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_532 ();
 DECAPx2_ASAP7_75t_R FILLER_129_551 ();
 DECAPx10_ASAP7_75t_R FILLER_129_573 ();
 DECAPx2_ASAP7_75t_R FILLER_129_595 ();
 FILLER_ASAP7_75t_R FILLER_129_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_603 ();
 DECAPx10_ASAP7_75t_R FILLER_129_611 ();
 DECAPx2_ASAP7_75t_R FILLER_129_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_639 ();
 DECAPx1_ASAP7_75t_R FILLER_129_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_694 ();
 DECAPx2_ASAP7_75t_R FILLER_129_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_708 ();
 DECAPx1_ASAP7_75t_R FILLER_129_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_738 ();
 DECAPx4_ASAP7_75t_R FILLER_129_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_758 ();
 DECAPx2_ASAP7_75t_R FILLER_129_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_792 ();
 FILLER_ASAP7_75t_R FILLER_129_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_807 ();
 DECAPx4_ASAP7_75t_R FILLER_129_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_835 ();
 DECAPx1_ASAP7_75t_R FILLER_129_844 ();
 DECAPx2_ASAP7_75t_R FILLER_129_855 ();
 FILLER_ASAP7_75t_R FILLER_129_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_863 ();
 DECAPx1_ASAP7_75t_R FILLER_129_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_880 ();
 DECAPx6_ASAP7_75t_R FILLER_129_893 ();
 DECAPx4_ASAP7_75t_R FILLER_129_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_923 ();
 FILLER_ASAP7_75t_R FILLER_129_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_934 ();
 DECAPx6_ASAP7_75t_R FILLER_129_942 ();
 DECAPx1_ASAP7_75t_R FILLER_129_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_960 ();
 DECAPx2_ASAP7_75t_R FILLER_129_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_998 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1030 ();
 FILLER_ASAP7_75t_R FILLER_129_1036 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_129_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_129_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1207 ();
 FILLER_ASAP7_75t_R FILLER_129_1213 ();
 FILLER_ASAP7_75t_R FILLER_129_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1239 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1250 ();
 FILLER_ASAP7_75t_R FILLER_129_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1272 ();
 FILLER_ASAP7_75t_R FILLER_129_1278 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1286 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1303 ();
 FILLER_ASAP7_75t_R FILLER_129_1314 ();
 FILLER_ASAP7_75t_R FILLER_129_1326 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1342 ();
 FILLER_ASAP7_75t_R FILLER_129_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1354 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_18 ();
 DECAPx10_ASAP7_75t_R FILLER_130_25 ();
 DECAPx2_ASAP7_75t_R FILLER_130_47 ();
 DECAPx2_ASAP7_75t_R FILLER_130_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_62 ();
 DECAPx10_ASAP7_75t_R FILLER_130_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_88 ();
 DECAPx10_ASAP7_75t_R FILLER_130_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_117 ();
 DECAPx1_ASAP7_75t_R FILLER_130_122 ();
 DECAPx4_ASAP7_75t_R FILLER_130_132 ();
 DECAPx6_ASAP7_75t_R FILLER_130_149 ();
 FILLER_ASAP7_75t_R FILLER_130_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_172 ();
 DECAPx4_ASAP7_75t_R FILLER_130_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_197 ();
 DECAPx4_ASAP7_75t_R FILLER_130_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_214 ();
 FILLER_ASAP7_75t_R FILLER_130_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_231 ();
 DECAPx6_ASAP7_75t_R FILLER_130_238 ();
 FILLER_ASAP7_75t_R FILLER_130_252 ();
 DECAPx2_ASAP7_75t_R FILLER_130_262 ();
 DECAPx1_ASAP7_75t_R FILLER_130_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_278 ();
 DECAPx2_ASAP7_75t_R FILLER_130_291 ();
 FILLER_ASAP7_75t_R FILLER_130_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_299 ();
 DECAPx1_ASAP7_75t_R FILLER_130_306 ();
 DECAPx10_ASAP7_75t_R FILLER_130_332 ();
 DECAPx2_ASAP7_75t_R FILLER_130_354 ();
 FILLER_ASAP7_75t_R FILLER_130_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_381 ();
 DECAPx1_ASAP7_75t_R FILLER_130_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_398 ();
 DECAPx4_ASAP7_75t_R FILLER_130_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_415 ();
 DECAPx2_ASAP7_75t_R FILLER_130_426 ();
 DECAPx6_ASAP7_75t_R FILLER_130_444 ();
 DECAPx1_ASAP7_75t_R FILLER_130_458 ();
 DECAPx4_ASAP7_75t_R FILLER_130_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_474 ();
 DECAPx1_ASAP7_75t_R FILLER_130_485 ();
 FILLER_ASAP7_75t_R FILLER_130_495 ();
 FILLER_ASAP7_75t_R FILLER_130_503 ();
 DECAPx4_ASAP7_75t_R FILLER_130_511 ();
 FILLER_ASAP7_75t_R FILLER_130_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_529 ();
 DECAPx1_ASAP7_75t_R FILLER_130_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_556 ();
 DECAPx6_ASAP7_75t_R FILLER_130_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_603 ();
 DECAPx4_ASAP7_75t_R FILLER_130_630 ();
 FILLER_ASAP7_75t_R FILLER_130_640 ();
 DECAPx4_ASAP7_75t_R FILLER_130_655 ();
 DECAPx1_ASAP7_75t_R FILLER_130_672 ();
 DECAPx4_ASAP7_75t_R FILLER_130_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_696 ();
 FILLER_ASAP7_75t_R FILLER_130_715 ();
 DECAPx6_ASAP7_75t_R FILLER_130_738 ();
 DECAPx10_ASAP7_75t_R FILLER_130_755 ();
 DECAPx2_ASAP7_75t_R FILLER_130_792 ();
 FILLER_ASAP7_75t_R FILLER_130_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_812 ();
 DECAPx1_ASAP7_75t_R FILLER_130_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_829 ();
 DECAPx4_ASAP7_75t_R FILLER_130_836 ();
 FILLER_ASAP7_75t_R FILLER_130_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_848 ();
 DECAPx2_ASAP7_75t_R FILLER_130_855 ();
 FILLER_ASAP7_75t_R FILLER_130_861 ();
 DECAPx4_ASAP7_75t_R FILLER_130_872 ();
 FILLER_ASAP7_75t_R FILLER_130_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_884 ();
 DECAPx6_ASAP7_75t_R FILLER_130_888 ();
 DECAPx1_ASAP7_75t_R FILLER_130_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_906 ();
 DECAPx10_ASAP7_75t_R FILLER_130_917 ();
 DECAPx6_ASAP7_75t_R FILLER_130_939 ();
 FILLER_ASAP7_75t_R FILLER_130_953 ();
 DECAPx6_ASAP7_75t_R FILLER_130_965 ();
 FILLER_ASAP7_75t_R FILLER_130_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_981 ();
 FILLER_ASAP7_75t_R FILLER_130_992 ();
 DECAPx4_ASAP7_75t_R FILLER_130_1000 ();
 FILLER_ASAP7_75t_R FILLER_130_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1048 ();
 FILLER_ASAP7_75t_R FILLER_130_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1081 ();
 FILLER_ASAP7_75t_R FILLER_130_1087 ();
 DECAPx4_ASAP7_75t_R FILLER_130_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1111 ();
 DECAPx4_ASAP7_75t_R FILLER_130_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1162 ();
 DECAPx4_ASAP7_75t_R FILLER_130_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1227 ();
 FILLER_ASAP7_75t_R FILLER_130_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1236 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1249 ();
 FILLER_ASAP7_75t_R FILLER_130_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1308 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1331 ();
 FILLER_ASAP7_75t_R FILLER_130_1343 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_131_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_45 ();
 DECAPx10_ASAP7_75t_R FILLER_131_52 ();
 DECAPx2_ASAP7_75t_R FILLER_131_74 ();
 FILLER_ASAP7_75t_R FILLER_131_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_82 ();
 FILLER_ASAP7_75t_R FILLER_131_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_117 ();
 DECAPx1_ASAP7_75t_R FILLER_131_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_151 ();
 FILLER_ASAP7_75t_R FILLER_131_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_172 ();
 FILLER_ASAP7_75t_R FILLER_131_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_197 ();
 DECAPx1_ASAP7_75t_R FILLER_131_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_214 ();
 DECAPx4_ASAP7_75t_R FILLER_131_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_245 ();
 FILLER_ASAP7_75t_R FILLER_131_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_260 ();
 FILLER_ASAP7_75t_R FILLER_131_269 ();
 FILLER_ASAP7_75t_R FILLER_131_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_279 ();
 DECAPx4_ASAP7_75t_R FILLER_131_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_313 ();
 DECAPx4_ASAP7_75t_R FILLER_131_326 ();
 FILLER_ASAP7_75t_R FILLER_131_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_346 ();
 DECAPx4_ASAP7_75t_R FILLER_131_353 ();
 FILLER_ASAP7_75t_R FILLER_131_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_365 ();
 DECAPx2_ASAP7_75t_R FILLER_131_374 ();
 DECAPx10_ASAP7_75t_R FILLER_131_388 ();
 FILLER_ASAP7_75t_R FILLER_131_410 ();
 DECAPx2_ASAP7_75t_R FILLER_131_422 ();
 DECAPx1_ASAP7_75t_R FILLER_131_436 ();
 DECAPx6_ASAP7_75t_R FILLER_131_448 ();
 FILLER_ASAP7_75t_R FILLER_131_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_464 ();
 FILLER_ASAP7_75t_R FILLER_131_483 ();
 DECAPx1_ASAP7_75t_R FILLER_131_493 ();
 DECAPx10_ASAP7_75t_R FILLER_131_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_535 ();
 DECAPx2_ASAP7_75t_R FILLER_131_548 ();
 DECAPx1_ASAP7_75t_R FILLER_131_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_577 ();
 DECAPx1_ASAP7_75t_R FILLER_131_604 ();
 DECAPx1_ASAP7_75t_R FILLER_131_614 ();
 DECAPx2_ASAP7_75t_R FILLER_131_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_627 ();
 DECAPx10_ASAP7_75t_R FILLER_131_635 ();
 DECAPx2_ASAP7_75t_R FILLER_131_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_663 ();
 DECAPx2_ASAP7_75t_R FILLER_131_670 ();
 DECAPx2_ASAP7_75t_R FILLER_131_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_721 ();
 DECAPx10_ASAP7_75t_R FILLER_131_728 ();
 DECAPx1_ASAP7_75t_R FILLER_131_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_778 ();
 DECAPx4_ASAP7_75t_R FILLER_131_788 ();
 FILLER_ASAP7_75t_R FILLER_131_798 ();
 FILLER_ASAP7_75t_R FILLER_131_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_805 ();
 DECAPx2_ASAP7_75t_R FILLER_131_833 ();
 DECAPx6_ASAP7_75t_R FILLER_131_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_864 ();
 DECAPx4_ASAP7_75t_R FILLER_131_874 ();
 DECAPx1_ASAP7_75t_R FILLER_131_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_900 ();
 DECAPx2_ASAP7_75t_R FILLER_131_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_962 ();
 DECAPx2_ASAP7_75t_R FILLER_131_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_975 ();
 DECAPx2_ASAP7_75t_R FILLER_131_979 ();
 FILLER_ASAP7_75t_R FILLER_131_985 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1011 ();
 FILLER_ASAP7_75t_R FILLER_131_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1087 ();
 FILLER_ASAP7_75t_R FILLER_131_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1101 ();
 FILLER_ASAP7_75t_R FILLER_131_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1130 ();
 FILLER_ASAP7_75t_R FILLER_131_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_131_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1241 ();
 DECAPx4_ASAP7_75t_R FILLER_131_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1262 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_131_1295 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1320 ();
 FILLER_ASAP7_75t_R FILLER_131_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1336 ();
 FILLER_ASAP7_75t_R FILLER_131_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1345 ();
 FILLER_ASAP7_75t_R FILLER_131_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1385 ();
 FILLER_ASAP7_75t_R FILLER_132_8 ();
 FILLER_ASAP7_75t_R FILLER_132_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_28 ();
 DECAPx4_ASAP7_75t_R FILLER_132_32 ();
 FILLER_ASAP7_75t_R FILLER_132_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_74 ();
 DECAPx1_ASAP7_75t_R FILLER_132_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_85 ();
 FILLER_ASAP7_75t_R FILLER_132_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_121 ();
 DECAPx1_ASAP7_75t_R FILLER_132_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_132 ();
 DECAPx10_ASAP7_75t_R FILLER_132_136 ();
 FILLER_ASAP7_75t_R FILLER_132_158 ();
 DECAPx2_ASAP7_75t_R FILLER_132_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_186 ();
 DECAPx4_ASAP7_75t_R FILLER_132_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_213 ();
 DECAPx2_ASAP7_75t_R FILLER_132_234 ();
 FILLER_ASAP7_75t_R FILLER_132_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_242 ();
 FILLER_ASAP7_75t_R FILLER_132_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_259 ();
 DECAPx1_ASAP7_75t_R FILLER_132_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_270 ();
 DECAPx2_ASAP7_75t_R FILLER_132_285 ();
 FILLER_ASAP7_75t_R FILLER_132_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_301 ();
 DECAPx6_ASAP7_75t_R FILLER_132_316 ();
 DECAPx1_ASAP7_75t_R FILLER_132_350 ();
 DECAPx2_ASAP7_75t_R FILLER_132_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_387 ();
 DECAPx6_ASAP7_75t_R FILLER_132_394 ();
 FILLER_ASAP7_75t_R FILLER_132_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_428 ();
 DECAPx1_ASAP7_75t_R FILLER_132_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_441 ();
 DECAPx2_ASAP7_75t_R FILLER_132_456 ();
 DECAPx6_ASAP7_75t_R FILLER_132_464 ();
 FILLER_ASAP7_75t_R FILLER_132_478 ();
 DECAPx1_ASAP7_75t_R FILLER_132_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_505 ();
 DECAPx4_ASAP7_75t_R FILLER_132_516 ();
 FILLER_ASAP7_75t_R FILLER_132_526 ();
 FILLER_ASAP7_75t_R FILLER_132_534 ();
 DECAPx6_ASAP7_75t_R FILLER_132_542 ();
 FILLER_ASAP7_75t_R FILLER_132_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_574 ();
 FILLER_ASAP7_75t_R FILLER_132_591 ();
 DECAPx1_ASAP7_75t_R FILLER_132_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_623 ();
 DECAPx2_ASAP7_75t_R FILLER_132_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_671 ();
 FILLER_ASAP7_75t_R FILLER_132_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_680 ();
 DECAPx10_ASAP7_75t_R FILLER_132_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_709 ();
 DECAPx6_ASAP7_75t_R FILLER_132_713 ();
 FILLER_ASAP7_75t_R FILLER_132_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_729 ();
 DECAPx2_ASAP7_75t_R FILLER_132_739 ();
 FILLER_ASAP7_75t_R FILLER_132_745 ();
 FILLER_ASAP7_75t_R FILLER_132_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_768 ();
 DECAPx6_ASAP7_75t_R FILLER_132_779 ();
 DECAPx1_ASAP7_75t_R FILLER_132_793 ();
 DECAPx4_ASAP7_75t_R FILLER_132_803 ();
 DECAPx2_ASAP7_75t_R FILLER_132_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_870 ();
 FILLER_ASAP7_75t_R FILLER_132_880 ();
 DECAPx2_ASAP7_75t_R FILLER_132_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_903 ();
 DECAPx2_ASAP7_75t_R FILLER_132_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_926 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1008 ();
 FILLER_ASAP7_75t_R FILLER_132_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1096 ();
 FILLER_ASAP7_75t_R FILLER_132_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1117 ();
 DECAPx4_ASAP7_75t_R FILLER_132_1128 ();
 FILLER_ASAP7_75t_R FILLER_132_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_132_1154 ();
 FILLER_ASAP7_75t_R FILLER_132_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1214 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1236 ();
 FILLER_ASAP7_75t_R FILLER_132_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1244 ();
 DECAPx4_ASAP7_75t_R FILLER_132_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1273 ();
 FILLER_ASAP7_75t_R FILLER_132_1295 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1297 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1306 ();
 FILLER_ASAP7_75t_R FILLER_132_1312 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1330 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1336 ();
 FILLER_ASAP7_75t_R FILLER_132_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1351 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1388 ();
 FILLER_ASAP7_75t_R FILLER_133_28 ();
 DECAPx2_ASAP7_75t_R FILLER_133_36 ();
 FILLER_ASAP7_75t_R FILLER_133_42 ();
 DECAPx2_ASAP7_75t_R FILLER_133_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_56 ();
 DECAPx2_ASAP7_75t_R FILLER_133_60 ();
 DECAPx2_ASAP7_75t_R FILLER_133_92 ();
 FILLER_ASAP7_75t_R FILLER_133_101 ();
 DECAPx1_ASAP7_75t_R FILLER_133_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_116 ();
 DECAPx6_ASAP7_75t_R FILLER_133_127 ();
 FILLER_ASAP7_75t_R FILLER_133_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_150 ();
 DECAPx2_ASAP7_75t_R FILLER_133_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_172 ();
 DECAPx6_ASAP7_75t_R FILLER_133_179 ();
 FILLER_ASAP7_75t_R FILLER_133_193 ();
 DECAPx4_ASAP7_75t_R FILLER_133_201 ();
 FILLER_ASAP7_75t_R FILLER_133_211 ();
 DECAPx4_ASAP7_75t_R FILLER_133_233 ();
 DECAPx2_ASAP7_75t_R FILLER_133_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_255 ();
 DECAPx6_ASAP7_75t_R FILLER_133_262 ();
 DECAPx4_ASAP7_75t_R FILLER_133_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_300 ();
 DECAPx6_ASAP7_75t_R FILLER_133_307 ();
 DECAPx2_ASAP7_75t_R FILLER_133_321 ();
 DECAPx6_ASAP7_75t_R FILLER_133_349 ();
 FILLER_ASAP7_75t_R FILLER_133_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_365 ();
 DECAPx2_ASAP7_75t_R FILLER_133_372 ();
 DECAPx10_ASAP7_75t_R FILLER_133_400 ();
 DECAPx2_ASAP7_75t_R FILLER_133_422 ();
 DECAPx1_ASAP7_75t_R FILLER_133_440 ();
 FILLER_ASAP7_75t_R FILLER_133_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_452 ();
 DECAPx2_ASAP7_75t_R FILLER_133_479 ();
 FILLER_ASAP7_75t_R FILLER_133_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_487 ();
 DECAPx6_ASAP7_75t_R FILLER_133_494 ();
 FILLER_ASAP7_75t_R FILLER_133_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_510 ();
 FILLER_ASAP7_75t_R FILLER_133_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_529 ();
 DECAPx2_ASAP7_75t_R FILLER_133_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_550 ();
 DECAPx10_ASAP7_75t_R FILLER_133_557 ();
 DECAPx4_ASAP7_75t_R FILLER_133_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_606 ();
 DECAPx6_ASAP7_75t_R FILLER_133_610 ();
 DECAPx1_ASAP7_75t_R FILLER_133_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_670 ();
 DECAPx10_ASAP7_75t_R FILLER_133_686 ();
 DECAPx4_ASAP7_75t_R FILLER_133_708 ();
 FILLER_ASAP7_75t_R FILLER_133_726 ();
 DECAPx4_ASAP7_75t_R FILLER_133_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_753 ();
 DECAPx4_ASAP7_75t_R FILLER_133_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_788 ();
 DECAPx2_ASAP7_75t_R FILLER_133_805 ();
 DECAPx6_ASAP7_75t_R FILLER_133_823 ();
 FILLER_ASAP7_75t_R FILLER_133_837 ();
 FILLER_ASAP7_75t_R FILLER_133_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_861 ();
 FILLER_ASAP7_75t_R FILLER_133_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_884 ();
 DECAPx4_ASAP7_75t_R FILLER_133_894 ();
 FILLER_ASAP7_75t_R FILLER_133_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_906 ();
 DECAPx4_ASAP7_75t_R FILLER_133_914 ();
 DECAPx10_ASAP7_75t_R FILLER_133_926 ();
 DECAPx6_ASAP7_75t_R FILLER_133_948 ();
 DECAPx1_ASAP7_75t_R FILLER_133_962 ();
 DECAPx1_ASAP7_75t_R FILLER_133_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_976 ();
 DECAPx2_ASAP7_75t_R FILLER_133_989 ();
 DECAPx4_ASAP7_75t_R FILLER_133_1001 ();
 FILLER_ASAP7_75t_R FILLER_133_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1049 ();
 DECAPx4_ASAP7_75t_R FILLER_133_1071 ();
 FILLER_ASAP7_75t_R FILLER_133_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1114 ();
 DECAPx6_ASAP7_75t_R FILLER_133_1144 ();
 FILLER_ASAP7_75t_R FILLER_133_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1180 ();
 FILLER_ASAP7_75t_R FILLER_133_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1204 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1221 ();
 DECAPx4_ASAP7_75t_R FILLER_133_1238 ();
 FILLER_ASAP7_75t_R FILLER_133_1296 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1298 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1327 ();
 DECAPx4_ASAP7_75t_R FILLER_133_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1359 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1369 ();
 DECAPx1_ASAP7_75t_R FILLER_134_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_6 ();
 FILLER_ASAP7_75t_R FILLER_134_13 ();
 DECAPx1_ASAP7_75t_R FILLER_134_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_52 ();
 FILLER_ASAP7_75t_R FILLER_134_59 ();
 FILLER_ASAP7_75t_R FILLER_134_64 ();
 DECAPx1_ASAP7_75t_R FILLER_134_76 ();
 DECAPx10_ASAP7_75t_R FILLER_134_83 ();
 DECAPx1_ASAP7_75t_R FILLER_134_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_162 ();
 DECAPx6_ASAP7_75t_R FILLER_134_177 ();
 DECAPx1_ASAP7_75t_R FILLER_134_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_195 ();
 DECAPx2_ASAP7_75t_R FILLER_134_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_208 ();
 DECAPx6_ASAP7_75t_R FILLER_134_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_252 ();
 DECAPx2_ASAP7_75t_R FILLER_134_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_265 ();
 FILLER_ASAP7_75t_R FILLER_134_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_280 ();
 DECAPx6_ASAP7_75t_R FILLER_134_287 ();
 DECAPx1_ASAP7_75t_R FILLER_134_301 ();
 DECAPx1_ASAP7_75t_R FILLER_134_313 ();
 DECAPx1_ASAP7_75t_R FILLER_134_323 ();
 DECAPx6_ASAP7_75t_R FILLER_134_345 ();
 DECAPx2_ASAP7_75t_R FILLER_134_359 ();
 DECAPx4_ASAP7_75t_R FILLER_134_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_385 ();
 DECAPx2_ASAP7_75t_R FILLER_134_392 ();
 FILLER_ASAP7_75t_R FILLER_134_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_400 ();
 DECAPx1_ASAP7_75t_R FILLER_134_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_412 ();
 DECAPx2_ASAP7_75t_R FILLER_134_416 ();
 FILLER_ASAP7_75t_R FILLER_134_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_445 ();
 FILLER_ASAP7_75t_R FILLER_134_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_461 ();
 DECAPx1_ASAP7_75t_R FILLER_134_464 ();
 DECAPx4_ASAP7_75t_R FILLER_134_471 ();
 FILLER_ASAP7_75t_R FILLER_134_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_483 ();
 DECAPx6_ASAP7_75t_R FILLER_134_496 ();
 DECAPx1_ASAP7_75t_R FILLER_134_510 ();
 DECAPx2_ASAP7_75t_R FILLER_134_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_526 ();
 DECAPx2_ASAP7_75t_R FILLER_134_543 ();
 FILLER_ASAP7_75t_R FILLER_134_549 ();
 DECAPx10_ASAP7_75t_R FILLER_134_558 ();
 DECAPx6_ASAP7_75t_R FILLER_134_580 ();
 FILLER_ASAP7_75t_R FILLER_134_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_596 ();
 DECAPx10_ASAP7_75t_R FILLER_134_603 ();
 DECAPx4_ASAP7_75t_R FILLER_134_625 ();
 FILLER_ASAP7_75t_R FILLER_134_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_637 ();
 DECAPx10_ASAP7_75t_R FILLER_134_645 ();
 DECAPx2_ASAP7_75t_R FILLER_134_667 ();
 DECAPx1_ASAP7_75t_R FILLER_134_688 ();
 FILLER_ASAP7_75t_R FILLER_134_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_708 ();
 FILLER_ASAP7_75t_R FILLER_134_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_732 ();
 DECAPx6_ASAP7_75t_R FILLER_134_758 ();
 DECAPx2_ASAP7_75t_R FILLER_134_772 ();
 FILLER_ASAP7_75t_R FILLER_134_788 ();
 DECAPx4_ASAP7_75t_R FILLER_134_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_810 ();
 DECAPx2_ASAP7_75t_R FILLER_134_824 ();
 FILLER_ASAP7_75t_R FILLER_134_830 ();
 DECAPx2_ASAP7_75t_R FILLER_134_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_848 ();
 DECAPx4_ASAP7_75t_R FILLER_134_858 ();
 DECAPx2_ASAP7_75t_R FILLER_134_880 ();
 FILLER_ASAP7_75t_R FILLER_134_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_896 ();
 DECAPx10_ASAP7_75t_R FILLER_134_903 ();
 DECAPx4_ASAP7_75t_R FILLER_134_925 ();
 DECAPx4_ASAP7_75t_R FILLER_134_942 ();
 DECAPx10_ASAP7_75t_R FILLER_134_970 ();
 FILLER_ASAP7_75t_R FILLER_134_992 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1000 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1022 ();
 DECAPx1_ASAP7_75t_R FILLER_134_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1058 ();
 FILLER_ASAP7_75t_R FILLER_134_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1103 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1113 ();
 FILLER_ASAP7_75t_R FILLER_134_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1165 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1172 ();
 FILLER_ASAP7_75t_R FILLER_134_1182 ();
 FILLER_ASAP7_75t_R FILLER_134_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_134_1235 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1247 ();
 FILLER_ASAP7_75t_R FILLER_134_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1277 ();
 FILLER_ASAP7_75t_R FILLER_134_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1315 ();
 DECAPx1_ASAP7_75t_R FILLER_134_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1347 ();
 FILLER_ASAP7_75t_R FILLER_134_1356 ();
 FILLER_ASAP7_75t_R FILLER_134_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_134_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_135_2 ();
 FILLER_ASAP7_75t_R FILLER_135_12 ();
 DECAPx1_ASAP7_75t_R FILLER_135_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_36 ();
 DECAPx2_ASAP7_75t_R FILLER_135_40 ();
 DECAPx1_ASAP7_75t_R FILLER_135_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_76 ();
 DECAPx1_ASAP7_75t_R FILLER_135_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_107 ();
 FILLER_ASAP7_75t_R FILLER_135_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_128 ();
 DECAPx2_ASAP7_75t_R FILLER_135_132 ();
 FILLER_ASAP7_75t_R FILLER_135_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_144 ();
 DECAPx4_ASAP7_75t_R FILLER_135_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_161 ();
 DECAPx1_ASAP7_75t_R FILLER_135_182 ();
 DECAPx2_ASAP7_75t_R FILLER_135_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_218 ();
 DECAPx1_ASAP7_75t_R FILLER_135_227 ();
 DECAPx2_ASAP7_75t_R FILLER_135_238 ();
 FILLER_ASAP7_75t_R FILLER_135_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_246 ();
 DECAPx1_ASAP7_75t_R FILLER_135_250 ();
 DECAPx1_ASAP7_75t_R FILLER_135_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_266 ();
 FILLER_ASAP7_75t_R FILLER_135_273 ();
 DECAPx1_ASAP7_75t_R FILLER_135_297 ();
 DECAPx10_ASAP7_75t_R FILLER_135_323 ();
 FILLER_ASAP7_75t_R FILLER_135_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_353 ();
 DECAPx10_ASAP7_75t_R FILLER_135_366 ();
 DECAPx4_ASAP7_75t_R FILLER_135_388 ();
 DECAPx1_ASAP7_75t_R FILLER_135_424 ();
 DECAPx1_ASAP7_75t_R FILLER_135_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_438 ();
 DECAPx2_ASAP7_75t_R FILLER_135_447 ();
 FILLER_ASAP7_75t_R FILLER_135_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_455 ();
 FILLER_ASAP7_75t_R FILLER_135_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_484 ();
 FILLER_ASAP7_75t_R FILLER_135_493 ();
 DECAPx2_ASAP7_75t_R FILLER_135_502 ();
 DECAPx1_ASAP7_75t_R FILLER_135_516 ();
 DECAPx1_ASAP7_75t_R FILLER_135_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_531 ();
 FILLER_ASAP7_75t_R FILLER_135_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_540 ();
 DECAPx1_ASAP7_75t_R FILLER_135_548 ();
 DECAPx2_ASAP7_75t_R FILLER_135_578 ();
 FILLER_ASAP7_75t_R FILLER_135_584 ();
 DECAPx2_ASAP7_75t_R FILLER_135_615 ();
 FILLER_ASAP7_75t_R FILLER_135_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_623 ();
 DECAPx1_ASAP7_75t_R FILLER_135_638 ();
 DECAPx6_ASAP7_75t_R FILLER_135_656 ();
 DECAPx1_ASAP7_75t_R FILLER_135_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_674 ();
 DECAPx10_ASAP7_75t_R FILLER_135_699 ();
 DECAPx10_ASAP7_75t_R FILLER_135_731 ();
 DECAPx2_ASAP7_75t_R FILLER_135_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_763 ();
 FILLER_ASAP7_75t_R FILLER_135_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_769 ();
 DECAPx10_ASAP7_75t_R FILLER_135_786 ();
 DECAPx2_ASAP7_75t_R FILLER_135_808 ();
 DECAPx10_ASAP7_75t_R FILLER_135_821 ();
 FILLER_ASAP7_75t_R FILLER_135_843 ();
 DECAPx2_ASAP7_75t_R FILLER_135_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_863 ();
 DECAPx6_ASAP7_75t_R FILLER_135_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_903 ();
 DECAPx1_ASAP7_75t_R FILLER_135_920 ();
 FILLER_ASAP7_75t_R FILLER_135_933 ();
 DECAPx2_ASAP7_75t_R FILLER_135_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_951 ();
 DECAPx2_ASAP7_75t_R FILLER_135_968 ();
 FILLER_ASAP7_75t_R FILLER_135_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_986 ();
 FILLER_ASAP7_75t_R FILLER_135_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1034 ();
 FILLER_ASAP7_75t_R FILLER_135_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1086 ();
 FILLER_ASAP7_75t_R FILLER_135_1092 ();
 DECAPx4_ASAP7_75t_R FILLER_135_1102 ();
 FILLER_ASAP7_75t_R FILLER_135_1112 ();
 DECAPx4_ASAP7_75t_R FILLER_135_1126 ();
 FILLER_ASAP7_75t_R FILLER_135_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1138 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1156 ();
 FILLER_ASAP7_75t_R FILLER_135_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1213 ();
 FILLER_ASAP7_75t_R FILLER_135_1219 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1233 ();
 FILLER_ASAP7_75t_R FILLER_135_1256 ();
 DECAPx4_ASAP7_75t_R FILLER_135_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1298 ();
 FILLER_ASAP7_75t_R FILLER_135_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_136_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_6 ();
 DECAPx4_ASAP7_75t_R FILLER_136_37 ();
 FILLER_ASAP7_75t_R FILLER_136_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_55 ();
 DECAPx6_ASAP7_75t_R FILLER_136_62 ();
 FILLER_ASAP7_75t_R FILLER_136_76 ();
 DECAPx10_ASAP7_75t_R FILLER_136_116 ();
 DECAPx1_ASAP7_75t_R FILLER_136_138 ();
 DECAPx1_ASAP7_75t_R FILLER_136_158 ();
 DECAPx1_ASAP7_75t_R FILLER_136_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_180 ();
 FILLER_ASAP7_75t_R FILLER_136_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_189 ();
 DECAPx1_ASAP7_75t_R FILLER_136_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_204 ();
 DECAPx2_ASAP7_75t_R FILLER_136_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_217 ();
 DECAPx2_ASAP7_75t_R FILLER_136_224 ();
 FILLER_ASAP7_75t_R FILLER_136_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_232 ();
 DECAPx6_ASAP7_75t_R FILLER_136_259 ();
 FILLER_ASAP7_75t_R FILLER_136_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_275 ();
 FILLER_ASAP7_75t_R FILLER_136_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_284 ();
 DECAPx4_ASAP7_75t_R FILLER_136_298 ();
 DECAPx2_ASAP7_75t_R FILLER_136_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_384 ();
 DECAPx2_ASAP7_75t_R FILLER_136_391 ();
 DECAPx2_ASAP7_75t_R FILLER_136_409 ();
 DECAPx2_ASAP7_75t_R FILLER_136_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_427 ();
 FILLER_ASAP7_75t_R FILLER_136_436 ();
 DECAPx4_ASAP7_75t_R FILLER_136_452 ();
 DECAPx2_ASAP7_75t_R FILLER_136_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_493 ();
 DECAPx1_ASAP7_75t_R FILLER_136_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_624 ();
 DECAPx4_ASAP7_75t_R FILLER_136_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_659 ();
 FILLER_ASAP7_75t_R FILLER_136_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_692 ();
 DECAPx6_ASAP7_75t_R FILLER_136_702 ();
 FILLER_ASAP7_75t_R FILLER_136_716 ();
 DECAPx2_ASAP7_75t_R FILLER_136_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_752 ();
 DECAPx2_ASAP7_75t_R FILLER_136_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_786 ();
 FILLER_ASAP7_75t_R FILLER_136_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_809 ();
 DECAPx1_ASAP7_75t_R FILLER_136_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_830 ();
 DECAPx1_ASAP7_75t_R FILLER_136_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_845 ();
 DECAPx1_ASAP7_75t_R FILLER_136_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_887 ();
 DECAPx1_ASAP7_75t_R FILLER_136_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_901 ();
 DECAPx1_ASAP7_75t_R FILLER_136_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_945 ();
 DECAPx2_ASAP7_75t_R FILLER_136_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_992 ();
 FILLER_ASAP7_75t_R FILLER_136_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1008 ();
 FILLER_ASAP7_75t_R FILLER_136_1019 ();
 FILLER_ASAP7_75t_R FILLER_136_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_136_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1093 ();
 FILLER_ASAP7_75t_R FILLER_136_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1155 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_136_1188 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1214 ();
 DECAPx6_ASAP7_75t_R FILLER_136_1221 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_136_1247 ();
 FILLER_ASAP7_75t_R FILLER_136_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_136_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_136_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_137_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_14 ();
 DECAPx6_ASAP7_75t_R FILLER_137_24 ();
 FILLER_ASAP7_75t_R FILLER_137_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_40 ();
 DECAPx2_ASAP7_75t_R FILLER_137_83 ();
 FILLER_ASAP7_75t_R FILLER_137_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_91 ();
 DECAPx1_ASAP7_75t_R FILLER_137_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_114 ();
 DECAPx2_ASAP7_75t_R FILLER_137_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_127 ();
 DECAPx2_ASAP7_75t_R FILLER_137_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_137 ();
 DECAPx1_ASAP7_75t_R FILLER_137_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_168 ();
 DECAPx10_ASAP7_75t_R FILLER_137_183 ();
 DECAPx6_ASAP7_75t_R FILLER_137_213 ();
 DECAPx2_ASAP7_75t_R FILLER_137_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_233 ();
 DECAPx4_ASAP7_75t_R FILLER_137_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_250 ();
 DECAPx2_ASAP7_75t_R FILLER_137_257 ();
 FILLER_ASAP7_75t_R FILLER_137_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_265 ();
 DECAPx1_ASAP7_75t_R FILLER_137_276 ();
 DECAPx1_ASAP7_75t_R FILLER_137_306 ();
 DECAPx2_ASAP7_75t_R FILLER_137_317 ();
 FILLER_ASAP7_75t_R FILLER_137_323 ();
 FILLER_ASAP7_75t_R FILLER_137_333 ();
 DECAPx2_ASAP7_75t_R FILLER_137_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_349 ();
 FILLER_ASAP7_75t_R FILLER_137_356 ();
 DECAPx2_ASAP7_75t_R FILLER_137_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_371 ();
 FILLER_ASAP7_75t_R FILLER_137_375 ();
 DECAPx4_ASAP7_75t_R FILLER_137_403 ();
 FILLER_ASAP7_75t_R FILLER_137_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_415 ();
 FILLER_ASAP7_75t_R FILLER_137_430 ();
 DECAPx2_ASAP7_75t_R FILLER_137_450 ();
 FILLER_ASAP7_75t_R FILLER_137_456 ();
 DECAPx10_ASAP7_75t_R FILLER_137_465 ();
 DECAPx4_ASAP7_75t_R FILLER_137_487 ();
 FILLER_ASAP7_75t_R FILLER_137_497 ();
 DECAPx1_ASAP7_75t_R FILLER_137_505 ();
 DECAPx2_ASAP7_75t_R FILLER_137_512 ();
 FILLER_ASAP7_75t_R FILLER_137_518 ();
 DECAPx2_ASAP7_75t_R FILLER_137_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_533 ();
 DECAPx2_ASAP7_75t_R FILLER_137_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_543 ();
 DECAPx2_ASAP7_75t_R FILLER_137_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_563 ();
 DECAPx6_ASAP7_75t_R FILLER_137_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_584 ();
 FILLER_ASAP7_75t_R FILLER_137_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_594 ();
 DECAPx10_ASAP7_75t_R FILLER_137_602 ();
 DECAPx6_ASAP7_75t_R FILLER_137_624 ();
 DECAPx1_ASAP7_75t_R FILLER_137_638 ();
 DECAPx6_ASAP7_75t_R FILLER_137_659 ();
 FILLER_ASAP7_75t_R FILLER_137_688 ();
 DECAPx1_ASAP7_75t_R FILLER_137_698 ();
 DECAPx4_ASAP7_75t_R FILLER_137_714 ();
 FILLER_ASAP7_75t_R FILLER_137_724 ();
 FILLER_ASAP7_75t_R FILLER_137_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_753 ();
 DECAPx4_ASAP7_75t_R FILLER_137_777 ();
 FILLER_ASAP7_75t_R FILLER_137_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_789 ();
 FILLER_ASAP7_75t_R FILLER_137_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_813 ();
 DECAPx2_ASAP7_75t_R FILLER_137_820 ();
 FILLER_ASAP7_75t_R FILLER_137_826 ();
 DECAPx2_ASAP7_75t_R FILLER_137_842 ();
 FILLER_ASAP7_75t_R FILLER_137_848 ();
 DECAPx1_ASAP7_75t_R FILLER_137_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_860 ();
 DECAPx1_ASAP7_75t_R FILLER_137_882 ();
 DECAPx2_ASAP7_75t_R FILLER_137_898 ();
 FILLER_ASAP7_75t_R FILLER_137_904 ();
 DECAPx2_ASAP7_75t_R FILLER_137_916 ();
 FILLER_ASAP7_75t_R FILLER_137_922 ();
 DECAPx2_ASAP7_75t_R FILLER_137_926 ();
 DECAPx4_ASAP7_75t_R FILLER_137_944 ();
 FILLER_ASAP7_75t_R FILLER_137_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_964 ();
 DECAPx4_ASAP7_75t_R FILLER_137_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_983 ();
 DECAPx2_ASAP7_75t_R FILLER_137_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1000 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1031 ();
 FILLER_ASAP7_75t_R FILLER_137_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1048 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1055 ();
 FILLER_ASAP7_75t_R FILLER_137_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1094 ();
 FILLER_ASAP7_75t_R FILLER_137_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_137_1146 ();
 FILLER_ASAP7_75t_R FILLER_137_1160 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1194 ();
 FILLER_ASAP7_75t_R FILLER_137_1200 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1225 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1234 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1268 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1282 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1296 ();
 FILLER_ASAP7_75t_R FILLER_137_1309 ();
 DECAPx6_ASAP7_75t_R FILLER_137_1325 ();
 FILLER_ASAP7_75t_R FILLER_137_1339 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1341 ();
 FILLER_ASAP7_75t_R FILLER_137_1349 ();
 DECAPx6_ASAP7_75t_R FILLER_137_1361 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_32 ();
 DECAPx1_ASAP7_75t_R FILLER_138_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_67 ();
 DECAPx1_ASAP7_75t_R FILLER_138_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_75 ();
 DECAPx6_ASAP7_75t_R FILLER_138_85 ();
 DECAPx1_ASAP7_75t_R FILLER_138_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_103 ();
 FILLER_ASAP7_75t_R FILLER_138_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_150 ();
 DECAPx4_ASAP7_75t_R FILLER_138_157 ();
 FILLER_ASAP7_75t_R FILLER_138_173 ();
 DECAPx6_ASAP7_75t_R FILLER_138_182 ();
 DECAPx2_ASAP7_75t_R FILLER_138_196 ();
 FILLER_ASAP7_75t_R FILLER_138_216 ();
 DECAPx2_ASAP7_75t_R FILLER_138_232 ();
 FILLER_ASAP7_75t_R FILLER_138_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_240 ();
 DECAPx2_ASAP7_75t_R FILLER_138_261 ();
 FILLER_ASAP7_75t_R FILLER_138_267 ();
 DECAPx6_ASAP7_75t_R FILLER_138_279 ();
 FILLER_ASAP7_75t_R FILLER_138_293 ();
 DECAPx2_ASAP7_75t_R FILLER_138_298 ();
 FILLER_ASAP7_75t_R FILLER_138_304 ();
 DECAPx1_ASAP7_75t_R FILLER_138_332 ();
 DECAPx2_ASAP7_75t_R FILLER_138_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_356 ();
 DECAPx6_ASAP7_75t_R FILLER_138_364 ();
 FILLER_ASAP7_75t_R FILLER_138_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_380 ();
 FILLER_ASAP7_75t_R FILLER_138_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_390 ();
 FILLER_ASAP7_75t_R FILLER_138_394 ();
 DECAPx2_ASAP7_75t_R FILLER_138_430 ();
 FILLER_ASAP7_75t_R FILLER_138_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_438 ();
 FILLER_ASAP7_75t_R FILLER_138_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_454 ();
 DECAPx1_ASAP7_75t_R FILLER_138_470 ();
 DECAPx2_ASAP7_75t_R FILLER_138_487 ();
 FILLER_ASAP7_75t_R FILLER_138_493 ();
 FILLER_ASAP7_75t_R FILLER_138_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_500 ();
 DECAPx6_ASAP7_75t_R FILLER_138_505 ();
 FILLER_ASAP7_75t_R FILLER_138_519 ();
 DECAPx10_ASAP7_75t_R FILLER_138_527 ();
 DECAPx1_ASAP7_75t_R FILLER_138_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_553 ();
 DECAPx6_ASAP7_75t_R FILLER_138_560 ();
 DECAPx2_ASAP7_75t_R FILLER_138_577 ();
 FILLER_ASAP7_75t_R FILLER_138_583 ();
 DECAPx4_ASAP7_75t_R FILLER_138_591 ();
 FILLER_ASAP7_75t_R FILLER_138_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_603 ();
 DECAPx2_ASAP7_75t_R FILLER_138_608 ();
 DECAPx1_ASAP7_75t_R FILLER_138_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_625 ();
 DECAPx10_ASAP7_75t_R FILLER_138_644 ();
 DECAPx1_ASAP7_75t_R FILLER_138_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_680 ();
 DECAPx6_ASAP7_75t_R FILLER_138_684 ();
 FILLER_ASAP7_75t_R FILLER_138_698 ();
 DECAPx6_ASAP7_75t_R FILLER_138_737 ();
 DECAPx2_ASAP7_75t_R FILLER_138_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_757 ();
 DECAPx2_ASAP7_75t_R FILLER_138_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_774 ();
 DECAPx1_ASAP7_75t_R FILLER_138_785 ();
 DECAPx2_ASAP7_75t_R FILLER_138_805 ();
 DECAPx1_ASAP7_75t_R FILLER_138_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_837 ();
 FILLER_ASAP7_75t_R FILLER_138_850 ();
 DECAPx10_ASAP7_75t_R FILLER_138_858 ();
 DECAPx2_ASAP7_75t_R FILLER_138_880 ();
 FILLER_ASAP7_75t_R FILLER_138_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_888 ();
 DECAPx6_ASAP7_75t_R FILLER_138_897 ();
 DECAPx1_ASAP7_75t_R FILLER_138_911 ();
 DECAPx2_ASAP7_75t_R FILLER_138_921 ();
 DECAPx1_ASAP7_75t_R FILLER_138_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_937 ();
 DECAPx6_ASAP7_75t_R FILLER_138_944 ();
 DECAPx1_ASAP7_75t_R FILLER_138_964 ();
 DECAPx10_ASAP7_75t_R FILLER_138_974 ();
 DECAPx6_ASAP7_75t_R FILLER_138_996 ();
 FILLER_ASAP7_75t_R FILLER_138_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1033 ();
 FILLER_ASAP7_75t_R FILLER_138_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1079 ();
 FILLER_ASAP7_75t_R FILLER_138_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1098 ();
 FILLER_ASAP7_75t_R FILLER_138_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1128 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1176 ();
 FILLER_ASAP7_75t_R FILLER_138_1185 ();
 FILLER_ASAP7_75t_R FILLER_138_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1222 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1249 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1272 ();
 FILLER_ASAP7_75t_R FILLER_138_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1284 ();
 FILLER_ASAP7_75t_R FILLER_138_1315 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1333 ();
 FILLER_ASAP7_75t_R FILLER_138_1351 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1363 ();
 FILLER_ASAP7_75t_R FILLER_138_1369 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1377 ();
 FILLER_ASAP7_75t_R FILLER_138_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_139_2 ();
 FILLER_ASAP7_75t_R FILLER_139_8 ();
 DECAPx6_ASAP7_75t_R FILLER_139_19 ();
 DECAPx1_ASAP7_75t_R FILLER_139_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_37 ();
 DECAPx1_ASAP7_75t_R FILLER_139_44 ();
 DECAPx6_ASAP7_75t_R FILLER_139_51 ();
 FILLER_ASAP7_75t_R FILLER_139_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_67 ();
 DECAPx4_ASAP7_75t_R FILLER_139_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_104 ();
 DECAPx2_ASAP7_75t_R FILLER_139_111 ();
 FILLER_ASAP7_75t_R FILLER_139_117 ();
 DECAPx4_ASAP7_75t_R FILLER_139_122 ();
 FILLER_ASAP7_75t_R FILLER_139_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_134 ();
 DECAPx4_ASAP7_75t_R FILLER_139_163 ();
 FILLER_ASAP7_75t_R FILLER_139_173 ();
 DECAPx2_ASAP7_75t_R FILLER_139_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_213 ();
 DECAPx2_ASAP7_75t_R FILLER_139_228 ();
 FILLER_ASAP7_75t_R FILLER_139_234 ();
 DECAPx2_ASAP7_75t_R FILLER_139_260 ();
 DECAPx1_ASAP7_75t_R FILLER_139_284 ();
 DECAPx1_ASAP7_75t_R FILLER_139_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_295 ();
 DECAPx2_ASAP7_75t_R FILLER_139_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_315 ();
 DECAPx1_ASAP7_75t_R FILLER_139_325 ();
 DECAPx2_ASAP7_75t_R FILLER_139_349 ();
 FILLER_ASAP7_75t_R FILLER_139_355 ();
 DECAPx1_ASAP7_75t_R FILLER_139_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_387 ();
 DECAPx1_ASAP7_75t_R FILLER_139_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_399 ();
 DECAPx2_ASAP7_75t_R FILLER_139_408 ();
 FILLER_ASAP7_75t_R FILLER_139_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_416 ();
 FILLER_ASAP7_75t_R FILLER_139_453 ();
 DECAPx2_ASAP7_75t_R FILLER_139_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_520 ();
 DECAPx2_ASAP7_75t_R FILLER_139_543 ();
 FILLER_ASAP7_75t_R FILLER_139_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_551 ();
 DECAPx1_ASAP7_75t_R FILLER_139_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_614 ();
 DECAPx2_ASAP7_75t_R FILLER_139_641 ();
 DECAPx6_ASAP7_75t_R FILLER_139_688 ();
 FILLER_ASAP7_75t_R FILLER_139_702 ();
 DECAPx2_ASAP7_75t_R FILLER_139_710 ();
 FILLER_ASAP7_75t_R FILLER_139_716 ();
 DECAPx6_ASAP7_75t_R FILLER_139_731 ();
 DECAPx10_ASAP7_75t_R FILLER_139_753 ();
 DECAPx1_ASAP7_75t_R FILLER_139_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_779 ();
 DECAPx4_ASAP7_75t_R FILLER_139_788 ();
 DECAPx4_ASAP7_75t_R FILLER_139_808 ();
 FILLER_ASAP7_75t_R FILLER_139_818 ();
 DECAPx2_ASAP7_75t_R FILLER_139_825 ();
 FILLER_ASAP7_75t_R FILLER_139_831 ();
 DECAPx10_ASAP7_75t_R FILLER_139_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_873 ();
 DECAPx2_ASAP7_75t_R FILLER_139_889 ();
 FILLER_ASAP7_75t_R FILLER_139_895 ();
 DECAPx2_ASAP7_75t_R FILLER_139_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_913 ();
 DECAPx1_ASAP7_75t_R FILLER_139_920 ();
 DECAPx2_ASAP7_75t_R FILLER_139_926 ();
 DECAPx6_ASAP7_75t_R FILLER_139_942 ();
 DECAPx1_ASAP7_75t_R FILLER_139_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_960 ();
 DECAPx4_ASAP7_75t_R FILLER_139_971 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1002 ();
 FILLER_ASAP7_75t_R FILLER_139_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1079 ();
 FILLER_ASAP7_75t_R FILLER_139_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1127 ();
 FILLER_ASAP7_75t_R FILLER_139_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1151 ();
 FILLER_ASAP7_75t_R FILLER_139_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1173 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1196 ();
 FILLER_ASAP7_75t_R FILLER_139_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1214 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1244 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1272 ();
 FILLER_ASAP7_75t_R FILLER_139_1286 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1300 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1307 ();
 FILLER_ASAP7_75t_R FILLER_139_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1345 ();
 FILLER_ASAP7_75t_R FILLER_139_1352 ();
 FILLER_ASAP7_75t_R FILLER_139_1384 ();
 DECAPx4_ASAP7_75t_R FILLER_140_2 ();
 FILLER_ASAP7_75t_R FILLER_140_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_14 ();
 DECAPx2_ASAP7_75t_R FILLER_140_21 ();
 FILLER_ASAP7_75t_R FILLER_140_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_41 ();
 DECAPx2_ASAP7_75t_R FILLER_140_48 ();
 FILLER_ASAP7_75t_R FILLER_140_54 ();
 DECAPx4_ASAP7_75t_R FILLER_140_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_70 ();
 DECAPx2_ASAP7_75t_R FILLER_140_77 ();
 FILLER_ASAP7_75t_R FILLER_140_83 ();
 DECAPx10_ASAP7_75t_R FILLER_140_115 ();
 DECAPx1_ASAP7_75t_R FILLER_140_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_141 ();
 DECAPx4_ASAP7_75t_R FILLER_140_168 ();
 FILLER_ASAP7_75t_R FILLER_140_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_180 ();
 FILLER_ASAP7_75t_R FILLER_140_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_189 ();
 DECAPx6_ASAP7_75t_R FILLER_140_193 ();
 FILLER_ASAP7_75t_R FILLER_140_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_215 ();
 DECAPx6_ASAP7_75t_R FILLER_140_228 ();
 DECAPx1_ASAP7_75t_R FILLER_140_242 ();
 DECAPx6_ASAP7_75t_R FILLER_140_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_266 ();
 DECAPx6_ASAP7_75t_R FILLER_140_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_333 ();
 DECAPx1_ASAP7_75t_R FILLER_140_342 ();
 DECAPx2_ASAP7_75t_R FILLER_140_352 ();
 DECAPx2_ASAP7_75t_R FILLER_140_364 ();
 FILLER_ASAP7_75t_R FILLER_140_370 ();
 DECAPx2_ASAP7_75t_R FILLER_140_375 ();
 FILLER_ASAP7_75t_R FILLER_140_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_383 ();
 DECAPx4_ASAP7_75t_R FILLER_140_410 ();
 FILLER_ASAP7_75t_R FILLER_140_420 ();
 DECAPx1_ASAP7_75t_R FILLER_140_432 ();
 DECAPx4_ASAP7_75t_R FILLER_140_470 ();
 DECAPx2_ASAP7_75t_R FILLER_140_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_503 ();
 FILLER_ASAP7_75t_R FILLER_140_553 ();
 DECAPx1_ASAP7_75t_R FILLER_140_581 ();
 FILLER_ASAP7_75t_R FILLER_140_611 ();
 DECAPx1_ASAP7_75t_R FILLER_140_619 ();
 DECAPx6_ASAP7_75t_R FILLER_140_659 ();
 DECAPx10_ASAP7_75t_R FILLER_140_695 ();
 DECAPx2_ASAP7_75t_R FILLER_140_725 ();
 DECAPx1_ASAP7_75t_R FILLER_140_739 ();
 DECAPx2_ASAP7_75t_R FILLER_140_763 ();
 DECAPx10_ASAP7_75t_R FILLER_140_779 ();
 DECAPx10_ASAP7_75t_R FILLER_140_801 ();
 DECAPx2_ASAP7_75t_R FILLER_140_823 ();
 FILLER_ASAP7_75t_R FILLER_140_829 ();
 DECAPx1_ASAP7_75t_R FILLER_140_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_853 ();
 DECAPx2_ASAP7_75t_R FILLER_140_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_896 ();
 DECAPx1_ASAP7_75t_R FILLER_140_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_911 ();
 FILLER_ASAP7_75t_R FILLER_140_934 ();
 DECAPx6_ASAP7_75t_R FILLER_140_947 ();
 FILLER_ASAP7_75t_R FILLER_140_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_963 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1014 ();
 FILLER_ASAP7_75t_R FILLER_140_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_140_1072 ();
 DECAPx4_ASAP7_75t_R FILLER_140_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1142 ();
 DECAPx4_ASAP7_75t_R FILLER_140_1170 ();
 FILLER_ASAP7_75t_R FILLER_140_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1182 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1190 ();
 FILLER_ASAP7_75t_R FILLER_140_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1248 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1284 ();
 DECAPx4_ASAP7_75t_R FILLER_140_1293 ();
 FILLER_ASAP7_75t_R FILLER_140_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1305 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1312 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1316 ();
 DECAPx4_ASAP7_75t_R FILLER_140_1323 ();
 FILLER_ASAP7_75t_R FILLER_140_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1341 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1363 ();
 FILLER_ASAP7_75t_R FILLER_140_1369 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1377 ();
 FILLER_ASAP7_75t_R FILLER_140_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1388 ();
 FILLER_ASAP7_75t_R FILLER_141_2 ();
 DECAPx1_ASAP7_75t_R FILLER_141_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_60 ();
 DECAPx4_ASAP7_75t_R FILLER_141_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_87 ();
 DECAPx2_ASAP7_75t_R FILLER_141_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_97 ();
 DECAPx4_ASAP7_75t_R FILLER_141_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_117 ();
 DECAPx4_ASAP7_75t_R FILLER_141_131 ();
 FILLER_ASAP7_75t_R FILLER_141_141 ();
 DECAPx4_ASAP7_75t_R FILLER_141_176 ();
 FILLER_ASAP7_75t_R FILLER_141_186 ();
 DECAPx2_ASAP7_75t_R FILLER_141_214 ();
 DECAPx10_ASAP7_75t_R FILLER_141_223 ();
 FILLER_ASAP7_75t_R FILLER_141_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_259 ();
 DECAPx2_ASAP7_75t_R FILLER_141_266 ();
 FILLER_ASAP7_75t_R FILLER_141_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_274 ();
 DECAPx6_ASAP7_75t_R FILLER_141_290 ();
 FILLER_ASAP7_75t_R FILLER_141_304 ();
 DECAPx6_ASAP7_75t_R FILLER_141_316 ();
 FILLER_ASAP7_75t_R FILLER_141_330 ();
 FILLER_ASAP7_75t_R FILLER_141_338 ();
 DECAPx2_ASAP7_75t_R FILLER_141_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_352 ();
 DECAPx4_ASAP7_75t_R FILLER_141_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_402 ();
 DECAPx4_ASAP7_75t_R FILLER_141_410 ();
 FILLER_ASAP7_75t_R FILLER_141_420 ();
 FILLER_ASAP7_75t_R FILLER_141_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_449 ();
 DECAPx10_ASAP7_75t_R FILLER_141_456 ();
 DECAPx4_ASAP7_75t_R FILLER_141_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_488 ();
 DECAPx2_ASAP7_75t_R FILLER_141_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_528 ();
 DECAPx2_ASAP7_75t_R FILLER_141_542 ();
 FILLER_ASAP7_75t_R FILLER_141_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_564 ();
 DECAPx1_ASAP7_75t_R FILLER_141_574 ();
 DECAPx2_ASAP7_75t_R FILLER_141_591 ();
 FILLER_ASAP7_75t_R FILLER_141_603 ();
 DECAPx6_ASAP7_75t_R FILLER_141_609 ();
 DECAPx2_ASAP7_75t_R FILLER_141_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_629 ();
 DECAPx4_ASAP7_75t_R FILLER_141_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_643 ();
 DECAPx2_ASAP7_75t_R FILLER_141_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_672 ();
 DECAPx1_ASAP7_75t_R FILLER_141_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_686 ();
 DECAPx6_ASAP7_75t_R FILLER_141_703 ();
 FILLER_ASAP7_75t_R FILLER_141_717 ();
 DECAPx1_ASAP7_75t_R FILLER_141_725 ();
 DECAPx2_ASAP7_75t_R FILLER_141_739 ();
 DECAPx6_ASAP7_75t_R FILLER_141_765 ();
 FILLER_ASAP7_75t_R FILLER_141_779 ();
 DECAPx1_ASAP7_75t_R FILLER_141_791 ();
 FILLER_ASAP7_75t_R FILLER_141_805 ();
 DECAPx2_ASAP7_75t_R FILLER_141_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_830 ();
 DECAPx2_ASAP7_75t_R FILLER_141_843 ();
 FILLER_ASAP7_75t_R FILLER_141_849 ();
 DECAPx1_ASAP7_75t_R FILLER_141_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_865 ();
 DECAPx1_ASAP7_75t_R FILLER_141_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_893 ();
 DECAPx6_ASAP7_75t_R FILLER_141_908 ();
 FILLER_ASAP7_75t_R FILLER_141_922 ();
 DECAPx1_ASAP7_75t_R FILLER_141_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_961 ();
 DECAPx2_ASAP7_75t_R FILLER_141_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_978 ();
 FILLER_ASAP7_75t_R FILLER_141_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1023 ();
 FILLER_ASAP7_75t_R FILLER_141_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_141_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1074 ();
 FILLER_ASAP7_75t_R FILLER_141_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1094 ();
 FILLER_ASAP7_75t_R FILLER_141_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_141_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1192 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1203 ();
 FILLER_ASAP7_75t_R FILLER_141_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1211 ();
 FILLER_ASAP7_75t_R FILLER_141_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1224 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1249 ();
 FILLER_ASAP7_75t_R FILLER_141_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1261 ();
 FILLER_ASAP7_75t_R FILLER_141_1302 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1318 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1335 ();
 DECAPx6_ASAP7_75t_R FILLER_141_1350 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_142_2 ();
 FILLER_ASAP7_75t_R FILLER_142_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_10 ();
 FILLER_ASAP7_75t_R FILLER_142_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_19 ();
 DECAPx6_ASAP7_75t_R FILLER_142_23 ();
 DECAPx2_ASAP7_75t_R FILLER_142_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_43 ();
 DECAPx4_ASAP7_75t_R FILLER_142_47 ();
 FILLER_ASAP7_75t_R FILLER_142_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_59 ();
 FILLER_ASAP7_75t_R FILLER_142_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_88 ();
 DECAPx4_ASAP7_75t_R FILLER_142_92 ();
 FILLER_ASAP7_75t_R FILLER_142_102 ();
 FILLER_ASAP7_75t_R FILLER_142_114 ();
 DECAPx1_ASAP7_75t_R FILLER_142_142 ();
 DECAPx1_ASAP7_75t_R FILLER_142_159 ();
 DECAPx2_ASAP7_75t_R FILLER_142_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_238 ();
 FILLER_ASAP7_75t_R FILLER_142_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_255 ();
 DECAPx10_ASAP7_75t_R FILLER_142_285 ();
 FILLER_ASAP7_75t_R FILLER_142_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_336 ();
 DECAPx2_ASAP7_75t_R FILLER_142_343 ();
 DECAPx1_ASAP7_75t_R FILLER_142_352 ();
 DECAPx1_ASAP7_75t_R FILLER_142_362 ();
 DECAPx10_ASAP7_75t_R FILLER_142_374 ();
 DECAPx1_ASAP7_75t_R FILLER_142_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_400 ();
 DECAPx2_ASAP7_75t_R FILLER_142_427 ();
 FILLER_ASAP7_75t_R FILLER_142_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_464 ();
 DECAPx2_ASAP7_75t_R FILLER_142_471 ();
 DECAPx4_ASAP7_75t_R FILLER_142_480 ();
 FILLER_ASAP7_75t_R FILLER_142_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_492 ();
 DECAPx2_ASAP7_75t_R FILLER_142_503 ();
 FILLER_ASAP7_75t_R FILLER_142_509 ();
 DECAPx10_ASAP7_75t_R FILLER_142_514 ();
 DECAPx6_ASAP7_75t_R FILLER_142_536 ();
 FILLER_ASAP7_75t_R FILLER_142_550 ();
 DECAPx10_ASAP7_75t_R FILLER_142_559 ();
 FILLER_ASAP7_75t_R FILLER_142_581 ();
 DECAPx6_ASAP7_75t_R FILLER_142_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_604 ();
 DECAPx10_ASAP7_75t_R FILLER_142_611 ();
 DECAPx10_ASAP7_75t_R FILLER_142_633 ();
 DECAPx10_ASAP7_75t_R FILLER_142_655 ();
 FILLER_ASAP7_75t_R FILLER_142_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_685 ();
 DECAPx2_ASAP7_75t_R FILLER_142_692 ();
 DECAPx6_ASAP7_75t_R FILLER_142_718 ();
 DECAPx4_ASAP7_75t_R FILLER_142_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_748 ();
 DECAPx1_ASAP7_75t_R FILLER_142_752 ();
 DECAPx2_ASAP7_75t_R FILLER_142_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_774 ();
 FILLER_ASAP7_75t_R FILLER_142_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_807 ();
 DECAPx2_ASAP7_75t_R FILLER_142_843 ();
 FILLER_ASAP7_75t_R FILLER_142_849 ();
 DECAPx1_ASAP7_75t_R FILLER_142_863 ();
 DECAPx10_ASAP7_75t_R FILLER_142_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_909 ();
 DECAPx4_ASAP7_75t_R FILLER_142_922 ();
 FILLER_ASAP7_75t_R FILLER_142_932 ();
 FILLER_ASAP7_75t_R FILLER_142_946 ();
 FILLER_ASAP7_75t_R FILLER_142_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_953 ();
 DECAPx4_ASAP7_75t_R FILLER_142_958 ();
 FILLER_ASAP7_75t_R FILLER_142_968 ();
 DECAPx2_ASAP7_75t_R FILLER_142_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_982 ();
 FILLER_ASAP7_75t_R FILLER_142_989 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1000 ();
 FILLER_ASAP7_75t_R FILLER_142_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1055 ();
 FILLER_ASAP7_75t_R FILLER_142_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1155 ();
 FILLER_ASAP7_75t_R FILLER_142_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1207 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1231 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1268 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1331 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1388 ();
 DECAPx1_ASAP7_75t_R FILLER_143_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_6 ();
 DECAPx1_ASAP7_75t_R FILLER_143_19 ();
 DECAPx1_ASAP7_75t_R FILLER_143_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_31 ();
 DECAPx1_ASAP7_75t_R FILLER_143_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_43 ();
 DECAPx4_ASAP7_75t_R FILLER_143_47 ();
 DECAPx2_ASAP7_75t_R FILLER_143_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_74 ();
 DECAPx2_ASAP7_75t_R FILLER_143_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_84 ();
 DECAPx2_ASAP7_75t_R FILLER_143_92 ();
 DECAPx6_ASAP7_75t_R FILLER_143_101 ();
 DECAPx2_ASAP7_75t_R FILLER_143_115 ();
 FILLER_ASAP7_75t_R FILLER_143_139 ();
 DECAPx2_ASAP7_75t_R FILLER_143_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_157 ();
 DECAPx2_ASAP7_75t_R FILLER_143_161 ();
 FILLER_ASAP7_75t_R FILLER_143_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_169 ();
 FILLER_ASAP7_75t_R FILLER_143_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_188 ();
 DECAPx4_ASAP7_75t_R FILLER_143_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_205 ();
 DECAPx4_ASAP7_75t_R FILLER_143_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_223 ();
 DECAPx4_ASAP7_75t_R FILLER_143_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_260 ();
 DECAPx1_ASAP7_75t_R FILLER_143_267 ();
 DECAPx4_ASAP7_75t_R FILLER_143_274 ();
 FILLER_ASAP7_75t_R FILLER_143_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_298 ();
 FILLER_ASAP7_75t_R FILLER_143_302 ();
 FILLER_ASAP7_75t_R FILLER_143_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_309 ();
 DECAPx2_ASAP7_75t_R FILLER_143_316 ();
 FILLER_ASAP7_75t_R FILLER_143_322 ();
 DECAPx2_ASAP7_75t_R FILLER_143_327 ();
 FILLER_ASAP7_75t_R FILLER_143_333 ();
 DECAPx4_ASAP7_75t_R FILLER_143_361 ();
 FILLER_ASAP7_75t_R FILLER_143_371 ();
 DECAPx2_ASAP7_75t_R FILLER_143_399 ();
 DECAPx1_ASAP7_75t_R FILLER_143_411 ();
 DECAPx2_ASAP7_75t_R FILLER_143_418 ();
 FILLER_ASAP7_75t_R FILLER_143_424 ();
 FILLER_ASAP7_75t_R FILLER_143_450 ();
 DECAPx4_ASAP7_75t_R FILLER_143_485 ();
 FILLER_ASAP7_75t_R FILLER_143_495 ();
 DECAPx4_ASAP7_75t_R FILLER_143_527 ();
 FILLER_ASAP7_75t_R FILLER_143_540 ();
 DECAPx1_ASAP7_75t_R FILLER_143_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_550 ();
 DECAPx6_ASAP7_75t_R FILLER_143_569 ();
 FILLER_ASAP7_75t_R FILLER_143_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_585 ();
 DECAPx1_ASAP7_75t_R FILLER_143_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_600 ();
 FILLER_ASAP7_75t_R FILLER_143_627 ();
 DECAPx1_ASAP7_75t_R FILLER_143_647 ();
 DECAPx10_ASAP7_75t_R FILLER_143_681 ();
 DECAPx1_ASAP7_75t_R FILLER_143_703 ();
 DECAPx10_ASAP7_75t_R FILLER_143_723 ();
 DECAPx2_ASAP7_75t_R FILLER_143_745 ();
 DECAPx2_ASAP7_75t_R FILLER_143_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_779 ();
 DECAPx6_ASAP7_75t_R FILLER_143_795 ();
 DECAPx1_ASAP7_75t_R FILLER_143_809 ();
 DECAPx10_ASAP7_75t_R FILLER_143_822 ();
 DECAPx10_ASAP7_75t_R FILLER_143_844 ();
 DECAPx4_ASAP7_75t_R FILLER_143_866 ();
 DECAPx6_ASAP7_75t_R FILLER_143_882 ();
 FILLER_ASAP7_75t_R FILLER_143_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_904 ();
 FILLER_ASAP7_75t_R FILLER_143_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_923 ();
 FILLER_ASAP7_75t_R FILLER_143_933 ();
 DECAPx4_ASAP7_75t_R FILLER_143_954 ();
 FILLER_ASAP7_75t_R FILLER_143_964 ();
 DECAPx2_ASAP7_75t_R FILLER_143_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_982 ();
 DECAPx2_ASAP7_75t_R FILLER_143_989 ();
 FILLER_ASAP7_75t_R FILLER_143_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1007 ();
 FILLER_ASAP7_75t_R FILLER_143_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1073 ();
 FILLER_ASAP7_75t_R FILLER_143_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1081 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1088 ();
 FILLER_ASAP7_75t_R FILLER_143_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1125 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1157 ();
 FILLER_ASAP7_75t_R FILLER_143_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1186 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1247 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1274 ();
 FILLER_ASAP7_75t_R FILLER_143_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1295 ();
 FILLER_ASAP7_75t_R FILLER_143_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1337 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1364 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_28 ();
 FILLER_ASAP7_75t_R FILLER_144_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_57 ();
 DECAPx4_ASAP7_75t_R FILLER_144_110 ();
 FILLER_ASAP7_75t_R FILLER_144_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_122 ();
 DECAPx2_ASAP7_75t_R FILLER_144_149 ();
 FILLER_ASAP7_75t_R FILLER_144_155 ();
 FILLER_ASAP7_75t_R FILLER_144_183 ();
 DECAPx6_ASAP7_75t_R FILLER_144_198 ();
 FILLER_ASAP7_75t_R FILLER_144_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_214 ();
 FILLER_ASAP7_75t_R FILLER_144_225 ();
 DECAPx1_ASAP7_75t_R FILLER_144_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_238 ();
 FILLER_ASAP7_75t_R FILLER_144_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_244 ();
 DECAPx6_ASAP7_75t_R FILLER_144_248 ();
 DECAPx2_ASAP7_75t_R FILLER_144_262 ();
 DECAPx1_ASAP7_75t_R FILLER_144_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_283 ();
 DECAPx1_ASAP7_75t_R FILLER_144_310 ();
 DECAPx4_ASAP7_75t_R FILLER_144_321 ();
 FILLER_ASAP7_75t_R FILLER_144_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_333 ();
 DECAPx4_ASAP7_75t_R FILLER_144_341 ();
 DECAPx2_ASAP7_75t_R FILLER_144_371 ();
 FILLER_ASAP7_75t_R FILLER_144_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_387 ();
 DECAPx10_ASAP7_75t_R FILLER_144_391 ();
 DECAPx10_ASAP7_75t_R FILLER_144_413 ();
 DECAPx2_ASAP7_75t_R FILLER_144_435 ();
 FILLER_ASAP7_75t_R FILLER_144_441 ();
 DECAPx4_ASAP7_75t_R FILLER_144_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_461 ();
 DECAPx2_ASAP7_75t_R FILLER_144_464 ();
 FILLER_ASAP7_75t_R FILLER_144_470 ();
 DECAPx2_ASAP7_75t_R FILLER_144_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_494 ();
 DECAPx2_ASAP7_75t_R FILLER_144_507 ();
 FILLER_ASAP7_75t_R FILLER_144_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_515 ();
 DECAPx6_ASAP7_75t_R FILLER_144_548 ();
 FILLER_ASAP7_75t_R FILLER_144_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_564 ();
 DECAPx2_ASAP7_75t_R FILLER_144_620 ();
 FILLER_ASAP7_75t_R FILLER_144_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_628 ();
 DECAPx4_ASAP7_75t_R FILLER_144_647 ();
 FILLER_ASAP7_75t_R FILLER_144_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_659 ();
 DECAPx1_ASAP7_75t_R FILLER_144_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_677 ();
 DECAPx2_ASAP7_75t_R FILLER_144_695 ();
 FILLER_ASAP7_75t_R FILLER_144_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_712 ();
 FILLER_ASAP7_75t_R FILLER_144_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_725 ();
 FILLER_ASAP7_75t_R FILLER_144_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_735 ();
 DECAPx6_ASAP7_75t_R FILLER_144_750 ();
 FILLER_ASAP7_75t_R FILLER_144_764 ();
 DECAPx4_ASAP7_75t_R FILLER_144_784 ();
 FILLER_ASAP7_75t_R FILLER_144_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_796 ();
 FILLER_ASAP7_75t_R FILLER_144_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_809 ();
 DECAPx2_ASAP7_75t_R FILLER_144_818 ();
 FILLER_ASAP7_75t_R FILLER_144_824 ();
 DECAPx1_ASAP7_75t_R FILLER_144_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_850 ();
 DECAPx4_ASAP7_75t_R FILLER_144_859 ();
 FILLER_ASAP7_75t_R FILLER_144_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_871 ();
 DECAPx4_ASAP7_75t_R FILLER_144_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_889 ();
 DECAPx4_ASAP7_75t_R FILLER_144_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_909 ();
 DECAPx4_ASAP7_75t_R FILLER_144_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_930 ();
 DECAPx6_ASAP7_75t_R FILLER_144_947 ();
 DECAPx6_ASAP7_75t_R FILLER_144_991 ();
 FILLER_ASAP7_75t_R FILLER_144_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1018 ();
 FILLER_ASAP7_75t_R FILLER_144_1024 ();
 FILLER_ASAP7_75t_R FILLER_144_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1045 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1071 ();
 FILLER_ASAP7_75t_R FILLER_144_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1116 ();
 FILLER_ASAP7_75t_R FILLER_144_1143 ();
 FILLER_ASAP7_75t_R FILLER_144_1148 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1168 ();
 FILLER_ASAP7_75t_R FILLER_144_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1220 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1227 ();
 FILLER_ASAP7_75t_R FILLER_144_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1254 ();
 DECAPx4_ASAP7_75t_R FILLER_144_1262 ();
 FILLER_ASAP7_75t_R FILLER_144_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1314 ();
 FILLER_ASAP7_75t_R FILLER_144_1320 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1322 ();
 DECAPx4_ASAP7_75t_R FILLER_144_1329 ();
 FILLER_ASAP7_75t_R FILLER_144_1339 ();
 FILLER_ASAP7_75t_R FILLER_144_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1349 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1356 ();
 FILLER_ASAP7_75t_R FILLER_144_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_145_2 ();
 FILLER_ASAP7_75t_R FILLER_145_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_14 ();
 DECAPx2_ASAP7_75t_R FILLER_145_18 ();
 FILLER_ASAP7_75t_R FILLER_145_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_37 ();
 FILLER_ASAP7_75t_R FILLER_145_44 ();
 DECAPx1_ASAP7_75t_R FILLER_145_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_57 ();
 DECAPx6_ASAP7_75t_R FILLER_145_68 ();
 DECAPx2_ASAP7_75t_R FILLER_145_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_94 ();
 DECAPx2_ASAP7_75t_R FILLER_145_121 ();
 FILLER_ASAP7_75t_R FILLER_145_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_129 ();
 DECAPx1_ASAP7_75t_R FILLER_145_133 ();
 DECAPx6_ASAP7_75t_R FILLER_145_167 ();
 FILLER_ASAP7_75t_R FILLER_145_181 ();
 FILLER_ASAP7_75t_R FILLER_145_216 ();
 DECAPx1_ASAP7_75t_R FILLER_145_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_248 ();
 FILLER_ASAP7_75t_R FILLER_145_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_287 ();
 FILLER_ASAP7_75t_R FILLER_145_294 ();
 DECAPx1_ASAP7_75t_R FILLER_145_310 ();
 DECAPx4_ASAP7_75t_R FILLER_145_340 ();
 FILLER_ASAP7_75t_R FILLER_145_350 ();
 DECAPx4_ASAP7_75t_R FILLER_145_366 ();
 DECAPx2_ASAP7_75t_R FILLER_145_386 ();
 DECAPx6_ASAP7_75t_R FILLER_145_420 ();
 FILLER_ASAP7_75t_R FILLER_145_434 ();
 FILLER_ASAP7_75t_R FILLER_145_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_477 ();
 DECAPx2_ASAP7_75t_R FILLER_145_507 ();
 FILLER_ASAP7_75t_R FILLER_145_513 ();
 FILLER_ASAP7_75t_R FILLER_145_518 ();
 DECAPx2_ASAP7_75t_R FILLER_145_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_572 ();
 DECAPx10_ASAP7_75t_R FILLER_145_600 ();
 DECAPx6_ASAP7_75t_R FILLER_145_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_636 ();
 DECAPx4_ASAP7_75t_R FILLER_145_675 ();
 FILLER_ASAP7_75t_R FILLER_145_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_687 ();
 DECAPx4_ASAP7_75t_R FILLER_145_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_715 ();
 FILLER_ASAP7_75t_R FILLER_145_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_737 ();
 DECAPx6_ASAP7_75t_R FILLER_145_755 ();
 FILLER_ASAP7_75t_R FILLER_145_769 ();
 DECAPx2_ASAP7_75t_R FILLER_145_784 ();
 FILLER_ASAP7_75t_R FILLER_145_790 ();
 FILLER_ASAP7_75t_R FILLER_145_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_807 ();
 DECAPx1_ASAP7_75t_R FILLER_145_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_818 ();
 DECAPx6_ASAP7_75t_R FILLER_145_825 ();
 FILLER_ASAP7_75t_R FILLER_145_839 ();
 FILLER_ASAP7_75t_R FILLER_145_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_864 ();
 DECAPx4_ASAP7_75t_R FILLER_145_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_914 ();
 FILLER_ASAP7_75t_R FILLER_145_922 ();
 DECAPx1_ASAP7_75t_R FILLER_145_926 ();
 DECAPx2_ASAP7_75t_R FILLER_145_944 ();
 FILLER_ASAP7_75t_R FILLER_145_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_952 ();
 DECAPx10_ASAP7_75t_R FILLER_145_971 ();
 DECAPx1_ASAP7_75t_R FILLER_145_993 ();
 FILLER_ASAP7_75t_R FILLER_145_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_145_1016 ();
 FILLER_ASAP7_75t_R FILLER_145_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1060 ();
 FILLER_ASAP7_75t_R FILLER_145_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1117 ();
 DECAPx6_ASAP7_75t_R FILLER_145_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1156 ();
 FILLER_ASAP7_75t_R FILLER_145_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1174 ();
 DECAPx6_ASAP7_75t_R FILLER_145_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_145_1224 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1244 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1303 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1328 ();
 FILLER_ASAP7_75t_R FILLER_145_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1353 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1360 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_146_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_32 ();
 DECAPx1_ASAP7_75t_R FILLER_146_59 ();
 DECAPx2_ASAP7_75t_R FILLER_146_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_76 ();
 DECAPx4_ASAP7_75t_R FILLER_146_80 ();
 FILLER_ASAP7_75t_R FILLER_146_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_96 ();
 DECAPx2_ASAP7_75t_R FILLER_146_113 ();
 FILLER_ASAP7_75t_R FILLER_146_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_141 ();
 DECAPx6_ASAP7_75t_R FILLER_146_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_162 ();
 DECAPx1_ASAP7_75t_R FILLER_146_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_174 ();
 DECAPx2_ASAP7_75t_R FILLER_146_181 ();
 FILLER_ASAP7_75t_R FILLER_146_187 ();
 DECAPx1_ASAP7_75t_R FILLER_146_215 ();
 DECAPx2_ASAP7_75t_R FILLER_146_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_231 ();
 DECAPx4_ASAP7_75t_R FILLER_146_235 ();
 FILLER_ASAP7_75t_R FILLER_146_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_247 ();
 DECAPx2_ASAP7_75t_R FILLER_146_258 ();
 FILLER_ASAP7_75t_R FILLER_146_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_266 ();
 FILLER_ASAP7_75t_R FILLER_146_273 ();
 DECAPx2_ASAP7_75t_R FILLER_146_278 ();
 FILLER_ASAP7_75t_R FILLER_146_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_286 ();
 DECAPx10_ASAP7_75t_R FILLER_146_295 ();
 DECAPx1_ASAP7_75t_R FILLER_146_323 ();
 DECAPx1_ASAP7_75t_R FILLER_146_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_360 ();
 DECAPx2_ASAP7_75t_R FILLER_146_371 ();
 DECAPx6_ASAP7_75t_R FILLER_146_383 ();
 FILLER_ASAP7_75t_R FILLER_146_397 ();
 DECAPx2_ASAP7_75t_R FILLER_146_417 ();
 FILLER_ASAP7_75t_R FILLER_146_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_425 ();
 DECAPx2_ASAP7_75t_R FILLER_146_453 ();
 FILLER_ASAP7_75t_R FILLER_146_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_461 ();
 DECAPx1_ASAP7_75t_R FILLER_146_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_494 ();
 DECAPx10_ASAP7_75t_R FILLER_146_498 ();
 DECAPx10_ASAP7_75t_R FILLER_146_520 ();
 DECAPx4_ASAP7_75t_R FILLER_146_542 ();
 DECAPx4_ASAP7_75t_R FILLER_146_572 ();
 FILLER_ASAP7_75t_R FILLER_146_582 ();
 DECAPx4_ASAP7_75t_R FILLER_146_592 ();
 FILLER_ASAP7_75t_R FILLER_146_602 ();
 DECAPx4_ASAP7_75t_R FILLER_146_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_624 ();
 DECAPx1_ASAP7_75t_R FILLER_146_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_639 ();
 DECAPx6_ASAP7_75t_R FILLER_146_658 ();
 DECAPx1_ASAP7_75t_R FILLER_146_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_676 ();
 DECAPx2_ASAP7_75t_R FILLER_146_695 ();
 FILLER_ASAP7_75t_R FILLER_146_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_703 ();
 FILLER_ASAP7_75t_R FILLER_146_722 ();
 FILLER_ASAP7_75t_R FILLER_146_730 ();
 FILLER_ASAP7_75t_R FILLER_146_735 ();
 DECAPx2_ASAP7_75t_R FILLER_146_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_755 ();
 DECAPx2_ASAP7_75t_R FILLER_146_759 ();
 FILLER_ASAP7_75t_R FILLER_146_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_767 ();
 DECAPx4_ASAP7_75t_R FILLER_146_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_781 ();
 DECAPx2_ASAP7_75t_R FILLER_146_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_811 ();
 DECAPx1_ASAP7_75t_R FILLER_146_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_839 ();
 FILLER_ASAP7_75t_R FILLER_146_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_876 ();
 DECAPx1_ASAP7_75t_R FILLER_146_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_888 ();
 DECAPx2_ASAP7_75t_R FILLER_146_907 ();
 DECAPx4_ASAP7_75t_R FILLER_146_943 ();
 FILLER_ASAP7_75t_R FILLER_146_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_955 ();
 DECAPx6_ASAP7_75t_R FILLER_146_981 ();
 DECAPx4_ASAP7_75t_R FILLER_146_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_146_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1111 ();
 FILLER_ASAP7_75t_R FILLER_146_1117 ();
 FILLER_ASAP7_75t_R FILLER_146_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_146_1159 ();
 DECAPx4_ASAP7_75t_R FILLER_146_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1191 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1214 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1237 ();
 FILLER_ASAP7_75t_R FILLER_146_1270 ();
 DECAPx4_ASAP7_75t_R FILLER_146_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1319 ();
 FILLER_ASAP7_75t_R FILLER_146_1333 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1353 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_147_2 ();
 FILLER_ASAP7_75t_R FILLER_147_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_18 ();
 DECAPx6_ASAP7_75t_R FILLER_147_31 ();
 FILLER_ASAP7_75t_R FILLER_147_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_47 ();
 DECAPx1_ASAP7_75t_R FILLER_147_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_61 ();
 DECAPx10_ASAP7_75t_R FILLER_147_88 ();
 DECAPx4_ASAP7_75t_R FILLER_147_110 ();
 FILLER_ASAP7_75t_R FILLER_147_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_122 ();
 DECAPx2_ASAP7_75t_R FILLER_147_130 ();
 FILLER_ASAP7_75t_R FILLER_147_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_171 ();
 DECAPx4_ASAP7_75t_R FILLER_147_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_185 ();
 FILLER_ASAP7_75t_R FILLER_147_189 ();
 DECAPx1_ASAP7_75t_R FILLER_147_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_201 ();
 DECAPx10_ASAP7_75t_R FILLER_147_208 ();
 DECAPx2_ASAP7_75t_R FILLER_147_230 ();
 FILLER_ASAP7_75t_R FILLER_147_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_238 ();
 DECAPx6_ASAP7_75t_R FILLER_147_271 ();
 DECAPx2_ASAP7_75t_R FILLER_147_285 ();
 DECAPx2_ASAP7_75t_R FILLER_147_297 ();
 FILLER_ASAP7_75t_R FILLER_147_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_305 ();
 DECAPx2_ASAP7_75t_R FILLER_147_324 ();
 FILLER_ASAP7_75t_R FILLER_147_330 ();
 DECAPx6_ASAP7_75t_R FILLER_147_348 ();
 FILLER_ASAP7_75t_R FILLER_147_362 ();
 DECAPx2_ASAP7_75t_R FILLER_147_371 ();
 FILLER_ASAP7_75t_R FILLER_147_380 ();
 DECAPx6_ASAP7_75t_R FILLER_147_403 ();
 FILLER_ASAP7_75t_R FILLER_147_417 ();
 DECAPx6_ASAP7_75t_R FILLER_147_437 ();
 FILLER_ASAP7_75t_R FILLER_147_451 ();
 DECAPx2_ASAP7_75t_R FILLER_147_471 ();
 FILLER_ASAP7_75t_R FILLER_147_477 ();
 DECAPx6_ASAP7_75t_R FILLER_147_482 ();
 FILLER_ASAP7_75t_R FILLER_147_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_498 ();
 DECAPx4_ASAP7_75t_R FILLER_147_505 ();
 FILLER_ASAP7_75t_R FILLER_147_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_517 ();
 DECAPx1_ASAP7_75t_R FILLER_147_521 ();
 DECAPx10_ASAP7_75t_R FILLER_147_529 ();
 DECAPx10_ASAP7_75t_R FILLER_147_551 ();
 DECAPx10_ASAP7_75t_R FILLER_147_573 ();
 DECAPx2_ASAP7_75t_R FILLER_147_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_601 ();
 DECAPx2_ASAP7_75t_R FILLER_147_634 ();
 FILLER_ASAP7_75t_R FILLER_147_640 ();
 DECAPx1_ASAP7_75t_R FILLER_147_662 ();
 DECAPx4_ASAP7_75t_R FILLER_147_684 ();
 DECAPx4_ASAP7_75t_R FILLER_147_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_714 ();
 DECAPx4_ASAP7_75t_R FILLER_147_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_733 ();
 DECAPx2_ASAP7_75t_R FILLER_147_744 ();
 DECAPx1_ASAP7_75t_R FILLER_147_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_774 ();
 DECAPx2_ASAP7_75t_R FILLER_147_783 ();
 DECAPx1_ASAP7_75t_R FILLER_147_804 ();
 FILLER_ASAP7_75t_R FILLER_147_834 ();
 DECAPx1_ASAP7_75t_R FILLER_147_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_861 ();
 DECAPx2_ASAP7_75t_R FILLER_147_884 ();
 DECAPx4_ASAP7_75t_R FILLER_147_905 ();
 FILLER_ASAP7_75t_R FILLER_147_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_923 ();
 DECAPx4_ASAP7_75t_R FILLER_147_926 ();
 FILLER_ASAP7_75t_R FILLER_147_936 ();
 DECAPx4_ASAP7_75t_R FILLER_147_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_954 ();
 DECAPx2_ASAP7_75t_R FILLER_147_961 ();
 DECAPx2_ASAP7_75t_R FILLER_147_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_996 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1023 ();
 FILLER_ASAP7_75t_R FILLER_147_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1037 ();
 FILLER_ASAP7_75t_R FILLER_147_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1052 ();
 FILLER_ASAP7_75t_R FILLER_147_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1088 ();
 FILLER_ASAP7_75t_R FILLER_147_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_147_1100 ();
 FILLER_ASAP7_75t_R FILLER_147_1116 ();
 FILLER_ASAP7_75t_R FILLER_147_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1158 ();
 FILLER_ASAP7_75t_R FILLER_147_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1202 ();
 FILLER_ASAP7_75t_R FILLER_147_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1210 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1315 ();
 FILLER_ASAP7_75t_R FILLER_147_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1346 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1372 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1391 ();
 DECAPx2_ASAP7_75t_R FILLER_148_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_40 ();
 FILLER_ASAP7_75t_R FILLER_148_48 ();
 DECAPx2_ASAP7_75t_R FILLER_148_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_60 ();
 DECAPx1_ASAP7_75t_R FILLER_148_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_77 ();
 DECAPx2_ASAP7_75t_R FILLER_148_82 ();
 FILLER_ASAP7_75t_R FILLER_148_88 ();
 DECAPx6_ASAP7_75t_R FILLER_148_116 ();
 FILLER_ASAP7_75t_R FILLER_148_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_132 ();
 FILLER_ASAP7_75t_R FILLER_148_139 ();
 DECAPx2_ASAP7_75t_R FILLER_148_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_157 ();
 FILLER_ASAP7_75t_R FILLER_148_184 ();
 DECAPx6_ASAP7_75t_R FILLER_148_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_208 ();
 DECAPx2_ASAP7_75t_R FILLER_148_229 ();
 DECAPx1_ASAP7_75t_R FILLER_148_242 ();
 DECAPx2_ASAP7_75t_R FILLER_148_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_259 ();
 DECAPx1_ASAP7_75t_R FILLER_148_263 ();
 FILLER_ASAP7_75t_R FILLER_148_273 ();
 FILLER_ASAP7_75t_R FILLER_148_281 ();
 DECAPx2_ASAP7_75t_R FILLER_148_298 ();
 DECAPx10_ASAP7_75t_R FILLER_148_314 ();
 DECAPx2_ASAP7_75t_R FILLER_148_336 ();
 FILLER_ASAP7_75t_R FILLER_148_342 ();
 DECAPx2_ASAP7_75t_R FILLER_148_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_356 ();
 DECAPx10_ASAP7_75t_R FILLER_148_389 ();
 DECAPx6_ASAP7_75t_R FILLER_148_411 ();
 DECAPx1_ASAP7_75t_R FILLER_148_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_429 ();
 DECAPx6_ASAP7_75t_R FILLER_148_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_464 ();
 FILLER_ASAP7_75t_R FILLER_148_495 ();
 DECAPx2_ASAP7_75t_R FILLER_148_530 ();
 FILLER_ASAP7_75t_R FILLER_148_544 ();
 DECAPx2_ASAP7_75t_R FILLER_148_559 ();
 FILLER_ASAP7_75t_R FILLER_148_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_567 ();
 DECAPx2_ASAP7_75t_R FILLER_148_586 ();
 DECAPx1_ASAP7_75t_R FILLER_148_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_622 ();
 DECAPx6_ASAP7_75t_R FILLER_148_626 ();
 FILLER_ASAP7_75t_R FILLER_148_640 ();
 DECAPx4_ASAP7_75t_R FILLER_148_648 ();
 FILLER_ASAP7_75t_R FILLER_148_658 ();
 DECAPx2_ASAP7_75t_R FILLER_148_680 ();
 FILLER_ASAP7_75t_R FILLER_148_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_699 ();
 FILLER_ASAP7_75t_R FILLER_148_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_729 ();
 FILLER_ASAP7_75t_R FILLER_148_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_746 ();
 FILLER_ASAP7_75t_R FILLER_148_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_755 ();
 FILLER_ASAP7_75t_R FILLER_148_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_772 ();
 DECAPx1_ASAP7_75t_R FILLER_148_784 ();
 DECAPx4_ASAP7_75t_R FILLER_148_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_808 ();
 DECAPx2_ASAP7_75t_R FILLER_148_841 ();
 DECAPx4_ASAP7_75t_R FILLER_148_854 ();
 DECAPx4_ASAP7_75t_R FILLER_148_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_893 ();
 DECAPx2_ASAP7_75t_R FILLER_148_905 ();
 FILLER_ASAP7_75t_R FILLER_148_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_913 ();
 FILLER_ASAP7_75t_R FILLER_148_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_930 ();
 DECAPx4_ASAP7_75t_R FILLER_148_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_948 ();
 DECAPx4_ASAP7_75t_R FILLER_148_961 ();
 DECAPx6_ASAP7_75t_R FILLER_148_983 ();
 DECAPx2_ASAP7_75t_R FILLER_148_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1016 ();
 FILLER_ASAP7_75t_R FILLER_148_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1040 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1061 ();
 FILLER_ASAP7_75t_R FILLER_148_1071 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1109 ();
 FILLER_ASAP7_75t_R FILLER_148_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1137 ();
 FILLER_ASAP7_75t_R FILLER_148_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1145 ();
 FILLER_ASAP7_75t_R FILLER_148_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1151 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1169 ();
 FILLER_ASAP7_75t_R FILLER_148_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1208 ();
 DECAPx1_ASAP7_75t_R FILLER_148_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1235 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1243 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1252 ();
 FILLER_ASAP7_75t_R FILLER_148_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1281 ();
 FILLER_ASAP7_75t_R FILLER_148_1287 ();
 FILLER_ASAP7_75t_R FILLER_148_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1301 ();
 FILLER_ASAP7_75t_R FILLER_148_1305 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1310 ();
 FILLER_ASAP7_75t_R FILLER_148_1316 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1318 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1378 ();
 FILLER_ASAP7_75t_R FILLER_148_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_148_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_149_2 ();
 FILLER_ASAP7_75t_R FILLER_149_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_14 ();
 FILLER_ASAP7_75t_R FILLER_149_18 ();
 FILLER_ASAP7_75t_R FILLER_149_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_52 ();
 DECAPx1_ASAP7_75t_R FILLER_149_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_157 ();
 DECAPx6_ASAP7_75t_R FILLER_149_165 ();
 DECAPx1_ASAP7_75t_R FILLER_149_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_209 ();
 FILLER_ASAP7_75t_R FILLER_149_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_226 ();
 DECAPx1_ASAP7_75t_R FILLER_149_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_263 ();
 DECAPx10_ASAP7_75t_R FILLER_149_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_300 ();
 FILLER_ASAP7_75t_R FILLER_149_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_339 ();
 DECAPx2_ASAP7_75t_R FILLER_149_366 ();
 FILLER_ASAP7_75t_R FILLER_149_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_408 ();
 FILLER_ASAP7_75t_R FILLER_149_412 ();
 FILLER_ASAP7_75t_R FILLER_149_432 ();
 DECAPx4_ASAP7_75t_R FILLER_149_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_450 ();
 DECAPx6_ASAP7_75t_R FILLER_149_469 ();
 DECAPx1_ASAP7_75t_R FILLER_149_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_558 ();
 DECAPx10_ASAP7_75t_R FILLER_149_633 ();
 DECAPx10_ASAP7_75t_R FILLER_149_655 ();
 DECAPx4_ASAP7_75t_R FILLER_149_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_687 ();
 FILLER_ASAP7_75t_R FILLER_149_698 ();
 DECAPx2_ASAP7_75t_R FILLER_149_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_721 ();
 DECAPx10_ASAP7_75t_R FILLER_149_728 ();
 DECAPx4_ASAP7_75t_R FILLER_149_762 ();
 FILLER_ASAP7_75t_R FILLER_149_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_774 ();
 DECAPx4_ASAP7_75t_R FILLER_149_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_793 ();
 DECAPx4_ASAP7_75t_R FILLER_149_804 ();
 FILLER_ASAP7_75t_R FILLER_149_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_822 ();
 DECAPx1_ASAP7_75t_R FILLER_149_829 ();
 DECAPx2_ASAP7_75t_R FILLER_149_843 ();
 DECAPx6_ASAP7_75t_R FILLER_149_858 ();
 FILLER_ASAP7_75t_R FILLER_149_872 ();
 FILLER_ASAP7_75t_R FILLER_149_886 ();
 DECAPx2_ASAP7_75t_R FILLER_149_905 ();
 DECAPx2_ASAP7_75t_R FILLER_149_918 ();
 DECAPx2_ASAP7_75t_R FILLER_149_933 ();
 DECAPx4_ASAP7_75t_R FILLER_149_946 ();
 DECAPx2_ASAP7_75t_R FILLER_149_962 ();
 FILLER_ASAP7_75t_R FILLER_149_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_970 ();
 DECAPx6_ASAP7_75t_R FILLER_149_977 ();
 DECAPx2_ASAP7_75t_R FILLER_149_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1024 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_149_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1055 ();
 DECAPx1_ASAP7_75t_R FILLER_149_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1154 ();
 FILLER_ASAP7_75t_R FILLER_149_1165 ();
 FILLER_ASAP7_75t_R FILLER_149_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_149_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1206 ();
 FILLER_ASAP7_75t_R FILLER_149_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1270 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1306 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1312 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1364 ();
 DECAPx4_ASAP7_75t_R FILLER_150_2 ();
 FILLER_ASAP7_75t_R FILLER_150_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_14 ();
 FILLER_ASAP7_75t_R FILLER_150_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_20 ();
 DECAPx2_ASAP7_75t_R FILLER_150_31 ();
 FILLER_ASAP7_75t_R FILLER_150_37 ();
 FILLER_ASAP7_75t_R FILLER_150_42 ();
 DECAPx2_ASAP7_75t_R FILLER_150_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_56 ();
 FILLER_ASAP7_75t_R FILLER_150_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_66 ();
 DECAPx6_ASAP7_75t_R FILLER_150_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_84 ();
 FILLER_ASAP7_75t_R FILLER_150_99 ();
 DECAPx1_ASAP7_75t_R FILLER_150_112 ();
 DECAPx4_ASAP7_75t_R FILLER_150_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_129 ();
 DECAPx4_ASAP7_75t_R FILLER_150_148 ();
 FILLER_ASAP7_75t_R FILLER_150_158 ();
 DECAPx2_ASAP7_75t_R FILLER_150_172 ();
 DECAPx2_ASAP7_75t_R FILLER_150_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_197 ();
 DECAPx2_ASAP7_75t_R FILLER_150_201 ();
 FILLER_ASAP7_75t_R FILLER_150_219 ();
 DECAPx2_ASAP7_75t_R FILLER_150_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_241 ();
 DECAPx6_ASAP7_75t_R FILLER_150_251 ();
 DECAPx2_ASAP7_75t_R FILLER_150_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_271 ();
 DECAPx2_ASAP7_75t_R FILLER_150_278 ();
 FILLER_ASAP7_75t_R FILLER_150_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_286 ();
 DECAPx6_ASAP7_75t_R FILLER_150_293 ();
 DECAPx2_ASAP7_75t_R FILLER_150_307 ();
 FILLER_ASAP7_75t_R FILLER_150_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_357 ();
 DECAPx4_ASAP7_75t_R FILLER_150_361 ();
 FILLER_ASAP7_75t_R FILLER_150_371 ();
 DECAPx6_ASAP7_75t_R FILLER_150_379 ();
 DECAPx6_ASAP7_75t_R FILLER_150_445 ();
 FILLER_ASAP7_75t_R FILLER_150_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_461 ();
 DECAPx2_ASAP7_75t_R FILLER_150_464 ();
 DECAPx1_ASAP7_75t_R FILLER_150_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_492 ();
 FILLER_ASAP7_75t_R FILLER_150_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_502 ();
 FILLER_ASAP7_75t_R FILLER_150_506 ();
 DECAPx6_ASAP7_75t_R FILLER_150_512 ();
 DECAPx1_ASAP7_75t_R FILLER_150_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_530 ();
 DECAPx2_ASAP7_75t_R FILLER_150_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_580 ();
 DECAPx1_ASAP7_75t_R FILLER_150_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_607 ();
 DECAPx2_ASAP7_75t_R FILLER_150_616 ();
 DECAPx6_ASAP7_75t_R FILLER_150_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_639 ();
 DECAPx2_ASAP7_75t_R FILLER_150_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_664 ();
 DECAPx1_ASAP7_75t_R FILLER_150_683 ();
 DECAPx1_ASAP7_75t_R FILLER_150_697 ();
 DECAPx1_ASAP7_75t_R FILLER_150_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_727 ();
 DECAPx6_ASAP7_75t_R FILLER_150_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_752 ();
 DECAPx2_ASAP7_75t_R FILLER_150_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_781 ();
 DECAPx2_ASAP7_75t_R FILLER_150_788 ();
 DECAPx2_ASAP7_75t_R FILLER_150_802 ();
 FILLER_ASAP7_75t_R FILLER_150_816 ();
 DECAPx2_ASAP7_75t_R FILLER_150_825 ();
 DECAPx1_ASAP7_75t_R FILLER_150_841 ();
 DECAPx1_ASAP7_75t_R FILLER_150_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_874 ();
 DECAPx2_ASAP7_75t_R FILLER_150_909 ();
 FILLER_ASAP7_75t_R FILLER_150_915 ();
 DECAPx1_ASAP7_75t_R FILLER_150_932 ();
 DECAPx2_ASAP7_75t_R FILLER_150_950 ();
 DECAPx1_ASAP7_75t_R FILLER_150_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_973 ();
 DECAPx4_ASAP7_75t_R FILLER_150_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_150_1015 ();
 FILLER_ASAP7_75t_R FILLER_150_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1027 ();
 FILLER_ASAP7_75t_R FILLER_150_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1052 ();
 DECAPx4_ASAP7_75t_R FILLER_150_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1096 ();
 FILLER_ASAP7_75t_R FILLER_150_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1112 ();
 DECAPx4_ASAP7_75t_R FILLER_150_1136 ();
 FILLER_ASAP7_75t_R FILLER_150_1146 ();
 FILLER_ASAP7_75t_R FILLER_150_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1162 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1184 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1229 ();
 FILLER_ASAP7_75t_R FILLER_150_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1250 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1272 ();
 DECAPx4_ASAP7_75t_R FILLER_150_1280 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1362 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_151_34 ();
 FILLER_ASAP7_75t_R FILLER_151_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_42 ();
 DECAPx2_ASAP7_75t_R FILLER_151_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_61 ();
 DECAPx2_ASAP7_75t_R FILLER_151_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_71 ();
 DECAPx2_ASAP7_75t_R FILLER_151_76 ();
 DECAPx1_ASAP7_75t_R FILLER_151_100 ();
 DECAPx10_ASAP7_75t_R FILLER_151_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_132 ();
 FILLER_ASAP7_75t_R FILLER_151_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_141 ();
 DECAPx6_ASAP7_75t_R FILLER_151_145 ();
 DECAPx1_ASAP7_75t_R FILLER_151_159 ();
 DECAPx10_ASAP7_75t_R FILLER_151_189 ();
 DECAPx2_ASAP7_75t_R FILLER_151_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_217 ();
 DECAPx6_ASAP7_75t_R FILLER_151_226 ();
 FILLER_ASAP7_75t_R FILLER_151_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_242 ();
 FILLER_ASAP7_75t_R FILLER_151_269 ();
 DECAPx1_ASAP7_75t_R FILLER_151_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_322 ();
 DECAPx1_ASAP7_75t_R FILLER_151_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_333 ();
 DECAPx1_ASAP7_75t_R FILLER_151_337 ();
 DECAPx4_ASAP7_75t_R FILLER_151_344 ();
 FILLER_ASAP7_75t_R FILLER_151_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_356 ();
 DECAPx4_ASAP7_75t_R FILLER_151_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_373 ();
 DECAPx2_ASAP7_75t_R FILLER_151_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_386 ();
 FILLER_ASAP7_75t_R FILLER_151_390 ();
 FILLER_ASAP7_75t_R FILLER_151_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_397 ();
 DECAPx4_ASAP7_75t_R FILLER_151_404 ();
 FILLER_ASAP7_75t_R FILLER_151_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_416 ();
 DECAPx10_ASAP7_75t_R FILLER_151_429 ();
 FILLER_ASAP7_75t_R FILLER_151_451 ();
 DECAPx4_ASAP7_75t_R FILLER_151_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_481 ();
 DECAPx6_ASAP7_75t_R FILLER_151_498 ();
 FILLER_ASAP7_75t_R FILLER_151_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_514 ();
 DECAPx10_ASAP7_75t_R FILLER_151_533 ();
 DECAPx2_ASAP7_75t_R FILLER_151_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_561 ();
 DECAPx1_ASAP7_75t_R FILLER_151_580 ();
 DECAPx1_ASAP7_75t_R FILLER_151_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_598 ();
 DECAPx4_ASAP7_75t_R FILLER_151_615 ();
 FILLER_ASAP7_75t_R FILLER_151_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_627 ();
 DECAPx2_ASAP7_75t_R FILLER_151_666 ();
 FILLER_ASAP7_75t_R FILLER_151_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_706 ();
 DECAPx6_ASAP7_75t_R FILLER_151_726 ();
 FILLER_ASAP7_75t_R FILLER_151_740 ();
 FILLER_ASAP7_75t_R FILLER_151_748 ();
 FILLER_ASAP7_75t_R FILLER_151_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_770 ();
 DECAPx1_ASAP7_75t_R FILLER_151_783 ();
 FILLER_ASAP7_75t_R FILLER_151_805 ();
 DECAPx2_ASAP7_75t_R FILLER_151_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_821 ();
 FILLER_ASAP7_75t_R FILLER_151_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_834 ();
 DECAPx6_ASAP7_75t_R FILLER_151_841 ();
 DECAPx4_ASAP7_75t_R FILLER_151_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_879 ();
 DECAPx1_ASAP7_75t_R FILLER_151_890 ();
 DECAPx2_ASAP7_75t_R FILLER_151_908 ();
 FILLER_ASAP7_75t_R FILLER_151_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_916 ();
 DECAPx4_ASAP7_75t_R FILLER_151_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_936 ();
 DECAPx4_ASAP7_75t_R FILLER_151_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_953 ();
 DECAPx1_ASAP7_75t_R FILLER_151_964 ();
 DECAPx1_ASAP7_75t_R FILLER_151_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_986 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1000 ();
 FILLER_ASAP7_75t_R FILLER_151_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1026 ();
 FILLER_ASAP7_75t_R FILLER_151_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1054 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1111 ();
 FILLER_ASAP7_75t_R FILLER_151_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1142 ();
 FILLER_ASAP7_75t_R FILLER_151_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1202 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1214 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1221 ();
 FILLER_ASAP7_75t_R FILLER_151_1231 ();
 FILLER_ASAP7_75t_R FILLER_151_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1305 ();
 FILLER_ASAP7_75t_R FILLER_151_1309 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1315 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1322 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_152_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_24 ();
 DECAPx6_ASAP7_75t_R FILLER_152_31 ();
 FILLER_ASAP7_75t_R FILLER_152_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_47 ();
 DECAPx4_ASAP7_75t_R FILLER_152_74 ();
 FILLER_ASAP7_75t_R FILLER_152_84 ();
 DECAPx2_ASAP7_75t_R FILLER_152_112 ();
 DECAPx6_ASAP7_75t_R FILLER_152_121 ();
 DECAPx2_ASAP7_75t_R FILLER_152_135 ();
 DECAPx2_ASAP7_75t_R FILLER_152_155 ();
 FILLER_ASAP7_75t_R FILLER_152_161 ();
 FILLER_ASAP7_75t_R FILLER_152_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_183 ();
 DECAPx2_ASAP7_75t_R FILLER_152_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_201 ();
 DECAPx4_ASAP7_75t_R FILLER_152_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_230 ();
 DECAPx1_ASAP7_75t_R FILLER_152_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_245 ();
 FILLER_ASAP7_75t_R FILLER_152_254 ();
 DECAPx1_ASAP7_75t_R FILLER_152_289 ();
 DECAPx10_ASAP7_75t_R FILLER_152_296 ();
 DECAPx6_ASAP7_75t_R FILLER_152_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_332 ();
 DECAPx2_ASAP7_75t_R FILLER_152_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_353 ();
 DECAPx2_ASAP7_75t_R FILLER_152_362 ();
 DECAPx10_ASAP7_75t_R FILLER_152_374 ();
 DECAPx6_ASAP7_75t_R FILLER_152_396 ();
 FILLER_ASAP7_75t_R FILLER_152_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_430 ();
 DECAPx4_ASAP7_75t_R FILLER_152_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_449 ();
 FILLER_ASAP7_75t_R FILLER_152_460 ();
 FILLER_ASAP7_75t_R FILLER_152_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_478 ();
 DECAPx2_ASAP7_75t_R FILLER_152_489 ();
 DECAPx2_ASAP7_75t_R FILLER_152_513 ();
 FILLER_ASAP7_75t_R FILLER_152_519 ();
 DECAPx10_ASAP7_75t_R FILLER_152_539 ();
 DECAPx2_ASAP7_75t_R FILLER_152_561 ();
 FILLER_ASAP7_75t_R FILLER_152_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_569 ();
 DECAPx2_ASAP7_75t_R FILLER_152_598 ();
 DECAPx10_ASAP7_75t_R FILLER_152_610 ();
 DECAPx6_ASAP7_75t_R FILLER_152_632 ();
 DECAPx2_ASAP7_75t_R FILLER_152_646 ();
 DECAPx2_ASAP7_75t_R FILLER_152_658 ();
 FILLER_ASAP7_75t_R FILLER_152_664 ();
 DECAPx1_ASAP7_75t_R FILLER_152_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_733 ();
 DECAPx2_ASAP7_75t_R FILLER_152_750 ();
 FILLER_ASAP7_75t_R FILLER_152_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_758 ();
 DECAPx2_ASAP7_75t_R FILLER_152_766 ();
 DECAPx10_ASAP7_75t_R FILLER_152_779 ();
 DECAPx2_ASAP7_75t_R FILLER_152_801 ();
 FILLER_ASAP7_75t_R FILLER_152_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_809 ();
 DECAPx4_ASAP7_75t_R FILLER_152_818 ();
 FILLER_ASAP7_75t_R FILLER_152_828 ();
 FILLER_ASAP7_75t_R FILLER_152_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_838 ();
 DECAPx6_ASAP7_75t_R FILLER_152_849 ();
 DECAPx2_ASAP7_75t_R FILLER_152_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_869 ();
 DECAPx6_ASAP7_75t_R FILLER_152_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_889 ();
 DECAPx1_ASAP7_75t_R FILLER_152_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_901 ();
 FILLER_ASAP7_75t_R FILLER_152_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_992 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1000 ();
 FILLER_ASAP7_75t_R FILLER_152_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1052 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1074 ();
 FILLER_ASAP7_75t_R FILLER_152_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1097 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1119 ();
 FILLER_ASAP7_75t_R FILLER_152_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1141 ();
 FILLER_ASAP7_75t_R FILLER_152_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1201 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1233 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1245 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1259 ();
 FILLER_ASAP7_75t_R FILLER_152_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1276 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1391 ();
 FILLER_ASAP7_75t_R FILLER_153_2 ();
 DECAPx2_ASAP7_75t_R FILLER_153_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_40 ();
 DECAPx6_ASAP7_75t_R FILLER_153_59 ();
 DECAPx2_ASAP7_75t_R FILLER_153_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_103 ();
 DECAPx6_ASAP7_75t_R FILLER_153_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_176 ();
 DECAPx1_ASAP7_75t_R FILLER_153_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_213 ();
 DECAPx6_ASAP7_75t_R FILLER_153_227 ();
 DECAPx1_ASAP7_75t_R FILLER_153_241 ();
 DECAPx2_ASAP7_75t_R FILLER_153_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_257 ();
 FILLER_ASAP7_75t_R FILLER_153_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_263 ();
 DECAPx4_ASAP7_75t_R FILLER_153_272 ();
 DECAPx6_ASAP7_75t_R FILLER_153_290 ();
 DECAPx1_ASAP7_75t_R FILLER_153_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_334 ();
 FILLER_ASAP7_75t_R FILLER_153_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_351 ();
 FILLER_ASAP7_75t_R FILLER_153_366 ();
 DECAPx2_ASAP7_75t_R FILLER_153_382 ();
 FILLER_ASAP7_75t_R FILLER_153_388 ();
 DECAPx4_ASAP7_75t_R FILLER_153_404 ();
 FILLER_ASAP7_75t_R FILLER_153_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_448 ();
 DECAPx6_ASAP7_75t_R FILLER_153_455 ();
 FILLER_ASAP7_75t_R FILLER_153_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_471 ();
 DECAPx6_ASAP7_75t_R FILLER_153_482 ();
 FILLER_ASAP7_75t_R FILLER_153_496 ();
 DECAPx2_ASAP7_75t_R FILLER_153_516 ();
 DECAPx10_ASAP7_75t_R FILLER_153_554 ();
 DECAPx4_ASAP7_75t_R FILLER_153_576 ();
 FILLER_ASAP7_75t_R FILLER_153_586 ();
 DECAPx1_ASAP7_75t_R FILLER_153_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_602 ();
 DECAPx6_ASAP7_75t_R FILLER_153_629 ();
 DECAPx1_ASAP7_75t_R FILLER_153_643 ();
 DECAPx2_ASAP7_75t_R FILLER_153_659 ();
 FILLER_ASAP7_75t_R FILLER_153_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_682 ();
 FILLER_ASAP7_75t_R FILLER_153_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_715 ();
 FILLER_ASAP7_75t_R FILLER_153_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_730 ();
 DECAPx6_ASAP7_75t_R FILLER_153_739 ();
 FILLER_ASAP7_75t_R FILLER_153_753 ();
 DECAPx6_ASAP7_75t_R FILLER_153_761 ();
 FILLER_ASAP7_75t_R FILLER_153_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_794 ();
 FILLER_ASAP7_75t_R FILLER_153_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_834 ();
 FILLER_ASAP7_75t_R FILLER_153_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_853 ();
 DECAPx4_ASAP7_75t_R FILLER_153_859 ();
 DECAPx2_ASAP7_75t_R FILLER_153_879 ();
 FILLER_ASAP7_75t_R FILLER_153_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_887 ();
 FILLER_ASAP7_75t_R FILLER_153_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_898 ();
 FILLER_ASAP7_75t_R FILLER_153_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_915 ();
 DECAPx1_ASAP7_75t_R FILLER_153_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_940 ();
 DECAPx6_ASAP7_75t_R FILLER_153_955 ();
 FILLER_ASAP7_75t_R FILLER_153_969 ();
 DECAPx2_ASAP7_75t_R FILLER_153_978 ();
 FILLER_ASAP7_75t_R FILLER_153_984 ();
 DECAPx4_ASAP7_75t_R FILLER_153_1000 ();
 FILLER_ASAP7_75t_R FILLER_153_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1032 ();
 DECAPx6_ASAP7_75t_R FILLER_153_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1074 ();
 DECAPx6_ASAP7_75t_R FILLER_153_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1124 ();
 FILLER_ASAP7_75t_R FILLER_153_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1159 ();
 FILLER_ASAP7_75t_R FILLER_153_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1204 ();
 FILLER_ASAP7_75t_R FILLER_153_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1213 ();
 DECAPx4_ASAP7_75t_R FILLER_153_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1285 ();
 DECAPx4_ASAP7_75t_R FILLER_153_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1324 ();
 FILLER_ASAP7_75t_R FILLER_153_1330 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1332 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_154_2 ();
 FILLER_ASAP7_75t_R FILLER_154_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_18 ();
 FILLER_ASAP7_75t_R FILLER_154_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_24 ();
 DECAPx6_ASAP7_75t_R FILLER_154_31 ();
 FILLER_ASAP7_75t_R FILLER_154_63 ();
 DECAPx4_ASAP7_75t_R FILLER_154_78 ();
 DECAPx1_ASAP7_75t_R FILLER_154_96 ();
 DECAPx2_ASAP7_75t_R FILLER_154_103 ();
 FILLER_ASAP7_75t_R FILLER_154_109 ();
 DECAPx1_ASAP7_75t_R FILLER_154_119 ();
 FILLER_ASAP7_75t_R FILLER_154_149 ();
 DECAPx4_ASAP7_75t_R FILLER_154_154 ();
 DECAPx6_ASAP7_75t_R FILLER_154_192 ();
 FILLER_ASAP7_75t_R FILLER_154_206 ();
 FILLER_ASAP7_75t_R FILLER_154_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_236 ();
 FILLER_ASAP7_75t_R FILLER_154_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_245 ();
 DECAPx4_ASAP7_75t_R FILLER_154_252 ();
 FILLER_ASAP7_75t_R FILLER_154_262 ();
 DECAPx1_ASAP7_75t_R FILLER_154_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_274 ();
 FILLER_ASAP7_75t_R FILLER_154_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_303 ();
 DECAPx1_ASAP7_75t_R FILLER_154_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_335 ();
 DECAPx2_ASAP7_75t_R FILLER_154_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_348 ();
 FILLER_ASAP7_75t_R FILLER_154_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_363 ();
 DECAPx1_ASAP7_75t_R FILLER_154_372 ();
 FILLER_ASAP7_75t_R FILLER_154_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_386 ();
 DECAPx2_ASAP7_75t_R FILLER_154_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_413 ();
 FILLER_ASAP7_75t_R FILLER_154_432 ();
 FILLER_ASAP7_75t_R FILLER_154_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_442 ();
 FILLER_ASAP7_75t_R FILLER_154_460 ();
 DECAPx4_ASAP7_75t_R FILLER_154_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_474 ();
 DECAPx4_ASAP7_75t_R FILLER_154_483 ();
 FILLER_ASAP7_75t_R FILLER_154_505 ();
 DECAPx2_ASAP7_75t_R FILLER_154_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_540 ();
 DECAPx1_ASAP7_75t_R FILLER_154_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_570 ();
 DECAPx4_ASAP7_75t_R FILLER_154_589 ();
 DECAPx2_ASAP7_75t_R FILLER_154_651 ();
 FILLER_ASAP7_75t_R FILLER_154_657 ();
 FILLER_ASAP7_75t_R FILLER_154_662 ();
 DECAPx2_ASAP7_75t_R FILLER_154_672 ();
 FILLER_ASAP7_75t_R FILLER_154_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_716 ();
 DECAPx4_ASAP7_75t_R FILLER_154_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_733 ();
 FILLER_ASAP7_75t_R FILLER_154_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_750 ();
 DECAPx1_ASAP7_75t_R FILLER_154_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_774 ();
 DECAPx2_ASAP7_75t_R FILLER_154_781 ();
 FILLER_ASAP7_75t_R FILLER_154_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_795 ();
 DECAPx2_ASAP7_75t_R FILLER_154_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_809 ();
 DECAPx6_ASAP7_75t_R FILLER_154_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_830 ();
 FILLER_ASAP7_75t_R FILLER_154_837 ();
 DECAPx2_ASAP7_75t_R FILLER_154_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_855 ();
 FILLER_ASAP7_75t_R FILLER_154_862 ();
 DECAPx6_ASAP7_75t_R FILLER_154_883 ();
 DECAPx2_ASAP7_75t_R FILLER_154_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_903 ();
 DECAPx6_ASAP7_75t_R FILLER_154_920 ();
 DECAPx1_ASAP7_75t_R FILLER_154_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_938 ();
 DECAPx1_ASAP7_75t_R FILLER_154_946 ();
 DECAPx6_ASAP7_75t_R FILLER_154_970 ();
 FILLER_ASAP7_75t_R FILLER_154_984 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1049 ();
 FILLER_ASAP7_75t_R FILLER_154_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1088 ();
 FILLER_ASAP7_75t_R FILLER_154_1094 ();
 FILLER_ASAP7_75t_R FILLER_154_1125 ();
 FILLER_ASAP7_75t_R FILLER_154_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1146 ();
 FILLER_ASAP7_75t_R FILLER_154_1152 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1171 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1232 ();
 FILLER_ASAP7_75t_R FILLER_154_1262 ();
 FILLER_ASAP7_75t_R FILLER_154_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1328 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1355 ();
 FILLER_ASAP7_75t_R FILLER_154_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1363 ();
 FILLER_ASAP7_75t_R FILLER_154_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_155_2 ();
 FILLER_ASAP7_75t_R FILLER_155_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_14 ();
 DECAPx4_ASAP7_75t_R FILLER_155_33 ();
 DECAPx2_ASAP7_75t_R FILLER_155_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_59 ();
 DECAPx4_ASAP7_75t_R FILLER_155_90 ();
 FILLER_ASAP7_75t_R FILLER_155_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_102 ();
 DECAPx1_ASAP7_75t_R FILLER_155_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_117 ();
 DECAPx2_ASAP7_75t_R FILLER_155_132 ();
 DECAPx10_ASAP7_75t_R FILLER_155_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_163 ();
 DECAPx10_ASAP7_75t_R FILLER_155_182 ();
 DECAPx1_ASAP7_75t_R FILLER_155_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_208 ();
 DECAPx1_ASAP7_75t_R FILLER_155_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_226 ();
 DECAPx2_ASAP7_75t_R FILLER_155_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_259 ();
 DECAPx6_ASAP7_75t_R FILLER_155_268 ();
 DECAPx1_ASAP7_75t_R FILLER_155_282 ();
 DECAPx6_ASAP7_75t_R FILLER_155_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_309 ();
 DECAPx6_ASAP7_75t_R FILLER_155_318 ();
 DECAPx1_ASAP7_75t_R FILLER_155_332 ();
 DECAPx2_ASAP7_75t_R FILLER_155_360 ();
 DECAPx6_ASAP7_75t_R FILLER_155_404 ();
 DECAPx2_ASAP7_75t_R FILLER_155_418 ();
 DECAPx10_ASAP7_75t_R FILLER_155_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_468 ();
 DECAPx10_ASAP7_75t_R FILLER_155_487 ();
 DECAPx2_ASAP7_75t_R FILLER_155_509 ();
 FILLER_ASAP7_75t_R FILLER_155_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_528 ();
 DECAPx2_ASAP7_75t_R FILLER_155_535 ();
 DECAPx1_ASAP7_75t_R FILLER_155_547 ();
 DECAPx6_ASAP7_75t_R FILLER_155_559 ();
 FILLER_ASAP7_75t_R FILLER_155_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_575 ();
 DECAPx1_ASAP7_75t_R FILLER_155_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_606 ();
 FILLER_ASAP7_75t_R FILLER_155_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_621 ();
 DECAPx6_ASAP7_75t_R FILLER_155_625 ();
 FILLER_ASAP7_75t_R FILLER_155_639 ();
 DECAPx1_ASAP7_75t_R FILLER_155_653 ();
 FILLER_ASAP7_75t_R FILLER_155_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_678 ();
 FILLER_ASAP7_75t_R FILLER_155_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_715 ();
 DECAPx2_ASAP7_75t_R FILLER_155_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_730 ();
 DECAPx1_ASAP7_75t_R FILLER_155_739 ();
 DECAPx6_ASAP7_75t_R FILLER_155_769 ();
 FILLER_ASAP7_75t_R FILLER_155_783 ();
 DECAPx4_ASAP7_75t_R FILLER_155_797 ();
 FILLER_ASAP7_75t_R FILLER_155_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_809 ();
 DECAPx4_ASAP7_75t_R FILLER_155_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_833 ();
 DECAPx2_ASAP7_75t_R FILLER_155_846 ();
 FILLER_ASAP7_75t_R FILLER_155_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_854 ();
 DECAPx10_ASAP7_75t_R FILLER_155_871 ();
 DECAPx6_ASAP7_75t_R FILLER_155_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_907 ();
 DECAPx4_ASAP7_75t_R FILLER_155_926 ();
 DECAPx2_ASAP7_75t_R FILLER_155_950 ();
 DECAPx1_ASAP7_75t_R FILLER_155_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_977 ();
 DECAPx2_ASAP7_75t_R FILLER_155_998 ();
 FILLER_ASAP7_75t_R FILLER_155_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_155_1028 ();
 FILLER_ASAP7_75t_R FILLER_155_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1139 ();
 FILLER_ASAP7_75t_R FILLER_155_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1162 ();
 FILLER_ASAP7_75t_R FILLER_155_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1178 ();
 FILLER_ASAP7_75t_R FILLER_155_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1192 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1196 ();
 FILLER_ASAP7_75t_R FILLER_155_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1215 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1222 ();
 FILLER_ASAP7_75t_R FILLER_155_1236 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1248 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1288 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1313 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1327 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1337 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1351 ();
 FILLER_ASAP7_75t_R FILLER_155_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1359 ();
 DECAPx10_ASAP7_75t_R FILLER_156_2 ();
 DECAPx10_ASAP7_75t_R FILLER_156_24 ();
 FILLER_ASAP7_75t_R FILLER_156_46 ();
 FILLER_ASAP7_75t_R FILLER_156_58 ();
 DECAPx10_ASAP7_75t_R FILLER_156_72 ();
 DECAPx2_ASAP7_75t_R FILLER_156_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_100 ();
 DECAPx1_ASAP7_75t_R FILLER_156_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_123 ();
 DECAPx6_ASAP7_75t_R FILLER_156_152 ();
 FILLER_ASAP7_75t_R FILLER_156_166 ();
 FILLER_ASAP7_75t_R FILLER_156_203 ();
 DECAPx6_ASAP7_75t_R FILLER_156_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_229 ();
 DECAPx1_ASAP7_75t_R FILLER_156_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_241 ();
 FILLER_ASAP7_75t_R FILLER_156_245 ();
 DECAPx10_ASAP7_75t_R FILLER_156_279 ();
 DECAPx2_ASAP7_75t_R FILLER_156_301 ();
 FILLER_ASAP7_75t_R FILLER_156_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_309 ();
 DECAPx6_ASAP7_75t_R FILLER_156_316 ();
 DECAPx2_ASAP7_75t_R FILLER_156_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_336 ();
 DECAPx1_ASAP7_75t_R FILLER_156_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_374 ();
 DECAPx2_ASAP7_75t_R FILLER_156_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_390 ();
 DECAPx10_ASAP7_75t_R FILLER_156_397 ();
 DECAPx4_ASAP7_75t_R FILLER_156_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_429 ();
 DECAPx6_ASAP7_75t_R FILLER_156_442 ();
 DECAPx2_ASAP7_75t_R FILLER_156_456 ();
 DECAPx1_ASAP7_75t_R FILLER_156_464 ();
 DECAPx1_ASAP7_75t_R FILLER_156_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_508 ();
 DECAPx10_ASAP7_75t_R FILLER_156_527 ();
 DECAPx6_ASAP7_75t_R FILLER_156_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_563 ();
 DECAPx1_ASAP7_75t_R FILLER_156_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_578 ();
 DECAPx1_ASAP7_75t_R FILLER_156_587 ();
 DECAPx4_ASAP7_75t_R FILLER_156_594 ();
 FILLER_ASAP7_75t_R FILLER_156_604 ();
 DECAPx4_ASAP7_75t_R FILLER_156_618 ();
 FILLER_ASAP7_75t_R FILLER_156_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_630 ();
 FILLER_ASAP7_75t_R FILLER_156_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_640 ();
 FILLER_ASAP7_75t_R FILLER_156_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_650 ();
 DECAPx1_ASAP7_75t_R FILLER_156_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_691 ();
 FILLER_ASAP7_75t_R FILLER_156_707 ();
 DECAPx6_ASAP7_75t_R FILLER_156_729 ();
 DECAPx1_ASAP7_75t_R FILLER_156_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_747 ();
 DECAPx10_ASAP7_75t_R FILLER_156_754 ();
 DECAPx4_ASAP7_75t_R FILLER_156_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_805 ();
 DECAPx6_ASAP7_75t_R FILLER_156_818 ();
 FILLER_ASAP7_75t_R FILLER_156_832 ();
 DECAPx4_ASAP7_75t_R FILLER_156_844 ();
 FILLER_ASAP7_75t_R FILLER_156_854 ();
 FILLER_ASAP7_75t_R FILLER_156_862 ();
 FILLER_ASAP7_75t_R FILLER_156_870 ();
 FILLER_ASAP7_75t_R FILLER_156_878 ();
 FILLER_ASAP7_75t_R FILLER_156_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_888 ();
 DECAPx10_ASAP7_75t_R FILLER_156_895 ();
 DECAPx1_ASAP7_75t_R FILLER_156_917 ();
 DECAPx10_ASAP7_75t_R FILLER_156_927 ();
 DECAPx1_ASAP7_75t_R FILLER_156_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_953 ();
 DECAPx2_ASAP7_75t_R FILLER_156_963 ();
 FILLER_ASAP7_75t_R FILLER_156_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_981 ();
 DECAPx2_ASAP7_75t_R FILLER_156_994 ();
 DECAPx6_ASAP7_75t_R FILLER_156_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_156_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1065 ();
 DECAPx6_ASAP7_75t_R FILLER_156_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1109 ();
 FILLER_ASAP7_75t_R FILLER_156_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1130 ();
 FILLER_ASAP7_75t_R FILLER_156_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1142 ();
 FILLER_ASAP7_75t_R FILLER_156_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1161 ();
 FILLER_ASAP7_75t_R FILLER_156_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1205 ();
 FILLER_ASAP7_75t_R FILLER_156_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1243 ();
 FILLER_ASAP7_75t_R FILLER_156_1249 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1261 ();
 FILLER_ASAP7_75t_R FILLER_156_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_156_1301 ();
 DECAPx6_ASAP7_75t_R FILLER_156_1323 ();
 FILLER_ASAP7_75t_R FILLER_156_1337 ();
 DECAPx6_ASAP7_75t_R FILLER_156_1349 ();
 FILLER_ASAP7_75t_R FILLER_156_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_157_2 ();
 FILLER_ASAP7_75t_R FILLER_157_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_26 ();
 DECAPx2_ASAP7_75t_R FILLER_157_39 ();
 FILLER_ASAP7_75t_R FILLER_157_45 ();
 DECAPx10_ASAP7_75t_R FILLER_157_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_91 ();
 DECAPx6_ASAP7_75t_R FILLER_157_106 ();
 FILLER_ASAP7_75t_R FILLER_157_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_148 ();
 FILLER_ASAP7_75t_R FILLER_157_155 ();
 FILLER_ASAP7_75t_R FILLER_157_160 ();
 FILLER_ASAP7_75t_R FILLER_157_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_176 ();
 DECAPx2_ASAP7_75t_R FILLER_157_183 ();
 FILLER_ASAP7_75t_R FILLER_157_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_194 ();
 FILLER_ASAP7_75t_R FILLER_157_201 ();
 DECAPx10_ASAP7_75t_R FILLER_157_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_248 ();
 DECAPx4_ASAP7_75t_R FILLER_157_255 ();
 FILLER_ASAP7_75t_R FILLER_157_280 ();
 DECAPx4_ASAP7_75t_R FILLER_157_289 ();
 DECAPx2_ASAP7_75t_R FILLER_157_317 ();
 DECAPx1_ASAP7_75t_R FILLER_157_347 ();
 FILLER_ASAP7_75t_R FILLER_157_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_361 ();
 DECAPx10_ASAP7_75t_R FILLER_157_365 ();
 DECAPx6_ASAP7_75t_R FILLER_157_387 ();
 DECAPx2_ASAP7_75t_R FILLER_157_401 ();
 DECAPx2_ASAP7_75t_R FILLER_157_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_431 ();
 DECAPx4_ASAP7_75t_R FILLER_157_441 ();
 FILLER_ASAP7_75t_R FILLER_157_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_453 ();
 DECAPx2_ASAP7_75t_R FILLER_157_472 ();
 FILLER_ASAP7_75t_R FILLER_157_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_520 ();
 DECAPx2_ASAP7_75t_R FILLER_157_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_563 ();
 FILLER_ASAP7_75t_R FILLER_157_582 ();
 DECAPx4_ASAP7_75t_R FILLER_157_590 ();
 FILLER_ASAP7_75t_R FILLER_157_618 ();
 FILLER_ASAP7_75t_R FILLER_157_623 ();
 DECAPx4_ASAP7_75t_R FILLER_157_635 ();
 FILLER_ASAP7_75t_R FILLER_157_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_699 ();
 FILLER_ASAP7_75t_R FILLER_157_706 ();
 FILLER_ASAP7_75t_R FILLER_157_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_732 ();
 FILLER_ASAP7_75t_R FILLER_157_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_742 ();
 FILLER_ASAP7_75t_R FILLER_157_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_751 ();
 DECAPx2_ASAP7_75t_R FILLER_157_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_765 ();
 DECAPx1_ASAP7_75t_R FILLER_157_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_808 ();
 DECAPx2_ASAP7_75t_R FILLER_157_825 ();
 FILLER_ASAP7_75t_R FILLER_157_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_833 ();
 FILLER_ASAP7_75t_R FILLER_157_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_846 ();
 DECAPx1_ASAP7_75t_R FILLER_157_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_863 ();
 DECAPx1_ASAP7_75t_R FILLER_157_870 ();
 FILLER_ASAP7_75t_R FILLER_157_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_888 ();
 DECAPx2_ASAP7_75t_R FILLER_157_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_917 ();
 DECAPx4_ASAP7_75t_R FILLER_157_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_936 ();
 DECAPx1_ASAP7_75t_R FILLER_157_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_949 ();
 DECAPx4_ASAP7_75t_R FILLER_157_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_967 ();
 DECAPx1_ASAP7_75t_R FILLER_157_987 ();
 DECAPx4_ASAP7_75t_R FILLER_157_997 ();
 DECAPx4_ASAP7_75t_R FILLER_157_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_157_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_157_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_157_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_157_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1105 ();
 FILLER_ASAP7_75t_R FILLER_157_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1121 ();
 FILLER_ASAP7_75t_R FILLER_157_1130 ();
 DECAPx4_ASAP7_75t_R FILLER_157_1138 ();
 FILLER_ASAP7_75t_R FILLER_157_1148 ();
 DECAPx4_ASAP7_75t_R FILLER_157_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1211 ();
 FILLER_ASAP7_75t_R FILLER_157_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1305 ();
 FILLER_ASAP7_75t_R FILLER_157_1378 ();
 DECAPx4_ASAP7_75t_R FILLER_158_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_30 ();
 DECAPx6_ASAP7_75t_R FILLER_158_49 ();
 DECAPx2_ASAP7_75t_R FILLER_158_75 ();
 FILLER_ASAP7_75t_R FILLER_158_81 ();
 DECAPx2_ASAP7_75t_R FILLER_158_119 ();
 DECAPx1_ASAP7_75t_R FILLER_158_139 ();
 FILLER_ASAP7_75t_R FILLER_158_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_195 ();
 FILLER_ASAP7_75t_R FILLER_158_212 ();
 DECAPx2_ASAP7_75t_R FILLER_158_220 ();
 FILLER_ASAP7_75t_R FILLER_158_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_234 ();
 DECAPx6_ASAP7_75t_R FILLER_158_249 ();
 FILLER_ASAP7_75t_R FILLER_158_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_265 ();
 DECAPx4_ASAP7_75t_R FILLER_158_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_345 ();
 DECAPx2_ASAP7_75t_R FILLER_158_354 ();
 DECAPx2_ASAP7_75t_R FILLER_158_378 ();
 DECAPx1_ASAP7_75t_R FILLER_158_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_395 ();
 FILLER_ASAP7_75t_R FILLER_158_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_416 ();
 FILLER_ASAP7_75t_R FILLER_158_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_445 ();
 DECAPx1_ASAP7_75t_R FILLER_158_458 ();
 DECAPx10_ASAP7_75t_R FILLER_158_464 ();
 DECAPx10_ASAP7_75t_R FILLER_158_486 ();
 DECAPx10_ASAP7_75t_R FILLER_158_508 ();
 DECAPx6_ASAP7_75t_R FILLER_158_530 ();
 DECAPx1_ASAP7_75t_R FILLER_158_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_548 ();
 DECAPx4_ASAP7_75t_R FILLER_158_567 ();
 FILLER_ASAP7_75t_R FILLER_158_577 ();
 DECAPx2_ASAP7_75t_R FILLER_158_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_648 ();
 DECAPx4_ASAP7_75t_R FILLER_158_655 ();
 DECAPx4_ASAP7_75t_R FILLER_158_674 ();
 FILLER_ASAP7_75t_R FILLER_158_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_686 ();
 FILLER_ASAP7_75t_R FILLER_158_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_707 ();
 FILLER_ASAP7_75t_R FILLER_158_714 ();
 DECAPx6_ASAP7_75t_R FILLER_158_724 ();
 DECAPx1_ASAP7_75t_R FILLER_158_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_742 ();
 DECAPx2_ASAP7_75t_R FILLER_158_759 ();
 FILLER_ASAP7_75t_R FILLER_158_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_767 ();
 DECAPx6_ASAP7_75t_R FILLER_158_790 ();
 FILLER_ASAP7_75t_R FILLER_158_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_806 ();
 DECAPx2_ASAP7_75t_R FILLER_158_813 ();
 DECAPx6_ASAP7_75t_R FILLER_158_831 ();
 FILLER_ASAP7_75t_R FILLER_158_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_847 ();
 DECAPx1_ASAP7_75t_R FILLER_158_858 ();
 DECAPx2_ASAP7_75t_R FILLER_158_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_878 ();
 DECAPx6_ASAP7_75t_R FILLER_158_889 ();
 FILLER_ASAP7_75t_R FILLER_158_903 ();
 DECAPx2_ASAP7_75t_R FILLER_158_923 ();
 DECAPx1_ASAP7_75t_R FILLER_158_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_949 ();
 DECAPx2_ASAP7_75t_R FILLER_158_961 ();
 DECAPx6_ASAP7_75t_R FILLER_158_973 ();
 FILLER_ASAP7_75t_R FILLER_158_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_989 ();
 FILLER_ASAP7_75t_R FILLER_158_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1029 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1097 ();
 FILLER_ASAP7_75t_R FILLER_158_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1149 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1185 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1192 ();
 FILLER_ASAP7_75t_R FILLER_158_1199 ();
 FILLER_ASAP7_75t_R FILLER_158_1211 ();
 FILLER_ASAP7_75t_R FILLER_158_1227 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1232 ();
 FILLER_ASAP7_75t_R FILLER_158_1242 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1254 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1272 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1313 ();
 FILLER_ASAP7_75t_R FILLER_158_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1365 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1369 ();
 FILLER_ASAP7_75t_R FILLER_158_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_159_2 ();
 FILLER_ASAP7_75t_R FILLER_159_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_10 ();
 DECAPx1_ASAP7_75t_R FILLER_159_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_27 ();
 DECAPx1_ASAP7_75t_R FILLER_159_38 ();
 DECAPx2_ASAP7_75t_R FILLER_159_58 ();
 FILLER_ASAP7_75t_R FILLER_159_64 ();
 DECAPx10_ASAP7_75t_R FILLER_159_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_110 ();
 FILLER_ASAP7_75t_R FILLER_159_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_136 ();
 DECAPx1_ASAP7_75t_R FILLER_159_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_144 ();
 DECAPx6_ASAP7_75t_R FILLER_159_153 ();
 FILLER_ASAP7_75t_R FILLER_159_167 ();
 DECAPx1_ASAP7_75t_R FILLER_159_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_219 ();
 DECAPx4_ASAP7_75t_R FILLER_159_228 ();
 FILLER_ASAP7_75t_R FILLER_159_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_240 ();
 DECAPx6_ASAP7_75t_R FILLER_159_253 ();
 FILLER_ASAP7_75t_R FILLER_159_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_269 ();
 FILLER_ASAP7_75t_R FILLER_159_278 ();
 DECAPx4_ASAP7_75t_R FILLER_159_286 ();
 DECAPx2_ASAP7_75t_R FILLER_159_306 ();
 DECAPx1_ASAP7_75t_R FILLER_159_324 ();
 FILLER_ASAP7_75t_R FILLER_159_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_348 ();
 DECAPx2_ASAP7_75t_R FILLER_159_355 ();
 FILLER_ASAP7_75t_R FILLER_159_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_363 ();
 DECAPx2_ASAP7_75t_R FILLER_159_396 ();
 FILLER_ASAP7_75t_R FILLER_159_402 ();
 DECAPx1_ASAP7_75t_R FILLER_159_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_420 ();
 DECAPx1_ASAP7_75t_R FILLER_159_427 ();
 DECAPx6_ASAP7_75t_R FILLER_159_434 ();
 FILLER_ASAP7_75t_R FILLER_159_448 ();
 DECAPx1_ASAP7_75t_R FILLER_159_468 ();
 DECAPx4_ASAP7_75t_R FILLER_159_490 ();
 FILLER_ASAP7_75t_R FILLER_159_500 ();
 DECAPx1_ASAP7_75t_R FILLER_159_556 ();
 DECAPx1_ASAP7_75t_R FILLER_159_577 ();
 DECAPx2_ASAP7_75t_R FILLER_159_588 ();
 DECAPx4_ASAP7_75t_R FILLER_159_597 ();
 DECAPx4_ASAP7_75t_R FILLER_159_615 ();
 FILLER_ASAP7_75t_R FILLER_159_625 ();
 DECAPx2_ASAP7_75t_R FILLER_159_637 ();
 DECAPx2_ASAP7_75t_R FILLER_159_675 ();
 FILLER_ASAP7_75t_R FILLER_159_681 ();
 DECAPx4_ASAP7_75t_R FILLER_159_695 ();
 DECAPx2_ASAP7_75t_R FILLER_159_711 ();
 DECAPx4_ASAP7_75t_R FILLER_159_725 ();
 DECAPx4_ASAP7_75t_R FILLER_159_753 ();
 FILLER_ASAP7_75t_R FILLER_159_763 ();
 DECAPx4_ASAP7_75t_R FILLER_159_781 ();
 FILLER_ASAP7_75t_R FILLER_159_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_793 ();
 DECAPx4_ASAP7_75t_R FILLER_159_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_810 ();
 DECAPx4_ASAP7_75t_R FILLER_159_827 ();
 FILLER_ASAP7_75t_R FILLER_159_849 ();
 DECAPx4_ASAP7_75t_R FILLER_159_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_880 ();
 DECAPx6_ASAP7_75t_R FILLER_159_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_912 ();
 DECAPx1_ASAP7_75t_R FILLER_159_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_941 ();
 DECAPx1_ASAP7_75t_R FILLER_159_954 ();
 FILLER_ASAP7_75t_R FILLER_159_973 ();
 DECAPx10_ASAP7_75t_R FILLER_159_997 ();
 FILLER_ASAP7_75t_R FILLER_159_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1103 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1122 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1135 ();
 FILLER_ASAP7_75t_R FILLER_159_1141 ();
 FILLER_ASAP7_75t_R FILLER_159_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1214 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1241 ();
 FILLER_ASAP7_75t_R FILLER_159_1247 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1262 ();
 FILLER_ASAP7_75t_R FILLER_159_1268 ();
 FILLER_ASAP7_75t_R FILLER_159_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1300 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1322 ();
 FILLER_ASAP7_75t_R FILLER_159_1332 ();
 FILLER_ASAP7_75t_R FILLER_159_1342 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1378 ();
 FILLER_ASAP7_75t_R FILLER_159_1384 ();
 DECAPx10_ASAP7_75t_R FILLER_160_2 ();
 FILLER_ASAP7_75t_R FILLER_160_24 ();
 FILLER_ASAP7_75t_R FILLER_160_42 ();
 DECAPx4_ASAP7_75t_R FILLER_160_54 ();
 DECAPx1_ASAP7_75t_R FILLER_160_74 ();
 DECAPx10_ASAP7_75t_R FILLER_160_96 ();
 DECAPx4_ASAP7_75t_R FILLER_160_118 ();
 DECAPx10_ASAP7_75t_R FILLER_160_138 ();
 DECAPx6_ASAP7_75t_R FILLER_160_160 ();
 FILLER_ASAP7_75t_R FILLER_160_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_176 ();
 DECAPx1_ASAP7_75t_R FILLER_160_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_214 ();
 DECAPx2_ASAP7_75t_R FILLER_160_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_251 ();
 DECAPx2_ASAP7_75t_R FILLER_160_260 ();
 DECAPx6_ASAP7_75t_R FILLER_160_280 ();
 DECAPx1_ASAP7_75t_R FILLER_160_294 ();
 DECAPx10_ASAP7_75t_R FILLER_160_308 ();
 DECAPx1_ASAP7_75t_R FILLER_160_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_334 ();
 DECAPx10_ASAP7_75t_R FILLER_160_347 ();
 FILLER_ASAP7_75t_R FILLER_160_369 ();
 DECAPx4_ASAP7_75t_R FILLER_160_377 ();
 FILLER_ASAP7_75t_R FILLER_160_387 ();
 DECAPx2_ASAP7_75t_R FILLER_160_405 ();
 FILLER_ASAP7_75t_R FILLER_160_411 ();
 DECAPx4_ASAP7_75t_R FILLER_160_425 ();
 DECAPx2_ASAP7_75t_R FILLER_160_453 ();
 FILLER_ASAP7_75t_R FILLER_160_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_461 ();
 DECAPx6_ASAP7_75t_R FILLER_160_474 ();
 DECAPx10_ASAP7_75t_R FILLER_160_512 ();
 DECAPx1_ASAP7_75t_R FILLER_160_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_538 ();
 DECAPx10_ASAP7_75t_R FILLER_160_589 ();
 DECAPx6_ASAP7_75t_R FILLER_160_611 ();
 DECAPx2_ASAP7_75t_R FILLER_160_625 ();
 DECAPx2_ASAP7_75t_R FILLER_160_662 ();
 FILLER_ASAP7_75t_R FILLER_160_668 ();
 DECAPx1_ASAP7_75t_R FILLER_160_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_678 ();
 DECAPx1_ASAP7_75t_R FILLER_160_682 ();
 DECAPx2_ASAP7_75t_R FILLER_160_694 ();
 FILLER_ASAP7_75t_R FILLER_160_712 ();
 DECAPx10_ASAP7_75t_R FILLER_160_724 ();
 DECAPx10_ASAP7_75t_R FILLER_160_752 ();
 FILLER_ASAP7_75t_R FILLER_160_774 ();
 DECAPx2_ASAP7_75t_R FILLER_160_782 ();
 FILLER_ASAP7_75t_R FILLER_160_788 ();
 DECAPx2_ASAP7_75t_R FILLER_160_802 ();
 DECAPx10_ASAP7_75t_R FILLER_160_814 ();
 FILLER_ASAP7_75t_R FILLER_160_836 ();
 DECAPx6_ASAP7_75t_R FILLER_160_844 ();
 DECAPx2_ASAP7_75t_R FILLER_160_858 ();
 DECAPx4_ASAP7_75t_R FILLER_160_874 ();
 DECAPx6_ASAP7_75t_R FILLER_160_887 ();
 DECAPx2_ASAP7_75t_R FILLER_160_913 ();
 FILLER_ASAP7_75t_R FILLER_160_919 ();
 DECAPx4_ASAP7_75t_R FILLER_160_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_940 ();
 DECAPx4_ASAP7_75t_R FILLER_160_949 ();
 DECAPx6_ASAP7_75t_R FILLER_160_978 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1008 ();
 FILLER_ASAP7_75t_R FILLER_160_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1060 ();
 FILLER_ASAP7_75t_R FILLER_160_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1081 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1112 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1154 ();
 FILLER_ASAP7_75t_R FILLER_160_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1236 ();
 FILLER_ASAP7_75t_R FILLER_160_1242 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1247 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1259 ();
 FILLER_ASAP7_75t_R FILLER_160_1269 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1307 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1347 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_161_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_12 ();
 DECAPx4_ASAP7_75t_R FILLER_161_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_33 ();
 DECAPx1_ASAP7_75t_R FILLER_161_44 ();
 DECAPx6_ASAP7_75t_R FILLER_161_58 ();
 DECAPx1_ASAP7_75t_R FILLER_161_72 ();
 DECAPx6_ASAP7_75t_R FILLER_161_118 ();
 FILLER_ASAP7_75t_R FILLER_161_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_134 ();
 FILLER_ASAP7_75t_R FILLER_161_145 ();
 DECAPx10_ASAP7_75t_R FILLER_161_157 ();
 DECAPx4_ASAP7_75t_R FILLER_161_179 ();
 FILLER_ASAP7_75t_R FILLER_161_189 ();
 DECAPx6_ASAP7_75t_R FILLER_161_194 ();
 FILLER_ASAP7_75t_R FILLER_161_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_223 ();
 DECAPx6_ASAP7_75t_R FILLER_161_230 ();
 FILLER_ASAP7_75t_R FILLER_161_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_272 ();
 DECAPx1_ASAP7_75t_R FILLER_161_307 ();
 DECAPx6_ASAP7_75t_R FILLER_161_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_331 ();
 DECAPx4_ASAP7_75t_R FILLER_161_358 ();
 FILLER_ASAP7_75t_R FILLER_161_368 ();
 DECAPx4_ASAP7_75t_R FILLER_161_388 ();
 DECAPx1_ASAP7_75t_R FILLER_161_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_439 ();
 DECAPx4_ASAP7_75t_R FILLER_161_458 ();
 DECAPx2_ASAP7_75t_R FILLER_161_492 ();
 FILLER_ASAP7_75t_R FILLER_161_498 ();
 DECAPx1_ASAP7_75t_R FILLER_161_516 ();
 DECAPx1_ASAP7_75t_R FILLER_161_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_542 ();
 DECAPx2_ASAP7_75t_R FILLER_161_569 ();
 FILLER_ASAP7_75t_R FILLER_161_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_577 ();
 DECAPx2_ASAP7_75t_R FILLER_161_581 ();
 DECAPx1_ASAP7_75t_R FILLER_161_593 ();
 DECAPx4_ASAP7_75t_R FILLER_161_600 ();
 DECAPx4_ASAP7_75t_R FILLER_161_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_638 ();
 DECAPx6_ASAP7_75t_R FILLER_161_656 ();
 DECAPx2_ASAP7_75t_R FILLER_161_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_676 ();
 DECAPx6_ASAP7_75t_R FILLER_161_693 ();
 DECAPx4_ASAP7_75t_R FILLER_161_713 ();
 FILLER_ASAP7_75t_R FILLER_161_723 ();
 DECAPx6_ASAP7_75t_R FILLER_161_741 ();
 DECAPx6_ASAP7_75t_R FILLER_161_762 ();
 FILLER_ASAP7_75t_R FILLER_161_776 ();
 FILLER_ASAP7_75t_R FILLER_161_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_792 ();
 FILLER_ASAP7_75t_R FILLER_161_806 ();
 DECAPx2_ASAP7_75t_R FILLER_161_824 ();
 FILLER_ASAP7_75t_R FILLER_161_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_832 ();
 FILLER_ASAP7_75t_R FILLER_161_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_862 ();
 DECAPx1_ASAP7_75t_R FILLER_161_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_873 ();
 DECAPx6_ASAP7_75t_R FILLER_161_886 ();
 DECAPx1_ASAP7_75t_R FILLER_161_900 ();
 FILLER_ASAP7_75t_R FILLER_161_916 ();
 DECAPx4_ASAP7_75t_R FILLER_161_936 ();
 FILLER_ASAP7_75t_R FILLER_161_946 ();
 DECAPx2_ASAP7_75t_R FILLER_161_955 ();
 FILLER_ASAP7_75t_R FILLER_161_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_963 ();
 FILLER_ASAP7_75t_R FILLER_161_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_970 ();
 FILLER_ASAP7_75t_R FILLER_161_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_997 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1042 ();
 FILLER_ASAP7_75t_R FILLER_161_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1122 ();
 FILLER_ASAP7_75t_R FILLER_161_1138 ();
 FILLER_ASAP7_75t_R FILLER_161_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1169 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1185 ();
 FILLER_ASAP7_75t_R FILLER_161_1199 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1223 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1289 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1324 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1328 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1332 ();
 FILLER_ASAP7_75t_R FILLER_161_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_162_2 ();
 DECAPx2_ASAP7_75t_R FILLER_162_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_36 ();
 DECAPx6_ASAP7_75t_R FILLER_162_47 ();
 DECAPx1_ASAP7_75t_R FILLER_162_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_65 ();
 FILLER_ASAP7_75t_R FILLER_162_76 ();
 FILLER_ASAP7_75t_R FILLER_162_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_96 ();
 DECAPx10_ASAP7_75t_R FILLER_162_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_122 ();
 DECAPx2_ASAP7_75t_R FILLER_162_141 ();
 DECAPx6_ASAP7_75t_R FILLER_162_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_187 ();
 DECAPx6_ASAP7_75t_R FILLER_162_206 ();
 DECAPx1_ASAP7_75t_R FILLER_162_220 ();
 DECAPx10_ASAP7_75t_R FILLER_162_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_252 ();
 FILLER_ASAP7_75t_R FILLER_162_262 ();
 DECAPx1_ASAP7_75t_R FILLER_162_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_282 ();
 DECAPx1_ASAP7_75t_R FILLER_162_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_300 ();
 DECAPx6_ASAP7_75t_R FILLER_162_327 ();
 DECAPx10_ASAP7_75t_R FILLER_162_350 ();
 DECAPx6_ASAP7_75t_R FILLER_162_372 ();
 DECAPx2_ASAP7_75t_R FILLER_162_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_416 ();
 DECAPx1_ASAP7_75t_R FILLER_162_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_427 ();
 DECAPx4_ASAP7_75t_R FILLER_162_431 ();
 FILLER_ASAP7_75t_R FILLER_162_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_443 ();
 DECAPx1_ASAP7_75t_R FILLER_162_474 ();
 FILLER_ASAP7_75t_R FILLER_162_514 ();
 FILLER_ASAP7_75t_R FILLER_162_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_536 ();
 DECAPx1_ASAP7_75t_R FILLER_162_553 ();
 DECAPx10_ASAP7_75t_R FILLER_162_560 ();
 DECAPx6_ASAP7_75t_R FILLER_162_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_658 ();
 DECAPx6_ASAP7_75t_R FILLER_162_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_683 ();
 FILLER_ASAP7_75t_R FILLER_162_690 ();
 FILLER_ASAP7_75t_R FILLER_162_708 ();
 FILLER_ASAP7_75t_R FILLER_162_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_736 ();
 DECAPx4_ASAP7_75t_R FILLER_162_743 ();
 FILLER_ASAP7_75t_R FILLER_162_753 ();
 FILLER_ASAP7_75t_R FILLER_162_771 ();
 DECAPx1_ASAP7_75t_R FILLER_162_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_789 ();
 DECAPx2_ASAP7_75t_R FILLER_162_802 ();
 FILLER_ASAP7_75t_R FILLER_162_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_810 ();
 FILLER_ASAP7_75t_R FILLER_162_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_819 ();
 DECAPx4_ASAP7_75t_R FILLER_162_836 ();
 FILLER_ASAP7_75t_R FILLER_162_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_848 ();
 DECAPx2_ASAP7_75t_R FILLER_162_865 ();
 FILLER_ASAP7_75t_R FILLER_162_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_890 ();
 DECAPx1_ASAP7_75t_R FILLER_162_929 ();
 DECAPx2_ASAP7_75t_R FILLER_162_953 ();
 DECAPx2_ASAP7_75t_R FILLER_162_975 ();
 FILLER_ASAP7_75t_R FILLER_162_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_983 ();
 DECAPx6_ASAP7_75t_R FILLER_162_991 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1024 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1034 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1065 ();
 FILLER_ASAP7_75t_R FILLER_162_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1100 ();
 FILLER_ASAP7_75t_R FILLER_162_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1125 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1176 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1187 ();
 FILLER_ASAP7_75t_R FILLER_162_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1217 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1231 ();
 FILLER_ASAP7_75t_R FILLER_162_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1282 ();
 FILLER_ASAP7_75t_R FILLER_162_1288 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1296 ();
 FILLER_ASAP7_75t_R FILLER_162_1306 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1317 ();
 FILLER_ASAP7_75t_R FILLER_162_1339 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1349 ();
 FILLER_ASAP7_75t_R FILLER_162_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1357 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1372 ();
 FILLER_ASAP7_75t_R FILLER_162_1378 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1388 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_2 ();
 DECAPx10_ASAP7_75t_R FILLER_163_29 ();
 FILLER_ASAP7_75t_R FILLER_163_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_53 ();
 FILLER_ASAP7_75t_R FILLER_163_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_66 ();
 FILLER_ASAP7_75t_R FILLER_163_97 ();
 DECAPx6_ASAP7_75t_R FILLER_163_111 ();
 FILLER_ASAP7_75t_R FILLER_163_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_162 ();
 FILLER_ASAP7_75t_R FILLER_163_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_202 ();
 DECAPx4_ASAP7_75t_R FILLER_163_211 ();
 FILLER_ASAP7_75t_R FILLER_163_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_223 ();
 FILLER_ASAP7_75t_R FILLER_163_230 ();
 DECAPx2_ASAP7_75t_R FILLER_163_246 ();
 DECAPx6_ASAP7_75t_R FILLER_163_258 ();
 DECAPx2_ASAP7_75t_R FILLER_163_272 ();
 FILLER_ASAP7_75t_R FILLER_163_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_294 ();
 DECAPx2_ASAP7_75t_R FILLER_163_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_304 ();
 FILLER_ASAP7_75t_R FILLER_163_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_318 ();
 DECAPx1_ASAP7_75t_R FILLER_163_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_329 ();
 FILLER_ASAP7_75t_R FILLER_163_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_380 ();
 FILLER_ASAP7_75t_R FILLER_163_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_386 ();
 FILLER_ASAP7_75t_R FILLER_163_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_407 ();
 DECAPx10_ASAP7_75t_R FILLER_163_422 ();
 DECAPx2_ASAP7_75t_R FILLER_163_444 ();
 DECAPx6_ASAP7_75t_R FILLER_163_511 ();
 DECAPx6_ASAP7_75t_R FILLER_163_549 ();
 DECAPx1_ASAP7_75t_R FILLER_163_563 ();
 DECAPx6_ASAP7_75t_R FILLER_163_591 ();
 FILLER_ASAP7_75t_R FILLER_163_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_625 ();
 DECAPx6_ASAP7_75t_R FILLER_163_644 ();
 DECAPx2_ASAP7_75t_R FILLER_163_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_677 ();
 DECAPx1_ASAP7_75t_R FILLER_163_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_692 ();
 DECAPx1_ASAP7_75t_R FILLER_163_700 ();
 DECAPx1_ASAP7_75t_R FILLER_163_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_731 ();
 DECAPx1_ASAP7_75t_R FILLER_163_751 ();
 FILLER_ASAP7_75t_R FILLER_163_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_793 ();
 DECAPx1_ASAP7_75t_R FILLER_163_806 ();
 DECAPx1_ASAP7_75t_R FILLER_163_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_820 ();
 FILLER_ASAP7_75t_R FILLER_163_837 ();
 DECAPx4_ASAP7_75t_R FILLER_163_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_855 ();
 DECAPx2_ASAP7_75t_R FILLER_163_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_874 ();
 DECAPx2_ASAP7_75t_R FILLER_163_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_903 ();
 DECAPx6_ASAP7_75t_R FILLER_163_910 ();
 DECAPx1_ASAP7_75t_R FILLER_163_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_930 ();
 DECAPx2_ASAP7_75t_R FILLER_163_958 ();
 FILLER_ASAP7_75t_R FILLER_163_964 ();
 DECAPx10_ASAP7_75t_R FILLER_163_976 ();
 DECAPx6_ASAP7_75t_R FILLER_163_998 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1012 ();
 FILLER_ASAP7_75t_R FILLER_163_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1062 ();
 FILLER_ASAP7_75t_R FILLER_163_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1070 ();
 FILLER_ASAP7_75t_R FILLER_163_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1103 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1124 ();
 FILLER_ASAP7_75t_R FILLER_163_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1132 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1162 ();
 FILLER_ASAP7_75t_R FILLER_163_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1168 ();
 DECAPx4_ASAP7_75t_R FILLER_163_1175 ();
 FILLER_ASAP7_75t_R FILLER_163_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1220 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1285 ();
 DECAPx4_ASAP7_75t_R FILLER_163_1296 ();
 FILLER_ASAP7_75t_R FILLER_163_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1326 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1337 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1351 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1365 ();
 DECAPx6_ASAP7_75t_R FILLER_164_2 ();
 FILLER_ASAP7_75t_R FILLER_164_16 ();
 FILLER_ASAP7_75t_R FILLER_164_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_23 ();
 DECAPx2_ASAP7_75t_R FILLER_164_34 ();
 FILLER_ASAP7_75t_R FILLER_164_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_42 ();
 DECAPx4_ASAP7_75t_R FILLER_164_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_59 ();
 DECAPx6_ASAP7_75t_R FILLER_164_78 ();
 DECAPx6_ASAP7_75t_R FILLER_164_130 ();
 FILLER_ASAP7_75t_R FILLER_164_144 ();
 FILLER_ASAP7_75t_R FILLER_164_165 ();
 DECAPx2_ASAP7_75t_R FILLER_164_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_188 ();
 DECAPx2_ASAP7_75t_R FILLER_164_217 ();
 FILLER_ASAP7_75t_R FILLER_164_223 ();
 DECAPx1_ASAP7_75t_R FILLER_164_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_253 ();
 DECAPx6_ASAP7_75t_R FILLER_164_268 ();
 DECAPx1_ASAP7_75t_R FILLER_164_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_286 ();
 DECAPx1_ASAP7_75t_R FILLER_164_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_301 ();
 DECAPx2_ASAP7_75t_R FILLER_164_308 ();
 FILLER_ASAP7_75t_R FILLER_164_314 ();
 DECAPx2_ASAP7_75t_R FILLER_164_329 ();
 FILLER_ASAP7_75t_R FILLER_164_335 ();
 FILLER_ASAP7_75t_R FILLER_164_359 ();
 DECAPx4_ASAP7_75t_R FILLER_164_393 ();
 DECAPx2_ASAP7_75t_R FILLER_164_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_423 ();
 DECAPx2_ASAP7_75t_R FILLER_164_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_439 ();
 DECAPx2_ASAP7_75t_R FILLER_164_443 ();
 FILLER_ASAP7_75t_R FILLER_164_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_461 ();
 DECAPx10_ASAP7_75t_R FILLER_164_464 ();
 DECAPx10_ASAP7_75t_R FILLER_164_516 ();
 DECAPx1_ASAP7_75t_R FILLER_164_538 ();
 DECAPx1_ASAP7_75t_R FILLER_164_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_558 ();
 FILLER_ASAP7_75t_R FILLER_164_562 ();
 DECAPx6_ASAP7_75t_R FILLER_164_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_582 ();
 DECAPx4_ASAP7_75t_R FILLER_164_595 ();
 DECAPx10_ASAP7_75t_R FILLER_164_615 ();
 DECAPx2_ASAP7_75t_R FILLER_164_637 ();
 FILLER_ASAP7_75t_R FILLER_164_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_663 ();
 DECAPx1_ASAP7_75t_R FILLER_164_682 ();
 DECAPx1_ASAP7_75t_R FILLER_164_702 ();
 DECAPx1_ASAP7_75t_R FILLER_164_718 ();
 DECAPx2_ASAP7_75t_R FILLER_164_728 ();
 FILLER_ASAP7_75t_R FILLER_164_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_736 ();
 FILLER_ASAP7_75t_R FILLER_164_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_746 ();
 DECAPx1_ASAP7_75t_R FILLER_164_759 ();
 DECAPx1_ASAP7_75t_R FILLER_164_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_783 ();
 DECAPx2_ASAP7_75t_R FILLER_164_808 ();
 FILLER_ASAP7_75t_R FILLER_164_814 ();
 DECAPx4_ASAP7_75t_R FILLER_164_822 ();
 FILLER_ASAP7_75t_R FILLER_164_832 ();
 DECAPx2_ASAP7_75t_R FILLER_164_850 ();
 FILLER_ASAP7_75t_R FILLER_164_856 ();
 DECAPx4_ASAP7_75t_R FILLER_164_868 ();
 FILLER_ASAP7_75t_R FILLER_164_878 ();
 DECAPx6_ASAP7_75t_R FILLER_164_886 ();
 DECAPx2_ASAP7_75t_R FILLER_164_900 ();
 DECAPx10_ASAP7_75t_R FILLER_164_912 ();
 DECAPx10_ASAP7_75t_R FILLER_164_934 ();
 DECAPx6_ASAP7_75t_R FILLER_164_962 ();
 DECAPx2_ASAP7_75t_R FILLER_164_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_982 ();
 FILLER_ASAP7_75t_R FILLER_164_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_997 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1020 ();
 FILLER_ASAP7_75t_R FILLER_164_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1040 ();
 FILLER_ASAP7_75t_R FILLER_164_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1063 ();
 FILLER_ASAP7_75t_R FILLER_164_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1143 ();
 DECAPx6_ASAP7_75t_R FILLER_164_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1197 ();
 FILLER_ASAP7_75t_R FILLER_164_1214 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1230 ();
 DECAPx6_ASAP7_75t_R FILLER_164_1239 ();
 FILLER_ASAP7_75t_R FILLER_164_1253 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1267 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1314 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1320 ();
 FILLER_ASAP7_75t_R FILLER_164_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1349 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1370 ();
 FILLER_ASAP7_75t_R FILLER_164_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_165_2 ();
 FILLER_ASAP7_75t_R FILLER_165_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_14 ();
 DECAPx2_ASAP7_75t_R FILLER_165_34 ();
 FILLER_ASAP7_75t_R FILLER_165_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_42 ();
 DECAPx2_ASAP7_75t_R FILLER_165_49 ();
 FILLER_ASAP7_75t_R FILLER_165_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_57 ();
 DECAPx10_ASAP7_75t_R FILLER_165_76 ();
 DECAPx2_ASAP7_75t_R FILLER_165_98 ();
 FILLER_ASAP7_75t_R FILLER_165_104 ();
 DECAPx6_ASAP7_75t_R FILLER_165_109 ();
 DECAPx1_ASAP7_75t_R FILLER_165_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_127 ();
 DECAPx2_ASAP7_75t_R FILLER_165_134 ();
 FILLER_ASAP7_75t_R FILLER_165_140 ();
 DECAPx10_ASAP7_75t_R FILLER_165_155 ();
 DECAPx6_ASAP7_75t_R FILLER_165_177 ();
 DECAPx2_ASAP7_75t_R FILLER_165_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_204 ();
 DECAPx1_ASAP7_75t_R FILLER_165_211 ();
 DECAPx1_ASAP7_75t_R FILLER_165_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_225 ();
 DECAPx2_ASAP7_75t_R FILLER_165_238 ();
 DECAPx1_ASAP7_75t_R FILLER_165_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_301 ();
 FILLER_ASAP7_75t_R FILLER_165_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_320 ();
 DECAPx2_ASAP7_75t_R FILLER_165_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_335 ();
 FILLER_ASAP7_75t_R FILLER_165_344 ();
 DECAPx6_ASAP7_75t_R FILLER_165_352 ();
 DECAPx1_ASAP7_75t_R FILLER_165_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_370 ();
 DECAPx2_ASAP7_75t_R FILLER_165_377 ();
 FILLER_ASAP7_75t_R FILLER_165_383 ();
 DECAPx1_ASAP7_75t_R FILLER_165_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_392 ();
 DECAPx1_ASAP7_75t_R FILLER_165_407 ();
 DECAPx1_ASAP7_75t_R FILLER_165_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_421 ();
 DECAPx2_ASAP7_75t_R FILLER_165_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_454 ();
 DECAPx4_ASAP7_75t_R FILLER_165_491 ();
 DECAPx2_ASAP7_75t_R FILLER_165_519 ();
 FILLER_ASAP7_75t_R FILLER_165_525 ();
 DECAPx4_ASAP7_75t_R FILLER_165_571 ();
 FILLER_ASAP7_75t_R FILLER_165_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_583 ();
 FILLER_ASAP7_75t_R FILLER_165_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_604 ();
 DECAPx2_ASAP7_75t_R FILLER_165_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_623 ();
 DECAPx2_ASAP7_75t_R FILLER_165_634 ();
 FILLER_ASAP7_75t_R FILLER_165_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_642 ();
 DECAPx1_ASAP7_75t_R FILLER_165_655 ();
 DECAPx4_ASAP7_75t_R FILLER_165_665 ();
 DECAPx6_ASAP7_75t_R FILLER_165_693 ();
 FILLER_ASAP7_75t_R FILLER_165_707 ();
 DECAPx2_ASAP7_75t_R FILLER_165_712 ();
 FILLER_ASAP7_75t_R FILLER_165_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_720 ();
 DECAPx2_ASAP7_75t_R FILLER_165_727 ();
 FILLER_ASAP7_75t_R FILLER_165_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_756 ();
 DECAPx2_ASAP7_75t_R FILLER_165_765 ();
 FILLER_ASAP7_75t_R FILLER_165_771 ();
 DECAPx2_ASAP7_75t_R FILLER_165_781 ();
 DECAPx1_ASAP7_75t_R FILLER_165_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_823 ();
 DECAPx1_ASAP7_75t_R FILLER_165_830 ();
 DECAPx10_ASAP7_75t_R FILLER_165_844 ();
 DECAPx10_ASAP7_75t_R FILLER_165_866 ();
 FILLER_ASAP7_75t_R FILLER_165_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_890 ();
 FILLER_ASAP7_75t_R FILLER_165_898 ();
 DECAPx1_ASAP7_75t_R FILLER_165_913 ();
 FILLER_ASAP7_75t_R FILLER_165_938 ();
 FILLER_ASAP7_75t_R FILLER_165_961 ();
 DECAPx1_ASAP7_75t_R FILLER_165_971 ();
 FILLER_ASAP7_75t_R FILLER_165_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1045 ();
 FILLER_ASAP7_75t_R FILLER_165_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1112 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1119 ();
 FILLER_ASAP7_75t_R FILLER_165_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_165_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1188 ();
 FILLER_ASAP7_75t_R FILLER_165_1194 ();
 DECAPx4_ASAP7_75t_R FILLER_165_1225 ();
 FILLER_ASAP7_75t_R FILLER_165_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1255 ();
 DECAPx1_ASAP7_75t_R FILLER_165_1277 ();
 DECAPx1_ASAP7_75t_R FILLER_165_1299 ();
 DECAPx4_ASAP7_75t_R FILLER_165_1306 ();
 FILLER_ASAP7_75t_R FILLER_165_1333 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1338 ();
 FILLER_ASAP7_75t_R FILLER_166_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_60 ();
 DECAPx6_ASAP7_75t_R FILLER_166_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_150 ();
 FILLER_ASAP7_75t_R FILLER_166_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_173 ();
 DECAPx4_ASAP7_75t_R FILLER_166_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_196 ();
 FILLER_ASAP7_75t_R FILLER_166_217 ();
 DECAPx10_ASAP7_75t_R FILLER_166_231 ();
 DECAPx6_ASAP7_75t_R FILLER_166_273 ();
 DECAPx2_ASAP7_75t_R FILLER_166_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_311 ();
 FILLER_ASAP7_75t_R FILLER_166_318 ();
 DECAPx1_ASAP7_75t_R FILLER_166_329 ();
 DECAPx2_ASAP7_75t_R FILLER_166_353 ();
 FILLER_ASAP7_75t_R FILLER_166_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_368 ();
 DECAPx6_ASAP7_75t_R FILLER_166_372 ();
 FILLER_ASAP7_75t_R FILLER_166_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_388 ();
 DECAPx2_ASAP7_75t_R FILLER_166_397 ();
 FILLER_ASAP7_75t_R FILLER_166_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_405 ();
 DECAPx4_ASAP7_75t_R FILLER_166_412 ();
 FILLER_ASAP7_75t_R FILLER_166_422 ();
 DECAPx10_ASAP7_75t_R FILLER_166_430 ();
 DECAPx4_ASAP7_75t_R FILLER_166_452 ();
 DECAPx4_ASAP7_75t_R FILLER_166_464 ();
 FILLER_ASAP7_75t_R FILLER_166_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_495 ();
 DECAPx1_ASAP7_75t_R FILLER_166_520 ();
 DECAPx1_ASAP7_75t_R FILLER_166_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_531 ();
 FILLER_ASAP7_75t_R FILLER_166_542 ();
 DECAPx6_ASAP7_75t_R FILLER_166_550 ();
 FILLER_ASAP7_75t_R FILLER_166_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_576 ();
 FILLER_ASAP7_75t_R FILLER_166_599 ();
 DECAPx2_ASAP7_75t_R FILLER_166_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_639 ();
 DECAPx4_ASAP7_75t_R FILLER_166_668 ();
 DECAPx2_ASAP7_75t_R FILLER_166_700 ();
 DECAPx2_ASAP7_75t_R FILLER_166_712 ();
 FILLER_ASAP7_75t_R FILLER_166_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_720 ();
 FILLER_ASAP7_75t_R FILLER_166_731 ();
 DECAPx1_ASAP7_75t_R FILLER_166_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_752 ();
 DECAPx4_ASAP7_75t_R FILLER_166_764 ();
 DECAPx2_ASAP7_75t_R FILLER_166_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_786 ();
 DECAPx6_ASAP7_75t_R FILLER_166_799 ();
 FILLER_ASAP7_75t_R FILLER_166_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_815 ();
 FILLER_ASAP7_75t_R FILLER_166_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_838 ();
 DECAPx2_ASAP7_75t_R FILLER_166_851 ();
 FILLER_ASAP7_75t_R FILLER_166_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_900 ();
 FILLER_ASAP7_75t_R FILLER_166_919 ();
 DECAPx1_ASAP7_75t_R FILLER_166_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_935 ();
 FILLER_ASAP7_75t_R FILLER_166_943 ();
 DECAPx1_ASAP7_75t_R FILLER_166_952 ();
 FILLER_ASAP7_75t_R FILLER_166_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_966 ();
 FILLER_ASAP7_75t_R FILLER_166_1000 ();
 FILLER_ASAP7_75t_R FILLER_166_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1066 ();
 DECAPx6_ASAP7_75t_R FILLER_166_1077 ();
 FILLER_ASAP7_75t_R FILLER_166_1091 ();
 FILLER_ASAP7_75t_R FILLER_166_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1124 ();
 FILLER_ASAP7_75t_R FILLER_166_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1184 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1210 ();
 FILLER_ASAP7_75t_R FILLER_166_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1216 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1237 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1268 ();
 FILLER_ASAP7_75t_R FILLER_166_1279 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1291 ();
 FILLER_ASAP7_75t_R FILLER_166_1360 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1369 ();
 FILLER_ASAP7_75t_R FILLER_166_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_167_2 ();
 DECAPx2_ASAP7_75t_R FILLER_167_16 ();
 DECAPx6_ASAP7_75t_R FILLER_167_28 ();
 DECAPx4_ASAP7_75t_R FILLER_167_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_61 ();
 DECAPx4_ASAP7_75t_R FILLER_167_92 ();
 FILLER_ASAP7_75t_R FILLER_167_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_166 ();
 FILLER_ASAP7_75t_R FILLER_167_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_203 ();
 DECAPx6_ASAP7_75t_R FILLER_167_212 ();
 DECAPx4_ASAP7_75t_R FILLER_167_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_242 ();
 DECAPx2_ASAP7_75t_R FILLER_167_246 ();
 DECAPx1_ASAP7_75t_R FILLER_167_258 ();
 DECAPx6_ASAP7_75t_R FILLER_167_268 ();
 FILLER_ASAP7_75t_R FILLER_167_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_284 ();
 DECAPx1_ASAP7_75t_R FILLER_167_295 ();
 DECAPx2_ASAP7_75t_R FILLER_167_325 ();
 FILLER_ASAP7_75t_R FILLER_167_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_333 ();
 DECAPx4_ASAP7_75t_R FILLER_167_340 ();
 FILLER_ASAP7_75t_R FILLER_167_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_352 ();
 FILLER_ASAP7_75t_R FILLER_167_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_399 ();
 DECAPx1_ASAP7_75t_R FILLER_167_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_418 ();
 DECAPx1_ASAP7_75t_R FILLER_167_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_429 ();
 DECAPx1_ASAP7_75t_R FILLER_167_446 ();
 DECAPx1_ASAP7_75t_R FILLER_167_468 ();
 DECAPx2_ASAP7_75t_R FILLER_167_496 ();
 DECAPx1_ASAP7_75t_R FILLER_167_505 ();
 DECAPx1_ASAP7_75t_R FILLER_167_535 ();
 DECAPx4_ASAP7_75t_R FILLER_167_571 ();
 FILLER_ASAP7_75t_R FILLER_167_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_583 ();
 DECAPx4_ASAP7_75t_R FILLER_167_594 ();
 FILLER_ASAP7_75t_R FILLER_167_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_641 ();
 DECAPx6_ASAP7_75t_R FILLER_167_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_678 ();
 FILLER_ASAP7_75t_R FILLER_167_685 ();
 DECAPx2_ASAP7_75t_R FILLER_167_699 ();
 FILLER_ASAP7_75t_R FILLER_167_705 ();
 FILLER_ASAP7_75t_R FILLER_167_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_717 ();
 DECAPx2_ASAP7_75t_R FILLER_167_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_730 ();
 DECAPx4_ASAP7_75t_R FILLER_167_738 ();
 FILLER_ASAP7_75t_R FILLER_167_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_750 ();
 DECAPx1_ASAP7_75t_R FILLER_167_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_761 ();
 DECAPx1_ASAP7_75t_R FILLER_167_774 ();
 DECAPx4_ASAP7_75t_R FILLER_167_784 ();
 FILLER_ASAP7_75t_R FILLER_167_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_796 ();
 DECAPx6_ASAP7_75t_R FILLER_167_804 ();
 FILLER_ASAP7_75t_R FILLER_167_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_820 ();
 DECAPx4_ASAP7_75t_R FILLER_167_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_845 ();
 DECAPx6_ASAP7_75t_R FILLER_167_888 ();
 FILLER_ASAP7_75t_R FILLER_167_902 ();
 FILLER_ASAP7_75t_R FILLER_167_910 ();
 DECAPx1_ASAP7_75t_R FILLER_167_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_923 ();
 DECAPx2_ASAP7_75t_R FILLER_167_934 ();
 FILLER_ASAP7_75t_R FILLER_167_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_942 ();
 DECAPx4_ASAP7_75t_R FILLER_167_961 ();
 FILLER_ASAP7_75t_R FILLER_167_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_980 ();
 DECAPx2_ASAP7_75t_R FILLER_167_991 ();
 FILLER_ASAP7_75t_R FILLER_167_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_999 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1018 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1035 ();
 FILLER_ASAP7_75t_R FILLER_167_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1064 ();
 DECAPx4_ASAP7_75t_R FILLER_167_1073 ();
 FILLER_ASAP7_75t_R FILLER_167_1083 ();
 FILLER_ASAP7_75t_R FILLER_167_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1103 ();
 FILLER_ASAP7_75t_R FILLER_167_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1120 ();
 FILLER_ASAP7_75t_R FILLER_167_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1146 ();
 FILLER_ASAP7_75t_R FILLER_167_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1172 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1206 ();
 FILLER_ASAP7_75t_R FILLER_167_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_167_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1236 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1247 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1258 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1272 ();
 FILLER_ASAP7_75t_R FILLER_167_1286 ();
 FILLER_ASAP7_75t_R FILLER_167_1304 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1364 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1391 ();
 DECAPx4_ASAP7_75t_R FILLER_168_2 ();
 FILLER_ASAP7_75t_R FILLER_168_12 ();
 FILLER_ASAP7_75t_R FILLER_168_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_31 ();
 DECAPx1_ASAP7_75t_R FILLER_168_62 ();
 DECAPx2_ASAP7_75t_R FILLER_168_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_90 ();
 FILLER_ASAP7_75t_R FILLER_168_97 ();
 DECAPx1_ASAP7_75t_R FILLER_168_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_109 ();
 DECAPx1_ASAP7_75t_R FILLER_168_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_144 ();
 FILLER_ASAP7_75t_R FILLER_168_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_186 ();
 FILLER_ASAP7_75t_R FILLER_168_201 ();
 DECAPx1_ASAP7_75t_R FILLER_168_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_213 ();
 DECAPx1_ASAP7_75t_R FILLER_168_224 ();
 DECAPx10_ASAP7_75t_R FILLER_168_272 ();
 FILLER_ASAP7_75t_R FILLER_168_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_296 ();
 DECAPx1_ASAP7_75t_R FILLER_168_309 ();
 DECAPx1_ASAP7_75t_R FILLER_168_316 ();
 DECAPx4_ASAP7_75t_R FILLER_168_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_348 ();
 DECAPx6_ASAP7_75t_R FILLER_168_370 ();
 DECAPx1_ASAP7_75t_R FILLER_168_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_388 ();
 DECAPx1_ASAP7_75t_R FILLER_168_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_399 ();
 DECAPx1_ASAP7_75t_R FILLER_168_412 ();
 DECAPx4_ASAP7_75t_R FILLER_168_442 ();
 DECAPx6_ASAP7_75t_R FILLER_168_464 ();
 DECAPx1_ASAP7_75t_R FILLER_168_478 ();
 DECAPx6_ASAP7_75t_R FILLER_168_520 ();
 DECAPx2_ASAP7_75t_R FILLER_168_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_540 ();
 DECAPx6_ASAP7_75t_R FILLER_168_544 ();
 FILLER_ASAP7_75t_R FILLER_168_558 ();
 DECAPx2_ASAP7_75t_R FILLER_168_563 ();
 DECAPx6_ASAP7_75t_R FILLER_168_587 ();
 FILLER_ASAP7_75t_R FILLER_168_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_603 ();
 DECAPx10_ASAP7_75t_R FILLER_168_614 ();
 DECAPx10_ASAP7_75t_R FILLER_168_636 ();
 DECAPx1_ASAP7_75t_R FILLER_168_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_694 ();
 DECAPx2_ASAP7_75t_R FILLER_168_737 ();
 FILLER_ASAP7_75t_R FILLER_168_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_745 ();
 DECAPx1_ASAP7_75t_R FILLER_168_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_763 ();
 FILLER_ASAP7_75t_R FILLER_168_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_776 ();
 DECAPx1_ASAP7_75t_R FILLER_168_783 ();
 FILLER_ASAP7_75t_R FILLER_168_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_816 ();
 DECAPx4_ASAP7_75t_R FILLER_168_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_833 ();
 DECAPx1_ASAP7_75t_R FILLER_168_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_856 ();
 DECAPx2_ASAP7_75t_R FILLER_168_863 ();
 FILLER_ASAP7_75t_R FILLER_168_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_871 ();
 DECAPx6_ASAP7_75t_R FILLER_168_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_905 ();
 DECAPx4_ASAP7_75t_R FILLER_168_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_927 ();
 DECAPx4_ASAP7_75t_R FILLER_168_935 ();
 DECAPx10_ASAP7_75t_R FILLER_168_965 ();
 DECAPx10_ASAP7_75t_R FILLER_168_987 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1009 ();
 FILLER_ASAP7_75t_R FILLER_168_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1048 ();
 FILLER_ASAP7_75t_R FILLER_168_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1060 ();
 FILLER_ASAP7_75t_R FILLER_168_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1102 ();
 FILLER_ASAP7_75t_R FILLER_168_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1126 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1156 ();
 FILLER_ASAP7_75t_R FILLER_168_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1263 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1272 ();
 FILLER_ASAP7_75t_R FILLER_168_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1311 ();
 FILLER_ASAP7_75t_R FILLER_168_1318 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_168_1324 ();
 FILLER_ASAP7_75t_R FILLER_168_1346 ();
 FILLER_ASAP7_75t_R FILLER_168_1358 ();
 DECAPx1_ASAP7_75t_R FILLER_168_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_169_32 ();
 FILLER_ASAP7_75t_R FILLER_169_42 ();
 DECAPx10_ASAP7_75t_R FILLER_169_53 ();
 DECAPx10_ASAP7_75t_R FILLER_169_75 ();
 DECAPx10_ASAP7_75t_R FILLER_169_123 ();
 DECAPx10_ASAP7_75t_R FILLER_169_145 ();
 DECAPx1_ASAP7_75t_R FILLER_169_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_171 ();
 DECAPx6_ASAP7_75t_R FILLER_169_175 ();
 FILLER_ASAP7_75t_R FILLER_169_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_191 ();
 DECAPx10_ASAP7_75t_R FILLER_169_204 ();
 FILLER_ASAP7_75t_R FILLER_169_226 ();
 DECAPx2_ASAP7_75t_R FILLER_169_260 ();
 DECAPx2_ASAP7_75t_R FILLER_169_272 ();
 DECAPx10_ASAP7_75t_R FILLER_169_281 ();
 DECAPx6_ASAP7_75t_R FILLER_169_303 ();
 FILLER_ASAP7_75t_R FILLER_169_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_319 ();
 DECAPx6_ASAP7_75t_R FILLER_169_338 ();
 DECAPx1_ASAP7_75t_R FILLER_169_352 ();
 DECAPx10_ASAP7_75t_R FILLER_169_366 ();
 DECAPx1_ASAP7_75t_R FILLER_169_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_418 ();
 DECAPx10_ASAP7_75t_R FILLER_169_425 ();
 DECAPx1_ASAP7_75t_R FILLER_169_447 ();
 DECAPx2_ASAP7_75t_R FILLER_169_477 ();
 FILLER_ASAP7_75t_R FILLER_169_483 ();
 DECAPx4_ASAP7_75t_R FILLER_169_495 ();
 FILLER_ASAP7_75t_R FILLER_169_505 ();
 FILLER_ASAP7_75t_R FILLER_169_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_512 ();
 DECAPx4_ASAP7_75t_R FILLER_169_519 ();
 FILLER_ASAP7_75t_R FILLER_169_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_531 ();
 DECAPx2_ASAP7_75t_R FILLER_169_538 ();
 DECAPx6_ASAP7_75t_R FILLER_169_562 ();
 DECAPx1_ASAP7_75t_R FILLER_169_576 ();
 DECAPx1_ASAP7_75t_R FILLER_169_596 ();
 DECAPx4_ASAP7_75t_R FILLER_169_603 ();
 DECAPx2_ASAP7_75t_R FILLER_169_619 ();
 FILLER_ASAP7_75t_R FILLER_169_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_627 ();
 DECAPx10_ASAP7_75t_R FILLER_169_635 ();
 DECAPx6_ASAP7_75t_R FILLER_169_697 ();
 FILLER_ASAP7_75t_R FILLER_169_711 ();
 DECAPx4_ASAP7_75t_R FILLER_169_726 ();
 FILLER_ASAP7_75t_R FILLER_169_736 ();
 DECAPx4_ASAP7_75t_R FILLER_169_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_754 ();
 DECAPx2_ASAP7_75t_R FILLER_169_768 ();
 FILLER_ASAP7_75t_R FILLER_169_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_795 ();
 DECAPx1_ASAP7_75t_R FILLER_169_802 ();
 DECAPx1_ASAP7_75t_R FILLER_169_812 ();
 DECAPx6_ASAP7_75t_R FILLER_169_822 ();
 FILLER_ASAP7_75t_R FILLER_169_836 ();
 DECAPx2_ASAP7_75t_R FILLER_169_848 ();
 FILLER_ASAP7_75t_R FILLER_169_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_856 ();
 DECAPx4_ASAP7_75t_R FILLER_169_863 ();
 FILLER_ASAP7_75t_R FILLER_169_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_875 ();
 DECAPx6_ASAP7_75t_R FILLER_169_895 ();
 DECAPx2_ASAP7_75t_R FILLER_169_909 ();
 FILLER_ASAP7_75t_R FILLER_169_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_923 ();
 DECAPx4_ASAP7_75t_R FILLER_169_941 ();
 FILLER_ASAP7_75t_R FILLER_169_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_953 ();
 DECAPx2_ASAP7_75t_R FILLER_169_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_977 ();
 DECAPx10_ASAP7_75t_R FILLER_169_981 ();
 FILLER_ASAP7_75t_R FILLER_169_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_169_1085 ();
 DECAPx4_ASAP7_75t_R FILLER_169_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1138 ();
 FILLER_ASAP7_75t_R FILLER_169_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1173 ();
 FILLER_ASAP7_75t_R FILLER_169_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1219 ();
 DECAPx6_ASAP7_75t_R FILLER_169_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_169_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1246 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1280 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1286 ();
 FILLER_ASAP7_75t_R FILLER_169_1294 ();
 DECAPx6_ASAP7_75t_R FILLER_169_1303 ();
 FILLER_ASAP7_75t_R FILLER_169_1317 ();
 DECAPx4_ASAP7_75t_R FILLER_169_1329 ();
 DECAPx4_ASAP7_75t_R FILLER_169_1365 ();
 FILLER_ASAP7_75t_R FILLER_169_1375 ();
 FILLER_ASAP7_75t_R FILLER_169_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_170_2 ();
 FILLER_ASAP7_75t_R FILLER_170_8 ();
 DECAPx4_ASAP7_75t_R FILLER_170_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_40 ();
 DECAPx6_ASAP7_75t_R FILLER_170_47 ();
 DECAPx1_ASAP7_75t_R FILLER_170_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_75 ();
 DECAPx1_ASAP7_75t_R FILLER_170_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_110 ();
 FILLER_ASAP7_75t_R FILLER_170_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_116 ();
 DECAPx1_ASAP7_75t_R FILLER_170_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_131 ();
 FILLER_ASAP7_75t_R FILLER_170_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_158 ();
 DECAPx1_ASAP7_75t_R FILLER_170_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_166 ();
 DECAPx1_ASAP7_75t_R FILLER_170_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_175 ();
 FILLER_ASAP7_75t_R FILLER_170_182 ();
 DECAPx2_ASAP7_75t_R FILLER_170_194 ();
 FILLER_ASAP7_75t_R FILLER_170_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_202 ();
 DECAPx1_ASAP7_75t_R FILLER_170_213 ();
 DECAPx2_ASAP7_75t_R FILLER_170_235 ();
 FILLER_ASAP7_75t_R FILLER_170_241 ();
 FILLER_ASAP7_75t_R FILLER_170_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_259 ();
 DECAPx1_ASAP7_75t_R FILLER_170_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_300 ();
 DECAPx6_ASAP7_75t_R FILLER_170_319 ();
 FILLER_ASAP7_75t_R FILLER_170_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_348 ();
 DECAPx6_ASAP7_75t_R FILLER_170_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_402 ();
 DECAPx6_ASAP7_75t_R FILLER_170_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_420 ();
 DECAPx4_ASAP7_75t_R FILLER_170_427 ();
 FILLER_ASAP7_75t_R FILLER_170_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_439 ();
 DECAPx1_ASAP7_75t_R FILLER_170_458 ();
 FILLER_ASAP7_75t_R FILLER_170_464 ();
 FILLER_ASAP7_75t_R FILLER_170_469 ();
 DECAPx4_ASAP7_75t_R FILLER_170_477 ();
 FILLER_ASAP7_75t_R FILLER_170_487 ();
 DECAPx4_ASAP7_75t_R FILLER_170_499 ();
 FILLER_ASAP7_75t_R FILLER_170_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_526 ();
 DECAPx1_ASAP7_75t_R FILLER_170_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_539 ();
 DECAPx10_ASAP7_75t_R FILLER_170_546 ();
 DECAPx6_ASAP7_75t_R FILLER_170_568 ();
 FILLER_ASAP7_75t_R FILLER_170_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_611 ();
 DECAPx2_ASAP7_75t_R FILLER_170_618 ();
 FILLER_ASAP7_75t_R FILLER_170_624 ();
 DECAPx6_ASAP7_75t_R FILLER_170_638 ();
 DECAPx1_ASAP7_75t_R FILLER_170_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_656 ();
 DECAPx10_ASAP7_75t_R FILLER_170_701 ();
 DECAPx2_ASAP7_75t_R FILLER_170_723 ();
 DECAPx1_ASAP7_75t_R FILLER_170_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_748 ();
 DECAPx4_ASAP7_75t_R FILLER_170_767 ();
 FILLER_ASAP7_75t_R FILLER_170_777 ();
 DECAPx1_ASAP7_75t_R FILLER_170_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_801 ();
 FILLER_ASAP7_75t_R FILLER_170_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_828 ();
 DECAPx4_ASAP7_75t_R FILLER_170_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_866 ();
 DECAPx4_ASAP7_75t_R FILLER_170_873 ();
 FILLER_ASAP7_75t_R FILLER_170_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_885 ();
 DECAPx1_ASAP7_75t_R FILLER_170_895 ();
 DECAPx4_ASAP7_75t_R FILLER_170_939 ();
 DECAPx2_ASAP7_75t_R FILLER_170_962 ();
 FILLER_ASAP7_75t_R FILLER_170_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_970 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1023 ();
 FILLER_ASAP7_75t_R FILLER_170_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1115 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1129 ();
 FILLER_ASAP7_75t_R FILLER_170_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1148 ();
 FILLER_ASAP7_75t_R FILLER_170_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1191 ();
 FILLER_ASAP7_75t_R FILLER_170_1205 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1210 ();
 FILLER_ASAP7_75t_R FILLER_170_1216 ();
 DECAPx1_ASAP7_75t_R FILLER_170_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1250 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1261 ();
 FILLER_ASAP7_75t_R FILLER_170_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1288 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1380 ();
 FILLER_ASAP7_75t_R FILLER_170_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_170_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_171_2 ();
 DECAPx1_ASAP7_75t_R FILLER_171_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_20 ();
 DECAPx1_ASAP7_75t_R FILLER_171_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_35 ();
 DECAPx1_ASAP7_75t_R FILLER_171_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_76 ();
 FILLER_ASAP7_75t_R FILLER_171_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_94 ();
 DECAPx4_ASAP7_75t_R FILLER_171_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_108 ();
 FILLER_ASAP7_75t_R FILLER_171_127 ();
 DECAPx1_ASAP7_75t_R FILLER_171_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_143 ();
 FILLER_ASAP7_75t_R FILLER_171_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_172 ();
 DECAPx1_ASAP7_75t_R FILLER_171_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_203 ();
 DECAPx2_ASAP7_75t_R FILLER_171_230 ();
 FILLER_ASAP7_75t_R FILLER_171_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_238 ();
 DECAPx2_ASAP7_75t_R FILLER_171_257 ();
 FILLER_ASAP7_75t_R FILLER_171_263 ();
 DECAPx1_ASAP7_75t_R FILLER_171_271 ();
 FILLER_ASAP7_75t_R FILLER_171_278 ();
 DECAPx2_ASAP7_75t_R FILLER_171_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_366 ();
 DECAPx4_ASAP7_75t_R FILLER_171_403 ();
 DECAPx4_ASAP7_75t_R FILLER_171_439 ();
 FILLER_ASAP7_75t_R FILLER_171_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_464 ();
 FILLER_ASAP7_75t_R FILLER_171_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_503 ();
 FILLER_ASAP7_75t_R FILLER_171_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_515 ();
 FILLER_ASAP7_75t_R FILLER_171_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_569 ();
 DECAPx6_ASAP7_75t_R FILLER_171_596 ();
 DECAPx1_ASAP7_75t_R FILLER_171_610 ();
 DECAPx1_ASAP7_75t_R FILLER_171_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_658 ();
 FILLER_ASAP7_75t_R FILLER_171_687 ();
 DECAPx2_ASAP7_75t_R FILLER_171_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_708 ();
 FILLER_ASAP7_75t_R FILLER_171_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_717 ();
 FILLER_ASAP7_75t_R FILLER_171_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_740 ();
 DECAPx2_ASAP7_75t_R FILLER_171_747 ();
 DECAPx6_ASAP7_75t_R FILLER_171_760 ();
 FILLER_ASAP7_75t_R FILLER_171_774 ();
 DECAPx4_ASAP7_75t_R FILLER_171_782 ();
 FILLER_ASAP7_75t_R FILLER_171_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_794 ();
 FILLER_ASAP7_75t_R FILLER_171_801 ();
 FILLER_ASAP7_75t_R FILLER_171_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_813 ();
 DECAPx6_ASAP7_75t_R FILLER_171_830 ();
 FILLER_ASAP7_75t_R FILLER_171_844 ();
 FILLER_ASAP7_75t_R FILLER_171_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_864 ();
 DECAPx4_ASAP7_75t_R FILLER_171_875 ();
 FILLER_ASAP7_75t_R FILLER_171_885 ();
 DECAPx2_ASAP7_75t_R FILLER_171_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_897 ();
 DECAPx6_ASAP7_75t_R FILLER_171_910 ();
 FILLER_ASAP7_75t_R FILLER_171_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_928 ();
 FILLER_ASAP7_75t_R FILLER_171_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_937 ();
 FILLER_ASAP7_75t_R FILLER_171_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_956 ();
 DECAPx4_ASAP7_75t_R FILLER_171_983 ();
 DECAPx2_ASAP7_75t_R FILLER_171_998 ();
 FILLER_ASAP7_75t_R FILLER_171_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1006 ();
 FILLER_ASAP7_75t_R FILLER_171_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1013 ();
 FILLER_ASAP7_75t_R FILLER_171_1025 ();
 FILLER_ASAP7_75t_R FILLER_171_1030 ();
 FILLER_ASAP7_75t_R FILLER_171_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1066 ();
 FILLER_ASAP7_75t_R FILLER_171_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1106 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1115 ();
 FILLER_ASAP7_75t_R FILLER_171_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1130 ();
 FILLER_ASAP7_75t_R FILLER_171_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1162 ();
 FILLER_ASAP7_75t_R FILLER_171_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1184 ();
 FILLER_ASAP7_75t_R FILLER_171_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1217 ();
 FILLER_ASAP7_75t_R FILLER_171_1239 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1296 ();
 FILLER_ASAP7_75t_R FILLER_171_1328 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_172_2 ();
 DECAPx2_ASAP7_75t_R FILLER_172_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_22 ();
 DECAPx1_ASAP7_75t_R FILLER_172_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_44 ();
 DECAPx1_ASAP7_75t_R FILLER_172_55 ();
 FILLER_ASAP7_75t_R FILLER_172_73 ();
 DECAPx1_ASAP7_75t_R FILLER_172_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_115 ();
 FILLER_ASAP7_75t_R FILLER_172_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_146 ();
 DECAPx10_ASAP7_75t_R FILLER_172_153 ();
 DECAPx1_ASAP7_75t_R FILLER_172_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_186 ();
 DECAPx6_ASAP7_75t_R FILLER_172_190 ();
 DECAPx1_ASAP7_75t_R FILLER_172_204 ();
 DECAPx1_ASAP7_75t_R FILLER_172_214 ();
 DECAPx1_ASAP7_75t_R FILLER_172_221 ();
 DECAPx6_ASAP7_75t_R FILLER_172_234 ();
 FILLER_ASAP7_75t_R FILLER_172_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_250 ();
 DECAPx4_ASAP7_75t_R FILLER_172_261 ();
 DECAPx10_ASAP7_75t_R FILLER_172_277 ();
 DECAPx10_ASAP7_75t_R FILLER_172_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_340 ();
 DECAPx10_ASAP7_75t_R FILLER_172_359 ();
 FILLER_ASAP7_75t_R FILLER_172_381 ();
 DECAPx2_ASAP7_75t_R FILLER_172_393 ();
 FILLER_ASAP7_75t_R FILLER_172_417 ();
 DECAPx6_ASAP7_75t_R FILLER_172_445 ();
 FILLER_ASAP7_75t_R FILLER_172_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_461 ();
 FILLER_ASAP7_75t_R FILLER_172_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_466 ();
 DECAPx2_ASAP7_75t_R FILLER_172_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_479 ();
 FILLER_ASAP7_75t_R FILLER_172_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_488 ();
 DECAPx2_ASAP7_75t_R FILLER_172_515 ();
 FILLER_ASAP7_75t_R FILLER_172_521 ();
 DECAPx1_ASAP7_75t_R FILLER_172_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_535 ();
 DECAPx1_ASAP7_75t_R FILLER_172_553 ();
 DECAPx4_ASAP7_75t_R FILLER_172_560 ();
 FILLER_ASAP7_75t_R FILLER_172_588 ();
 FILLER_ASAP7_75t_R FILLER_172_604 ();
 DECAPx1_ASAP7_75t_R FILLER_172_624 ();
 FILLER_ASAP7_75t_R FILLER_172_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_633 ();
 DECAPx1_ASAP7_75t_R FILLER_172_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_664 ();
 DECAPx2_ASAP7_75t_R FILLER_172_671 ();
 FILLER_ASAP7_75t_R FILLER_172_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_679 ();
 DECAPx1_ASAP7_75t_R FILLER_172_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_711 ();
 FILLER_ASAP7_75t_R FILLER_172_719 ();
 DECAPx1_ASAP7_75t_R FILLER_172_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_739 ();
 DECAPx10_ASAP7_75t_R FILLER_172_748 ();
 DECAPx2_ASAP7_75t_R FILLER_172_770 ();
 DECAPx6_ASAP7_75t_R FILLER_172_782 ();
 DECAPx4_ASAP7_75t_R FILLER_172_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_812 ();
 DECAPx4_ASAP7_75t_R FILLER_172_819 ();
 FILLER_ASAP7_75t_R FILLER_172_829 ();
 DECAPx2_ASAP7_75t_R FILLER_172_846 ();
 FILLER_ASAP7_75t_R FILLER_172_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_864 ();
 DECAPx4_ASAP7_75t_R FILLER_172_871 ();
 DECAPx1_ASAP7_75t_R FILLER_172_893 ();
 FILLER_ASAP7_75t_R FILLER_172_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_908 ();
 DECAPx2_ASAP7_75t_R FILLER_172_915 ();
 FILLER_ASAP7_75t_R FILLER_172_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_923 ();
 DECAPx2_ASAP7_75t_R FILLER_172_941 ();
 DECAPx4_ASAP7_75t_R FILLER_172_959 ();
 FILLER_ASAP7_75t_R FILLER_172_969 ();
 DECAPx10_ASAP7_75t_R FILLER_172_974 ();
 DECAPx2_ASAP7_75t_R FILLER_172_996 ();
 FILLER_ASAP7_75t_R FILLER_172_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1025 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1054 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1068 ();
 FILLER_ASAP7_75t_R FILLER_172_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1094 ();
 FILLER_ASAP7_75t_R FILLER_172_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1102 ();
 FILLER_ASAP7_75t_R FILLER_172_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1155 ();
 FILLER_ASAP7_75t_R FILLER_172_1161 ();
 FILLER_ASAP7_75t_R FILLER_172_1177 ();
 DECAPx4_ASAP7_75t_R FILLER_172_1187 ();
 FILLER_ASAP7_75t_R FILLER_172_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1199 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1240 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1265 ();
 FILLER_ASAP7_75t_R FILLER_172_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1281 ();
 FILLER_ASAP7_75t_R FILLER_172_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1310 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1321 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1335 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1355 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1373 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_173_2 ();
 FILLER_ASAP7_75t_R FILLER_173_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_18 ();
 DECAPx2_ASAP7_75t_R FILLER_173_29 ();
 FILLER_ASAP7_75t_R FILLER_173_35 ();
 DECAPx2_ASAP7_75t_R FILLER_173_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_49 ();
 DECAPx10_ASAP7_75t_R FILLER_173_53 ();
 DECAPx2_ASAP7_75t_R FILLER_173_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_81 ();
 DECAPx10_ASAP7_75t_R FILLER_173_88 ();
 DECAPx10_ASAP7_75t_R FILLER_173_110 ();
 DECAPx6_ASAP7_75t_R FILLER_173_132 ();
 DECAPx1_ASAP7_75t_R FILLER_173_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_150 ();
 DECAPx10_ASAP7_75t_R FILLER_173_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_183 ();
 DECAPx10_ASAP7_75t_R FILLER_173_196 ();
 DECAPx10_ASAP7_75t_R FILLER_173_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_240 ();
 FILLER_ASAP7_75t_R FILLER_173_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_246 ();
 DECAPx6_ASAP7_75t_R FILLER_173_253 ();
 FILLER_ASAP7_75t_R FILLER_173_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_269 ();
 DECAPx1_ASAP7_75t_R FILLER_173_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_283 ();
 DECAPx1_ASAP7_75t_R FILLER_173_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_291 ();
 DECAPx1_ASAP7_75t_R FILLER_173_302 ();
 DECAPx10_ASAP7_75t_R FILLER_173_324 ();
 DECAPx4_ASAP7_75t_R FILLER_173_346 ();
 DECAPx10_ASAP7_75t_R FILLER_173_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_407 ();
 DECAPx2_ASAP7_75t_R FILLER_173_420 ();
 DECAPx6_ASAP7_75t_R FILLER_173_441 ();
 DECAPx2_ASAP7_75t_R FILLER_173_455 ();
 DECAPx4_ASAP7_75t_R FILLER_173_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_489 ();
 DECAPx2_ASAP7_75t_R FILLER_173_496 ();
 FILLER_ASAP7_75t_R FILLER_173_502 ();
 DECAPx4_ASAP7_75t_R FILLER_173_507 ();
 FILLER_ASAP7_75t_R FILLER_173_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_519 ();
 DECAPx4_ASAP7_75t_R FILLER_173_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_538 ();
 DECAPx4_ASAP7_75t_R FILLER_173_546 ();
 DECAPx10_ASAP7_75t_R FILLER_173_562 ();
 DECAPx1_ASAP7_75t_R FILLER_173_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_588 ();
 DECAPx6_ASAP7_75t_R FILLER_173_595 ();
 DECAPx1_ASAP7_75t_R FILLER_173_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_623 ();
 DECAPx4_ASAP7_75t_R FILLER_173_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_670 ();
 DECAPx6_ASAP7_75t_R FILLER_173_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_692 ();
 DECAPx2_ASAP7_75t_R FILLER_173_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_718 ();
 FILLER_ASAP7_75t_R FILLER_173_729 ();
 DECAPx2_ASAP7_75t_R FILLER_173_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_743 ();
 DECAPx1_ASAP7_75t_R FILLER_173_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_759 ();
 FILLER_ASAP7_75t_R FILLER_173_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_778 ();
 FILLER_ASAP7_75t_R FILLER_173_785 ();
 FILLER_ASAP7_75t_R FILLER_173_793 ();
 DECAPx4_ASAP7_75t_R FILLER_173_813 ();
 DECAPx10_ASAP7_75t_R FILLER_173_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_861 ();
 FILLER_ASAP7_75t_R FILLER_173_872 ();
 DECAPx2_ASAP7_75t_R FILLER_173_890 ();
 FILLER_ASAP7_75t_R FILLER_173_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_898 ();
 FILLER_ASAP7_75t_R FILLER_173_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_908 ();
 DECAPx1_ASAP7_75t_R FILLER_173_920 ();
 DECAPx2_ASAP7_75t_R FILLER_173_942 ();
 DECAPx6_ASAP7_75t_R FILLER_173_960 ();
 FILLER_ASAP7_75t_R FILLER_173_974 ();
 FILLER_ASAP7_75t_R FILLER_173_988 ();
 DECAPx6_ASAP7_75t_R FILLER_173_1008 ();
 FILLER_ASAP7_75t_R FILLER_173_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1024 ();
 DECAPx6_ASAP7_75t_R FILLER_173_1032 ();
 FILLER_ASAP7_75t_R FILLER_173_1046 ();
 FILLER_ASAP7_75t_R FILLER_173_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_173_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1087 ();
 FILLER_ASAP7_75t_R FILLER_173_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1111 ();
 FILLER_ASAP7_75t_R FILLER_173_1164 ();
 DECAPx4_ASAP7_75t_R FILLER_173_1192 ();
 FILLER_ASAP7_75t_R FILLER_173_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1204 ();
 FILLER_ASAP7_75t_R FILLER_173_1213 ();
 FILLER_ASAP7_75t_R FILLER_173_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1220 ();
 DECAPx1_ASAP7_75t_R FILLER_173_1249 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1263 ();
 FILLER_ASAP7_75t_R FILLER_173_1269 ();
 FILLER_ASAP7_75t_R FILLER_173_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1319 ();
 FILLER_ASAP7_75t_R FILLER_173_1341 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1359 ();
 DECAPx6_ASAP7_75t_R FILLER_174_2 ();
 FILLER_ASAP7_75t_R FILLER_174_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_18 ();
 DECAPx2_ASAP7_75t_R FILLER_174_29 ();
 DECAPx1_ASAP7_75t_R FILLER_174_45 ();
 DECAPx6_ASAP7_75t_R FILLER_174_52 ();
 DECAPx1_ASAP7_75t_R FILLER_174_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_70 ();
 DECAPx2_ASAP7_75t_R FILLER_174_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_83 ();
 DECAPx6_ASAP7_75t_R FILLER_174_93 ();
 FILLER_ASAP7_75t_R FILLER_174_107 ();
 FILLER_ASAP7_75t_R FILLER_174_127 ();
 FILLER_ASAP7_75t_R FILLER_174_147 ();
 DECAPx6_ASAP7_75t_R FILLER_174_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_210 ();
 FILLER_ASAP7_75t_R FILLER_174_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_225 ();
 DECAPx4_ASAP7_75t_R FILLER_174_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_265 ();
 DECAPx6_ASAP7_75t_R FILLER_174_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_306 ();
 DECAPx2_ASAP7_75t_R FILLER_174_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_347 ();
 DECAPx4_ASAP7_75t_R FILLER_174_351 ();
 FILLER_ASAP7_75t_R FILLER_174_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_363 ();
 DECAPx2_ASAP7_75t_R FILLER_174_400 ();
 FILLER_ASAP7_75t_R FILLER_174_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_423 ();
 DECAPx2_ASAP7_75t_R FILLER_174_428 ();
 DECAPx1_ASAP7_75t_R FILLER_174_437 ();
 DECAPx4_ASAP7_75t_R FILLER_174_449 ();
 FILLER_ASAP7_75t_R FILLER_174_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_461 ();
 DECAPx2_ASAP7_75t_R FILLER_174_492 ();
 FILLER_ASAP7_75t_R FILLER_174_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_500 ();
 DECAPx1_ASAP7_75t_R FILLER_174_505 ();
 DECAPx1_ASAP7_75t_R FILLER_174_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_524 ();
 DECAPx2_ASAP7_75t_R FILLER_174_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_539 ();
 DECAPx4_ASAP7_75t_R FILLER_174_547 ();
 FILLER_ASAP7_75t_R FILLER_174_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_559 ();
 DECAPx2_ASAP7_75t_R FILLER_174_578 ();
 FILLER_ASAP7_75t_R FILLER_174_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_586 ();
 DECAPx4_ASAP7_75t_R FILLER_174_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_607 ();
 DECAPx1_ASAP7_75t_R FILLER_174_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_622 ();
 FILLER_ASAP7_75t_R FILLER_174_651 ();
 DECAPx4_ASAP7_75t_R FILLER_174_660 ();
 FILLER_ASAP7_75t_R FILLER_174_670 ();
 DECAPx1_ASAP7_75t_R FILLER_174_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_682 ();
 FILLER_ASAP7_75t_R FILLER_174_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_695 ();
 DECAPx2_ASAP7_75t_R FILLER_174_702 ();
 DECAPx2_ASAP7_75t_R FILLER_174_714 ();
 FILLER_ASAP7_75t_R FILLER_174_730 ();
 DECAPx1_ASAP7_75t_R FILLER_174_738 ();
 DECAPx4_ASAP7_75t_R FILLER_174_750 ();
 FILLER_ASAP7_75t_R FILLER_174_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_778 ();
 DECAPx1_ASAP7_75t_R FILLER_174_809 ();
 DECAPx2_ASAP7_75t_R FILLER_174_835 ();
 DECAPx10_ASAP7_75t_R FILLER_174_847 ();
 FILLER_ASAP7_75t_R FILLER_174_869 ();
 DECAPx2_ASAP7_75t_R FILLER_174_889 ();
 FILLER_ASAP7_75t_R FILLER_174_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_897 ();
 DECAPx10_ASAP7_75t_R FILLER_174_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_945 ();
 DECAPx2_ASAP7_75t_R FILLER_174_960 ();
 FILLER_ASAP7_75t_R FILLER_174_966 ();
 DECAPx2_ASAP7_75t_R FILLER_174_986 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1086 ();
 DECAPx4_ASAP7_75t_R FILLER_174_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1151 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1223 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1245 ();
 DECAPx4_ASAP7_75t_R FILLER_174_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1311 ();
 FILLER_ASAP7_75t_R FILLER_174_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1337 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_175_2 ();
 FILLER_ASAP7_75t_R FILLER_175_16 ();
 DECAPx2_ASAP7_75t_R FILLER_175_28 ();
 DECAPx1_ASAP7_75t_R FILLER_175_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_68 ();
 DECAPx2_ASAP7_75t_R FILLER_175_99 ();
 FILLER_ASAP7_75t_R FILLER_175_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_126 ();
 FILLER_ASAP7_75t_R FILLER_175_135 ();
 FILLER_ASAP7_75t_R FILLER_175_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_168 ();
 DECAPx1_ASAP7_75t_R FILLER_175_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_213 ();
 FILLER_ASAP7_75t_R FILLER_175_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_224 ();
 DECAPx2_ASAP7_75t_R FILLER_175_241 ();
 DECAPx4_ASAP7_75t_R FILLER_175_279 ();
 DECAPx6_ASAP7_75t_R FILLER_175_359 ();
 FILLER_ASAP7_75t_R FILLER_175_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_375 ();
 DECAPx1_ASAP7_75t_R FILLER_175_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_424 ();
 FILLER_ASAP7_75t_R FILLER_175_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_443 ();
 DECAPx4_ASAP7_75t_R FILLER_175_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_472 ();
 FILLER_ASAP7_75t_R FILLER_175_493 ();
 FILLER_ASAP7_75t_R FILLER_175_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_531 ();
 DECAPx2_ASAP7_75t_R FILLER_175_550 ();
 DECAPx2_ASAP7_75t_R FILLER_175_598 ();
 FILLER_ASAP7_75t_R FILLER_175_604 ();
 DECAPx4_ASAP7_75t_R FILLER_175_624 ();
 DECAPx4_ASAP7_75t_R FILLER_175_677 ();
 FILLER_ASAP7_75t_R FILLER_175_687 ();
 FILLER_ASAP7_75t_R FILLER_175_699 ();
 DECAPx2_ASAP7_75t_R FILLER_175_721 ();
 FILLER_ASAP7_75t_R FILLER_175_727 ();
 FILLER_ASAP7_75t_R FILLER_175_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_737 ();
 DECAPx2_ASAP7_75t_R FILLER_175_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_762 ();
 DECAPx6_ASAP7_75t_R FILLER_175_769 ();
 FILLER_ASAP7_75t_R FILLER_175_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_785 ();
 DECAPx4_ASAP7_75t_R FILLER_175_792 ();
 FILLER_ASAP7_75t_R FILLER_175_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_804 ();
 FILLER_ASAP7_75t_R FILLER_175_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_815 ();
 DECAPx2_ASAP7_75t_R FILLER_175_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_853 ();
 DECAPx1_ASAP7_75t_R FILLER_175_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_876 ();
 DECAPx2_ASAP7_75t_R FILLER_175_897 ();
 FILLER_ASAP7_75t_R FILLER_175_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_905 ();
 DECAPx4_ASAP7_75t_R FILLER_175_914 ();
 DECAPx6_ASAP7_75t_R FILLER_175_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_940 ();
 DECAPx6_ASAP7_75t_R FILLER_175_978 ();
 DECAPx1_ASAP7_75t_R FILLER_175_992 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1014 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1086 ();
 DECAPx4_ASAP7_75t_R FILLER_175_1129 ();
 FILLER_ASAP7_75t_R FILLER_175_1139 ();
 FILLER_ASAP7_75t_R FILLER_175_1149 ();
 FILLER_ASAP7_75t_R FILLER_175_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1192 ();
 FILLER_ASAP7_75t_R FILLER_175_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1211 ();
 DECAPx4_ASAP7_75t_R FILLER_175_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1272 ();
 FILLER_ASAP7_75t_R FILLER_175_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1288 ();
 FILLER_ASAP7_75t_R FILLER_175_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1365 ();
 DECAPx4_ASAP7_75t_R FILLER_176_2 ();
 FILLER_ASAP7_75t_R FILLER_176_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_14 ();
 DECAPx2_ASAP7_75t_R FILLER_176_27 ();
 FILLER_ASAP7_75t_R FILLER_176_33 ();
 FILLER_ASAP7_75t_R FILLER_176_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_43 ();
 DECAPx10_ASAP7_75t_R FILLER_176_74 ();
 FILLER_ASAP7_75t_R FILLER_176_96 ();
 DECAPx6_ASAP7_75t_R FILLER_176_106 ();
 FILLER_ASAP7_75t_R FILLER_176_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_122 ();
 FILLER_ASAP7_75t_R FILLER_176_149 ();
 DECAPx1_ASAP7_75t_R FILLER_176_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_164 ();
 FILLER_ASAP7_75t_R FILLER_176_168 ();
 DECAPx4_ASAP7_75t_R FILLER_176_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_209 ();
 DECAPx10_ASAP7_75t_R FILLER_176_230 ();
 DECAPx4_ASAP7_75t_R FILLER_176_252 ();
 DECAPx6_ASAP7_75t_R FILLER_176_276 ();
 DECAPx2_ASAP7_75t_R FILLER_176_290 ();
 DECAPx2_ASAP7_75t_R FILLER_176_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_364 ();
 DECAPx10_ASAP7_75t_R FILLER_176_372 ();
 DECAPx2_ASAP7_75t_R FILLER_176_394 ();
 FILLER_ASAP7_75t_R FILLER_176_400 ();
 DECAPx4_ASAP7_75t_R FILLER_176_422 ();
 FILLER_ASAP7_75t_R FILLER_176_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_434 ();
 DECAPx6_ASAP7_75t_R FILLER_176_443 ();
 DECAPx1_ASAP7_75t_R FILLER_176_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_461 ();
 DECAPx2_ASAP7_75t_R FILLER_176_464 ();
 FILLER_ASAP7_75t_R FILLER_176_470 ();
 DECAPx6_ASAP7_75t_R FILLER_176_488 ();
 DECAPx1_ASAP7_75t_R FILLER_176_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_512 ();
 DECAPx1_ASAP7_75t_R FILLER_176_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_539 ();
 DECAPx4_ASAP7_75t_R FILLER_176_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_558 ();
 DECAPx1_ASAP7_75t_R FILLER_176_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_590 ();
 DECAPx10_ASAP7_75t_R FILLER_176_594 ();
 DECAPx10_ASAP7_75t_R FILLER_176_616 ();
 DECAPx10_ASAP7_75t_R FILLER_176_638 ();
 DECAPx10_ASAP7_75t_R FILLER_176_660 ();
 DECAPx4_ASAP7_75t_R FILLER_176_682 ();
 FILLER_ASAP7_75t_R FILLER_176_692 ();
 DECAPx4_ASAP7_75t_R FILLER_176_704 ();
 FILLER_ASAP7_75t_R FILLER_176_714 ();
 FILLER_ASAP7_75t_R FILLER_176_726 ();
 DECAPx1_ASAP7_75t_R FILLER_176_740 ();
 DECAPx1_ASAP7_75t_R FILLER_176_752 ();
 DECAPx6_ASAP7_75t_R FILLER_176_778 ();
 FILLER_ASAP7_75t_R FILLER_176_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_794 ();
 DECAPx4_ASAP7_75t_R FILLER_176_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_821 ();
 DECAPx1_ASAP7_75t_R FILLER_176_838 ();
 DECAPx4_ASAP7_75t_R FILLER_176_848 ();
 DECAPx2_ASAP7_75t_R FILLER_176_876 ();
 FILLER_ASAP7_75t_R FILLER_176_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_884 ();
 DECAPx4_ASAP7_75t_R FILLER_176_891 ();
 FILLER_ASAP7_75t_R FILLER_176_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_903 ();
 DECAPx6_ASAP7_75t_R FILLER_176_915 ();
 DECAPx1_ASAP7_75t_R FILLER_176_929 ();
 DECAPx1_ASAP7_75t_R FILLER_176_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_962 ();
 DECAPx10_ASAP7_75t_R FILLER_176_970 ();
 DECAPx10_ASAP7_75t_R FILLER_176_992 ();
 DECAPx6_ASAP7_75t_R FILLER_176_1014 ();
 FILLER_ASAP7_75t_R FILLER_176_1028 ();
 FILLER_ASAP7_75t_R FILLER_176_1033 ();
 FILLER_ASAP7_75t_R FILLER_176_1041 ();
 FILLER_ASAP7_75t_R FILLER_176_1057 ();
 FILLER_ASAP7_75t_R FILLER_176_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1127 ();
 FILLER_ASAP7_75t_R FILLER_176_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1135 ();
 FILLER_ASAP7_75t_R FILLER_176_1172 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1187 ();
 FILLER_ASAP7_75t_R FILLER_176_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1226 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1282 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1293 ();
 FILLER_ASAP7_75t_R FILLER_176_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1301 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_176_1353 ();
 FILLER_ASAP7_75t_R FILLER_176_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1388 ();
 FILLER_ASAP7_75t_R FILLER_177_32 ();
 DECAPx1_ASAP7_75t_R FILLER_177_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_48 ();
 DECAPx2_ASAP7_75t_R FILLER_177_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_70 ();
 FILLER_ASAP7_75t_R FILLER_177_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_81 ();
 DECAPx2_ASAP7_75t_R FILLER_177_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_91 ();
 DECAPx2_ASAP7_75t_R FILLER_177_118 ();
 FILLER_ASAP7_75t_R FILLER_177_124 ();
 DECAPx10_ASAP7_75t_R FILLER_177_132 ();
 DECAPx10_ASAP7_75t_R FILLER_177_154 ();
 DECAPx2_ASAP7_75t_R FILLER_177_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_182 ();
 DECAPx2_ASAP7_75t_R FILLER_177_186 ();
 FILLER_ASAP7_75t_R FILLER_177_192 ();
 DECAPx1_ASAP7_75t_R FILLER_177_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_212 ();
 DECAPx6_ASAP7_75t_R FILLER_177_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_267 ();
 FILLER_ASAP7_75t_R FILLER_177_271 ();
 DECAPx4_ASAP7_75t_R FILLER_177_279 ();
 FILLER_ASAP7_75t_R FILLER_177_289 ();
 DECAPx2_ASAP7_75t_R FILLER_177_309 ();
 FILLER_ASAP7_75t_R FILLER_177_315 ();
 FILLER_ASAP7_75t_R FILLER_177_354 ();
 DECAPx2_ASAP7_75t_R FILLER_177_364 ();
 DECAPx2_ASAP7_75t_R FILLER_177_396 ();
 FILLER_ASAP7_75t_R FILLER_177_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_424 ();
 FILLER_ASAP7_75t_R FILLER_177_437 ();
 DECAPx2_ASAP7_75t_R FILLER_177_445 ();
 FILLER_ASAP7_75t_R FILLER_177_451 ();
 FILLER_ASAP7_75t_R FILLER_177_479 ();
 FILLER_ASAP7_75t_R FILLER_177_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_489 ();
 FILLER_ASAP7_75t_R FILLER_177_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_515 ();
 FILLER_ASAP7_75t_R FILLER_177_538 ();
 DECAPx4_ASAP7_75t_R FILLER_177_546 ();
 FILLER_ASAP7_75t_R FILLER_177_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_558 ();
 DECAPx4_ASAP7_75t_R FILLER_177_567 ();
 DECAPx4_ASAP7_75t_R FILLER_177_586 ();
 DECAPx6_ASAP7_75t_R FILLER_177_599 ();
 DECAPx10_ASAP7_75t_R FILLER_177_621 ();
 FILLER_ASAP7_75t_R FILLER_177_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_645 ();
 DECAPx6_ASAP7_75t_R FILLER_177_682 ();
 DECAPx2_ASAP7_75t_R FILLER_177_696 ();
 DECAPx1_ASAP7_75t_R FILLER_177_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_726 ();
 FILLER_ASAP7_75t_R FILLER_177_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_750 ();
 FILLER_ASAP7_75t_R FILLER_177_767 ();
 DECAPx2_ASAP7_75t_R FILLER_177_797 ();
 FILLER_ASAP7_75t_R FILLER_177_803 ();
 DECAPx10_ASAP7_75t_R FILLER_177_813 ();
 DECAPx1_ASAP7_75t_R FILLER_177_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_839 ();
 DECAPx6_ASAP7_75t_R FILLER_177_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_860 ();
 DECAPx6_ASAP7_75t_R FILLER_177_877 ();
 FILLER_ASAP7_75t_R FILLER_177_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_893 ();
 DECAPx1_ASAP7_75t_R FILLER_177_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_905 ();
 DECAPx2_ASAP7_75t_R FILLER_177_912 ();
 DECAPx4_ASAP7_75t_R FILLER_177_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_942 ();
 DECAPx10_ASAP7_75t_R FILLER_177_951 ();
 DECAPx2_ASAP7_75t_R FILLER_177_973 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1103 ();
 DECAPx4_ASAP7_75t_R FILLER_177_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1133 ();
 FILLER_ASAP7_75t_R FILLER_177_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_177_1196 ();
 FILLER_ASAP7_75t_R FILLER_177_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1244 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1271 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1295 ();
 FILLER_ASAP7_75t_R FILLER_177_1314 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1333 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1337 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1348 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1365 ();
 FILLER_ASAP7_75t_R FILLER_177_1372 ();
 DECAPx4_ASAP7_75t_R FILLER_178_2 ();
 FILLER_ASAP7_75t_R FILLER_178_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_14 ();
 DECAPx10_ASAP7_75t_R FILLER_178_18 ();
 FILLER_ASAP7_75t_R FILLER_178_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_49 ();
 DECAPx6_ASAP7_75t_R FILLER_178_53 ();
 DECAPx1_ASAP7_75t_R FILLER_178_93 ();
 DECAPx1_ASAP7_75t_R FILLER_178_103 ();
 DECAPx4_ASAP7_75t_R FILLER_178_110 ();
 DECAPx1_ASAP7_75t_R FILLER_178_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_176 ();
 DECAPx6_ASAP7_75t_R FILLER_178_183 ();
 DECAPx2_ASAP7_75t_R FILLER_178_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_209 ();
 DECAPx6_ASAP7_75t_R FILLER_178_224 ();
 FILLER_ASAP7_75t_R FILLER_178_238 ();
 DECAPx1_ASAP7_75t_R FILLER_178_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_267 ();
 FILLER_ASAP7_75t_R FILLER_178_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_358 ();
 FILLER_ASAP7_75t_R FILLER_178_367 ();
 DECAPx10_ASAP7_75t_R FILLER_178_414 ();
 FILLER_ASAP7_75t_R FILLER_178_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_466 ();
 FILLER_ASAP7_75t_R FILLER_178_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_490 ();
 DECAPx2_ASAP7_75t_R FILLER_178_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_504 ();
 DECAPx2_ASAP7_75t_R FILLER_178_508 ();
 FILLER_ASAP7_75t_R FILLER_178_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_526 ();
 DECAPx4_ASAP7_75t_R FILLER_178_533 ();
 FILLER_ASAP7_75t_R FILLER_178_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_545 ();
 DECAPx1_ASAP7_75t_R FILLER_178_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_607 ();
 DECAPx2_ASAP7_75t_R FILLER_178_640 ();
 FILLER_ASAP7_75t_R FILLER_178_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_660 ();
 FILLER_ASAP7_75t_R FILLER_178_664 ();
 FILLER_ASAP7_75t_R FILLER_178_692 ();
 DECAPx2_ASAP7_75t_R FILLER_178_704 ();
 FILLER_ASAP7_75t_R FILLER_178_710 ();
 FILLER_ASAP7_75t_R FILLER_178_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_724 ();
 DECAPx10_ASAP7_75t_R FILLER_178_740 ();
 DECAPx2_ASAP7_75t_R FILLER_178_762 ();
 FILLER_ASAP7_75t_R FILLER_178_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_770 ();
 DECAPx6_ASAP7_75t_R FILLER_178_787 ();
 DECAPx1_ASAP7_75t_R FILLER_178_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_805 ();
 FILLER_ASAP7_75t_R FILLER_178_812 ();
 DECAPx4_ASAP7_75t_R FILLER_178_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_841 ();
 DECAPx6_ASAP7_75t_R FILLER_178_848 ();
 DECAPx2_ASAP7_75t_R FILLER_178_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_868 ();
 DECAPx6_ASAP7_75t_R FILLER_178_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_930 ();
 FILLER_ASAP7_75t_R FILLER_178_943 ();
 DECAPx6_ASAP7_75t_R FILLER_178_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_969 ();
 FILLER_ASAP7_75t_R FILLER_178_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1214 ();
 FILLER_ASAP7_75t_R FILLER_178_1220 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1241 ();
 FILLER_ASAP7_75t_R FILLER_178_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1286 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1306 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1324 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1333 ();
 FILLER_ASAP7_75t_R FILLER_178_1343 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1373 ();
 DECAPx1_ASAP7_75t_R FILLER_178_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_179_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_12 ();
 DECAPx2_ASAP7_75t_R FILLER_179_29 ();
 FILLER_ASAP7_75t_R FILLER_179_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_37 ();
 DECAPx1_ASAP7_75t_R FILLER_179_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_68 ();
 DECAPx4_ASAP7_75t_R FILLER_179_75 ();
 FILLER_ASAP7_75t_R FILLER_179_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_87 ();
 DECAPx4_ASAP7_75t_R FILLER_179_98 ();
 DECAPx2_ASAP7_75t_R FILLER_179_114 ();
 FILLER_ASAP7_75t_R FILLER_179_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_122 ();
 FILLER_ASAP7_75t_R FILLER_179_163 ();
 DECAPx1_ASAP7_75t_R FILLER_179_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_195 ();
 DECAPx2_ASAP7_75t_R FILLER_179_210 ();
 DECAPx2_ASAP7_75t_R FILLER_179_230 ();
 FILLER_ASAP7_75t_R FILLER_179_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_238 ();
 FILLER_ASAP7_75t_R FILLER_179_247 ();
 DECAPx4_ASAP7_75t_R FILLER_179_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_274 ();
 DECAPx6_ASAP7_75t_R FILLER_179_289 ();
 FILLER_ASAP7_75t_R FILLER_179_303 ();
 FILLER_ASAP7_75t_R FILLER_179_355 ();
 DECAPx6_ASAP7_75t_R FILLER_179_370 ();
 DECAPx2_ASAP7_75t_R FILLER_179_394 ();
 FILLER_ASAP7_75t_R FILLER_179_400 ();
 DECAPx6_ASAP7_75t_R FILLER_179_405 ();
 DECAPx2_ASAP7_75t_R FILLER_179_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_444 ();
 FILLER_ASAP7_75t_R FILLER_179_466 ();
 FILLER_ASAP7_75t_R FILLER_179_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_473 ();
 DECAPx6_ASAP7_75t_R FILLER_179_477 ();
 FILLER_ASAP7_75t_R FILLER_179_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_519 ();
 DECAPx2_ASAP7_75t_R FILLER_179_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_547 ();
 FILLER_ASAP7_75t_R FILLER_179_558 ();
 DECAPx2_ASAP7_75t_R FILLER_179_568 ();
 DECAPx2_ASAP7_75t_R FILLER_179_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_592 ();
 DECAPx1_ASAP7_75t_R FILLER_179_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_660 ();
 FILLER_ASAP7_75t_R FILLER_179_678 ();
 DECAPx1_ASAP7_75t_R FILLER_179_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_690 ();
 DECAPx10_ASAP7_75t_R FILLER_179_698 ();
 DECAPx2_ASAP7_75t_R FILLER_179_720 ();
 FILLER_ASAP7_75t_R FILLER_179_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_728 ();
 FILLER_ASAP7_75t_R FILLER_179_742 ();
 DECAPx6_ASAP7_75t_R FILLER_179_750 ();
 FILLER_ASAP7_75t_R FILLER_179_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_766 ();
 DECAPx2_ASAP7_75t_R FILLER_179_773 ();
 DECAPx2_ASAP7_75t_R FILLER_179_789 ();
 FILLER_ASAP7_75t_R FILLER_179_809 ();
 FILLER_ASAP7_75t_R FILLER_179_827 ();
 DECAPx1_ASAP7_75t_R FILLER_179_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_893 ();
 FILLER_ASAP7_75t_R FILLER_179_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_902 ();
 DECAPx2_ASAP7_75t_R FILLER_179_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_923 ();
 DECAPx4_ASAP7_75t_R FILLER_179_932 ();
 FILLER_ASAP7_75t_R FILLER_179_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_944 ();
 DECAPx2_ASAP7_75t_R FILLER_179_951 ();
 FILLER_ASAP7_75t_R FILLER_179_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_959 ();
 FILLER_ASAP7_75t_R FILLER_179_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_984 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1013 ();
 FILLER_ASAP7_75t_R FILLER_179_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1062 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1083 ();
 FILLER_ASAP7_75t_R FILLER_179_1089 ();
 FILLER_ASAP7_75t_R FILLER_179_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_179_1106 ();
 FILLER_ASAP7_75t_R FILLER_179_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1122 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1176 ();
 FILLER_ASAP7_75t_R FILLER_179_1200 ();
 FILLER_ASAP7_75t_R FILLER_179_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1216 ();
 FILLER_ASAP7_75t_R FILLER_179_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_179_1256 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1309 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1317 ();
 FILLER_ASAP7_75t_R FILLER_179_1333 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1342 ();
 FILLER_ASAP7_75t_R FILLER_179_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1391 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_39 ();
 DECAPx2_ASAP7_75t_R FILLER_180_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_52 ();
 DECAPx1_ASAP7_75t_R FILLER_180_56 ();
 DECAPx6_ASAP7_75t_R FILLER_180_92 ();
 FILLER_ASAP7_75t_R FILLER_180_139 ();
 DECAPx2_ASAP7_75t_R FILLER_180_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_164 ();
 DECAPx1_ASAP7_75t_R FILLER_180_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_172 ();
 DECAPx1_ASAP7_75t_R FILLER_180_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_197 ();
 DECAPx1_ASAP7_75t_R FILLER_180_204 ();
 DECAPx1_ASAP7_75t_R FILLER_180_216 ();
 FILLER_ASAP7_75t_R FILLER_180_233 ();
 FILLER_ASAP7_75t_R FILLER_180_249 ();
 FILLER_ASAP7_75t_R FILLER_180_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_259 ();
 DECAPx4_ASAP7_75t_R FILLER_180_266 ();
 DECAPx6_ASAP7_75t_R FILLER_180_284 ();
 DECAPx1_ASAP7_75t_R FILLER_180_298 ();
 DECAPx2_ASAP7_75t_R FILLER_180_320 ();
 FILLER_ASAP7_75t_R FILLER_180_326 ();
 DECAPx1_ASAP7_75t_R FILLER_180_368 ();
 DECAPx6_ASAP7_75t_R FILLER_180_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_404 ();
 DECAPx4_ASAP7_75t_R FILLER_180_411 ();
 FILLER_ASAP7_75t_R FILLER_180_421 ();
 DECAPx6_ASAP7_75t_R FILLER_180_441 ();
 DECAPx2_ASAP7_75t_R FILLER_180_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_461 ();
 DECAPx2_ASAP7_75t_R FILLER_180_464 ();
 DECAPx6_ASAP7_75t_R FILLER_180_478 ();
 FILLER_ASAP7_75t_R FILLER_180_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_494 ();
 DECAPx6_ASAP7_75t_R FILLER_180_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_515 ();
 FILLER_ASAP7_75t_R FILLER_180_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_532 ();
 DECAPx6_ASAP7_75t_R FILLER_180_539 ();
 DECAPx2_ASAP7_75t_R FILLER_180_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_559 ();
 DECAPx2_ASAP7_75t_R FILLER_180_566 ();
 FILLER_ASAP7_75t_R FILLER_180_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_574 ();
 DECAPx6_ASAP7_75t_R FILLER_180_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_627 ();
 DECAPx10_ASAP7_75t_R FILLER_180_631 ();
 DECAPx6_ASAP7_75t_R FILLER_180_653 ();
 DECAPx2_ASAP7_75t_R FILLER_180_685 ();
 FILLER_ASAP7_75t_R FILLER_180_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_704 ();
 DECAPx4_ASAP7_75t_R FILLER_180_713 ();
 FILLER_ASAP7_75t_R FILLER_180_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_725 ();
 FILLER_ASAP7_75t_R FILLER_180_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_775 ();
 DECAPx4_ASAP7_75t_R FILLER_180_812 ();
 FILLER_ASAP7_75t_R FILLER_180_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_844 ();
 DECAPx2_ASAP7_75t_R FILLER_180_855 ();
 FILLER_ASAP7_75t_R FILLER_180_861 ();
 DECAPx1_ASAP7_75t_R FILLER_180_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_891 ();
 DECAPx1_ASAP7_75t_R FILLER_180_902 ();
 DECAPx2_ASAP7_75t_R FILLER_180_938 ();
 DECAPx10_ASAP7_75t_R FILLER_180_952 ();
 DECAPx2_ASAP7_75t_R FILLER_180_974 ();
 FILLER_ASAP7_75t_R FILLER_180_980 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1000 ();
 FILLER_ASAP7_75t_R FILLER_180_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1014 ();
 FILLER_ASAP7_75t_R FILLER_180_1024 ();
 FILLER_ASAP7_75t_R FILLER_180_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1135 ();
 DECAPx6_ASAP7_75t_R FILLER_180_1162 ();
 FILLER_ASAP7_75t_R FILLER_180_1176 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1248 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1264 ();
 FILLER_ASAP7_75t_R FILLER_180_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1314 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1341 ();
 FILLER_ASAP7_75t_R FILLER_180_1351 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1367 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_181_2 ();
 FILLER_ASAP7_75t_R FILLER_181_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_14 ();
 FILLER_ASAP7_75t_R FILLER_181_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_57 ();
 DECAPx1_ASAP7_75t_R FILLER_181_70 ();
 FILLER_ASAP7_75t_R FILLER_181_77 ();
 FILLER_ASAP7_75t_R FILLER_181_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_111 ();
 DECAPx1_ASAP7_75t_R FILLER_181_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_119 ();
 DECAPx1_ASAP7_75t_R FILLER_181_123 ();
 DECAPx10_ASAP7_75t_R FILLER_181_133 ();
 DECAPx10_ASAP7_75t_R FILLER_181_155 ();
 DECAPx2_ASAP7_75t_R FILLER_181_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_183 ();
 DECAPx2_ASAP7_75t_R FILLER_181_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_196 ();
 FILLER_ASAP7_75t_R FILLER_181_203 ();
 DECAPx1_ASAP7_75t_R FILLER_181_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_225 ();
 FILLER_ASAP7_75t_R FILLER_181_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_235 ();
 DECAPx2_ASAP7_75t_R FILLER_181_242 ();
 FILLER_ASAP7_75t_R FILLER_181_248 ();
 DECAPx1_ASAP7_75t_R FILLER_181_257 ();
 FILLER_ASAP7_75t_R FILLER_181_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_271 ();
 DECAPx10_ASAP7_75t_R FILLER_181_286 ();
 DECAPx1_ASAP7_75t_R FILLER_181_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_312 ();
 FILLER_ASAP7_75t_R FILLER_181_323 ();
 FILLER_ASAP7_75t_R FILLER_181_343 ();
 DECAPx6_ASAP7_75t_R FILLER_181_363 ();
 DECAPx2_ASAP7_75t_R FILLER_181_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_383 ();
 DECAPx6_ASAP7_75t_R FILLER_181_416 ();
 DECAPx1_ASAP7_75t_R FILLER_181_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_434 ();
 DECAPx2_ASAP7_75t_R FILLER_181_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_491 ();
 DECAPx1_ASAP7_75t_R FILLER_181_507 ();
 DECAPx4_ASAP7_75t_R FILLER_181_524 ();
 FILLER_ASAP7_75t_R FILLER_181_534 ();
 DECAPx4_ASAP7_75t_R FILLER_181_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_560 ();
 DECAPx1_ASAP7_75t_R FILLER_181_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_571 ();
 DECAPx10_ASAP7_75t_R FILLER_181_578 ();
 DECAPx2_ASAP7_75t_R FILLER_181_600 ();
 FILLER_ASAP7_75t_R FILLER_181_606 ();
 DECAPx2_ASAP7_75t_R FILLER_181_614 ();
 FILLER_ASAP7_75t_R FILLER_181_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_622 ();
 FILLER_ASAP7_75t_R FILLER_181_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_631 ();
 DECAPx10_ASAP7_75t_R FILLER_181_638 ();
 DECAPx4_ASAP7_75t_R FILLER_181_660 ();
 DECAPx10_ASAP7_75t_R FILLER_181_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_705 ();
 DECAPx2_ASAP7_75t_R FILLER_181_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_729 ();
 DECAPx2_ASAP7_75t_R FILLER_181_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_744 ();
 DECAPx6_ASAP7_75t_R FILLER_181_773 ();
 DECAPx1_ASAP7_75t_R FILLER_181_787 ();
 DECAPx10_ASAP7_75t_R FILLER_181_811 ();
 DECAPx10_ASAP7_75t_R FILLER_181_833 ();
 DECAPx1_ASAP7_75t_R FILLER_181_855 ();
 FILLER_ASAP7_75t_R FILLER_181_877 ();
 DECAPx6_ASAP7_75t_R FILLER_181_891 ();
 DECAPx1_ASAP7_75t_R FILLER_181_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_923 ();
 DECAPx4_ASAP7_75t_R FILLER_181_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_943 ();
 DECAPx2_ASAP7_75t_R FILLER_181_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_983 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1036 ();
 DECAPx1_ASAP7_75t_R FILLER_181_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1056 ();
 FILLER_ASAP7_75t_R FILLER_181_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1072 ();
 FILLER_ASAP7_75t_R FILLER_181_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_181_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1170 ();
 FILLER_ASAP7_75t_R FILLER_181_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1242 ();
 FILLER_ASAP7_75t_R FILLER_181_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1283 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1300 ();
 FILLER_ASAP7_75t_R FILLER_181_1316 ();
 FILLER_ASAP7_75t_R FILLER_181_1325 ();
 FILLER_ASAP7_75t_R FILLER_181_1336 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1344 ();
 FILLER_ASAP7_75t_R FILLER_181_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_182_2 ();
 DECAPx2_ASAP7_75t_R FILLER_182_24 ();
 FILLER_ASAP7_75t_R FILLER_182_30 ();
 DECAPx1_ASAP7_75t_R FILLER_182_38 ();
 DECAPx2_ASAP7_75t_R FILLER_182_45 ();
 DECAPx10_ASAP7_75t_R FILLER_182_59 ();
 DECAPx2_ASAP7_75t_R FILLER_182_87 ();
 DECAPx2_ASAP7_75t_R FILLER_182_96 ();
 FILLER_ASAP7_75t_R FILLER_182_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_104 ();
 DECAPx10_ASAP7_75t_R FILLER_182_117 ();
 DECAPx6_ASAP7_75t_R FILLER_182_139 ();
 FILLER_ASAP7_75t_R FILLER_182_153 ();
 DECAPx2_ASAP7_75t_R FILLER_182_171 ();
 FILLER_ASAP7_75t_R FILLER_182_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_197 ();
 FILLER_ASAP7_75t_R FILLER_182_204 ();
 FILLER_ASAP7_75t_R FILLER_182_214 ();
 FILLER_ASAP7_75t_R FILLER_182_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_226 ();
 DECAPx10_ASAP7_75t_R FILLER_182_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_282 ();
 DECAPx1_ASAP7_75t_R FILLER_182_290 ();
 DECAPx6_ASAP7_75t_R FILLER_182_328 ();
 DECAPx1_ASAP7_75t_R FILLER_182_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_346 ();
 DECAPx2_ASAP7_75t_R FILLER_182_359 ();
 FILLER_ASAP7_75t_R FILLER_182_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_367 ();
 FILLER_ASAP7_75t_R FILLER_182_386 ();
 DECAPx2_ASAP7_75t_R FILLER_182_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_426 ();
 DECAPx1_ASAP7_75t_R FILLER_182_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_443 ();
 FILLER_ASAP7_75t_R FILLER_182_464 ();
 DECAPx2_ASAP7_75t_R FILLER_182_484 ();
 FILLER_ASAP7_75t_R FILLER_182_530 ();
 DECAPx1_ASAP7_75t_R FILLER_182_544 ();
 FILLER_ASAP7_75t_R FILLER_182_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_662 ();
 DECAPx2_ASAP7_75t_R FILLER_182_681 ();
 FILLER_ASAP7_75t_R FILLER_182_687 ();
 DECAPx6_ASAP7_75t_R FILLER_182_707 ();
 DECAPx2_ASAP7_75t_R FILLER_182_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_727 ();
 DECAPx10_ASAP7_75t_R FILLER_182_734 ();
 DECAPx10_ASAP7_75t_R FILLER_182_762 ();
 DECAPx4_ASAP7_75t_R FILLER_182_784 ();
 FILLER_ASAP7_75t_R FILLER_182_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_796 ();
 FILLER_ASAP7_75t_R FILLER_182_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_811 ();
 DECAPx4_ASAP7_75t_R FILLER_182_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_838 ();
 DECAPx6_ASAP7_75t_R FILLER_182_851 ();
 DECAPx1_ASAP7_75t_R FILLER_182_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_869 ();
 DECAPx1_ASAP7_75t_R FILLER_182_875 ();
 DECAPx4_ASAP7_75t_R FILLER_182_893 ();
 FILLER_ASAP7_75t_R FILLER_182_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_905 ();
 DECAPx2_ASAP7_75t_R FILLER_182_924 ();
 FILLER_ASAP7_75t_R FILLER_182_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_942 ();
 DECAPx4_ASAP7_75t_R FILLER_182_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_182_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1018 ();
 DECAPx4_ASAP7_75t_R FILLER_182_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1060 ();
 FILLER_ASAP7_75t_R FILLER_182_1066 ();
 DECAPx6_ASAP7_75t_R FILLER_182_1074 ();
 FILLER_ASAP7_75t_R FILLER_182_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1090 ();
 FILLER_ASAP7_75t_R FILLER_182_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_182_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1203 ();
 FILLER_ASAP7_75t_R FILLER_182_1225 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1253 ();
 DECAPx4_ASAP7_75t_R FILLER_182_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1270 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1277 ();
 DECAPx6_ASAP7_75t_R FILLER_182_1290 ();
 DECAPx6_ASAP7_75t_R FILLER_182_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1324 ();
 FILLER_ASAP7_75t_R FILLER_182_1354 ();
 DECAPx6_ASAP7_75t_R FILLER_182_1362 ();
 FILLER_ASAP7_75t_R FILLER_182_1376 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1378 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_183_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_12 ();
 FILLER_ASAP7_75t_R FILLER_183_33 ();
 DECAPx1_ASAP7_75t_R FILLER_183_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_65 ();
 FILLER_ASAP7_75t_R FILLER_183_78 ();
 DECAPx1_ASAP7_75t_R FILLER_183_83 ();
 DECAPx1_ASAP7_75t_R FILLER_183_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_152 ();
 DECAPx6_ASAP7_75t_R FILLER_183_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_212 ();
 DECAPx10_ASAP7_75t_R FILLER_183_225 ();
 DECAPx2_ASAP7_75t_R FILLER_183_247 ();
 FILLER_ASAP7_75t_R FILLER_183_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_255 ();
 FILLER_ASAP7_75t_R FILLER_183_274 ();
 FILLER_ASAP7_75t_R FILLER_183_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_284 ();
 DECAPx2_ASAP7_75t_R FILLER_183_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_301 ();
 DECAPx10_ASAP7_75t_R FILLER_183_320 ();
 DECAPx2_ASAP7_75t_R FILLER_183_342 ();
 FILLER_ASAP7_75t_R FILLER_183_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_350 ();
 DECAPx10_ASAP7_75t_R FILLER_183_361 ();
 FILLER_ASAP7_75t_R FILLER_183_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_385 ();
 FILLER_ASAP7_75t_R FILLER_183_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_401 ();
 DECAPx4_ASAP7_75t_R FILLER_183_414 ();
 DECAPx6_ASAP7_75t_R FILLER_183_444 ();
 DECAPx2_ASAP7_75t_R FILLER_183_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_464 ();
 DECAPx2_ASAP7_75t_R FILLER_183_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_477 ();
 FILLER_ASAP7_75t_R FILLER_183_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_487 ();
 DECAPx2_ASAP7_75t_R FILLER_183_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_508 ();
 DECAPx4_ASAP7_75t_R FILLER_183_512 ();
 FILLER_ASAP7_75t_R FILLER_183_522 ();
 DECAPx1_ASAP7_75t_R FILLER_183_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_565 ();
 DECAPx1_ASAP7_75t_R FILLER_183_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_582 ();
 DECAPx4_ASAP7_75t_R FILLER_183_618 ();
 FILLER_ASAP7_75t_R FILLER_183_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_630 ();
 DECAPx4_ASAP7_75t_R FILLER_183_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_667 ();
 FILLER_ASAP7_75t_R FILLER_183_679 ();
 FILLER_ASAP7_75t_R FILLER_183_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_689 ();
 FILLER_ASAP7_75t_R FILLER_183_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_703 ();
 DECAPx2_ASAP7_75t_R FILLER_183_710 ();
 FILLER_ASAP7_75t_R FILLER_183_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_725 ();
 FILLER_ASAP7_75t_R FILLER_183_739 ();
 DECAPx2_ASAP7_75t_R FILLER_183_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_766 ();
 DECAPx2_ASAP7_75t_R FILLER_183_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_779 ();
 FILLER_ASAP7_75t_R FILLER_183_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_796 ();
 DECAPx2_ASAP7_75t_R FILLER_183_804 ();
 FILLER_ASAP7_75t_R FILLER_183_810 ();
 DECAPx2_ASAP7_75t_R FILLER_183_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_834 ();
 DECAPx2_ASAP7_75t_R FILLER_183_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_861 ();
 DECAPx1_ASAP7_75t_R FILLER_183_868 ();
 DECAPx4_ASAP7_75t_R FILLER_183_879 ();
 DECAPx1_ASAP7_75t_R FILLER_183_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_960 ();
 DECAPx1_ASAP7_75t_R FILLER_183_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_968 ();
 DECAPx4_ASAP7_75t_R FILLER_183_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_988 ();
 DECAPx1_ASAP7_75t_R FILLER_183_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1003 ();
 FILLER_ASAP7_75t_R FILLER_183_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_183_1059 ();
 FILLER_ASAP7_75t_R FILLER_183_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_183_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_183_1137 ();
 FILLER_ASAP7_75t_R FILLER_183_1143 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1155 ();
 FILLER_ASAP7_75t_R FILLER_183_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1171 ();
 DECAPx4_ASAP7_75t_R FILLER_183_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1185 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1213 ();
 DECAPx2_ASAP7_75t_R FILLER_183_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1241 ();
 FILLER_ASAP7_75t_R FILLER_183_1245 ();
 DECAPx1_ASAP7_75t_R FILLER_183_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1268 ();
 DECAPx4_ASAP7_75t_R FILLER_183_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1318 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1329 ();
 DECAPx1_ASAP7_75t_R FILLER_183_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_183_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1361 ();
 DECAPx1_ASAP7_75t_R FILLER_183_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_184_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_16 ();
 DECAPx2_ASAP7_75t_R FILLER_184_23 ();
 FILLER_ASAP7_75t_R FILLER_184_29 ();
 DECAPx4_ASAP7_75t_R FILLER_184_37 ();
 FILLER_ASAP7_75t_R FILLER_184_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_49 ();
 DECAPx2_ASAP7_75t_R FILLER_184_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_65 ();
 DECAPx4_ASAP7_75t_R FILLER_184_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_102 ();
 DECAPx6_ASAP7_75t_R FILLER_184_106 ();
 FILLER_ASAP7_75t_R FILLER_184_120 ();
 FILLER_ASAP7_75t_R FILLER_184_132 ();
 DECAPx2_ASAP7_75t_R FILLER_184_160 ();
 DECAPx4_ASAP7_75t_R FILLER_184_172 ();
 FILLER_ASAP7_75t_R FILLER_184_182 ();
 DECAPx2_ASAP7_75t_R FILLER_184_196 ();
 FILLER_ASAP7_75t_R FILLER_184_202 ();
 DECAPx6_ASAP7_75t_R FILLER_184_218 ();
 DECAPx1_ASAP7_75t_R FILLER_184_232 ();
 DECAPx6_ASAP7_75t_R FILLER_184_254 ();
 FILLER_ASAP7_75t_R FILLER_184_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_270 ();
 DECAPx2_ASAP7_75t_R FILLER_184_274 ();
 FILLER_ASAP7_75t_R FILLER_184_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_282 ();
 DECAPx2_ASAP7_75t_R FILLER_184_315 ();
 FILLER_ASAP7_75t_R FILLER_184_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_328 ();
 DECAPx2_ASAP7_75t_R FILLER_184_347 ();
 FILLER_ASAP7_75t_R FILLER_184_353 ();
 DECAPx4_ASAP7_75t_R FILLER_184_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_373 ();
 DECAPx10_ASAP7_75t_R FILLER_184_392 ();
 DECAPx6_ASAP7_75t_R FILLER_184_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_428 ();
 DECAPx10_ASAP7_75t_R FILLER_184_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_461 ();
 DECAPx10_ASAP7_75t_R FILLER_184_464 ();
 DECAPx4_ASAP7_75t_R FILLER_184_486 ();
 DECAPx10_ASAP7_75t_R FILLER_184_502 ();
 FILLER_ASAP7_75t_R FILLER_184_524 ();
 FILLER_ASAP7_75t_R FILLER_184_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_554 ();
 DECAPx1_ASAP7_75t_R FILLER_184_567 ();
 DECAPx4_ASAP7_75t_R FILLER_184_577 ();
 DECAPx2_ASAP7_75t_R FILLER_184_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_606 ();
 DECAPx10_ASAP7_75t_R FILLER_184_614 ();
 DECAPx2_ASAP7_75t_R FILLER_184_636 ();
 FILLER_ASAP7_75t_R FILLER_184_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_644 ();
 FILLER_ASAP7_75t_R FILLER_184_648 ();
 DECAPx1_ASAP7_75t_R FILLER_184_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_697 ();
 DECAPx2_ASAP7_75t_R FILLER_184_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_720 ();
 FILLER_ASAP7_75t_R FILLER_184_737 ();
 DECAPx2_ASAP7_75t_R FILLER_184_754 ();
 FILLER_ASAP7_75t_R FILLER_184_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_781 ();
 DECAPx2_ASAP7_75t_R FILLER_184_806 ();
 FILLER_ASAP7_75t_R FILLER_184_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_814 ();
 DECAPx2_ASAP7_75t_R FILLER_184_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_860 ();
 DECAPx4_ASAP7_75t_R FILLER_184_878 ();
 FILLER_ASAP7_75t_R FILLER_184_888 ();
 DECAPx4_ASAP7_75t_R FILLER_184_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_911 ();
 DECAPx4_ASAP7_75t_R FILLER_184_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_934 ();
 FILLER_ASAP7_75t_R FILLER_184_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_947 ();
 DECAPx10_ASAP7_75t_R FILLER_184_954 ();
 DECAPx10_ASAP7_75t_R FILLER_184_976 ();
 DECAPx6_ASAP7_75t_R FILLER_184_998 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_184_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1168 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1193 ();
 DECAPx4_ASAP7_75t_R FILLER_184_1209 ();
 FILLER_ASAP7_75t_R FILLER_184_1219 ();
 FILLER_ASAP7_75t_R FILLER_184_1239 ();
 FILLER_ASAP7_75t_R FILLER_184_1251 ();
 FILLER_ASAP7_75t_R FILLER_184_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1297 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1312 ();
 FILLER_ASAP7_75t_R FILLER_184_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1369 ();
 FILLER_ASAP7_75t_R FILLER_184_1381 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_185_2 ();
 FILLER_ASAP7_75t_R FILLER_185_8 ();
 FILLER_ASAP7_75t_R FILLER_185_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_44 ();
 DECAPx2_ASAP7_75t_R FILLER_185_48 ();
 DECAPx6_ASAP7_75t_R FILLER_185_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_77 ();
 FILLER_ASAP7_75t_R FILLER_185_110 ();
 DECAPx2_ASAP7_75t_R FILLER_185_118 ();
 FILLER_ASAP7_75t_R FILLER_185_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_126 ();
 DECAPx6_ASAP7_75t_R FILLER_185_133 ();
 FILLER_ASAP7_75t_R FILLER_185_147 ();
 DECAPx4_ASAP7_75t_R FILLER_185_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_165 ();
 DECAPx2_ASAP7_75t_R FILLER_185_172 ();
 FILLER_ASAP7_75t_R FILLER_185_178 ();
 DECAPx6_ASAP7_75t_R FILLER_185_186 ();
 DECAPx1_ASAP7_75t_R FILLER_185_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_204 ();
 DECAPx2_ASAP7_75t_R FILLER_185_211 ();
 FILLER_ASAP7_75t_R FILLER_185_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_225 ();
 DECAPx1_ASAP7_75t_R FILLER_185_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_252 ();
 DECAPx2_ASAP7_75t_R FILLER_185_259 ();
 DECAPx2_ASAP7_75t_R FILLER_185_276 ();
 FILLER_ASAP7_75t_R FILLER_185_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_284 ();
 DECAPx2_ASAP7_75t_R FILLER_185_298 ();
 FILLER_ASAP7_75t_R FILLER_185_304 ();
 FILLER_ASAP7_75t_R FILLER_185_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_314 ();
 FILLER_ASAP7_75t_R FILLER_185_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_329 ();
 FILLER_ASAP7_75t_R FILLER_185_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_360 ();
 DECAPx6_ASAP7_75t_R FILLER_185_367 ();
 FILLER_ASAP7_75t_R FILLER_185_381 ();
 DECAPx1_ASAP7_75t_R FILLER_185_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_405 ();
 DECAPx1_ASAP7_75t_R FILLER_185_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_425 ();
 DECAPx6_ASAP7_75t_R FILLER_185_429 ();
 FILLER_ASAP7_75t_R FILLER_185_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_457 ();
 DECAPx2_ASAP7_75t_R FILLER_185_476 ();
 DECAPx2_ASAP7_75t_R FILLER_185_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_506 ();
 FILLER_ASAP7_75t_R FILLER_185_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_527 ();
 DECAPx2_ASAP7_75t_R FILLER_185_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_543 ();
 DECAPx10_ASAP7_75t_R FILLER_185_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_569 ();
 DECAPx10_ASAP7_75t_R FILLER_185_578 ();
 DECAPx2_ASAP7_75t_R FILLER_185_600 ();
 FILLER_ASAP7_75t_R FILLER_185_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_608 ();
 DECAPx10_ASAP7_75t_R FILLER_185_635 ();
 DECAPx2_ASAP7_75t_R FILLER_185_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_663 ();
 DECAPx6_ASAP7_75t_R FILLER_185_685 ();
 DECAPx10_ASAP7_75t_R FILLER_185_706 ();
 DECAPx4_ASAP7_75t_R FILLER_185_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_748 ();
 DECAPx6_ASAP7_75t_R FILLER_185_755 ();
 FILLER_ASAP7_75t_R FILLER_185_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_771 ();
 DECAPx1_ASAP7_75t_R FILLER_185_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_784 ();
 DECAPx6_ASAP7_75t_R FILLER_185_797 ();
 DECAPx2_ASAP7_75t_R FILLER_185_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_833 ();
 DECAPx1_ASAP7_75t_R FILLER_185_846 ();
 FILLER_ASAP7_75t_R FILLER_185_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_859 ();
 DECAPx2_ASAP7_75t_R FILLER_185_875 ();
 FILLER_ASAP7_75t_R FILLER_185_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_883 ();
 DECAPx10_ASAP7_75t_R FILLER_185_890 ();
 FILLER_ASAP7_75t_R FILLER_185_912 ();
 DECAPx1_ASAP7_75t_R FILLER_185_920 ();
 DECAPx4_ASAP7_75t_R FILLER_185_926 ();
 FILLER_ASAP7_75t_R FILLER_185_936 ();
 DECAPx6_ASAP7_75t_R FILLER_185_944 ();
 DECAPx10_ASAP7_75t_R FILLER_185_974 ();
 DECAPx2_ASAP7_75t_R FILLER_185_996 ();
 FILLER_ASAP7_75t_R FILLER_185_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1025 ();
 DECAPx4_ASAP7_75t_R FILLER_185_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1055 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1079 ();
 DECAPx6_ASAP7_75t_R FILLER_185_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1113 ();
 FILLER_ASAP7_75t_R FILLER_185_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1121 ();
 FILLER_ASAP7_75t_R FILLER_185_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1215 ();
 FILLER_ASAP7_75t_R FILLER_185_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1229 ();
 DECAPx4_ASAP7_75t_R FILLER_185_1262 ();
 FILLER_ASAP7_75t_R FILLER_185_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1277 ();
 FILLER_ASAP7_75t_R FILLER_185_1283 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1311 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1323 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1330 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1352 ();
 FILLER_ASAP7_75t_R FILLER_185_1358 ();
 DECAPx4_ASAP7_75t_R FILLER_186_2 ();
 FILLER_ASAP7_75t_R FILLER_186_12 ();
 DECAPx1_ASAP7_75t_R FILLER_186_20 ();
 DECAPx1_ASAP7_75t_R FILLER_186_27 ();
 DECAPx1_ASAP7_75t_R FILLER_186_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_80 ();
 DECAPx1_ASAP7_75t_R FILLER_186_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_88 ();
 FILLER_ASAP7_75t_R FILLER_186_121 ();
 DECAPx2_ASAP7_75t_R FILLER_186_129 ();
 FILLER_ASAP7_75t_R FILLER_186_135 ();
 DECAPx1_ASAP7_75t_R FILLER_186_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_147 ();
 DECAPx1_ASAP7_75t_R FILLER_186_154 ();
 DECAPx2_ASAP7_75t_R FILLER_186_172 ();
 FILLER_ASAP7_75t_R FILLER_186_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_180 ();
 FILLER_ASAP7_75t_R FILLER_186_189 ();
 DECAPx1_ASAP7_75t_R FILLER_186_197 ();
 DECAPx4_ASAP7_75t_R FILLER_186_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_281 ();
 DECAPx4_ASAP7_75t_R FILLER_186_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_329 ();
 DECAPx1_ASAP7_75t_R FILLER_186_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_352 ();
 DECAPx6_ASAP7_75t_R FILLER_186_369 ();
 FILLER_ASAP7_75t_R FILLER_186_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_391 ();
 DECAPx2_ASAP7_75t_R FILLER_186_438 ();
 FILLER_ASAP7_75t_R FILLER_186_464 ();
 DECAPx2_ASAP7_75t_R FILLER_186_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_490 ();
 DECAPx6_ASAP7_75t_R FILLER_186_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_542 ();
 FILLER_ASAP7_75t_R FILLER_186_561 ();
 DECAPx2_ASAP7_75t_R FILLER_186_586 ();
 DECAPx2_ASAP7_75t_R FILLER_186_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_622 ();
 DECAPx1_ASAP7_75t_R FILLER_186_626 ();
 DECAPx6_ASAP7_75t_R FILLER_186_652 ();
 DECAPx1_ASAP7_75t_R FILLER_186_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_670 ();
 DECAPx4_ASAP7_75t_R FILLER_186_683 ();
 FILLER_ASAP7_75t_R FILLER_186_693 ();
 DECAPx10_ASAP7_75t_R FILLER_186_704 ();
 DECAPx2_ASAP7_75t_R FILLER_186_726 ();
 FILLER_ASAP7_75t_R FILLER_186_732 ();
 DECAPx4_ASAP7_75t_R FILLER_186_769 ();
 FILLER_ASAP7_75t_R FILLER_186_779 ();
 DECAPx10_ASAP7_75t_R FILLER_186_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_811 ();
 DECAPx1_ASAP7_75t_R FILLER_186_828 ();
 DECAPx2_ASAP7_75t_R FILLER_186_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_850 ();
 FILLER_ASAP7_75t_R FILLER_186_857 ();
 DECAPx2_ASAP7_75t_R FILLER_186_868 ();
 FILLER_ASAP7_75t_R FILLER_186_874 ();
 DECAPx4_ASAP7_75t_R FILLER_186_904 ();
 FILLER_ASAP7_75t_R FILLER_186_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_938 ();
 DECAPx1_ASAP7_75t_R FILLER_186_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_963 ();
 DECAPx4_ASAP7_75t_R FILLER_186_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1051 ();
 FILLER_ASAP7_75t_R FILLER_186_1091 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1101 ();
 FILLER_ASAP7_75t_R FILLER_186_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1117 ();
 FILLER_ASAP7_75t_R FILLER_186_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1194 ();
 FILLER_ASAP7_75t_R FILLER_186_1201 ();
 FILLER_ASAP7_75t_R FILLER_186_1216 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1250 ();
 FILLER_ASAP7_75t_R FILLER_186_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1256 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1263 ();
 FILLER_ASAP7_75t_R FILLER_186_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1278 ();
 DECAPx1_ASAP7_75t_R FILLER_186_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1307 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1316 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1330 ();
 FILLER_ASAP7_75t_R FILLER_186_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_186_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_187_2 ();
 DECAPx4_ASAP7_75t_R FILLER_187_24 ();
 DECAPx6_ASAP7_75t_R FILLER_187_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_52 ();
 DECAPx6_ASAP7_75t_R FILLER_187_79 ();
 DECAPx1_ASAP7_75t_R FILLER_187_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_100 ();
 DECAPx1_ASAP7_75t_R FILLER_187_111 ();
 FILLER_ASAP7_75t_R FILLER_187_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_121 ();
 FILLER_ASAP7_75t_R FILLER_187_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_178 ();
 FILLER_ASAP7_75t_R FILLER_187_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_189 ();
 DECAPx6_ASAP7_75t_R FILLER_187_196 ();
 DECAPx1_ASAP7_75t_R FILLER_187_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_214 ();
 FILLER_ASAP7_75t_R FILLER_187_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_241 ();
 DECAPx1_ASAP7_75t_R FILLER_187_256 ();
 FILLER_ASAP7_75t_R FILLER_187_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_282 ();
 DECAPx6_ASAP7_75t_R FILLER_187_291 ();
 DECAPx1_ASAP7_75t_R FILLER_187_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_309 ();
 FILLER_ASAP7_75t_R FILLER_187_319 ();
 DECAPx6_ASAP7_75t_R FILLER_187_327 ();
 DECAPx1_ASAP7_75t_R FILLER_187_341 ();
 FILLER_ASAP7_75t_R FILLER_187_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_360 ();
 DECAPx4_ASAP7_75t_R FILLER_187_375 ();
 DECAPx1_ASAP7_75t_R FILLER_187_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_397 ();
 FILLER_ASAP7_75t_R FILLER_187_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_408 ();
 DECAPx6_ASAP7_75t_R FILLER_187_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_435 ();
 DECAPx10_ASAP7_75t_R FILLER_187_454 ();
 DECAPx2_ASAP7_75t_R FILLER_187_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_482 ();
 DECAPx2_ASAP7_75t_R FILLER_187_501 ();
 FILLER_ASAP7_75t_R FILLER_187_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_527 ();
 DECAPx4_ASAP7_75t_R FILLER_187_535 ();
 FILLER_ASAP7_75t_R FILLER_187_545 ();
 FILLER_ASAP7_75t_R FILLER_187_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_573 ();
 DECAPx1_ASAP7_75t_R FILLER_187_618 ();
 FILLER_ASAP7_75t_R FILLER_187_644 ();
 DECAPx1_ASAP7_75t_R FILLER_187_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_668 ();
 FILLER_ASAP7_75t_R FILLER_187_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_692 ();
 DECAPx1_ASAP7_75t_R FILLER_187_728 ();
 DECAPx6_ASAP7_75t_R FILLER_187_738 ();
 FILLER_ASAP7_75t_R FILLER_187_752 ();
 DECAPx6_ASAP7_75t_R FILLER_187_767 ();
 FILLER_ASAP7_75t_R FILLER_187_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_801 ();
 DECAPx10_ASAP7_75t_R FILLER_187_812 ();
 DECAPx10_ASAP7_75t_R FILLER_187_834 ();
 DECAPx1_ASAP7_75t_R FILLER_187_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_860 ();
 DECAPx6_ASAP7_75t_R FILLER_187_874 ();
 DECAPx2_ASAP7_75t_R FILLER_187_888 ();
 FILLER_ASAP7_75t_R FILLER_187_912 ();
 DECAPx4_ASAP7_75t_R FILLER_187_926 ();
 DECAPx10_ASAP7_75t_R FILLER_187_950 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1030 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1037 ();
 FILLER_ASAP7_75t_R FILLER_187_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1051 ();
 FILLER_ASAP7_75t_R FILLER_187_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1083 ();
 FILLER_ASAP7_75t_R FILLER_187_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1091 ();
 FILLER_ASAP7_75t_R FILLER_187_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1111 ();
 DECAPx6_ASAP7_75t_R FILLER_187_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_187_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1224 ();
 FILLER_ASAP7_75t_R FILLER_187_1230 ();
 DECAPx6_ASAP7_75t_R FILLER_187_1235 ();
 FILLER_ASAP7_75t_R FILLER_187_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1251 ();
 FILLER_ASAP7_75t_R FILLER_187_1262 ();
 DECAPx6_ASAP7_75t_R FILLER_187_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1297 ();
 FILLER_ASAP7_75t_R FILLER_187_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1352 ();
 FILLER_ASAP7_75t_R FILLER_187_1364 ();
 DECAPx6_ASAP7_75t_R FILLER_188_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_16 ();
 DECAPx2_ASAP7_75t_R FILLER_188_27 ();
 DECAPx4_ASAP7_75t_R FILLER_188_49 ();
 FILLER_ASAP7_75t_R FILLER_188_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_61 ();
 DECAPx2_ASAP7_75t_R FILLER_188_72 ();
 FILLER_ASAP7_75t_R FILLER_188_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_80 ();
 DECAPx4_ASAP7_75t_R FILLER_188_91 ();
 FILLER_ASAP7_75t_R FILLER_188_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_103 ();
 DECAPx6_ASAP7_75t_R FILLER_188_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_121 ();
 DECAPx4_ASAP7_75t_R FILLER_188_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_169 ();
 DECAPx1_ASAP7_75t_R FILLER_188_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_188 ();
 FILLER_ASAP7_75t_R FILLER_188_195 ();
 DECAPx1_ASAP7_75t_R FILLER_188_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_225 ();
 DECAPx10_ASAP7_75t_R FILLER_188_234 ();
 FILLER_ASAP7_75t_R FILLER_188_256 ();
 DECAPx4_ASAP7_75t_R FILLER_188_267 ();
 FILLER_ASAP7_75t_R FILLER_188_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_279 ();
 DECAPx2_ASAP7_75t_R FILLER_188_300 ();
 DECAPx10_ASAP7_75t_R FILLER_188_312 ();
 DECAPx4_ASAP7_75t_R FILLER_188_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_362 ();
 FILLER_ASAP7_75t_R FILLER_188_369 ();
 FILLER_ASAP7_75t_R FILLER_188_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_380 ();
 DECAPx1_ASAP7_75t_R FILLER_188_399 ();
 DECAPx10_ASAP7_75t_R FILLER_188_412 ();
 FILLER_ASAP7_75t_R FILLER_188_434 ();
 DECAPx2_ASAP7_75t_R FILLER_188_454 ();
 FILLER_ASAP7_75t_R FILLER_188_460 ();
 DECAPx4_ASAP7_75t_R FILLER_188_464 ();
 FILLER_ASAP7_75t_R FILLER_188_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_507 ();
 DECAPx10_ASAP7_75t_R FILLER_188_534 ();
 FILLER_ASAP7_75t_R FILLER_188_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_558 ();
 DECAPx10_ASAP7_75t_R FILLER_188_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_593 ();
 DECAPx2_ASAP7_75t_R FILLER_188_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_610 ();
 FILLER_ASAP7_75t_R FILLER_188_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_626 ();
 DECAPx10_ASAP7_75t_R FILLER_188_630 ();
 DECAPx2_ASAP7_75t_R FILLER_188_652 ();
 FILLER_ASAP7_75t_R FILLER_188_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_692 ();
 DECAPx1_ASAP7_75t_R FILLER_188_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_705 ();
 DECAPx2_ASAP7_75t_R FILLER_188_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_715 ();
 FILLER_ASAP7_75t_R FILLER_188_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_721 ();
 DECAPx6_ASAP7_75t_R FILLER_188_743 ();
 FILLER_ASAP7_75t_R FILLER_188_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_759 ();
 DECAPx4_ASAP7_75t_R FILLER_188_770 ();
 FILLER_ASAP7_75t_R FILLER_188_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_794 ();
 FILLER_ASAP7_75t_R FILLER_188_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_805 ();
 DECAPx4_ASAP7_75t_R FILLER_188_816 ();
 DECAPx4_ASAP7_75t_R FILLER_188_845 ();
 FILLER_ASAP7_75t_R FILLER_188_855 ();
 FILLER_ASAP7_75t_R FILLER_188_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_865 ();
 FILLER_ASAP7_75t_R FILLER_188_875 ();
 DECAPx4_ASAP7_75t_R FILLER_188_883 ();
 FILLER_ASAP7_75t_R FILLER_188_893 ();
 DECAPx1_ASAP7_75t_R FILLER_188_913 ();
 DECAPx2_ASAP7_75t_R FILLER_188_929 ();
 FILLER_ASAP7_75t_R FILLER_188_935 ();
 DECAPx2_ASAP7_75t_R FILLER_188_943 ();
 FILLER_ASAP7_75t_R FILLER_188_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_951 ();
 DECAPx2_ASAP7_75t_R FILLER_188_970 ();
 FILLER_ASAP7_75t_R FILLER_188_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_978 ();
 DECAPx1_ASAP7_75t_R FILLER_188_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_990 ();
 FILLER_ASAP7_75t_R FILLER_188_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1011 ();
 DECAPx4_ASAP7_75t_R FILLER_188_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1066 ();
 FILLER_ASAP7_75t_R FILLER_188_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1096 ();
 FILLER_ASAP7_75t_R FILLER_188_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1112 ();
 FILLER_ASAP7_75t_R FILLER_188_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1133 ();
 FILLER_ASAP7_75t_R FILLER_188_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_188_1147 ();
 FILLER_ASAP7_75t_R FILLER_188_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1226 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1262 ();
 FILLER_ASAP7_75t_R FILLER_188_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1299 ();
 FILLER_ASAP7_75t_R FILLER_188_1305 ();
 FILLER_ASAP7_75t_R FILLER_188_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1315 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1329 ();
 FILLER_ASAP7_75t_R FILLER_188_1343 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_189_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_16 ();
 DECAPx2_ASAP7_75t_R FILLER_189_23 ();
 DECAPx6_ASAP7_75t_R FILLER_189_59 ();
 DECAPx1_ASAP7_75t_R FILLER_189_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_77 ();
 DECAPx1_ASAP7_75t_R FILLER_189_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_85 ();
 DECAPx4_ASAP7_75t_R FILLER_189_92 ();
 DECAPx4_ASAP7_75t_R FILLER_189_112 ();
 DECAPx4_ASAP7_75t_R FILLER_189_125 ();
 FILLER_ASAP7_75t_R FILLER_189_135 ();
 DECAPx4_ASAP7_75t_R FILLER_189_140 ();
 FILLER_ASAP7_75t_R FILLER_189_150 ();
 DECAPx6_ASAP7_75t_R FILLER_189_159 ();
 DECAPx2_ASAP7_75t_R FILLER_189_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_179 ();
 DECAPx1_ASAP7_75t_R FILLER_189_186 ();
 DECAPx10_ASAP7_75t_R FILLER_189_196 ();
 DECAPx1_ASAP7_75t_R FILLER_189_218 ();
 FILLER_ASAP7_75t_R FILLER_189_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_238 ();
 DECAPx10_ASAP7_75t_R FILLER_189_245 ();
 DECAPx6_ASAP7_75t_R FILLER_189_267 ();
 FILLER_ASAP7_75t_R FILLER_189_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_283 ();
 DECAPx6_ASAP7_75t_R FILLER_189_292 ();
 FILLER_ASAP7_75t_R FILLER_189_306 ();
 DECAPx6_ASAP7_75t_R FILLER_189_316 ();
 DECAPx1_ASAP7_75t_R FILLER_189_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_346 ();
 DECAPx4_ASAP7_75t_R FILLER_189_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_369 ();
 DECAPx2_ASAP7_75t_R FILLER_189_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_383 ();
 FILLER_ASAP7_75t_R FILLER_189_417 ();
 DECAPx10_ASAP7_75t_R FILLER_189_427 ();
 DECAPx4_ASAP7_75t_R FILLER_189_449 ();
 FILLER_ASAP7_75t_R FILLER_189_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_461 ();
 DECAPx2_ASAP7_75t_R FILLER_189_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_486 ();
 DECAPx6_ASAP7_75t_R FILLER_189_503 ();
 DECAPx1_ASAP7_75t_R FILLER_189_517 ();
 DECAPx2_ASAP7_75t_R FILLER_189_531 ();
 DECAPx1_ASAP7_75t_R FILLER_189_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_559 ();
 FILLER_ASAP7_75t_R FILLER_189_570 ();
 DECAPx1_ASAP7_75t_R FILLER_189_590 ();
 DECAPx4_ASAP7_75t_R FILLER_189_600 ();
 FILLER_ASAP7_75t_R FILLER_189_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_612 ();
 DECAPx10_ASAP7_75t_R FILLER_189_639 ();
 DECAPx10_ASAP7_75t_R FILLER_189_661 ();
 DECAPx2_ASAP7_75t_R FILLER_189_683 ();
 FILLER_ASAP7_75t_R FILLER_189_689 ();
 DECAPx4_ASAP7_75t_R FILLER_189_717 ();
 FILLER_ASAP7_75t_R FILLER_189_727 ();
 DECAPx6_ASAP7_75t_R FILLER_189_741 ();
 FILLER_ASAP7_75t_R FILLER_189_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_767 ();
 DECAPx1_ASAP7_75t_R FILLER_189_778 ();
 DECAPx1_ASAP7_75t_R FILLER_189_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_810 ();
 FILLER_ASAP7_75t_R FILLER_189_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_837 ();
 DECAPx1_ASAP7_75t_R FILLER_189_852 ();
 FILLER_ASAP7_75t_R FILLER_189_876 ();
 DECAPx10_ASAP7_75t_R FILLER_189_893 ();
 DECAPx2_ASAP7_75t_R FILLER_189_915 ();
 FILLER_ASAP7_75t_R FILLER_189_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_923 ();
 DECAPx2_ASAP7_75t_R FILLER_189_926 ();
 FILLER_ASAP7_75t_R FILLER_189_932 ();
 DECAPx2_ASAP7_75t_R FILLER_189_944 ();
 FILLER_ASAP7_75t_R FILLER_189_950 ();
 DECAPx10_ASAP7_75t_R FILLER_189_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_997 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1004 ();
 FILLER_ASAP7_75t_R FILLER_189_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1082 ();
 FILLER_ASAP7_75t_R FILLER_189_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1111 ();
 FILLER_ASAP7_75t_R FILLER_189_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1146 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1186 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1213 ();
 FILLER_ASAP7_75t_R FILLER_189_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1221 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1261 ();
 FILLER_ASAP7_75t_R FILLER_189_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1310 ();
 FILLER_ASAP7_75t_R FILLER_189_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1329 ();
 DECAPx4_ASAP7_75t_R FILLER_189_1373 ();
 DECAPx1_ASAP7_75t_R FILLER_190_2 ();
 FILLER_ASAP7_75t_R FILLER_190_38 ();
 FILLER_ASAP7_75t_R FILLER_190_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_130 ();
 FILLER_ASAP7_75t_R FILLER_190_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_163 ();
 DECAPx4_ASAP7_75t_R FILLER_190_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_188 ();
 DECAPx1_ASAP7_75t_R FILLER_190_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_201 ();
 DECAPx1_ASAP7_75t_R FILLER_190_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_230 ();
 FILLER_ASAP7_75t_R FILLER_190_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_241 ();
 DECAPx2_ASAP7_75t_R FILLER_190_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_265 ();
 DECAPx2_ASAP7_75t_R FILLER_190_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_282 ();
 DECAPx1_ASAP7_75t_R FILLER_190_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_327 ();
 DECAPx1_ASAP7_75t_R FILLER_190_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_350 ();
 DECAPx10_ASAP7_75t_R FILLER_190_368 ();
 DECAPx1_ASAP7_75t_R FILLER_190_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_410 ();
 DECAPx2_ASAP7_75t_R FILLER_190_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_437 ();
 DECAPx2_ASAP7_75t_R FILLER_190_456 ();
 DECAPx2_ASAP7_75t_R FILLER_190_464 ();
 DECAPx10_ASAP7_75t_R FILLER_190_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_510 ();
 DECAPx4_ASAP7_75t_R FILLER_190_525 ();
 FILLER_ASAP7_75t_R FILLER_190_535 ();
 DECAPx2_ASAP7_75t_R FILLER_190_573 ();
 FILLER_ASAP7_75t_R FILLER_190_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_581 ();
 DECAPx1_ASAP7_75t_R FILLER_190_600 ();
 DECAPx6_ASAP7_75t_R FILLER_190_610 ();
 DECAPx1_ASAP7_75t_R FILLER_190_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_628 ();
 DECAPx2_ASAP7_75t_R FILLER_190_636 ();
 FILLER_ASAP7_75t_R FILLER_190_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_644 ();
 DECAPx2_ASAP7_75t_R FILLER_190_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_654 ();
 DECAPx6_ASAP7_75t_R FILLER_190_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_687 ();
 DECAPx6_ASAP7_75t_R FILLER_190_700 ();
 FILLER_ASAP7_75t_R FILLER_190_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_724 ();
 DECAPx2_ASAP7_75t_R FILLER_190_728 ();
 DECAPx6_ASAP7_75t_R FILLER_190_741 ();
 DECAPx1_ASAP7_75t_R FILLER_190_755 ();
 DECAPx4_ASAP7_75t_R FILLER_190_769 ();
 DECAPx4_ASAP7_75t_R FILLER_190_785 ();
 FILLER_ASAP7_75t_R FILLER_190_795 ();
 FILLER_ASAP7_75t_R FILLER_190_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_809 ();
 DECAPx6_ASAP7_75t_R FILLER_190_822 ();
 DECAPx2_ASAP7_75t_R FILLER_190_836 ();
 DECAPx6_ASAP7_75t_R FILLER_190_860 ();
 DECAPx2_ASAP7_75t_R FILLER_190_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_880 ();
 DECAPx10_ASAP7_75t_R FILLER_190_899 ();
 DECAPx2_ASAP7_75t_R FILLER_190_930 ();
 DECAPx4_ASAP7_75t_R FILLER_190_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_959 ();
 DECAPx6_ASAP7_75t_R FILLER_190_972 ();
 DECAPx2_ASAP7_75t_R FILLER_190_986 ();
 FILLER_ASAP7_75t_R FILLER_190_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1020 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1064 ();
 DECAPx4_ASAP7_75t_R FILLER_190_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1097 ();
 FILLER_ASAP7_75t_R FILLER_190_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1105 ();
 FILLER_ASAP7_75t_R FILLER_190_1116 ();
 DECAPx4_ASAP7_75t_R FILLER_190_1124 ();
 FILLER_ASAP7_75t_R FILLER_190_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1136 ();
 DECAPx4_ASAP7_75t_R FILLER_190_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1192 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1228 ();
 DECAPx4_ASAP7_75t_R FILLER_190_1273 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1283 ();
 FILLER_ASAP7_75t_R FILLER_190_1287 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1315 ();
 FILLER_ASAP7_75t_R FILLER_190_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1349 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_191_2 ();
 FILLER_ASAP7_75t_R FILLER_191_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_20 ();
 DECAPx4_ASAP7_75t_R FILLER_191_35 ();
 FILLER_ASAP7_75t_R FILLER_191_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_47 ();
 DECAPx4_ASAP7_75t_R FILLER_191_54 ();
 FILLER_ASAP7_75t_R FILLER_191_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_80 ();
 FILLER_ASAP7_75t_R FILLER_191_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_89 ();
 DECAPx1_ASAP7_75t_R FILLER_191_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_97 ();
 FILLER_ASAP7_75t_R FILLER_191_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_126 ();
 DECAPx1_ASAP7_75t_R FILLER_191_139 ();
 FILLER_ASAP7_75t_R FILLER_191_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_186 ();
 DECAPx2_ASAP7_75t_R FILLER_191_193 ();
 FILLER_ASAP7_75t_R FILLER_191_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_201 ();
 DECAPx1_ASAP7_75t_R FILLER_191_230 ();
 DECAPx4_ASAP7_75t_R FILLER_191_248 ();
 FILLER_ASAP7_75t_R FILLER_191_258 ();
 DECAPx1_ASAP7_75t_R FILLER_191_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_282 ();
 DECAPx10_ASAP7_75t_R FILLER_191_309 ();
 DECAPx4_ASAP7_75t_R FILLER_191_331 ();
 DECAPx1_ASAP7_75t_R FILLER_191_355 ();
 FILLER_ASAP7_75t_R FILLER_191_377 ();
 DECAPx1_ASAP7_75t_R FILLER_191_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_401 ();
 DECAPx6_ASAP7_75t_R FILLER_191_408 ();
 FILLER_ASAP7_75t_R FILLER_191_422 ();
 DECAPx2_ASAP7_75t_R FILLER_191_434 ();
 FILLER_ASAP7_75t_R FILLER_191_440 ();
 DECAPx1_ASAP7_75t_R FILLER_191_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_525 ();
 FILLER_ASAP7_75t_R FILLER_191_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_546 ();
 DECAPx4_ASAP7_75t_R FILLER_191_565 ();
 FILLER_ASAP7_75t_R FILLER_191_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_585 ();
 DECAPx1_ASAP7_75t_R FILLER_191_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_629 ();
 DECAPx2_ASAP7_75t_R FILLER_191_656 ();
 FILLER_ASAP7_75t_R FILLER_191_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_664 ();
 DECAPx4_ASAP7_75t_R FILLER_191_683 ();
 DECAPx4_ASAP7_75t_R FILLER_191_700 ();
 FILLER_ASAP7_75t_R FILLER_191_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_738 ();
 FILLER_ASAP7_75t_R FILLER_191_745 ();
 DECAPx6_ASAP7_75t_R FILLER_191_757 ();
 FILLER_ASAP7_75t_R FILLER_191_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_773 ();
 DECAPx10_ASAP7_75t_R FILLER_191_800 ();
 DECAPx10_ASAP7_75t_R FILLER_191_822 ();
 DECAPx6_ASAP7_75t_R FILLER_191_844 ();
 FILLER_ASAP7_75t_R FILLER_191_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_860 ();
 DECAPx2_ASAP7_75t_R FILLER_191_871 ();
 FILLER_ASAP7_75t_R FILLER_191_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_879 ();
 FILLER_ASAP7_75t_R FILLER_191_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_908 ();
 DECAPx2_ASAP7_75t_R FILLER_191_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_941 ();
 DECAPx4_ASAP7_75t_R FILLER_191_951 ();
 FILLER_ASAP7_75t_R FILLER_191_961 ();
 DECAPx2_ASAP7_75t_R FILLER_191_989 ();
 FILLER_ASAP7_75t_R FILLER_191_995 ();
 FILLER_ASAP7_75t_R FILLER_191_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1066 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1162 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1207 ();
 FILLER_ASAP7_75t_R FILLER_191_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1219 ();
 FILLER_ASAP7_75t_R FILLER_191_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_191_1265 ();
 FILLER_ASAP7_75t_R FILLER_191_1275 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1285 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1299 ();
 FILLER_ASAP7_75t_R FILLER_191_1306 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1308 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1331 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1340 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1391 ();
 DECAPx6_ASAP7_75t_R FILLER_192_2 ();
 DECAPx1_ASAP7_75t_R FILLER_192_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_20 ();
 DECAPx6_ASAP7_75t_R FILLER_192_24 ();
 FILLER_ASAP7_75t_R FILLER_192_38 ();
 DECAPx6_ASAP7_75t_R FILLER_192_46 ();
 DECAPx1_ASAP7_75t_R FILLER_192_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_64 ();
 DECAPx4_ASAP7_75t_R FILLER_192_71 ();
 FILLER_ASAP7_75t_R FILLER_192_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_101 ();
 DECAPx1_ASAP7_75t_R FILLER_192_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_112 ();
 DECAPx6_ASAP7_75t_R FILLER_192_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_130 ();
 DECAPx4_ASAP7_75t_R FILLER_192_149 ();
 FILLER_ASAP7_75t_R FILLER_192_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_165 ();
 DECAPx10_ASAP7_75t_R FILLER_192_172 ();
 DECAPx10_ASAP7_75t_R FILLER_192_194 ();
 DECAPx2_ASAP7_75t_R FILLER_192_216 ();
 FILLER_ASAP7_75t_R FILLER_192_222 ();
 FILLER_ASAP7_75t_R FILLER_192_230 ();
 DECAPx6_ASAP7_75t_R FILLER_192_238 ();
 FILLER_ASAP7_75t_R FILLER_192_252 ();
 DECAPx2_ASAP7_75t_R FILLER_192_264 ();
 FILLER_ASAP7_75t_R FILLER_192_270 ();
 DECAPx6_ASAP7_75t_R FILLER_192_282 ();
 FILLER_ASAP7_75t_R FILLER_192_296 ();
 DECAPx4_ASAP7_75t_R FILLER_192_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_311 ();
 DECAPx1_ASAP7_75t_R FILLER_192_324 ();
 DECAPx10_ASAP7_75t_R FILLER_192_346 ();
 DECAPx10_ASAP7_75t_R FILLER_192_368 ();
 DECAPx1_ASAP7_75t_R FILLER_192_390 ();
 DECAPx10_ASAP7_75t_R FILLER_192_415 ();
 DECAPx10_ASAP7_75t_R FILLER_192_437 ();
 FILLER_ASAP7_75t_R FILLER_192_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_461 ();
 DECAPx6_ASAP7_75t_R FILLER_192_464 ();
 FILLER_ASAP7_75t_R FILLER_192_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_480 ();
 DECAPx1_ASAP7_75t_R FILLER_192_489 ();
 DECAPx4_ASAP7_75t_R FILLER_192_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_506 ();
 FILLER_ASAP7_75t_R FILLER_192_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_515 ();
 DECAPx10_ASAP7_75t_R FILLER_192_523 ();
 DECAPx6_ASAP7_75t_R FILLER_192_545 ();
 DECAPx1_ASAP7_75t_R FILLER_192_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_588 ();
 FILLER_ASAP7_75t_R FILLER_192_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_603 ();
 DECAPx2_ASAP7_75t_R FILLER_192_610 ();
 FILLER_ASAP7_75t_R FILLER_192_616 ();
 DECAPx2_ASAP7_75t_R FILLER_192_621 ();
 FILLER_ASAP7_75t_R FILLER_192_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_629 ();
 DECAPx10_ASAP7_75t_R FILLER_192_636 ();
 DECAPx6_ASAP7_75t_R FILLER_192_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_672 ();
 FILLER_ASAP7_75t_R FILLER_192_691 ();
 DECAPx6_ASAP7_75t_R FILLER_192_719 ();
 DECAPx1_ASAP7_75t_R FILLER_192_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_751 ();
 DECAPx2_ASAP7_75t_R FILLER_192_760 ();
 DECAPx2_ASAP7_75t_R FILLER_192_776 ();
 FILLER_ASAP7_75t_R FILLER_192_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_784 ();
 DECAPx4_ASAP7_75t_R FILLER_192_802 ();
 FILLER_ASAP7_75t_R FILLER_192_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_814 ();
 DECAPx1_ASAP7_75t_R FILLER_192_823 ();
 DECAPx4_ASAP7_75t_R FILLER_192_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_843 ();
 DECAPx2_ASAP7_75t_R FILLER_192_848 ();
 DECAPx2_ASAP7_75t_R FILLER_192_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_886 ();
 DECAPx1_ASAP7_75t_R FILLER_192_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_920 ();
 DECAPx4_ASAP7_75t_R FILLER_192_936 ();
 FILLER_ASAP7_75t_R FILLER_192_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_952 ();
 DECAPx1_ASAP7_75t_R FILLER_192_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_964 ();
 FILLER_ASAP7_75t_R FILLER_192_971 ();
 DECAPx6_ASAP7_75t_R FILLER_192_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1056 ();
 FILLER_ASAP7_75t_R FILLER_192_1086 ();
 FILLER_ASAP7_75t_R FILLER_192_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_192_1187 ();
 FILLER_ASAP7_75t_R FILLER_192_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1251 ();
 FILLER_ASAP7_75t_R FILLER_192_1273 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1302 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1306 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1333 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1342 ();
 FILLER_ASAP7_75t_R FILLER_192_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1391 ();
 DECAPx6_ASAP7_75t_R FILLER_193_2 ();
 FILLER_ASAP7_75t_R FILLER_193_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_25 ();
 FILLER_ASAP7_75t_R FILLER_193_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_104 ();
 DECAPx1_ASAP7_75t_R FILLER_193_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_112 ();
 DECAPx2_ASAP7_75t_R FILLER_193_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_163 ();
 DECAPx2_ASAP7_75t_R FILLER_193_170 ();
 FILLER_ASAP7_75t_R FILLER_193_176 ();
 DECAPx4_ASAP7_75t_R FILLER_193_186 ();
 DECAPx4_ASAP7_75t_R FILLER_193_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_220 ();
 DECAPx2_ASAP7_75t_R FILLER_193_235 ();
 FILLER_ASAP7_75t_R FILLER_193_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_243 ();
 DECAPx10_ASAP7_75t_R FILLER_193_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_272 ();
 DECAPx4_ASAP7_75t_R FILLER_193_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_308 ();
 DECAPx2_ASAP7_75t_R FILLER_193_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_325 ();
 FILLER_ASAP7_75t_R FILLER_193_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_346 ();
 DECAPx2_ASAP7_75t_R FILLER_193_361 ();
 FILLER_ASAP7_75t_R FILLER_193_367 ();
 DECAPx2_ASAP7_75t_R FILLER_193_375 ();
 DECAPx2_ASAP7_75t_R FILLER_193_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_411 ();
 DECAPx6_ASAP7_75t_R FILLER_193_420 ();
 DECAPx10_ASAP7_75t_R FILLER_193_452 ();
 FILLER_ASAP7_75t_R FILLER_193_474 ();
 DECAPx10_ASAP7_75t_R FILLER_193_488 ();
 DECAPx2_ASAP7_75t_R FILLER_193_510 ();
 FILLER_ASAP7_75t_R FILLER_193_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_518 ();
 DECAPx10_ASAP7_75t_R FILLER_193_526 ();
 DECAPx4_ASAP7_75t_R FILLER_193_548 ();
 FILLER_ASAP7_75t_R FILLER_193_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_586 ();
 DECAPx6_ASAP7_75t_R FILLER_193_607 ();
 FILLER_ASAP7_75t_R FILLER_193_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_623 ();
 DECAPx10_ASAP7_75t_R FILLER_193_657 ();
 DECAPx2_ASAP7_75t_R FILLER_193_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_685 ();
 DECAPx2_ASAP7_75t_R FILLER_193_702 ();
 DECAPx1_ASAP7_75t_R FILLER_193_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_715 ();
 FILLER_ASAP7_75t_R FILLER_193_733 ();
 DECAPx4_ASAP7_75t_R FILLER_193_749 ();
 DECAPx10_ASAP7_75t_R FILLER_193_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_828 ();
 FILLER_ASAP7_75t_R FILLER_193_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_867 ();
 DECAPx2_ASAP7_75t_R FILLER_193_878 ();
 DECAPx10_ASAP7_75t_R FILLER_193_894 ();
 DECAPx2_ASAP7_75t_R FILLER_193_916 ();
 FILLER_ASAP7_75t_R FILLER_193_922 ();
 DECAPx2_ASAP7_75t_R FILLER_193_926 ();
 FILLER_ASAP7_75t_R FILLER_193_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_934 ();
 FILLER_ASAP7_75t_R FILLER_193_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_950 ();
 DECAPx4_ASAP7_75t_R FILLER_193_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_978 ();
 DECAPx1_ASAP7_75t_R FILLER_193_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_986 ();
 FILLER_ASAP7_75t_R FILLER_193_990 ();
 DECAPx6_ASAP7_75t_R FILLER_193_1000 ();
 FILLER_ASAP7_75t_R FILLER_193_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_193_1025 ();
 FILLER_ASAP7_75t_R FILLER_193_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1074 ();
 FILLER_ASAP7_75t_R FILLER_193_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1090 ();
 FILLER_ASAP7_75t_R FILLER_193_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1122 ();
 FILLER_ASAP7_75t_R FILLER_193_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1179 ();
 FILLER_ASAP7_75t_R FILLER_193_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1187 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1211 ();
 FILLER_ASAP7_75t_R FILLER_193_1223 ();
 FILLER_ASAP7_75t_R FILLER_193_1251 ();
 FILLER_ASAP7_75t_R FILLER_193_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1310 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1317 ();
 DECAPx6_ASAP7_75t_R FILLER_193_1358 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1379 ();
 DECAPx4_ASAP7_75t_R FILLER_194_2 ();
 FILLER_ASAP7_75t_R FILLER_194_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_18 ();
 DECAPx1_ASAP7_75t_R FILLER_194_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_29 ();
 FILLER_ASAP7_75t_R FILLER_194_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_61 ();
 DECAPx6_ASAP7_75t_R FILLER_194_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_89 ();
 DECAPx4_ASAP7_75t_R FILLER_194_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_129 ();
 FILLER_ASAP7_75t_R FILLER_194_143 ();
 DECAPx1_ASAP7_75t_R FILLER_194_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_189 ();
 DECAPx1_ASAP7_75t_R FILLER_194_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_202 ();
 FILLER_ASAP7_75t_R FILLER_194_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_239 ();
 DECAPx2_ASAP7_75t_R FILLER_194_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_267 ();
 FILLER_ASAP7_75t_R FILLER_194_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_298 ();
 FILLER_ASAP7_75t_R FILLER_194_307 ();
 DECAPx6_ASAP7_75t_R FILLER_194_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_333 ();
 DECAPx1_ASAP7_75t_R FILLER_194_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_368 ();
 DECAPx1_ASAP7_75t_R FILLER_194_395 ();
 DECAPx4_ASAP7_75t_R FILLER_194_431 ();
 FILLER_ASAP7_75t_R FILLER_194_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_461 ();
 DECAPx2_ASAP7_75t_R FILLER_194_464 ();
 DECAPx2_ASAP7_75t_R FILLER_194_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_494 ();
 FILLER_ASAP7_75t_R FILLER_194_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_518 ();
 FILLER_ASAP7_75t_R FILLER_194_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_539 ();
 DECAPx4_ASAP7_75t_R FILLER_194_558 ();
 DECAPx2_ASAP7_75t_R FILLER_194_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_627 ();
 DECAPx4_ASAP7_75t_R FILLER_194_634 ();
 FILLER_ASAP7_75t_R FILLER_194_644 ();
 DECAPx1_ASAP7_75t_R FILLER_194_649 ();
 DECAPx10_ASAP7_75t_R FILLER_194_659 ();
 DECAPx2_ASAP7_75t_R FILLER_194_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_687 ();
 FILLER_ASAP7_75t_R FILLER_194_695 ();
 DECAPx4_ASAP7_75t_R FILLER_194_707 ();
 FILLER_ASAP7_75t_R FILLER_194_717 ();
 DECAPx6_ASAP7_75t_R FILLER_194_725 ();
 DECAPx2_ASAP7_75t_R FILLER_194_739 ();
 FILLER_ASAP7_75t_R FILLER_194_755 ();
 DECAPx2_ASAP7_75t_R FILLER_194_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_773 ();
 DECAPx1_ASAP7_75t_R FILLER_194_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_781 ();
 DECAPx6_ASAP7_75t_R FILLER_194_792 ();
 DECAPx1_ASAP7_75t_R FILLER_194_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_810 ();
 DECAPx1_ASAP7_75t_R FILLER_194_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_846 ();
 DECAPx2_ASAP7_75t_R FILLER_194_860 ();
 DECAPx6_ASAP7_75t_R FILLER_194_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_892 ();
 DECAPx4_ASAP7_75t_R FILLER_194_911 ();
 DECAPx2_ASAP7_75t_R FILLER_194_926 ();
 FILLER_ASAP7_75t_R FILLER_194_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_934 ();
 FILLER_ASAP7_75t_R FILLER_194_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_943 ();
 DECAPx2_ASAP7_75t_R FILLER_194_962 ();
 FILLER_ASAP7_75t_R FILLER_194_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_970 ();
 FILLER_ASAP7_75t_R FILLER_194_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_194_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1061 ();
 FILLER_ASAP7_75t_R FILLER_194_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1107 ();
 FILLER_ASAP7_75t_R FILLER_194_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1141 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1176 ();
 FILLER_ASAP7_75t_R FILLER_194_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1276 ();
 FILLER_ASAP7_75t_R FILLER_194_1298 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1356 ();
 FILLER_ASAP7_75t_R FILLER_194_1378 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1388 ();
 FILLER_ASAP7_75t_R FILLER_195_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_34 ();
 FILLER_ASAP7_75t_R FILLER_195_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_43 ();
 DECAPx6_ASAP7_75t_R FILLER_195_47 ();
 DECAPx1_ASAP7_75t_R FILLER_195_61 ();
 DECAPx2_ASAP7_75t_R FILLER_195_75 ();
 FILLER_ASAP7_75t_R FILLER_195_81 ();
 FILLER_ASAP7_75t_R FILLER_195_109 ();
 DECAPx10_ASAP7_75t_R FILLER_195_117 ();
 DECAPx10_ASAP7_75t_R FILLER_195_142 ();
 DECAPx2_ASAP7_75t_R FILLER_195_164 ();
 FILLER_ASAP7_75t_R FILLER_195_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_172 ();
 FILLER_ASAP7_75t_R FILLER_195_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_215 ();
 DECAPx1_ASAP7_75t_R FILLER_195_231 ();
 DECAPx2_ASAP7_75t_R FILLER_195_249 ();
 DECAPx1_ASAP7_75t_R FILLER_195_265 ();
 DECAPx4_ASAP7_75t_R FILLER_195_275 ();
 FILLER_ASAP7_75t_R FILLER_195_285 ();
 DECAPx1_ASAP7_75t_R FILLER_195_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_309 ();
 DECAPx10_ASAP7_75t_R FILLER_195_319 ();
 DECAPx6_ASAP7_75t_R FILLER_195_341 ();
 FILLER_ASAP7_75t_R FILLER_195_355 ();
 DECAPx1_ASAP7_75t_R FILLER_195_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_367 ();
 DECAPx4_ASAP7_75t_R FILLER_195_374 ();
 DECAPx2_ASAP7_75t_R FILLER_195_387 ();
 DECAPx4_ASAP7_75t_R FILLER_195_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_406 ();
 DECAPx4_ASAP7_75t_R FILLER_195_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_429 ();
 FILLER_ASAP7_75t_R FILLER_195_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_486 ();
 DECAPx6_ASAP7_75t_R FILLER_195_513 ();
 DECAPx6_ASAP7_75t_R FILLER_195_545 ();
 DECAPx2_ASAP7_75t_R FILLER_195_591 ();
 FILLER_ASAP7_75t_R FILLER_195_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_599 ();
 DECAPx2_ASAP7_75t_R FILLER_195_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_609 ();
 DECAPx2_ASAP7_75t_R FILLER_195_626 ();
 FILLER_ASAP7_75t_R FILLER_195_632 ();
 DECAPx1_ASAP7_75t_R FILLER_195_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_664 ();
 DECAPx2_ASAP7_75t_R FILLER_195_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_685 ();
 FILLER_ASAP7_75t_R FILLER_195_693 ();
 DECAPx2_ASAP7_75t_R FILLER_195_725 ();
 DECAPx6_ASAP7_75t_R FILLER_195_737 ();
 FILLER_ASAP7_75t_R FILLER_195_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_753 ();
 DECAPx10_ASAP7_75t_R FILLER_195_766 ();
 DECAPx1_ASAP7_75t_R FILLER_195_788 ();
 DECAPx6_ASAP7_75t_R FILLER_195_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_816 ();
 DECAPx10_ASAP7_75t_R FILLER_195_824 ();
 FILLER_ASAP7_75t_R FILLER_195_846 ();
 FILLER_ASAP7_75t_R FILLER_195_863 ();
 FILLER_ASAP7_75t_R FILLER_195_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_883 ();
 FILLER_ASAP7_75t_R FILLER_195_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_894 ();
 DECAPx4_ASAP7_75t_R FILLER_195_911 ();
 FILLER_ASAP7_75t_R FILLER_195_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_923 ();
 FILLER_ASAP7_75t_R FILLER_195_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_928 ();
 DECAPx6_ASAP7_75t_R FILLER_195_933 ();
 FILLER_ASAP7_75t_R FILLER_195_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_969 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1006 ();
 FILLER_ASAP7_75t_R FILLER_195_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_195_1031 ();
 FILLER_ASAP7_75t_R FILLER_195_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1167 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1180 ();
 FILLER_ASAP7_75t_R FILLER_195_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1225 ();
 FILLER_ASAP7_75t_R FILLER_195_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1274 ();
 FILLER_ASAP7_75t_R FILLER_195_1280 ();
 DECAPx4_ASAP7_75t_R FILLER_195_1285 ();
 FILLER_ASAP7_75t_R FILLER_195_1307 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1309 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1343 ();
 FILLER_ASAP7_75t_R FILLER_195_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1359 ();
 DECAPx10_ASAP7_75t_R FILLER_196_2 ();
 DECAPx2_ASAP7_75t_R FILLER_196_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_30 ();
 DECAPx10_ASAP7_75t_R FILLER_196_37 ();
 DECAPx2_ASAP7_75t_R FILLER_196_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_97 ();
 DECAPx4_ASAP7_75t_R FILLER_196_101 ();
 FILLER_ASAP7_75t_R FILLER_196_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_125 ();
 DECAPx6_ASAP7_75t_R FILLER_196_130 ();
 FILLER_ASAP7_75t_R FILLER_196_144 ();
 DECAPx1_ASAP7_75t_R FILLER_196_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_157 ();
 DECAPx2_ASAP7_75t_R FILLER_196_184 ();
 DECAPx2_ASAP7_75t_R FILLER_196_196 ();
 DECAPx10_ASAP7_75t_R FILLER_196_208 ();
 DECAPx4_ASAP7_75t_R FILLER_196_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_240 ();
 DECAPx2_ASAP7_75t_R FILLER_196_247 ();
 FILLER_ASAP7_75t_R FILLER_196_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_255 ();
 DECAPx6_ASAP7_75t_R FILLER_196_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_296 ();
 DECAPx2_ASAP7_75t_R FILLER_196_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_340 ();
 DECAPx10_ASAP7_75t_R FILLER_196_361 ();
 DECAPx2_ASAP7_75t_R FILLER_196_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_389 ();
 DECAPx2_ASAP7_75t_R FILLER_196_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_423 ();
 DECAPx1_ASAP7_75t_R FILLER_196_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_446 ();
 DECAPx1_ASAP7_75t_R FILLER_196_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_461 ();
 FILLER_ASAP7_75t_R FILLER_196_482 ();
 DECAPx2_ASAP7_75t_R FILLER_196_495 ();
 FILLER_ASAP7_75t_R FILLER_196_504 ();
 DECAPx6_ASAP7_75t_R FILLER_196_518 ();
 DECAPx1_ASAP7_75t_R FILLER_196_564 ();
 FILLER_ASAP7_75t_R FILLER_196_574 ();
 FILLER_ASAP7_75t_R FILLER_196_623 ();
 DECAPx2_ASAP7_75t_R FILLER_196_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_648 ();
 DECAPx6_ASAP7_75t_R FILLER_196_652 ();
 FILLER_ASAP7_75t_R FILLER_196_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_668 ();
 DECAPx1_ASAP7_75t_R FILLER_196_687 ();
 DECAPx4_ASAP7_75t_R FILLER_196_697 ();
 FILLER_ASAP7_75t_R FILLER_196_707 ();
 DECAPx2_ASAP7_75t_R FILLER_196_712 ();
 FILLER_ASAP7_75t_R FILLER_196_718 ();
 DECAPx1_ASAP7_75t_R FILLER_196_756 ();
 FILLER_ASAP7_75t_R FILLER_196_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_768 ();
 FILLER_ASAP7_75t_R FILLER_196_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_778 ();
 DECAPx4_ASAP7_75t_R FILLER_196_789 ();
 FILLER_ASAP7_75t_R FILLER_196_809 ();
 DECAPx2_ASAP7_75t_R FILLER_196_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_836 ();
 DECAPx4_ASAP7_75t_R FILLER_196_843 ();
 FILLER_ASAP7_75t_R FILLER_196_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_855 ();
 DECAPx2_ASAP7_75t_R FILLER_196_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_872 ();
 DECAPx2_ASAP7_75t_R FILLER_196_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_904 ();
 DECAPx1_ASAP7_75t_R FILLER_196_933 ();
 DECAPx2_ASAP7_75t_R FILLER_196_947 ();
 FILLER_ASAP7_75t_R FILLER_196_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_955 ();
 DECAPx6_ASAP7_75t_R FILLER_196_966 ();
 FILLER_ASAP7_75t_R FILLER_196_980 ();
 FILLER_ASAP7_75t_R FILLER_196_988 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1030 ();
 FILLER_ASAP7_75t_R FILLER_196_1062 ();
 DECAPx4_ASAP7_75t_R FILLER_196_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_196_1135 ();
 FILLER_ASAP7_75t_R FILLER_196_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1155 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1184 ();
 FILLER_ASAP7_75t_R FILLER_196_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1219 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1255 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1268 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1272 ();
 FILLER_ASAP7_75t_R FILLER_196_1286 ();
 FILLER_ASAP7_75t_R FILLER_196_1314 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1323 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1336 ();
 FILLER_ASAP7_75t_R FILLER_196_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1347 ();
 FILLER_ASAP7_75t_R FILLER_196_1360 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1391 ();
 DECAPx6_ASAP7_75t_R FILLER_197_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_16 ();
 DECAPx1_ASAP7_75t_R FILLER_197_56 ();
 DECAPx2_ASAP7_75t_R FILLER_197_95 ();
 FILLER_ASAP7_75t_R FILLER_197_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_129 ();
 FILLER_ASAP7_75t_R FILLER_197_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_139 ();
 FILLER_ASAP7_75t_R FILLER_197_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_185 ();
 DECAPx1_ASAP7_75t_R FILLER_197_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_197 ();
 DECAPx6_ASAP7_75t_R FILLER_197_206 ();
 DECAPx2_ASAP7_75t_R FILLER_197_238 ();
 FILLER_ASAP7_75t_R FILLER_197_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_246 ();
 DECAPx4_ASAP7_75t_R FILLER_197_253 ();
 DECAPx4_ASAP7_75t_R FILLER_197_274 ();
 FILLER_ASAP7_75t_R FILLER_197_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_286 ();
 DECAPx4_ASAP7_75t_R FILLER_197_295 ();
 FILLER_ASAP7_75t_R FILLER_197_305 ();
 DECAPx2_ASAP7_75t_R FILLER_197_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_319 ();
 DECAPx2_ASAP7_75t_R FILLER_197_327 ();
 DECAPx1_ASAP7_75t_R FILLER_197_362 ();
 DECAPx6_ASAP7_75t_R FILLER_197_380 ();
 DECAPx2_ASAP7_75t_R FILLER_197_394 ();
 DECAPx6_ASAP7_75t_R FILLER_197_414 ();
 DECAPx10_ASAP7_75t_R FILLER_197_446 ();
 DECAPx2_ASAP7_75t_R FILLER_197_468 ();
 DECAPx1_ASAP7_75t_R FILLER_197_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_498 ();
 DECAPx6_ASAP7_75t_R FILLER_197_511 ();
 DECAPx2_ASAP7_75t_R FILLER_197_533 ();
 DECAPx2_ASAP7_75t_R FILLER_197_547 ();
 DECAPx10_ASAP7_75t_R FILLER_197_556 ();
 DECAPx4_ASAP7_75t_R FILLER_197_578 ();
 DECAPx6_ASAP7_75t_R FILLER_197_596 ();
 FILLER_ASAP7_75t_R FILLER_197_610 ();
 DECAPx10_ASAP7_75t_R FILLER_197_638 ();
 DECAPx10_ASAP7_75t_R FILLER_197_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_682 ();
 FILLER_ASAP7_75t_R FILLER_197_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_691 ();
 DECAPx2_ASAP7_75t_R FILLER_197_707 ();
 FILLER_ASAP7_75t_R FILLER_197_713 ();
 FILLER_ASAP7_75t_R FILLER_197_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_742 ();
 DECAPx2_ASAP7_75t_R FILLER_197_786 ();
 FILLER_ASAP7_75t_R FILLER_197_792 ();
 DECAPx1_ASAP7_75t_R FILLER_197_822 ();
 DECAPx2_ASAP7_75t_R FILLER_197_862 ();
 FILLER_ASAP7_75t_R FILLER_197_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_870 ();
 FILLER_ASAP7_75t_R FILLER_197_881 ();
 DECAPx2_ASAP7_75t_R FILLER_197_891 ();
 FILLER_ASAP7_75t_R FILLER_197_897 ();
 DECAPx6_ASAP7_75t_R FILLER_197_907 ();
 FILLER_ASAP7_75t_R FILLER_197_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_923 ();
 DECAPx1_ASAP7_75t_R FILLER_197_926 ();
 DECAPx2_ASAP7_75t_R FILLER_197_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_945 ();
 DECAPx1_ASAP7_75t_R FILLER_197_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_973 ();
 DECAPx10_ASAP7_75t_R FILLER_197_977 ();
 DECAPx2_ASAP7_75t_R FILLER_197_999 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1057 ();
 FILLER_ASAP7_75t_R FILLER_197_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1067 ();
 DECAPx6_ASAP7_75t_R FILLER_197_1071 ();
 FILLER_ASAP7_75t_R FILLER_197_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1101 ();
 FILLER_ASAP7_75t_R FILLER_197_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1109 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1134 ();
 FILLER_ASAP7_75t_R FILLER_197_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_197_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1168 ();
 FILLER_ASAP7_75t_R FILLER_197_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1211 ();
 FILLER_ASAP7_75t_R FILLER_197_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1241 ();
 DECAPx4_ASAP7_75t_R FILLER_197_1280 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1307 ();
 FILLER_ASAP7_75t_R FILLER_197_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1341 ();
 FILLER_ASAP7_75t_R FILLER_197_1347 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1365 ();
 DECAPx4_ASAP7_75t_R FILLER_198_2 ();
 FILLER_ASAP7_75t_R FILLER_198_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_36 ();
 FILLER_ASAP7_75t_R FILLER_198_48 ();
 DECAPx4_ASAP7_75t_R FILLER_198_53 ();
 FILLER_ASAP7_75t_R FILLER_198_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_65 ();
 FILLER_ASAP7_75t_R FILLER_198_72 ();
 DECAPx4_ASAP7_75t_R FILLER_198_77 ();
 DECAPx10_ASAP7_75t_R FILLER_198_93 ();
 FILLER_ASAP7_75t_R FILLER_198_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_120 ();
 DECAPx2_ASAP7_75t_R FILLER_198_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_153 ();
 DECAPx2_ASAP7_75t_R FILLER_198_157 ();
 DECAPx6_ASAP7_75t_R FILLER_198_177 ();
 DECAPx1_ASAP7_75t_R FILLER_198_191 ();
 DECAPx4_ASAP7_75t_R FILLER_198_209 ();
 FILLER_ASAP7_75t_R FILLER_198_219 ();
 DECAPx2_ASAP7_75t_R FILLER_198_254 ();
 FILLER_ASAP7_75t_R FILLER_198_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_262 ();
 DECAPx6_ASAP7_75t_R FILLER_198_269 ();
 FILLER_ASAP7_75t_R FILLER_198_283 ();
 DECAPx2_ASAP7_75t_R FILLER_198_297 ();
 FILLER_ASAP7_75t_R FILLER_198_303 ();
 DECAPx2_ASAP7_75t_R FILLER_198_311 ();
 FILLER_ASAP7_75t_R FILLER_198_317 ();
 DECAPx6_ASAP7_75t_R FILLER_198_325 ();
 DECAPx1_ASAP7_75t_R FILLER_198_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_343 ();
 DECAPx6_ASAP7_75t_R FILLER_198_384 ();
 FILLER_ASAP7_75t_R FILLER_198_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_400 ();
 DECAPx10_ASAP7_75t_R FILLER_198_409 ();
 DECAPx2_ASAP7_75t_R FILLER_198_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_437 ();
 DECAPx2_ASAP7_75t_R FILLER_198_456 ();
 DECAPx6_ASAP7_75t_R FILLER_198_464 ();
 DECAPx4_ASAP7_75t_R FILLER_198_490 ();
 FILLER_ASAP7_75t_R FILLER_198_500 ();
 DECAPx4_ASAP7_75t_R FILLER_198_508 ();
 FILLER_ASAP7_75t_R FILLER_198_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_552 ();
 DECAPx2_ASAP7_75t_R FILLER_198_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_565 ();
 DECAPx2_ASAP7_75t_R FILLER_198_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_580 ();
 DECAPx10_ASAP7_75t_R FILLER_198_597 ();
 DECAPx2_ASAP7_75t_R FILLER_198_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_625 ();
 DECAPx2_ASAP7_75t_R FILLER_198_640 ();
 FILLER_ASAP7_75t_R FILLER_198_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_648 ();
 DECAPx1_ASAP7_75t_R FILLER_198_652 ();
 DECAPx2_ASAP7_75t_R FILLER_198_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_680 ();
 DECAPx1_ASAP7_75t_R FILLER_198_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_697 ();
 DECAPx1_ASAP7_75t_R FILLER_198_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_709 ();
 DECAPx4_ASAP7_75t_R FILLER_198_717 ();
 DECAPx10_ASAP7_75t_R FILLER_198_730 ();
 FILLER_ASAP7_75t_R FILLER_198_752 ();
 DECAPx4_ASAP7_75t_R FILLER_198_764 ();
 FILLER_ASAP7_75t_R FILLER_198_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_779 ();
 DECAPx2_ASAP7_75t_R FILLER_198_790 ();
 DECAPx10_ASAP7_75t_R FILLER_198_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_836 ();
 DECAPx10_ASAP7_75t_R FILLER_198_843 ();
 DECAPx6_ASAP7_75t_R FILLER_198_865 ();
 DECAPx1_ASAP7_75t_R FILLER_198_879 ();
 DECAPx10_ASAP7_75t_R FILLER_198_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_929 ();
 DECAPx6_ASAP7_75t_R FILLER_198_944 ();
 DECAPx4_ASAP7_75t_R FILLER_198_984 ();
 FILLER_ASAP7_75t_R FILLER_198_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_996 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1036 ();
 DECAPx6_ASAP7_75t_R FILLER_198_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1061 ();
 FILLER_ASAP7_75t_R FILLER_198_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_198_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1166 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1203 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1223 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1250 ();
 FILLER_ASAP7_75t_R FILLER_198_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1324 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1333 ();
 FILLER_ASAP7_75t_R FILLER_198_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1345 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1358 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1370 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_199_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_61 ();
 DECAPx4_ASAP7_75t_R FILLER_199_65 ();
 FILLER_ASAP7_75t_R FILLER_199_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_77 ();
 FILLER_ASAP7_75t_R FILLER_199_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_106 ();
 DECAPx6_ASAP7_75t_R FILLER_199_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_131 ();
 DECAPx6_ASAP7_75t_R FILLER_199_148 ();
 FILLER_ASAP7_75t_R FILLER_199_162 ();
 DECAPx4_ASAP7_75t_R FILLER_199_176 ();
 FILLER_ASAP7_75t_R FILLER_199_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_188 ();
 DECAPx1_ASAP7_75t_R FILLER_199_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_213 ();
 DECAPx2_ASAP7_75t_R FILLER_199_228 ();
 FILLER_ASAP7_75t_R FILLER_199_234 ();
 DECAPx1_ASAP7_75t_R FILLER_199_239 ();
 DECAPx2_ASAP7_75t_R FILLER_199_250 ();
 FILLER_ASAP7_75t_R FILLER_199_262 ();
 FILLER_ASAP7_75t_R FILLER_199_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_274 ();
 DECAPx2_ASAP7_75t_R FILLER_199_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_317 ();
 DECAPx1_ASAP7_75t_R FILLER_199_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_336 ();
 FILLER_ASAP7_75t_R FILLER_199_345 ();
 DECAPx1_ASAP7_75t_R FILLER_199_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_354 ();
 DECAPx4_ASAP7_75t_R FILLER_199_361 ();
 FILLER_ASAP7_75t_R FILLER_199_371 ();
 DECAPx2_ASAP7_75t_R FILLER_199_387 ();
 FILLER_ASAP7_75t_R FILLER_199_393 ();
 DECAPx2_ASAP7_75t_R FILLER_199_413 ();
 DECAPx1_ASAP7_75t_R FILLER_199_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_441 ();
 FILLER_ASAP7_75t_R FILLER_199_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_500 ();
 DECAPx4_ASAP7_75t_R FILLER_199_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_537 ();
 DECAPx4_ASAP7_75t_R FILLER_199_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_551 ();
 FILLER_ASAP7_75t_R FILLER_199_558 ();
 DECAPx2_ASAP7_75t_R FILLER_199_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_624 ();
 DECAPx6_ASAP7_75t_R FILLER_199_661 ();
 FILLER_ASAP7_75t_R FILLER_199_675 ();
 DECAPx10_ASAP7_75t_R FILLER_199_691 ();
 DECAPx1_ASAP7_75t_R FILLER_199_713 ();
 DECAPx2_ASAP7_75t_R FILLER_199_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_733 ();
 FILLER_ASAP7_75t_R FILLER_199_737 ();
 DECAPx4_ASAP7_75t_R FILLER_199_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_756 ();
 DECAPx6_ASAP7_75t_R FILLER_199_765 ();
 DECAPx1_ASAP7_75t_R FILLER_199_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_783 ();
 DECAPx10_ASAP7_75t_R FILLER_199_794 ();
 FILLER_ASAP7_75t_R FILLER_199_816 ();
 FILLER_ASAP7_75t_R FILLER_199_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_838 ();
 DECAPx2_ASAP7_75t_R FILLER_199_849 ();
 DECAPx1_ASAP7_75t_R FILLER_199_869 ();
 DECAPx2_ASAP7_75t_R FILLER_199_883 ();
 DECAPx2_ASAP7_75t_R FILLER_199_895 ();
 FILLER_ASAP7_75t_R FILLER_199_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_926 ();
 DECAPx10_ASAP7_75t_R FILLER_199_935 ();
 DECAPx2_ASAP7_75t_R FILLER_199_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_963 ();
 FILLER_ASAP7_75t_R FILLER_199_985 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1013 ();
 FILLER_ASAP7_75t_R FILLER_199_1019 ();
 DECAPx4_ASAP7_75t_R FILLER_199_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1038 ();
 FILLER_ASAP7_75t_R FILLER_199_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1059 ();
 FILLER_ASAP7_75t_R FILLER_199_1065 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1104 ();
 FILLER_ASAP7_75t_R FILLER_199_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1120 ();
 DECAPx4_ASAP7_75t_R FILLER_199_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1171 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1186 ();
 FILLER_ASAP7_75t_R FILLER_199_1200 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1222 ();
 FILLER_ASAP7_75t_R FILLER_199_1236 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1244 ();
 DECAPx1_ASAP7_75t_R FILLER_199_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_199_1298 ();
 FILLER_ASAP7_75t_R FILLER_199_1308 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1344 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1357 ();
 FILLER_ASAP7_75t_R FILLER_199_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1391 ();
 DECAPx4_ASAP7_75t_R FILLER_200_2 ();
 FILLER_ASAP7_75t_R FILLER_200_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_14 ();
 DECAPx2_ASAP7_75t_R FILLER_200_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_24 ();
 FILLER_ASAP7_75t_R FILLER_200_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_35 ();
 DECAPx2_ASAP7_75t_R FILLER_200_40 ();
 DECAPx4_ASAP7_75t_R FILLER_200_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_62 ();
 DECAPx1_ASAP7_75t_R FILLER_200_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_81 ();
 DECAPx1_ASAP7_75t_R FILLER_200_88 ();
 DECAPx1_ASAP7_75t_R FILLER_200_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_99 ();
 DECAPx4_ASAP7_75t_R FILLER_200_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_139 ();
 DECAPx4_ASAP7_75t_R FILLER_200_166 ();
 FILLER_ASAP7_75t_R FILLER_200_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_182 ();
 FILLER_ASAP7_75t_R FILLER_200_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_193 ();
 DECAPx1_ASAP7_75t_R FILLER_200_208 ();
 DECAPx4_ASAP7_75t_R FILLER_200_220 ();
 FILLER_ASAP7_75t_R FILLER_200_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_232 ();
 DECAPx1_ASAP7_75t_R FILLER_200_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_263 ();
 DECAPx1_ASAP7_75t_R FILLER_200_270 ();
 DECAPx1_ASAP7_75t_R FILLER_200_294 ();
 DECAPx2_ASAP7_75t_R FILLER_200_324 ();
 FILLER_ASAP7_75t_R FILLER_200_330 ();
 FILLER_ASAP7_75t_R FILLER_200_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_360 ();
 DECAPx2_ASAP7_75t_R FILLER_200_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_375 ();
 DECAPx2_ASAP7_75t_R FILLER_200_388 ();
 FILLER_ASAP7_75t_R FILLER_200_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_396 ();
 DECAPx6_ASAP7_75t_R FILLER_200_411 ();
 DECAPx1_ASAP7_75t_R FILLER_200_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_429 ();
 DECAPx6_ASAP7_75t_R FILLER_200_448 ();
 FILLER_ASAP7_75t_R FILLER_200_490 ();
 DECAPx2_ASAP7_75t_R FILLER_200_508 ();
 FILLER_ASAP7_75t_R FILLER_200_514 ();
 FILLER_ASAP7_75t_R FILLER_200_519 ();
 DECAPx2_ASAP7_75t_R FILLER_200_537 ();
 FILLER_ASAP7_75t_R FILLER_200_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_545 ();
 DECAPx2_ASAP7_75t_R FILLER_200_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_555 ();
 FILLER_ASAP7_75t_R FILLER_200_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_564 ();
 DECAPx1_ASAP7_75t_R FILLER_200_575 ();
 DECAPx1_ASAP7_75t_R FILLER_200_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_586 ();
 DECAPx1_ASAP7_75t_R FILLER_200_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_599 ();
 DECAPx6_ASAP7_75t_R FILLER_200_637 ();
 DECAPx1_ASAP7_75t_R FILLER_200_651 ();
 DECAPx2_ASAP7_75t_R FILLER_200_662 ();
 DECAPx2_ASAP7_75t_R FILLER_200_671 ();
 FILLER_ASAP7_75t_R FILLER_200_693 ();
 DECAPx4_ASAP7_75t_R FILLER_200_702 ();
 DECAPx6_ASAP7_75t_R FILLER_200_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_732 ();
 FILLER_ASAP7_75t_R FILLER_200_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_743 ();
 DECAPx2_ASAP7_75t_R FILLER_200_750 ();
 FILLER_ASAP7_75t_R FILLER_200_756 ();
 DECAPx2_ASAP7_75t_R FILLER_200_764 ();
 FILLER_ASAP7_75t_R FILLER_200_770 ();
 DECAPx10_ASAP7_75t_R FILLER_200_780 ();
 DECAPx4_ASAP7_75t_R FILLER_200_802 ();
 FILLER_ASAP7_75t_R FILLER_200_812 ();
 DECAPx4_ASAP7_75t_R FILLER_200_820 ();
 FILLER_ASAP7_75t_R FILLER_200_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_860 ();
 DECAPx4_ASAP7_75t_R FILLER_200_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_927 ();
 DECAPx4_ASAP7_75t_R FILLER_200_934 ();
 DECAPx6_ASAP7_75t_R FILLER_200_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_982 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1009 ();
 FILLER_ASAP7_75t_R FILLER_200_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1069 ();
 FILLER_ASAP7_75t_R FILLER_200_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1111 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1152 ();
 FILLER_ASAP7_75t_R FILLER_200_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1176 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_200_1197 ();
 FILLER_ASAP7_75t_R FILLER_200_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1233 ();
 DECAPx4_ASAP7_75t_R FILLER_200_1259 ();
 FILLER_ASAP7_75t_R FILLER_200_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1279 ();
 FILLER_ASAP7_75t_R FILLER_200_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1296 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1305 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1376 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1391 ();
 DECAPx1_ASAP7_75t_R FILLER_201_2 ();
 DECAPx6_ASAP7_75t_R FILLER_201_38 ();
 DECAPx1_ASAP7_75t_R FILLER_201_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_90 ();
 DECAPx4_ASAP7_75t_R FILLER_201_94 ();
 FILLER_ASAP7_75t_R FILLER_201_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_113 ();
 DECAPx6_ASAP7_75t_R FILLER_201_123 ();
 FILLER_ASAP7_75t_R FILLER_201_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_153 ();
 DECAPx2_ASAP7_75t_R FILLER_201_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_163 ();
 DECAPx6_ASAP7_75t_R FILLER_201_196 ();
 DECAPx2_ASAP7_75t_R FILLER_201_210 ();
 DECAPx6_ASAP7_75t_R FILLER_201_229 ();
 DECAPx1_ASAP7_75t_R FILLER_201_243 ();
 DECAPx1_ASAP7_75t_R FILLER_201_250 ();
 DECAPx6_ASAP7_75t_R FILLER_201_260 ();
 DECAPx2_ASAP7_75t_R FILLER_201_294 ();
 FILLER_ASAP7_75t_R FILLER_201_300 ();
 DECAPx4_ASAP7_75t_R FILLER_201_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_318 ();
 DECAPx6_ASAP7_75t_R FILLER_201_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_341 ();
 DECAPx2_ASAP7_75t_R FILLER_201_351 ();
 DECAPx1_ASAP7_75t_R FILLER_201_360 ();
 DECAPx1_ASAP7_75t_R FILLER_201_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_376 ();
 DECAPx1_ASAP7_75t_R FILLER_201_391 ();
 DECAPx10_ASAP7_75t_R FILLER_201_421 ();
 DECAPx10_ASAP7_75t_R FILLER_201_443 ();
 DECAPx2_ASAP7_75t_R FILLER_201_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_500 ();
 DECAPx10_ASAP7_75t_R FILLER_201_507 ();
 FILLER_ASAP7_75t_R FILLER_201_529 ();
 FILLER_ASAP7_75t_R FILLER_201_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_565 ();
 DECAPx10_ASAP7_75t_R FILLER_201_572 ();
 DECAPx4_ASAP7_75t_R FILLER_201_594 ();
 FILLER_ASAP7_75t_R FILLER_201_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_606 ();
 FILLER_ASAP7_75t_R FILLER_201_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_617 ();
 DECAPx2_ASAP7_75t_R FILLER_201_621 ();
 FILLER_ASAP7_75t_R FILLER_201_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_712 ();
 DECAPx1_ASAP7_75t_R FILLER_201_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_729 ();
 FILLER_ASAP7_75t_R FILLER_201_746 ();
 DECAPx1_ASAP7_75t_R FILLER_201_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_772 ();
 DECAPx10_ASAP7_75t_R FILLER_201_793 ();
 DECAPx2_ASAP7_75t_R FILLER_201_815 ();
 DECAPx4_ASAP7_75t_R FILLER_201_827 ();
 FILLER_ASAP7_75t_R FILLER_201_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_839 ();
 FILLER_ASAP7_75t_R FILLER_201_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_860 ();
 DECAPx1_ASAP7_75t_R FILLER_201_868 ();
 DECAPx2_ASAP7_75t_R FILLER_201_880 ();
 DECAPx2_ASAP7_75t_R FILLER_201_900 ();
 FILLER_ASAP7_75t_R FILLER_201_906 ();
 DECAPx2_ASAP7_75t_R FILLER_201_915 ();
 FILLER_ASAP7_75t_R FILLER_201_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_923 ();
 DECAPx1_ASAP7_75t_R FILLER_201_956 ();
 DECAPx2_ASAP7_75t_R FILLER_201_980 ();
 FILLER_ASAP7_75t_R FILLER_201_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_997 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1021 ();
 FILLER_ASAP7_75t_R FILLER_201_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1029 ();
 FILLER_ASAP7_75t_R FILLER_201_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1045 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1053 ();
 DECAPx4_ASAP7_75t_R FILLER_201_1060 ();
 FILLER_ASAP7_75t_R FILLER_201_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1099 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1126 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1158 ();
 FILLER_ASAP7_75t_R FILLER_201_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1164 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1187 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1255 ();
 FILLER_ASAP7_75t_R FILLER_201_1261 ();
 FILLER_ASAP7_75t_R FILLER_201_1280 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1282 ();
 FILLER_ASAP7_75t_R FILLER_201_1289 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1302 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1323 ();
 FILLER_ASAP7_75t_R FILLER_201_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1335 ();
 FILLER_ASAP7_75t_R FILLER_201_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1359 ();
 DECAPx6_ASAP7_75t_R FILLER_202_2 ();
 DECAPx1_ASAP7_75t_R FILLER_202_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_24 ();
 DECAPx4_ASAP7_75t_R FILLER_202_33 ();
 FILLER_ASAP7_75t_R FILLER_202_43 ();
 FILLER_ASAP7_75t_R FILLER_202_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_55 ();
 DECAPx4_ASAP7_75t_R FILLER_202_59 ();
 FILLER_ASAP7_75t_R FILLER_202_69 ();
 FILLER_ASAP7_75t_R FILLER_202_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_76 ();
 DECAPx4_ASAP7_75t_R FILLER_202_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_113 ();
 DECAPx2_ASAP7_75t_R FILLER_202_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_134 ();
 DECAPx2_ASAP7_75t_R FILLER_202_161 ();
 FILLER_ASAP7_75t_R FILLER_202_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_169 ();
 DECAPx6_ASAP7_75t_R FILLER_202_188 ();
 FILLER_ASAP7_75t_R FILLER_202_202 ();
 FILLER_ASAP7_75t_R FILLER_202_230 ();
 FILLER_ASAP7_75t_R FILLER_202_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_254 ();
 DECAPx4_ASAP7_75t_R FILLER_202_269 ();
 FILLER_ASAP7_75t_R FILLER_202_279 ();
 DECAPx2_ASAP7_75t_R FILLER_202_287 ();
 FILLER_ASAP7_75t_R FILLER_202_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_295 ();
 DECAPx2_ASAP7_75t_R FILLER_202_311 ();
 DECAPx10_ASAP7_75t_R FILLER_202_331 ();
 FILLER_ASAP7_75t_R FILLER_202_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_355 ();
 DECAPx4_ASAP7_75t_R FILLER_202_368 ();
 FILLER_ASAP7_75t_R FILLER_202_378 ();
 FILLER_ASAP7_75t_R FILLER_202_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_394 ();
 FILLER_ASAP7_75t_R FILLER_202_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_409 ();
 DECAPx1_ASAP7_75t_R FILLER_202_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_417 ();
 DECAPx6_ASAP7_75t_R FILLER_202_424 ();
 DECAPx1_ASAP7_75t_R FILLER_202_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_461 ();
 DECAPx2_ASAP7_75t_R FILLER_202_464 ();
 FILLER_ASAP7_75t_R FILLER_202_470 ();
 DECAPx6_ASAP7_75t_R FILLER_202_489 ();
 DECAPx2_ASAP7_75t_R FILLER_202_503 ();
 DECAPx1_ASAP7_75t_R FILLER_202_517 ();
 FILLER_ASAP7_75t_R FILLER_202_527 ();
 DECAPx10_ASAP7_75t_R FILLER_202_537 ();
 DECAPx2_ASAP7_75t_R FILLER_202_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_565 ();
 FILLER_ASAP7_75t_R FILLER_202_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_576 ();
 DECAPx1_ASAP7_75t_R FILLER_202_580 ();
 DECAPx2_ASAP7_75t_R FILLER_202_595 ();
 FILLER_ASAP7_75t_R FILLER_202_601 ();
 DECAPx10_ASAP7_75t_R FILLER_202_606 ();
 DECAPx2_ASAP7_75t_R FILLER_202_634 ();
 FILLER_ASAP7_75t_R FILLER_202_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_642 ();
 DECAPx1_ASAP7_75t_R FILLER_202_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_650 ();
 DECAPx4_ASAP7_75t_R FILLER_202_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_675 ();
 FILLER_ASAP7_75t_R FILLER_202_693 ();
 DECAPx1_ASAP7_75t_R FILLER_202_703 ();
 FILLER_ASAP7_75t_R FILLER_202_719 ();
 DECAPx6_ASAP7_75t_R FILLER_202_735 ();
 FILLER_ASAP7_75t_R FILLER_202_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_761 ();
 DECAPx1_ASAP7_75t_R FILLER_202_768 ();
 DECAPx6_ASAP7_75t_R FILLER_202_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_798 ();
 DECAPx4_ASAP7_75t_R FILLER_202_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_816 ();
 DECAPx4_ASAP7_75t_R FILLER_202_835 ();
 FILLER_ASAP7_75t_R FILLER_202_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_856 ();
 DECAPx2_ASAP7_75t_R FILLER_202_867 ();
 DECAPx4_ASAP7_75t_R FILLER_202_879 ();
 FILLER_ASAP7_75t_R FILLER_202_889 ();
 DECAPx4_ASAP7_75t_R FILLER_202_898 ();
 FILLER_ASAP7_75t_R FILLER_202_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_910 ();
 FILLER_ASAP7_75t_R FILLER_202_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_927 ();
 DECAPx1_ASAP7_75t_R FILLER_202_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_938 ();
 DECAPx6_ASAP7_75t_R FILLER_202_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_967 ();
 DECAPx6_ASAP7_75t_R FILLER_202_975 ();
 DECAPx6_ASAP7_75t_R FILLER_202_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_202_1054 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1072 ();
 FILLER_ASAP7_75t_R FILLER_202_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1088 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1114 ();
 FILLER_ASAP7_75t_R FILLER_202_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1127 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1171 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1186 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1209 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1217 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1228 ();
 DECAPx4_ASAP7_75t_R FILLER_202_1252 ();
 FILLER_ASAP7_75t_R FILLER_202_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1290 ();
 FILLER_ASAP7_75t_R FILLER_202_1296 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1306 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1328 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1348 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1356 ();
 FILLER_ASAP7_75t_R FILLER_202_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1364 ();
 FILLER_ASAP7_75t_R FILLER_202_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1373 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_203_2 ();
 FILLER_ASAP7_75t_R FILLER_203_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_14 ();
 DECAPx10_ASAP7_75t_R FILLER_203_67 ();
 DECAPx4_ASAP7_75t_R FILLER_203_95 ();
 FILLER_ASAP7_75t_R FILLER_203_105 ();
 DECAPx4_ASAP7_75t_R FILLER_203_133 ();
 DECAPx10_ASAP7_75t_R FILLER_203_152 ();
 DECAPx6_ASAP7_75t_R FILLER_203_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_188 ();
 DECAPx4_ASAP7_75t_R FILLER_203_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_217 ();
 DECAPx6_ASAP7_75t_R FILLER_203_221 ();
 FILLER_ASAP7_75t_R FILLER_203_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_237 ();
 FILLER_ASAP7_75t_R FILLER_203_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_248 ();
 DECAPx1_ASAP7_75t_R FILLER_203_263 ();
 FILLER_ASAP7_75t_R FILLER_203_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_277 ();
 DECAPx1_ASAP7_75t_R FILLER_203_289 ();
 FILLER_ASAP7_75t_R FILLER_203_319 ();
 DECAPx6_ASAP7_75t_R FILLER_203_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_361 ();
 DECAPx2_ASAP7_75t_R FILLER_203_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_400 ();
 DECAPx4_ASAP7_75t_R FILLER_203_404 ();
 FILLER_ASAP7_75t_R FILLER_203_414 ();
 FILLER_ASAP7_75t_R FILLER_203_424 ();
 FILLER_ASAP7_75t_R FILLER_203_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_462 ();
 DECAPx4_ASAP7_75t_R FILLER_203_481 ();
 FILLER_ASAP7_75t_R FILLER_203_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_502 ();
 FILLER_ASAP7_75t_R FILLER_203_517 ();
 FILLER_ASAP7_75t_R FILLER_203_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_539 ();
 DECAPx2_ASAP7_75t_R FILLER_203_546 ();
 FILLER_ASAP7_75t_R FILLER_203_552 ();
 FILLER_ASAP7_75t_R FILLER_203_560 ();
 DECAPx6_ASAP7_75t_R FILLER_203_614 ();
 DECAPx2_ASAP7_75t_R FILLER_203_636 ();
 DECAPx2_ASAP7_75t_R FILLER_203_645 ();
 DECAPx2_ASAP7_75t_R FILLER_203_667 ();
 FILLER_ASAP7_75t_R FILLER_203_673 ();
 FILLER_ASAP7_75t_R FILLER_203_681 ();
 DECAPx1_ASAP7_75t_R FILLER_203_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_695 ();
 FILLER_ASAP7_75t_R FILLER_203_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_704 ();
 DECAPx6_ASAP7_75t_R FILLER_203_709 ();
 DECAPx1_ASAP7_75t_R FILLER_203_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_727 ();
 DECAPx10_ASAP7_75t_R FILLER_203_734 ();
 FILLER_ASAP7_75t_R FILLER_203_756 ();
 DECAPx1_ASAP7_75t_R FILLER_203_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_770 ();
 DECAPx10_ASAP7_75t_R FILLER_203_779 ();
 DECAPx10_ASAP7_75t_R FILLER_203_801 ();
 DECAPx2_ASAP7_75t_R FILLER_203_823 ();
 FILLER_ASAP7_75t_R FILLER_203_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_831 ();
 DECAPx1_ASAP7_75t_R FILLER_203_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_841 ();
 DECAPx4_ASAP7_75t_R FILLER_203_858 ();
 DECAPx6_ASAP7_75t_R FILLER_203_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_895 ();
 FILLER_ASAP7_75t_R FILLER_203_912 ();
 DECAPx10_ASAP7_75t_R FILLER_203_926 ();
 DECAPx6_ASAP7_75t_R FILLER_203_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_962 ();
 DECAPx4_ASAP7_75t_R FILLER_203_970 ();
 FILLER_ASAP7_75t_R FILLER_203_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_982 ();
 FILLER_ASAP7_75t_R FILLER_203_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1028 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1044 ();
 FILLER_ASAP7_75t_R FILLER_203_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1072 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1140 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1160 ();
 FILLER_ASAP7_75t_R FILLER_203_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1168 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1187 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1206 ();
 DECAPx6_ASAP7_75t_R FILLER_203_1219 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1255 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1276 ();
 FILLER_ASAP7_75t_R FILLER_203_1287 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1307 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1318 ();
 FILLER_ASAP7_75t_R FILLER_203_1327 ();
 FILLER_ASAP7_75t_R FILLER_203_1364 ();
 DECAPx10_ASAP7_75t_R FILLER_204_2 ();
 FILLER_ASAP7_75t_R FILLER_204_24 ();
 DECAPx6_ASAP7_75t_R FILLER_204_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_49 ();
 DECAPx4_ASAP7_75t_R FILLER_204_56 ();
 DECAPx4_ASAP7_75t_R FILLER_204_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_120 ();
 DECAPx10_ASAP7_75t_R FILLER_204_124 ();
 DECAPx10_ASAP7_75t_R FILLER_204_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_168 ();
 DECAPx4_ASAP7_75t_R FILLER_204_187 ();
 FILLER_ASAP7_75t_R FILLER_204_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_199 ();
 DECAPx2_ASAP7_75t_R FILLER_204_206 ();
 FILLER_ASAP7_75t_R FILLER_204_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_214 ();
 DECAPx6_ASAP7_75t_R FILLER_204_222 ();
 FILLER_ASAP7_75t_R FILLER_204_242 ();
 DECAPx2_ASAP7_75t_R FILLER_204_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_258 ();
 FILLER_ASAP7_75t_R FILLER_204_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_268 ();
 DECAPx1_ASAP7_75t_R FILLER_204_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_290 ();
 DECAPx1_ASAP7_75t_R FILLER_204_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_298 ();
 DECAPx2_ASAP7_75t_R FILLER_204_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_319 ();
 DECAPx10_ASAP7_75t_R FILLER_204_328 ();
 FILLER_ASAP7_75t_R FILLER_204_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_370 ();
 DECAPx1_ASAP7_75t_R FILLER_204_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_410 ();
 DECAPx6_ASAP7_75t_R FILLER_204_437 ();
 FILLER_ASAP7_75t_R FILLER_204_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_453 ();
 DECAPx4_ASAP7_75t_R FILLER_204_464 ();
 FILLER_ASAP7_75t_R FILLER_204_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_500 ();
 FILLER_ASAP7_75t_R FILLER_204_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_513 ();
 DECAPx2_ASAP7_75t_R FILLER_204_520 ();
 DECAPx6_ASAP7_75t_R FILLER_204_549 ();
 DECAPx1_ASAP7_75t_R FILLER_204_563 ();
 DECAPx2_ASAP7_75t_R FILLER_204_573 ();
 FILLER_ASAP7_75t_R FILLER_204_579 ();
 DECAPx2_ASAP7_75t_R FILLER_204_619 ();
 FILLER_ASAP7_75t_R FILLER_204_625 ();
 DECAPx10_ASAP7_75t_R FILLER_204_653 ();
 FILLER_ASAP7_75t_R FILLER_204_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_686 ();
 DECAPx2_ASAP7_75t_R FILLER_204_699 ();
 FILLER_ASAP7_75t_R FILLER_204_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_728 ();
 DECAPx4_ASAP7_75t_R FILLER_204_735 ();
 DECAPx2_ASAP7_75t_R FILLER_204_755 ();
 FILLER_ASAP7_75t_R FILLER_204_767 ();
 DECAPx10_ASAP7_75t_R FILLER_204_775 ();
 DECAPx6_ASAP7_75t_R FILLER_204_797 ();
 DECAPx2_ASAP7_75t_R FILLER_204_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_817 ();
 FILLER_ASAP7_75t_R FILLER_204_836 ();
 DECAPx10_ASAP7_75t_R FILLER_204_850 ();
 DECAPx2_ASAP7_75t_R FILLER_204_872 ();
 DECAPx1_ASAP7_75t_R FILLER_204_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_898 ();
 DECAPx2_ASAP7_75t_R FILLER_204_909 ();
 DECAPx4_ASAP7_75t_R FILLER_204_937 ();
 FILLER_ASAP7_75t_R FILLER_204_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_949 ();
 DECAPx2_ASAP7_75t_R FILLER_204_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_985 ();
 DECAPx4_ASAP7_75t_R FILLER_204_1000 ();
 FILLER_ASAP7_75t_R FILLER_204_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1102 ();
 DECAPx6_ASAP7_75t_R FILLER_204_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1157 ();
 FILLER_ASAP7_75t_R FILLER_204_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1178 ();
 DECAPx4_ASAP7_75t_R FILLER_204_1195 ();
 FILLER_ASAP7_75t_R FILLER_204_1205 ();
 DECAPx4_ASAP7_75t_R FILLER_204_1230 ();
 FILLER_ASAP7_75t_R FILLER_204_1240 ();
 FILLER_ASAP7_75t_R FILLER_204_1249 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1267 ();
 DECAPx6_ASAP7_75t_R FILLER_204_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1301 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1309 ();
 FILLER_ASAP7_75t_R FILLER_204_1315 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1347 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1360 ();
 FILLER_ASAP7_75t_R FILLER_204_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1373 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_205_2 ();
 DECAPx6_ASAP7_75t_R FILLER_205_27 ();
 FILLER_ASAP7_75t_R FILLER_205_41 ();
 FILLER_ASAP7_75t_R FILLER_205_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_71 ();
 DECAPx1_ASAP7_75t_R FILLER_205_87 ();
 DECAPx2_ASAP7_75t_R FILLER_205_117 ();
 FILLER_ASAP7_75t_R FILLER_205_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_125 ();
 FILLER_ASAP7_75t_R FILLER_205_136 ();
 DECAPx2_ASAP7_75t_R FILLER_205_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_166 ();
 DECAPx4_ASAP7_75t_R FILLER_205_173 ();
 DECAPx1_ASAP7_75t_R FILLER_205_227 ();
 DECAPx1_ASAP7_75t_R FILLER_205_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_259 ();
 DECAPx4_ASAP7_75t_R FILLER_205_266 ();
 FILLER_ASAP7_75t_R FILLER_205_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_278 ();
 DECAPx10_ASAP7_75t_R FILLER_205_291 ();
 DECAPx2_ASAP7_75t_R FILLER_205_313 ();
 FILLER_ASAP7_75t_R FILLER_205_319 ();
 DECAPx4_ASAP7_75t_R FILLER_205_327 ();
 FILLER_ASAP7_75t_R FILLER_205_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_339 ();
 DECAPx10_ASAP7_75t_R FILLER_205_358 ();
 DECAPx2_ASAP7_75t_R FILLER_205_380 ();
 DECAPx2_ASAP7_75t_R FILLER_205_389 ();
 FILLER_ASAP7_75t_R FILLER_205_395 ();
 DECAPx6_ASAP7_75t_R FILLER_205_415 ();
 DECAPx2_ASAP7_75t_R FILLER_205_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_453 ();
 DECAPx6_ASAP7_75t_R FILLER_205_469 ();
 DECAPx2_ASAP7_75t_R FILLER_205_483 ();
 DECAPx2_ASAP7_75t_R FILLER_205_516 ();
 FILLER_ASAP7_75t_R FILLER_205_522 ();
 FILLER_ASAP7_75t_R FILLER_205_530 ();
 DECAPx4_ASAP7_75t_R FILLER_205_540 ();
 FILLER_ASAP7_75t_R FILLER_205_550 ();
 DECAPx6_ASAP7_75t_R FILLER_205_576 ();
 FILLER_ASAP7_75t_R FILLER_205_590 ();
 DECAPx2_ASAP7_75t_R FILLER_205_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_606 ();
 DECAPx2_ASAP7_75t_R FILLER_205_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_627 ();
 DECAPx6_ASAP7_75t_R FILLER_205_652 ();
 FILLER_ASAP7_75t_R FILLER_205_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_699 ();
 DECAPx6_ASAP7_75t_R FILLER_205_707 ();
 FILLER_ASAP7_75t_R FILLER_205_721 ();
 DECAPx6_ASAP7_75t_R FILLER_205_734 ();
 FILLER_ASAP7_75t_R FILLER_205_748 ();
 FILLER_ASAP7_75t_R FILLER_205_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_768 ();
 DECAPx6_ASAP7_75t_R FILLER_205_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_789 ();
 DECAPx10_ASAP7_75t_R FILLER_205_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_822 ();
 DECAPx1_ASAP7_75t_R FILLER_205_843 ();
 DECAPx1_ASAP7_75t_R FILLER_205_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_858 ();
 DECAPx1_ASAP7_75t_R FILLER_205_888 ();
 DECAPx4_ASAP7_75t_R FILLER_205_911 ();
 FILLER_ASAP7_75t_R FILLER_205_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_968 ();
 DECAPx2_ASAP7_75t_R FILLER_205_981 ();
 FILLER_ASAP7_75t_R FILLER_205_987 ();
 FILLER_ASAP7_75t_R FILLER_205_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1020 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_205_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1127 ();
 FILLER_ASAP7_75t_R FILLER_205_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1142 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1254 ();
 FILLER_ASAP7_75t_R FILLER_205_1260 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1282 ();
 FILLER_ASAP7_75t_R FILLER_205_1296 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1308 ();
 FILLER_ASAP7_75t_R FILLER_205_1314 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1316 ();
 FILLER_ASAP7_75t_R FILLER_205_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1331 ();
 DECAPx4_ASAP7_75t_R FILLER_205_1339 ();
 FILLER_ASAP7_75t_R FILLER_205_1349 ();
 FILLER_ASAP7_75t_R FILLER_205_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_206_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_59 ();
 DECAPx6_ASAP7_75t_R FILLER_206_92 ();
 DECAPx2_ASAP7_75t_R FILLER_206_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_141 ();
 FILLER_ASAP7_75t_R FILLER_206_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_170 ();
 DECAPx4_ASAP7_75t_R FILLER_206_179 ();
 DECAPx2_ASAP7_75t_R FILLER_206_207 ();
 FILLER_ASAP7_75t_R FILLER_206_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_219 ();
 DECAPx6_ASAP7_75t_R FILLER_206_226 ();
 FILLER_ASAP7_75t_R FILLER_206_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_242 ();
 FILLER_ASAP7_75t_R FILLER_206_257 ();
 DECAPx6_ASAP7_75t_R FILLER_206_271 ();
 DECAPx1_ASAP7_75t_R FILLER_206_285 ();
 DECAPx2_ASAP7_75t_R FILLER_206_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_302 ();
 DECAPx4_ASAP7_75t_R FILLER_206_309 ();
 FILLER_ASAP7_75t_R FILLER_206_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_321 ();
 DECAPx2_ASAP7_75t_R FILLER_206_328 ();
 DECAPx4_ASAP7_75t_R FILLER_206_344 ();
 FILLER_ASAP7_75t_R FILLER_206_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_362 ();
 DECAPx2_ASAP7_75t_R FILLER_206_370 ();
 FILLER_ASAP7_75t_R FILLER_206_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_378 ();
 FILLER_ASAP7_75t_R FILLER_206_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_399 ();
 DECAPx1_ASAP7_75t_R FILLER_206_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_412 ();
 DECAPx6_ASAP7_75t_R FILLER_206_425 ();
 DECAPx1_ASAP7_75t_R FILLER_206_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_443 ();
 DECAPx4_ASAP7_75t_R FILLER_206_452 ();
 DECAPx2_ASAP7_75t_R FILLER_206_470 ();
 FILLER_ASAP7_75t_R FILLER_206_476 ();
 DECAPx10_ASAP7_75t_R FILLER_206_484 ();
 FILLER_ASAP7_75t_R FILLER_206_516 ();
 FILLER_ASAP7_75t_R FILLER_206_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_534 ();
 FILLER_ASAP7_75t_R FILLER_206_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_545 ();
 DECAPx2_ASAP7_75t_R FILLER_206_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_584 ();
 DECAPx1_ASAP7_75t_R FILLER_206_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_592 ();
 DECAPx6_ASAP7_75t_R FILLER_206_599 ();
 DECAPx6_ASAP7_75t_R FILLER_206_639 ();
 DECAPx1_ASAP7_75t_R FILLER_206_653 ();
 FILLER_ASAP7_75t_R FILLER_206_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_685 ();
 DECAPx1_ASAP7_75t_R FILLER_206_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_696 ();
 DECAPx4_ASAP7_75t_R FILLER_206_710 ();
 DECAPx4_ASAP7_75t_R FILLER_206_739 ();
 FILLER_ASAP7_75t_R FILLER_206_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_757 ();
 FILLER_ASAP7_75t_R FILLER_206_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_775 ();
 FILLER_ASAP7_75t_R FILLER_206_784 ();
 DECAPx10_ASAP7_75t_R FILLER_206_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_818 ();
 FILLER_ASAP7_75t_R FILLER_206_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_838 ();
 FILLER_ASAP7_75t_R FILLER_206_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_847 ();
 DECAPx1_ASAP7_75t_R FILLER_206_866 ();
 FILLER_ASAP7_75t_R FILLER_206_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_881 ();
 DECAPx4_ASAP7_75t_R FILLER_206_889 ();
 FILLER_ASAP7_75t_R FILLER_206_899 ();
 DECAPx10_ASAP7_75t_R FILLER_206_907 ();
 DECAPx4_ASAP7_75t_R FILLER_206_929 ();
 FILLER_ASAP7_75t_R FILLER_206_939 ();
 DECAPx4_ASAP7_75t_R FILLER_206_951 ();
 FILLER_ASAP7_75t_R FILLER_206_961 ();
 DECAPx4_ASAP7_75t_R FILLER_206_991 ();
 FILLER_ASAP7_75t_R FILLER_206_1001 ();
 DECAPx6_ASAP7_75t_R FILLER_206_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1020 ();
 FILLER_ASAP7_75t_R FILLER_206_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1035 ();
 FILLER_ASAP7_75t_R FILLER_206_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1041 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1050 ();
 FILLER_ASAP7_75t_R FILLER_206_1060 ();
 FILLER_ASAP7_75t_R FILLER_206_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1143 ();
 FILLER_ASAP7_75t_R FILLER_206_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1173 ();
 FILLER_ASAP7_75t_R FILLER_206_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1209 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1232 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1255 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1264 ();
 FILLER_ASAP7_75t_R FILLER_206_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1309 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1313 ();
 FILLER_ASAP7_75t_R FILLER_206_1324 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1338 ();
 FILLER_ASAP7_75t_R FILLER_206_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1346 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1373 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_207_2 ();
 DECAPx6_ASAP7_75t_R FILLER_207_24 ();
 DECAPx1_ASAP7_75t_R FILLER_207_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_57 ();
 DECAPx2_ASAP7_75t_R FILLER_207_61 ();
 FILLER_ASAP7_75t_R FILLER_207_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_69 ();
 DECAPx1_ASAP7_75t_R FILLER_207_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_80 ();
 DECAPx6_ASAP7_75t_R FILLER_207_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_98 ();
 DECAPx10_ASAP7_75t_R FILLER_207_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_128 ();
 FILLER_ASAP7_75t_R FILLER_207_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_134 ();
 DECAPx2_ASAP7_75t_R FILLER_207_149 ();
 FILLER_ASAP7_75t_R FILLER_207_155 ();
 FILLER_ASAP7_75t_R FILLER_207_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_162 ();
 DECAPx2_ASAP7_75t_R FILLER_207_173 ();
 FILLER_ASAP7_75t_R FILLER_207_179 ();
 DECAPx4_ASAP7_75t_R FILLER_207_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_216 ();
 DECAPx2_ASAP7_75t_R FILLER_207_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_229 ();
 DECAPx2_ASAP7_75t_R FILLER_207_244 ();
 FILLER_ASAP7_75t_R FILLER_207_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_252 ();
 DECAPx2_ASAP7_75t_R FILLER_207_265 ();
 FILLER_ASAP7_75t_R FILLER_207_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_285 ();
 DECAPx1_ASAP7_75t_R FILLER_207_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_298 ();
 DECAPx2_ASAP7_75t_R FILLER_207_306 ();
 DECAPx2_ASAP7_75t_R FILLER_207_319 ();
 FILLER_ASAP7_75t_R FILLER_207_325 ();
 DECAPx2_ASAP7_75t_R FILLER_207_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_343 ();
 FILLER_ASAP7_75t_R FILLER_207_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_360 ();
 DECAPx6_ASAP7_75t_R FILLER_207_369 ();
 DECAPx2_ASAP7_75t_R FILLER_207_383 ();
 DECAPx4_ASAP7_75t_R FILLER_207_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_405 ();
 DECAPx2_ASAP7_75t_R FILLER_207_412 ();
 DECAPx4_ASAP7_75t_R FILLER_207_426 ();
 FILLER_ASAP7_75t_R FILLER_207_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_464 ();
 FILLER_ASAP7_75t_R FILLER_207_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_481 ();
 DECAPx1_ASAP7_75t_R FILLER_207_499 ();
 DECAPx2_ASAP7_75t_R FILLER_207_517 ();
 FILLER_ASAP7_75t_R FILLER_207_523 ();
 DECAPx10_ASAP7_75t_R FILLER_207_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_553 ();
 FILLER_ASAP7_75t_R FILLER_207_562 ();
 DECAPx2_ASAP7_75t_R FILLER_207_602 ();
 FILLER_ASAP7_75t_R FILLER_207_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_613 ();
 DECAPx2_ASAP7_75t_R FILLER_207_620 ();
 FILLER_ASAP7_75t_R FILLER_207_626 ();
 DECAPx10_ASAP7_75t_R FILLER_207_631 ();
 DECAPx10_ASAP7_75t_R FILLER_207_653 ();
 DECAPx1_ASAP7_75t_R FILLER_207_675 ();
 DECAPx10_ASAP7_75t_R FILLER_207_687 ();
 DECAPx2_ASAP7_75t_R FILLER_207_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_715 ();
 DECAPx4_ASAP7_75t_R FILLER_207_744 ();
 FILLER_ASAP7_75t_R FILLER_207_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_756 ();
 DECAPx10_ASAP7_75t_R FILLER_207_786 ();
 DECAPx10_ASAP7_75t_R FILLER_207_808 ();
 DECAPx4_ASAP7_75t_R FILLER_207_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_852 ();
 FILLER_ASAP7_75t_R FILLER_207_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_861 ();
 DECAPx6_ASAP7_75t_R FILLER_207_869 ();
 FILLER_ASAP7_75t_R FILLER_207_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_901 ();
 DECAPx1_ASAP7_75t_R FILLER_207_909 ();
 FILLER_ASAP7_75t_R FILLER_207_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_923 ();
 FILLER_ASAP7_75t_R FILLER_207_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_935 ();
 FILLER_ASAP7_75t_R FILLER_207_943 ();
 DECAPx6_ASAP7_75t_R FILLER_207_953 ();
 DECAPx2_ASAP7_75t_R FILLER_207_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_973 ();
 DECAPx10_ASAP7_75t_R FILLER_207_980 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1002 ();
 FILLER_ASAP7_75t_R FILLER_207_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_207_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1050 ();
 FILLER_ASAP7_75t_R FILLER_207_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1138 ();
 DECAPx4_ASAP7_75t_R FILLER_207_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1208 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1245 ();
 FILLER_ASAP7_75t_R FILLER_207_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1286 ();
 DECAPx4_ASAP7_75t_R FILLER_207_1311 ();
 FILLER_ASAP7_75t_R FILLER_207_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1323 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1330 ();
 FILLER_ASAP7_75t_R FILLER_207_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1346 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_208_2 ();
 FILLER_ASAP7_75t_R FILLER_208_24 ();
 DECAPx10_ASAP7_75t_R FILLER_208_56 ();
 DECAPx4_ASAP7_75t_R FILLER_208_78 ();
 FILLER_ASAP7_75t_R FILLER_208_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_90 ();
 FILLER_ASAP7_75t_R FILLER_208_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_119 ();
 DECAPx2_ASAP7_75t_R FILLER_208_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_132 ();
 FILLER_ASAP7_75t_R FILLER_208_166 ();
 DECAPx6_ASAP7_75t_R FILLER_208_176 ();
 DECAPx2_ASAP7_75t_R FILLER_208_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_196 ();
 FILLER_ASAP7_75t_R FILLER_208_209 ();
 DECAPx1_ASAP7_75t_R FILLER_208_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_244 ();
 FILLER_ASAP7_75t_R FILLER_208_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_253 ();
 DECAPx2_ASAP7_75t_R FILLER_208_287 ();
 FILLER_ASAP7_75t_R FILLER_208_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_295 ();
 DECAPx2_ASAP7_75t_R FILLER_208_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_310 ();
 DECAPx2_ASAP7_75t_R FILLER_208_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_361 ();
 DECAPx2_ASAP7_75t_R FILLER_208_368 ();
 FILLER_ASAP7_75t_R FILLER_208_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_376 ();
 FILLER_ASAP7_75t_R FILLER_208_391 ();
 DECAPx4_ASAP7_75t_R FILLER_208_400 ();
 FILLER_ASAP7_75t_R FILLER_208_410 ();
 DECAPx4_ASAP7_75t_R FILLER_208_421 ();
 FILLER_ASAP7_75t_R FILLER_208_431 ();
 DECAPx2_ASAP7_75t_R FILLER_208_441 ();
 DECAPx2_ASAP7_75t_R FILLER_208_456 ();
 FILLER_ASAP7_75t_R FILLER_208_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_466 ();
 DECAPx10_ASAP7_75t_R FILLER_208_491 ();
 DECAPx1_ASAP7_75t_R FILLER_208_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_517 ();
 DECAPx2_ASAP7_75t_R FILLER_208_530 ();
 FILLER_ASAP7_75t_R FILLER_208_536 ();
 DECAPx6_ASAP7_75t_R FILLER_208_546 ();
 DECAPx2_ASAP7_75t_R FILLER_208_560 ();
 FILLER_ASAP7_75t_R FILLER_208_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_581 ();
 DECAPx1_ASAP7_75t_R FILLER_208_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_592 ();
 DECAPx2_ASAP7_75t_R FILLER_208_619 ();
 FILLER_ASAP7_75t_R FILLER_208_625 ();
 DECAPx10_ASAP7_75t_R FILLER_208_634 ();
 DECAPx6_ASAP7_75t_R FILLER_208_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_670 ();
 DECAPx10_ASAP7_75t_R FILLER_208_681 ();
 FILLER_ASAP7_75t_R FILLER_208_703 ();
 DECAPx2_ASAP7_75t_R FILLER_208_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_722 ();
 FILLER_ASAP7_75t_R FILLER_208_737 ();
 FILLER_ASAP7_75t_R FILLER_208_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_773 ();
 FILLER_ASAP7_75t_R FILLER_208_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_790 ();
 DECAPx6_ASAP7_75t_R FILLER_208_801 ();
 DECAPx2_ASAP7_75t_R FILLER_208_815 ();
 DECAPx10_ASAP7_75t_R FILLER_208_833 ();
 DECAPx4_ASAP7_75t_R FILLER_208_855 ();
 FILLER_ASAP7_75t_R FILLER_208_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_880 ();
 FILLER_ASAP7_75t_R FILLER_208_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_901 ();
 FILLER_ASAP7_75t_R FILLER_208_945 ();
 FILLER_ASAP7_75t_R FILLER_208_961 ();
 FILLER_ASAP7_75t_R FILLER_208_973 ();
 DECAPx4_ASAP7_75t_R FILLER_208_986 ();
 FILLER_ASAP7_75t_R FILLER_208_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_998 ();
 DECAPx1_ASAP7_75t_R FILLER_208_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1071 ();
 FILLER_ASAP7_75t_R FILLER_208_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1109 ();
 FILLER_ASAP7_75t_R FILLER_208_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_208_1125 ();
 DECAPx4_ASAP7_75t_R FILLER_208_1155 ();
 FILLER_ASAP7_75t_R FILLER_208_1165 ();
 FILLER_ASAP7_75t_R FILLER_208_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1181 ();
 FILLER_ASAP7_75t_R FILLER_208_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_208_1220 ();
 FILLER_ASAP7_75t_R FILLER_208_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1233 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1285 ();
 FILLER_ASAP7_75t_R FILLER_208_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_208_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1370 ();
 DECAPx1_ASAP7_75t_R FILLER_208_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_209_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_41 ();
 DECAPx6_ASAP7_75t_R FILLER_209_48 ();
 DECAPx1_ASAP7_75t_R FILLER_209_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_66 ();
 DECAPx2_ASAP7_75t_R FILLER_209_93 ();
 FILLER_ASAP7_75t_R FILLER_209_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_108 ();
 FILLER_ASAP7_75t_R FILLER_209_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_137 ();
 DECAPx4_ASAP7_75t_R FILLER_209_171 ();
 FILLER_ASAP7_75t_R FILLER_209_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_183 ();
 DECAPx1_ASAP7_75t_R FILLER_209_190 ();
 DECAPx1_ASAP7_75t_R FILLER_209_226 ();
 DECAPx1_ASAP7_75t_R FILLER_209_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_240 ();
 DECAPx4_ASAP7_75t_R FILLER_209_247 ();
 DECAPx4_ASAP7_75t_R FILLER_209_271 ();
 DECAPx2_ASAP7_75t_R FILLER_209_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_307 ();
 DECAPx1_ASAP7_75t_R FILLER_209_322 ();
 DECAPx6_ASAP7_75t_R FILLER_209_335 ();
 DECAPx2_ASAP7_75t_R FILLER_209_394 ();
 FILLER_ASAP7_75t_R FILLER_209_400 ();
 DECAPx4_ASAP7_75t_R FILLER_209_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_451 ();
 DECAPx4_ASAP7_75t_R FILLER_209_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_472 ();
 DECAPx1_ASAP7_75t_R FILLER_209_483 ();
 FILLER_ASAP7_75t_R FILLER_209_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_561 ();
 DECAPx2_ASAP7_75t_R FILLER_209_572 ();
 FILLER_ASAP7_75t_R FILLER_209_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_580 ();
 DECAPx2_ASAP7_75t_R FILLER_209_607 ();
 DECAPx1_ASAP7_75t_R FILLER_209_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_621 ();
 DECAPx10_ASAP7_75t_R FILLER_209_654 ();
 DECAPx1_ASAP7_75t_R FILLER_209_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_680 ();
 DECAPx1_ASAP7_75t_R FILLER_209_709 ();
 FILLER_ASAP7_75t_R FILLER_209_721 ();
 DECAPx1_ASAP7_75t_R FILLER_209_729 ();
 DECAPx6_ASAP7_75t_R FILLER_209_739 ();
 FILLER_ASAP7_75t_R FILLER_209_753 ();
 DECAPx2_ASAP7_75t_R FILLER_209_761 ();
 FILLER_ASAP7_75t_R FILLER_209_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_769 ();
 DECAPx2_ASAP7_75t_R FILLER_209_782 ();
 FILLER_ASAP7_75t_R FILLER_209_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_790 ();
 DECAPx4_ASAP7_75t_R FILLER_209_801 ();
 FILLER_ASAP7_75t_R FILLER_209_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_850 ();
 DECAPx6_ASAP7_75t_R FILLER_209_858 ();
 DECAPx1_ASAP7_75t_R FILLER_209_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_904 ();
 DECAPx1_ASAP7_75t_R FILLER_209_920 ();
 DECAPx6_ASAP7_75t_R FILLER_209_926 ();
 DECAPx2_ASAP7_75t_R FILLER_209_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_946 ();
 DECAPx6_ASAP7_75t_R FILLER_209_954 ();
 DECAPx1_ASAP7_75t_R FILLER_209_968 ();
 DECAPx2_ASAP7_75t_R FILLER_209_1005 ();
 FILLER_ASAP7_75t_R FILLER_209_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1013 ();
 DECAPx4_ASAP7_75t_R FILLER_209_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1077 ();
 FILLER_ASAP7_75t_R FILLER_209_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_209_1092 ();
 FILLER_ASAP7_75t_R FILLER_209_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1100 ();
 DECAPx4_ASAP7_75t_R FILLER_209_1107 ();
 FILLER_ASAP7_75t_R FILLER_209_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1119 ();
 FILLER_ASAP7_75t_R FILLER_209_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_209_1174 ();
 FILLER_ASAP7_75t_R FILLER_209_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1194 ();
 FILLER_ASAP7_75t_R FILLER_209_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1211 ();
 DECAPx1_ASAP7_75t_R FILLER_209_1225 ();
 FILLER_ASAP7_75t_R FILLER_209_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_209_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1271 ();
 FILLER_ASAP7_75t_R FILLER_209_1275 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1280 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1294 ();
 DECAPx4_ASAP7_75t_R FILLER_209_1302 ();
 DECAPx4_ASAP7_75t_R FILLER_209_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1391 ();
 DECAPx6_ASAP7_75t_R FILLER_210_2 ();
 DECAPx1_ASAP7_75t_R FILLER_210_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_20 ();
 DECAPx1_ASAP7_75t_R FILLER_210_32 ();
 DECAPx1_ASAP7_75t_R FILLER_210_40 ();
 DECAPx2_ASAP7_75t_R FILLER_210_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_65 ();
 FILLER_ASAP7_75t_R FILLER_210_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_80 ();
 FILLER_ASAP7_75t_R FILLER_210_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_86 ();
 DECAPx2_ASAP7_75t_R FILLER_210_96 ();
 FILLER_ASAP7_75t_R FILLER_210_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_108 ();
 DECAPx1_ASAP7_75t_R FILLER_210_155 ();
 FILLER_ASAP7_75t_R FILLER_210_162 ();
 DECAPx2_ASAP7_75t_R FILLER_210_170 ();
 FILLER_ASAP7_75t_R FILLER_210_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_178 ();
 DECAPx1_ASAP7_75t_R FILLER_210_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_197 ();
 DECAPx1_ASAP7_75t_R FILLER_210_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_208 ();
 DECAPx10_ASAP7_75t_R FILLER_210_212 ();
 DECAPx2_ASAP7_75t_R FILLER_210_234 ();
 DECAPx1_ASAP7_75t_R FILLER_210_252 ();
 DECAPx6_ASAP7_75t_R FILLER_210_262 ();
 FILLER_ASAP7_75t_R FILLER_210_276 ();
 DECAPx1_ASAP7_75t_R FILLER_210_292 ();
 DECAPx2_ASAP7_75t_R FILLER_210_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_310 ();
 DECAPx2_ASAP7_75t_R FILLER_210_317 ();
 FILLER_ASAP7_75t_R FILLER_210_323 ();
 DECAPx2_ASAP7_75t_R FILLER_210_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_339 ();
 DECAPx2_ASAP7_75t_R FILLER_210_350 ();
 FILLER_ASAP7_75t_R FILLER_210_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_358 ();
 DECAPx2_ASAP7_75t_R FILLER_210_399 ();
 DECAPx2_ASAP7_75t_R FILLER_210_421 ();
 DECAPx4_ASAP7_75t_R FILLER_210_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_451 ();
 DECAPx1_ASAP7_75t_R FILLER_210_458 ();
 FILLER_ASAP7_75t_R FILLER_210_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_466 ();
 DECAPx6_ASAP7_75t_R FILLER_210_477 ();
 DECAPx1_ASAP7_75t_R FILLER_210_491 ();
 DECAPx2_ASAP7_75t_R FILLER_210_513 ();
 DECAPx2_ASAP7_75t_R FILLER_210_529 ();
 DECAPx1_ASAP7_75t_R FILLER_210_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_560 ();
 DECAPx6_ASAP7_75t_R FILLER_210_569 ();
 DECAPx2_ASAP7_75t_R FILLER_210_589 ();
 FILLER_ASAP7_75t_R FILLER_210_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_600 ();
 DECAPx2_ASAP7_75t_R FILLER_210_605 ();
 FILLER_ASAP7_75t_R FILLER_210_611 ();
 DECAPx4_ASAP7_75t_R FILLER_210_657 ();
 FILLER_ASAP7_75t_R FILLER_210_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_669 ();
 FILLER_ASAP7_75t_R FILLER_210_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_698 ();
 DECAPx2_ASAP7_75t_R FILLER_210_724 ();
 FILLER_ASAP7_75t_R FILLER_210_730 ();
 FILLER_ASAP7_75t_R FILLER_210_740 ();
 DECAPx2_ASAP7_75t_R FILLER_210_745 ();
 FILLER_ASAP7_75t_R FILLER_210_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_753 ();
 DECAPx2_ASAP7_75t_R FILLER_210_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_776 ();
 FILLER_ASAP7_75t_R FILLER_210_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_789 ();
 DECAPx6_ASAP7_75t_R FILLER_210_800 ();
 DECAPx1_ASAP7_75t_R FILLER_210_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_818 ();
 DECAPx2_ASAP7_75t_R FILLER_210_840 ();
 FILLER_ASAP7_75t_R FILLER_210_846 ();
 DECAPx1_ASAP7_75t_R FILLER_210_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_864 ();
 DECAPx10_ASAP7_75t_R FILLER_210_875 ();
 DECAPx2_ASAP7_75t_R FILLER_210_897 ();
 DECAPx4_ASAP7_75t_R FILLER_210_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_919 ();
 DECAPx2_ASAP7_75t_R FILLER_210_934 ();
 DECAPx6_ASAP7_75t_R FILLER_210_953 ();
 FILLER_ASAP7_75t_R FILLER_210_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_969 ();
 FILLER_ASAP7_75t_R FILLER_210_978 ();
 FILLER_ASAP7_75t_R FILLER_210_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1036 ();
 FILLER_ASAP7_75t_R FILLER_210_1055 ();
 FILLER_ASAP7_75t_R FILLER_210_1072 ();
 FILLER_ASAP7_75t_R FILLER_210_1112 ();
 DECAPx6_ASAP7_75t_R FILLER_210_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1140 ();
 FILLER_ASAP7_75t_R FILLER_210_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1159 ();
 DECAPx4_ASAP7_75t_R FILLER_210_1173 ();
 FILLER_ASAP7_75t_R FILLER_210_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1227 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1297 ();
 FILLER_ASAP7_75t_R FILLER_210_1303 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1311 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1324 ();
 FILLER_ASAP7_75t_R FILLER_210_1330 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1332 ();
 DECAPx6_ASAP7_75t_R FILLER_210_1336 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1350 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1354 ();
 FILLER_ASAP7_75t_R FILLER_210_1358 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_211_2 ();
 DECAPx6_ASAP7_75t_R FILLER_211_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_38 ();
 FILLER_ASAP7_75t_R FILLER_211_73 ();
 DECAPx1_ASAP7_75t_R FILLER_211_127 ();
 DECAPx4_ASAP7_75t_R FILLER_211_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_165 ();
 DECAPx2_ASAP7_75t_R FILLER_211_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_178 ();
 DECAPx1_ASAP7_75t_R FILLER_211_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_218 ();
 FILLER_ASAP7_75t_R FILLER_211_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_227 ();
 DECAPx4_ASAP7_75t_R FILLER_211_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_244 ();
 DECAPx1_ASAP7_75t_R FILLER_211_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_255 ();
 DECAPx4_ASAP7_75t_R FILLER_211_262 ();
 DECAPx2_ASAP7_75t_R FILLER_211_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_292 ();
 DECAPx6_ASAP7_75t_R FILLER_211_307 ();
 DECAPx2_ASAP7_75t_R FILLER_211_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_327 ();
 DECAPx10_ASAP7_75t_R FILLER_211_334 ();
 FILLER_ASAP7_75t_R FILLER_211_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_358 ();
 DECAPx2_ASAP7_75t_R FILLER_211_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_387 ();
 FILLER_ASAP7_75t_R FILLER_211_396 ();
 DECAPx4_ASAP7_75t_R FILLER_211_412 ();
 DECAPx2_ASAP7_75t_R FILLER_211_432 ();
 DECAPx4_ASAP7_75t_R FILLER_211_444 ();
 FILLER_ASAP7_75t_R FILLER_211_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_456 ();
 DECAPx1_ASAP7_75t_R FILLER_211_475 ();
 DECAPx10_ASAP7_75t_R FILLER_211_485 ();
 DECAPx10_ASAP7_75t_R FILLER_211_507 ();
 DECAPx2_ASAP7_75t_R FILLER_211_529 ();
 FILLER_ASAP7_75t_R FILLER_211_535 ();
 FILLER_ASAP7_75t_R FILLER_211_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_554 ();
 DECAPx4_ASAP7_75t_R FILLER_211_567 ();
 DECAPx6_ASAP7_75t_R FILLER_211_603 ();
 DECAPx2_ASAP7_75t_R FILLER_211_617 ();
 DECAPx2_ASAP7_75t_R FILLER_211_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_642 ();
 DECAPx10_ASAP7_75t_R FILLER_211_649 ();
 DECAPx2_ASAP7_75t_R FILLER_211_671 ();
 FILLER_ASAP7_75t_R FILLER_211_677 ();
 DECAPx2_ASAP7_75t_R FILLER_211_695 ();
 DECAPx4_ASAP7_75t_R FILLER_211_721 ();
 FILLER_ASAP7_75t_R FILLER_211_731 ();
 DECAPx2_ASAP7_75t_R FILLER_211_741 ();
 FILLER_ASAP7_75t_R FILLER_211_747 ();
 DECAPx10_ASAP7_75t_R FILLER_211_764 ();
 DECAPx1_ASAP7_75t_R FILLER_211_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_790 ();
 DECAPx10_ASAP7_75t_R FILLER_211_801 ();
 DECAPx6_ASAP7_75t_R FILLER_211_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_837 ();
 FILLER_ASAP7_75t_R FILLER_211_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_848 ();
 DECAPx6_ASAP7_75t_R FILLER_211_857 ();
 DECAPx1_ASAP7_75t_R FILLER_211_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_875 ();
 DECAPx1_ASAP7_75t_R FILLER_211_888 ();
 FILLER_ASAP7_75t_R FILLER_211_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_912 ();
 DECAPx4_ASAP7_75t_R FILLER_211_926 ();
 FILLER_ASAP7_75t_R FILLER_211_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_938 ();
 DECAPx2_ASAP7_75t_R FILLER_211_954 ();
 DECAPx10_ASAP7_75t_R FILLER_211_978 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1000 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1021 ();
 FILLER_ASAP7_75t_R FILLER_211_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_211_1077 ();
 FILLER_ASAP7_75t_R FILLER_211_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1096 ();
 FILLER_ASAP7_75t_R FILLER_211_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_211_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1186 ();
 DECAPx1_ASAP7_75t_R FILLER_211_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1256 ();
 FILLER_ASAP7_75t_R FILLER_211_1278 ();
 FILLER_ASAP7_75t_R FILLER_211_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1292 ();
 DECAPx1_ASAP7_75t_R FILLER_211_1296 ();
 DECAPx4_ASAP7_75t_R FILLER_211_1317 ();
 FILLER_ASAP7_75t_R FILLER_211_1327 ();
 DECAPx4_ASAP7_75t_R FILLER_211_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1367 ();
 DECAPx10_ASAP7_75t_R FILLER_212_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_24 ();
 FILLER_ASAP7_75t_R FILLER_212_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_53 ();
 DECAPx4_ASAP7_75t_R FILLER_212_60 ();
 DECAPx2_ASAP7_75t_R FILLER_212_74 ();
 FILLER_ASAP7_75t_R FILLER_212_80 ();
 DECAPx1_ASAP7_75t_R FILLER_212_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_92 ();
 DECAPx2_ASAP7_75t_R FILLER_212_96 ();
 FILLER_ASAP7_75t_R FILLER_212_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_104 ();
 DECAPx1_ASAP7_75t_R FILLER_212_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_115 ();
 DECAPx4_ASAP7_75t_R FILLER_212_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_129 ();
 DECAPx2_ASAP7_75t_R FILLER_212_140 ();
 FILLER_ASAP7_75t_R FILLER_212_146 ();
 DECAPx4_ASAP7_75t_R FILLER_212_151 ();
 DECAPx6_ASAP7_75t_R FILLER_212_187 ();
 FILLER_ASAP7_75t_R FILLER_212_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_203 ();
 FILLER_ASAP7_75t_R FILLER_212_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_246 ();
 FILLER_ASAP7_75t_R FILLER_212_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_275 ();
 DECAPx6_ASAP7_75t_R FILLER_212_290 ();
 DECAPx1_ASAP7_75t_R FILLER_212_304 ();
 FILLER_ASAP7_75t_R FILLER_212_323 ();
 DECAPx1_ASAP7_75t_R FILLER_212_347 ();
 DECAPx6_ASAP7_75t_R FILLER_212_357 ();
 FILLER_ASAP7_75t_R FILLER_212_371 ();
 DECAPx10_ASAP7_75t_R FILLER_212_384 ();
 DECAPx2_ASAP7_75t_R FILLER_212_406 ();
 FILLER_ASAP7_75t_R FILLER_212_412 ();
 DECAPx6_ASAP7_75t_R FILLER_212_420 ();
 FILLER_ASAP7_75t_R FILLER_212_434 ();
 FILLER_ASAP7_75t_R FILLER_212_442 ();
 DECAPx4_ASAP7_75t_R FILLER_212_450 ();
 FILLER_ASAP7_75t_R FILLER_212_460 ();
 DECAPx2_ASAP7_75t_R FILLER_212_464 ();
 FILLER_ASAP7_75t_R FILLER_212_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_472 ();
 FILLER_ASAP7_75t_R FILLER_212_489 ();
 DECAPx4_ASAP7_75t_R FILLER_212_509 ();
 DECAPx6_ASAP7_75t_R FILLER_212_529 ();
 DECAPx1_ASAP7_75t_R FILLER_212_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_547 ();
 DECAPx2_ASAP7_75t_R FILLER_212_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_576 ();
 FILLER_ASAP7_75t_R FILLER_212_589 ();
 DECAPx10_ASAP7_75t_R FILLER_212_623 ();
 DECAPx6_ASAP7_75t_R FILLER_212_659 ();
 DECAPx1_ASAP7_75t_R FILLER_212_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_677 ();
 DECAPx6_ASAP7_75t_R FILLER_212_686 ();
 DECAPx1_ASAP7_75t_R FILLER_212_700 ();
 DECAPx4_ASAP7_75t_R FILLER_212_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_726 ();
 DECAPx1_ASAP7_75t_R FILLER_212_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_749 ();
 DECAPx10_ASAP7_75t_R FILLER_212_764 ();
 DECAPx1_ASAP7_75t_R FILLER_212_786 ();
 DECAPx2_ASAP7_75t_R FILLER_212_796 ();
 FILLER_ASAP7_75t_R FILLER_212_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_841 ();
 FILLER_ASAP7_75t_R FILLER_212_860 ();
 FILLER_ASAP7_75t_R FILLER_212_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_883 ();
 DECAPx1_ASAP7_75t_R FILLER_212_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_915 ();
 DECAPx1_ASAP7_75t_R FILLER_212_933 ();
 DECAPx6_ASAP7_75t_R FILLER_212_954 ();
 FILLER_ASAP7_75t_R FILLER_212_988 ();
 FILLER_ASAP7_75t_R FILLER_212_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1043 ();
 FILLER_ASAP7_75t_R FILLER_212_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1055 ();
 FILLER_ASAP7_75t_R FILLER_212_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1102 ();
 FILLER_ASAP7_75t_R FILLER_212_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1126 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1134 ();
 FILLER_ASAP7_75t_R FILLER_212_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_212_1145 ();
 FILLER_ASAP7_75t_R FILLER_212_1155 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1166 ();
 FILLER_ASAP7_75t_R FILLER_212_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1192 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1211 ();
 FILLER_ASAP7_75t_R FILLER_212_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1224 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1228 ();
 FILLER_ASAP7_75t_R FILLER_212_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1280 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1294 ();
 FILLER_ASAP7_75t_R FILLER_212_1323 ();
 FILLER_ASAP7_75t_R FILLER_212_1341 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1367 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_213_2 ();
 DECAPx2_ASAP7_75t_R FILLER_213_16 ();
 FILLER_ASAP7_75t_R FILLER_213_38 ();
 DECAPx10_ASAP7_75t_R FILLER_213_43 ();
 FILLER_ASAP7_75t_R FILLER_213_65 ();
 FILLER_ASAP7_75t_R FILLER_213_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_77 ();
 DECAPx6_ASAP7_75t_R FILLER_213_81 ();
 DECAPx6_ASAP7_75t_R FILLER_213_98 ();
 FILLER_ASAP7_75t_R FILLER_213_112 ();
 DECAPx1_ASAP7_75t_R FILLER_213_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_132 ();
 DECAPx2_ASAP7_75t_R FILLER_213_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_145 ();
 DECAPx6_ASAP7_75t_R FILLER_213_149 ();
 FILLER_ASAP7_75t_R FILLER_213_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_165 ();
 DECAPx10_ASAP7_75t_R FILLER_213_181 ();
 DECAPx6_ASAP7_75t_R FILLER_213_203 ();
 FILLER_ASAP7_75t_R FILLER_213_217 ();
 DECAPx4_ASAP7_75t_R FILLER_213_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_232 ();
 FILLER_ASAP7_75t_R FILLER_213_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_241 ();
 FILLER_ASAP7_75t_R FILLER_213_268 ();
 DECAPx1_ASAP7_75t_R FILLER_213_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_286 ();
 DECAPx4_ASAP7_75t_R FILLER_213_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_303 ();
 DECAPx2_ASAP7_75t_R FILLER_213_310 ();
 FILLER_ASAP7_75t_R FILLER_213_316 ();
 FILLER_ASAP7_75t_R FILLER_213_338 ();
 DECAPx10_ASAP7_75t_R FILLER_213_356 ();
 DECAPx6_ASAP7_75t_R FILLER_213_378 ();
 DECAPx4_ASAP7_75t_R FILLER_213_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_408 ();
 DECAPx2_ASAP7_75t_R FILLER_213_429 ();
 FILLER_ASAP7_75t_R FILLER_213_435 ();
 DECAPx2_ASAP7_75t_R FILLER_213_451 ();
 DECAPx4_ASAP7_75t_R FILLER_213_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_477 ();
 FILLER_ASAP7_75t_R FILLER_213_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_511 ();
 FILLER_ASAP7_75t_R FILLER_213_529 ();
 FILLER_ASAP7_75t_R FILLER_213_541 ();
 DECAPx2_ASAP7_75t_R FILLER_213_555 ();
 FILLER_ASAP7_75t_R FILLER_213_561 ();
 DECAPx10_ASAP7_75t_R FILLER_213_569 ();
 DECAPx1_ASAP7_75t_R FILLER_213_594 ();
 DECAPx1_ASAP7_75t_R FILLER_213_604 ();
 DECAPx1_ASAP7_75t_R FILLER_213_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_647 ();
 DECAPx2_ASAP7_75t_R FILLER_213_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_691 ();
 DECAPx1_ASAP7_75t_R FILLER_213_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_709 ();
 DECAPx1_ASAP7_75t_R FILLER_213_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_727 ();
 DECAPx1_ASAP7_75t_R FILLER_213_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_749 ();
 DECAPx2_ASAP7_75t_R FILLER_213_767 ();
 FILLER_ASAP7_75t_R FILLER_213_773 ();
 DECAPx4_ASAP7_75t_R FILLER_213_798 ();
 FILLER_ASAP7_75t_R FILLER_213_808 ();
 DECAPx4_ASAP7_75t_R FILLER_213_826 ();
 DECAPx6_ASAP7_75t_R FILLER_213_849 ();
 FILLER_ASAP7_75t_R FILLER_213_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_865 ();
 FILLER_ASAP7_75t_R FILLER_213_872 ();
 DECAPx1_ASAP7_75t_R FILLER_213_882 ();
 DECAPx1_ASAP7_75t_R FILLER_213_906 ();
 DECAPx2_ASAP7_75t_R FILLER_213_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_926 ();
 FILLER_ASAP7_75t_R FILLER_213_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_945 ();
 DECAPx6_ASAP7_75t_R FILLER_213_966 ();
 FILLER_ASAP7_75t_R FILLER_213_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1019 ();
 DECAPx4_ASAP7_75t_R FILLER_213_1051 ();
 FILLER_ASAP7_75t_R FILLER_213_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1063 ();
 DECAPx6_ASAP7_75t_R FILLER_213_1074 ();
 FILLER_ASAP7_75t_R FILLER_213_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1116 ();
 FILLER_ASAP7_75t_R FILLER_213_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1156 ();
 FILLER_ASAP7_75t_R FILLER_213_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1188 ();
 FILLER_ASAP7_75t_R FILLER_213_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1200 ();
 DECAPx6_ASAP7_75t_R FILLER_213_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1243 ();
 DECAPx6_ASAP7_75t_R FILLER_213_1250 ();
 FILLER_ASAP7_75t_R FILLER_213_1264 ();
 DECAPx4_ASAP7_75t_R FILLER_213_1269 ();
 FILLER_ASAP7_75t_R FILLER_213_1282 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1287 ();
 FILLER_ASAP7_75t_R FILLER_213_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1295 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1309 ();
 DECAPx6_ASAP7_75t_R FILLER_213_1317 ();
 DECAPx4_ASAP7_75t_R FILLER_213_1337 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1367 ();
 DECAPx2_ASAP7_75t_R FILLER_214_2 ();
 DECAPx4_ASAP7_75t_R FILLER_214_34 ();
 FILLER_ASAP7_75t_R FILLER_214_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_46 ();
 DECAPx2_ASAP7_75t_R FILLER_214_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_95 ();
 DECAPx2_ASAP7_75t_R FILLER_214_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_157 ();
 FILLER_ASAP7_75t_R FILLER_214_168 ();
 FILLER_ASAP7_75t_R FILLER_214_184 ();
 FILLER_ASAP7_75t_R FILLER_214_201 ();
 DECAPx2_ASAP7_75t_R FILLER_214_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_215 ();
 DECAPx6_ASAP7_75t_R FILLER_214_236 ();
 DECAPx1_ASAP7_75t_R FILLER_214_250 ();
 DECAPx2_ASAP7_75t_R FILLER_214_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_271 ();
 DECAPx4_ASAP7_75t_R FILLER_214_278 ();
 FILLER_ASAP7_75t_R FILLER_214_288 ();
 FILLER_ASAP7_75t_R FILLER_214_303 ();
 DECAPx6_ASAP7_75t_R FILLER_214_319 ();
 FILLER_ASAP7_75t_R FILLER_214_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_335 ();
 DECAPx1_ASAP7_75t_R FILLER_214_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_371 ();
 DECAPx1_ASAP7_75t_R FILLER_214_379 ();
 DECAPx2_ASAP7_75t_R FILLER_214_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_410 ();
 DECAPx4_ASAP7_75t_R FILLER_214_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_451 ();
 DECAPx2_ASAP7_75t_R FILLER_214_464 ();
 FILLER_ASAP7_75t_R FILLER_214_470 ();
 FILLER_ASAP7_75t_R FILLER_214_513 ();
 DECAPx2_ASAP7_75t_R FILLER_214_531 ();
 DECAPx1_ASAP7_75t_R FILLER_214_555 ();
 DECAPx6_ASAP7_75t_R FILLER_214_569 ();
 FILLER_ASAP7_75t_R FILLER_214_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_585 ();
 DECAPx10_ASAP7_75t_R FILLER_214_592 ();
 DECAPx1_ASAP7_75t_R FILLER_214_614 ();
 FILLER_ASAP7_75t_R FILLER_214_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_627 ();
 DECAPx10_ASAP7_75t_R FILLER_214_637 ();
 DECAPx4_ASAP7_75t_R FILLER_214_659 ();
 DECAPx1_ASAP7_75t_R FILLER_214_685 ();
 DECAPx1_ASAP7_75t_R FILLER_214_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_712 ();
 DECAPx2_ASAP7_75t_R FILLER_214_721 ();
 FILLER_ASAP7_75t_R FILLER_214_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_729 ();
 FILLER_ASAP7_75t_R FILLER_214_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_746 ();
 DECAPx1_ASAP7_75t_R FILLER_214_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_771 ();
 DECAPx2_ASAP7_75t_R FILLER_214_806 ();
 DECAPx4_ASAP7_75t_R FILLER_214_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_830 ();
 DECAPx2_ASAP7_75t_R FILLER_214_854 ();
 DECAPx1_ASAP7_75t_R FILLER_214_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_870 ();
 DECAPx2_ASAP7_75t_R FILLER_214_887 ();
 FILLER_ASAP7_75t_R FILLER_214_893 ();
 DECAPx4_ASAP7_75t_R FILLER_214_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_937 ();
 DECAPx6_ASAP7_75t_R FILLER_214_950 ();
 DECAPx10_ASAP7_75t_R FILLER_214_984 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1076 ();
 FILLER_ASAP7_75t_R FILLER_214_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1091 ();
 DECAPx6_ASAP7_75t_R FILLER_214_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_214_1143 ();
 FILLER_ASAP7_75t_R FILLER_214_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1171 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1214 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1222 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1258 ();
 FILLER_ASAP7_75t_R FILLER_214_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1289 ();
 DECAPx6_ASAP7_75t_R FILLER_214_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1332 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1342 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1346 ();
 FILLER_ASAP7_75t_R FILLER_214_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1361 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_215_2 ();
 DECAPx2_ASAP7_75t_R FILLER_215_16 ();
 DECAPx2_ASAP7_75t_R FILLER_215_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_74 ();
 FILLER_ASAP7_75t_R FILLER_215_107 ();
 DECAPx4_ASAP7_75t_R FILLER_215_112 ();
 DECAPx1_ASAP7_75t_R FILLER_215_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_129 ();
 DECAPx2_ASAP7_75t_R FILLER_215_136 ();
 FILLER_ASAP7_75t_R FILLER_215_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_144 ();
 DECAPx4_ASAP7_75t_R FILLER_215_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_181 ();
 DECAPx4_ASAP7_75t_R FILLER_215_214 ();
 DECAPx2_ASAP7_75t_R FILLER_215_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_238 ();
 DECAPx10_ASAP7_75t_R FILLER_215_246 ();
 DECAPx1_ASAP7_75t_R FILLER_215_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_272 ();
 DECAPx6_ASAP7_75t_R FILLER_215_281 ();
 DECAPx4_ASAP7_75t_R FILLER_215_315 ();
 FILLER_ASAP7_75t_R FILLER_215_325 ();
 DECAPx4_ASAP7_75t_R FILLER_215_334 ();
 FILLER_ASAP7_75t_R FILLER_215_344 ();
 FILLER_ASAP7_75t_R FILLER_215_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_370 ();
 FILLER_ASAP7_75t_R FILLER_215_382 ();
 FILLER_ASAP7_75t_R FILLER_215_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_398 ();
 FILLER_ASAP7_75t_R FILLER_215_413 ();
 DECAPx6_ASAP7_75t_R FILLER_215_422 ();
 DECAPx1_ASAP7_75t_R FILLER_215_436 ();
 DECAPx2_ASAP7_75t_R FILLER_215_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_454 ();
 DECAPx10_ASAP7_75t_R FILLER_215_461 ();
 FILLER_ASAP7_75t_R FILLER_215_483 ();
 FILLER_ASAP7_75t_R FILLER_215_491 ();
 DECAPx6_ASAP7_75t_R FILLER_215_499 ();
 FILLER_ASAP7_75t_R FILLER_215_513 ();
 DECAPx1_ASAP7_75t_R FILLER_215_522 ();
 DECAPx1_ASAP7_75t_R FILLER_215_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_536 ();
 DECAPx2_ASAP7_75t_R FILLER_215_545 ();
 FILLER_ASAP7_75t_R FILLER_215_551 ();
 FILLER_ASAP7_75t_R FILLER_215_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_567 ();
 DECAPx1_ASAP7_75t_R FILLER_215_574 ();
 DECAPx6_ASAP7_75t_R FILLER_215_610 ();
 DECAPx1_ASAP7_75t_R FILLER_215_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_628 ();
 DECAPx4_ASAP7_75t_R FILLER_215_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_668 ();
 DECAPx6_ASAP7_75t_R FILLER_215_692 ();
 DECAPx4_ASAP7_75t_R FILLER_215_716 ();
 FILLER_ASAP7_75t_R FILLER_215_726 ();
 DECAPx4_ASAP7_75t_R FILLER_215_740 ();
 FILLER_ASAP7_75t_R FILLER_215_750 ();
 DECAPx2_ASAP7_75t_R FILLER_215_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_772 ();
 FILLER_ASAP7_75t_R FILLER_215_779 ();
 DECAPx6_ASAP7_75t_R FILLER_215_799 ();
 FILLER_ASAP7_75t_R FILLER_215_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_822 ();
 DECAPx6_ASAP7_75t_R FILLER_215_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_861 ();
 DECAPx2_ASAP7_75t_R FILLER_215_880 ();
 FILLER_ASAP7_75t_R FILLER_215_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_888 ();
 DECAPx2_ASAP7_75t_R FILLER_215_897 ();
 FILLER_ASAP7_75t_R FILLER_215_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_905 ();
 FILLER_ASAP7_75t_R FILLER_215_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_914 ();
 FILLER_ASAP7_75t_R FILLER_215_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_923 ();
 DECAPx6_ASAP7_75t_R FILLER_215_926 ();
 DECAPx1_ASAP7_75t_R FILLER_215_940 ();
 DECAPx4_ASAP7_75t_R FILLER_215_951 ();
 DECAPx4_ASAP7_75t_R FILLER_215_967 ();
 FILLER_ASAP7_75t_R FILLER_215_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_985 ();
 DECAPx6_ASAP7_75t_R FILLER_215_996 ();
 DECAPx6_ASAP7_75t_R FILLER_215_1036 ();
 FILLER_ASAP7_75t_R FILLER_215_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1062 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1073 ();
 FILLER_ASAP7_75t_R FILLER_215_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_215_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1097 ();
 FILLER_ASAP7_75t_R FILLER_215_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_215_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_215_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1195 ();
 FILLER_ASAP7_75t_R FILLER_215_1211 ();
 FILLER_ASAP7_75t_R FILLER_215_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1222 ();
 DECAPx4_ASAP7_75t_R FILLER_215_1233 ();
 FILLER_ASAP7_75t_R FILLER_215_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1245 ();
 DECAPx4_ASAP7_75t_R FILLER_215_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1272 ();
 FILLER_ASAP7_75t_R FILLER_215_1278 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_215_1310 ();
 FILLER_ASAP7_75t_R FILLER_215_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1343 ();
 DECAPx10_ASAP7_75t_R FILLER_216_2 ();
 DECAPx1_ASAP7_75t_R FILLER_216_50 ();
 DECAPx6_ASAP7_75t_R FILLER_216_63 ();
 FILLER_ASAP7_75t_R FILLER_216_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_79 ();
 DECAPx2_ASAP7_75t_R FILLER_216_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_92 ();
 DECAPx6_ASAP7_75t_R FILLER_216_99 ();
 DECAPx2_ASAP7_75t_R FILLER_216_119 ();
 FILLER_ASAP7_75t_R FILLER_216_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_127 ();
 DECAPx4_ASAP7_75t_R FILLER_216_134 ();
 FILLER_ASAP7_75t_R FILLER_216_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_146 ();
 DECAPx6_ASAP7_75t_R FILLER_216_163 ();
 DECAPx1_ASAP7_75t_R FILLER_216_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_187 ();
 DECAPx4_ASAP7_75t_R FILLER_216_206 ();
 FILLER_ASAP7_75t_R FILLER_216_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_218 ();
 FILLER_ASAP7_75t_R FILLER_216_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_241 ();
 FILLER_ASAP7_75t_R FILLER_216_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_254 ();
 FILLER_ASAP7_75t_R FILLER_216_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_275 ();
 FILLER_ASAP7_75t_R FILLER_216_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_286 ();
 FILLER_ASAP7_75t_R FILLER_216_299 ();
 DECAPx6_ASAP7_75t_R FILLER_216_309 ();
 DECAPx1_ASAP7_75t_R FILLER_216_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_327 ();
 DECAPx4_ASAP7_75t_R FILLER_216_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_348 ();
 DECAPx2_ASAP7_75t_R FILLER_216_356 ();
 DECAPx6_ASAP7_75t_R FILLER_216_388 ();
 FILLER_ASAP7_75t_R FILLER_216_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_404 ();
 DECAPx1_ASAP7_75t_R FILLER_216_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_426 ();
 FILLER_ASAP7_75t_R FILLER_216_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_435 ();
 DECAPx1_ASAP7_75t_R FILLER_216_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_461 ();
 DECAPx4_ASAP7_75t_R FILLER_216_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_474 ();
 DECAPx2_ASAP7_75t_R FILLER_216_501 ();
 FILLER_ASAP7_75t_R FILLER_216_519 ();
 DECAPx4_ASAP7_75t_R FILLER_216_527 ();
 FILLER_ASAP7_75t_R FILLER_216_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_539 ();
 DECAPx1_ASAP7_75t_R FILLER_216_546 ();
 FILLER_ASAP7_75t_R FILLER_216_566 ();
 DECAPx1_ASAP7_75t_R FILLER_216_594 ();
 FILLER_ASAP7_75t_R FILLER_216_601 ();
 DECAPx1_ASAP7_75t_R FILLER_216_609 ();
 DECAPx4_ASAP7_75t_R FILLER_216_657 ();
 DECAPx6_ASAP7_75t_R FILLER_216_693 ();
 DECAPx1_ASAP7_75t_R FILLER_216_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_717 ();
 DECAPx2_ASAP7_75t_R FILLER_216_728 ();
 DECAPx2_ASAP7_75t_R FILLER_216_746 ();
 FILLER_ASAP7_75t_R FILLER_216_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_754 ();
 DECAPx2_ASAP7_75t_R FILLER_216_765 ();
 FILLER_ASAP7_75t_R FILLER_216_771 ();
 DECAPx4_ASAP7_75t_R FILLER_216_779 ();
 FILLER_ASAP7_75t_R FILLER_216_789 ();
 DECAPx10_ASAP7_75t_R FILLER_216_803 ();
 DECAPx6_ASAP7_75t_R FILLER_216_825 ();
 DECAPx1_ASAP7_75t_R FILLER_216_839 ();
 DECAPx6_ASAP7_75t_R FILLER_216_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_873 ();
 DECAPx4_ASAP7_75t_R FILLER_216_902 ();
 FILLER_ASAP7_75t_R FILLER_216_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_914 ();
 DECAPx6_ASAP7_75t_R FILLER_216_925 ();
 DECAPx1_ASAP7_75t_R FILLER_216_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_943 ();
 DECAPx6_ASAP7_75t_R FILLER_216_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_965 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1002 ();
 FILLER_ASAP7_75t_R FILLER_216_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1017 ();
 FILLER_ASAP7_75t_R FILLER_216_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1028 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1063 ();
 FILLER_ASAP7_75t_R FILLER_216_1074 ();
 FILLER_ASAP7_75t_R FILLER_216_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1107 ();
 FILLER_ASAP7_75t_R FILLER_216_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1167 ();
 DECAPx4_ASAP7_75t_R FILLER_216_1180 ();
 FILLER_ASAP7_75t_R FILLER_216_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1192 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1203 ();
 DECAPx6_ASAP7_75t_R FILLER_216_1210 ();
 FILLER_ASAP7_75t_R FILLER_216_1224 ();
 DECAPx6_ASAP7_75t_R FILLER_216_1239 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1253 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1272 ();
 DECAPx4_ASAP7_75t_R FILLER_216_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1298 ();
 DECAPx4_ASAP7_75t_R FILLER_216_1305 ();
 FILLER_ASAP7_75t_R FILLER_216_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1353 ();
 FILLER_ASAP7_75t_R FILLER_216_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_217_2 ();
 DECAPx2_ASAP7_75t_R FILLER_217_16 ();
 DECAPx1_ASAP7_75t_R FILLER_217_34 ();
 DECAPx6_ASAP7_75t_R FILLER_217_41 ();
 DECAPx1_ASAP7_75t_R FILLER_217_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_59 ();
 DECAPx2_ASAP7_75t_R FILLER_217_66 ();
 FILLER_ASAP7_75t_R FILLER_217_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_80 ();
 DECAPx2_ASAP7_75t_R FILLER_217_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_90 ();
 FILLER_ASAP7_75t_R FILLER_217_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_101 ();
 DECAPx1_ASAP7_75t_R FILLER_217_105 ();
 FILLER_ASAP7_75t_R FILLER_217_149 ();
 DECAPx2_ASAP7_75t_R FILLER_217_165 ();
 FILLER_ASAP7_75t_R FILLER_217_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_173 ();
 DECAPx4_ASAP7_75t_R FILLER_217_202 ();
 DECAPx1_ASAP7_75t_R FILLER_217_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_228 ();
 DECAPx4_ASAP7_75t_R FILLER_217_237 ();
 FILLER_ASAP7_75t_R FILLER_217_247 ();
 DECAPx4_ASAP7_75t_R FILLER_217_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_273 ();
 FILLER_ASAP7_75t_R FILLER_217_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_282 ();
 FILLER_ASAP7_75t_R FILLER_217_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_299 ();
 DECAPx6_ASAP7_75t_R FILLER_217_306 ();
 DECAPx1_ASAP7_75t_R FILLER_217_326 ();
 DECAPx2_ASAP7_75t_R FILLER_217_340 ();
 FILLER_ASAP7_75t_R FILLER_217_346 ();
 DECAPx10_ASAP7_75t_R FILLER_217_354 ();
 DECAPx1_ASAP7_75t_R FILLER_217_376 ();
 DECAPx1_ASAP7_75t_R FILLER_217_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_393 ();
 DECAPx10_ASAP7_75t_R FILLER_217_400 ();
 FILLER_ASAP7_75t_R FILLER_217_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_439 ();
 DECAPx1_ASAP7_75t_R FILLER_217_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_452 ();
 DECAPx10_ASAP7_75t_R FILLER_217_459 ();
 DECAPx4_ASAP7_75t_R FILLER_217_481 ();
 DECAPx6_ASAP7_75t_R FILLER_217_515 ();
 DECAPx1_ASAP7_75t_R FILLER_217_529 ();
 DECAPx6_ASAP7_75t_R FILLER_217_539 ();
 DECAPx2_ASAP7_75t_R FILLER_217_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_581 ();
 DECAPx6_ASAP7_75t_R FILLER_217_585 ();
 FILLER_ASAP7_75t_R FILLER_217_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_601 ();
 FILLER_ASAP7_75t_R FILLER_217_628 ();
 DECAPx4_ASAP7_75t_R FILLER_217_643 ();
 FILLER_ASAP7_75t_R FILLER_217_653 ();
 DECAPx6_ASAP7_75t_R FILLER_217_658 ();
 DECAPx1_ASAP7_75t_R FILLER_217_692 ();
 DECAPx4_ASAP7_75t_R FILLER_217_708 ();
 FILLER_ASAP7_75t_R FILLER_217_718 ();
 DECAPx10_ASAP7_75t_R FILLER_217_757 ();
 DECAPx2_ASAP7_75t_R FILLER_217_779 ();
 FILLER_ASAP7_75t_R FILLER_217_785 ();
 DECAPx10_ASAP7_75t_R FILLER_217_790 ();
 DECAPx2_ASAP7_75t_R FILLER_217_812 ();
 FILLER_ASAP7_75t_R FILLER_217_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_820 ();
 FILLER_ASAP7_75t_R FILLER_217_839 ();
 DECAPx2_ASAP7_75t_R FILLER_217_853 ();
 FILLER_ASAP7_75t_R FILLER_217_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_861 ();
 DECAPx1_ASAP7_75t_R FILLER_217_876 ();
 DECAPx2_ASAP7_75t_R FILLER_217_894 ();
 FILLER_ASAP7_75t_R FILLER_217_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_902 ();
 DECAPx6_ASAP7_75t_R FILLER_217_910 ();
 DECAPx1_ASAP7_75t_R FILLER_217_926 ();
 FILLER_ASAP7_75t_R FILLER_217_938 ();
 DECAPx10_ASAP7_75t_R FILLER_217_960 ();
 DECAPx2_ASAP7_75t_R FILLER_217_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_988 ();
 DECAPx4_ASAP7_75t_R FILLER_217_1017 ();
 FILLER_ASAP7_75t_R FILLER_217_1027 ();
 FILLER_ASAP7_75t_R FILLER_217_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1064 ();
 DECAPx6_ASAP7_75t_R FILLER_217_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_217_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1121 ();
 DECAPx4_ASAP7_75t_R FILLER_217_1125 ();
 FILLER_ASAP7_75t_R FILLER_217_1153 ();
 DECAPx4_ASAP7_75t_R FILLER_217_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1224 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1249 ();
 DECAPx4_ASAP7_75t_R FILLER_217_1265 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1316 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1320 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1327 ();
 FILLER_ASAP7_75t_R FILLER_217_1333 ();
 FILLER_ASAP7_75t_R FILLER_217_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1385 ();
 FILLER_ASAP7_75t_R FILLER_218_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_35 ();
 DECAPx2_ASAP7_75t_R FILLER_218_114 ();
 FILLER_ASAP7_75t_R FILLER_218_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_122 ();
 DECAPx6_ASAP7_75t_R FILLER_218_126 ();
 DECAPx2_ASAP7_75t_R FILLER_218_140 ();
 DECAPx4_ASAP7_75t_R FILLER_218_172 ();
 FILLER_ASAP7_75t_R FILLER_218_182 ();
 DECAPx2_ASAP7_75t_R FILLER_218_202 ();
 DECAPx1_ASAP7_75t_R FILLER_218_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_218 ();
 DECAPx10_ASAP7_75t_R FILLER_218_227 ();
 FILLER_ASAP7_75t_R FILLER_218_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_267 ();
 DECAPx2_ASAP7_75t_R FILLER_218_288 ();
 DECAPx2_ASAP7_75t_R FILLER_218_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_316 ();
 FILLER_ASAP7_75t_R FILLER_218_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_330 ();
 FILLER_ASAP7_75t_R FILLER_218_343 ();
 DECAPx1_ASAP7_75t_R FILLER_218_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_363 ();
 DECAPx2_ASAP7_75t_R FILLER_218_380 ();
 FILLER_ASAP7_75t_R FILLER_218_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_388 ();
 DECAPx6_ASAP7_75t_R FILLER_218_411 ();
 DECAPx2_ASAP7_75t_R FILLER_218_431 ();
 FILLER_ASAP7_75t_R FILLER_218_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_439 ();
 DECAPx6_ASAP7_75t_R FILLER_218_446 ();
 FILLER_ASAP7_75t_R FILLER_218_460 ();
 DECAPx1_ASAP7_75t_R FILLER_218_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_468 ();
 FILLER_ASAP7_75t_R FILLER_218_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_489 ();
 DECAPx4_ASAP7_75t_R FILLER_218_496 ();
 FILLER_ASAP7_75t_R FILLER_218_506 ();
 DECAPx2_ASAP7_75t_R FILLER_218_514 ();
 DECAPx1_ASAP7_75t_R FILLER_218_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_530 ();
 DECAPx10_ASAP7_75t_R FILLER_218_557 ();
 DECAPx2_ASAP7_75t_R FILLER_218_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_585 ();
 DECAPx4_ASAP7_75t_R FILLER_218_592 ();
 DECAPx1_ASAP7_75t_R FILLER_218_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_612 ();
 DECAPx1_ASAP7_75t_R FILLER_218_622 ();
 DECAPx2_ASAP7_75t_R FILLER_218_632 ();
 FILLER_ASAP7_75t_R FILLER_218_638 ();
 DECAPx6_ASAP7_75t_R FILLER_218_666 ();
 FILLER_ASAP7_75t_R FILLER_218_680 ();
 DECAPx6_ASAP7_75t_R FILLER_218_688 ();
 DECAPx1_ASAP7_75t_R FILLER_218_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_716 ();
 DECAPx1_ASAP7_75t_R FILLER_218_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_767 ();
 FILLER_ASAP7_75t_R FILLER_218_790 ();
 FILLER_ASAP7_75t_R FILLER_218_818 ();
 DECAPx2_ASAP7_75t_R FILLER_218_838 ();
 DECAPx4_ASAP7_75t_R FILLER_218_854 ();
 DECAPx2_ASAP7_75t_R FILLER_218_872 ();
 FILLER_ASAP7_75t_R FILLER_218_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_880 ();
 DECAPx1_ASAP7_75t_R FILLER_218_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_908 ();
 FILLER_ASAP7_75t_R FILLER_218_916 ();
 DECAPx6_ASAP7_75t_R FILLER_218_928 ();
 FILLER_ASAP7_75t_R FILLER_218_942 ();
 FILLER_ASAP7_75t_R FILLER_218_956 ();
 FILLER_ASAP7_75t_R FILLER_218_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_972 ();
 DECAPx1_ASAP7_75t_R FILLER_218_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_995 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1110 ();
 FILLER_ASAP7_75t_R FILLER_218_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1120 ();
 DECAPx4_ASAP7_75t_R FILLER_218_1127 ();
 FILLER_ASAP7_75t_R FILLER_218_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1151 ();
 FILLER_ASAP7_75t_R FILLER_218_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1186 ();
 FILLER_ASAP7_75t_R FILLER_218_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1194 ();
 FILLER_ASAP7_75t_R FILLER_218_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1211 ();
 DECAPx4_ASAP7_75t_R FILLER_218_1218 ();
 FILLER_ASAP7_75t_R FILLER_218_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1230 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1267 ();
 FILLER_ASAP7_75t_R FILLER_218_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1281 ();
 FILLER_ASAP7_75t_R FILLER_218_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1308 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1330 ();
 FILLER_ASAP7_75t_R FILLER_218_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1338 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1354 ();
 FILLER_ASAP7_75t_R FILLER_218_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_219_2 ();
 DECAPx1_ASAP7_75t_R FILLER_219_16 ();
 DECAPx2_ASAP7_75t_R FILLER_219_31 ();
 FILLER_ASAP7_75t_R FILLER_219_37 ();
 DECAPx2_ASAP7_75t_R FILLER_219_42 ();
 FILLER_ASAP7_75t_R FILLER_219_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_50 ();
 FILLER_ASAP7_75t_R FILLER_219_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_63 ();
 DECAPx10_ASAP7_75t_R FILLER_219_78 ();
 DECAPx2_ASAP7_75t_R FILLER_219_100 ();
 FILLER_ASAP7_75t_R FILLER_219_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_108 ();
 DECAPx1_ASAP7_75t_R FILLER_219_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_119 ();
 DECAPx1_ASAP7_75t_R FILLER_219_123 ();
 DECAPx4_ASAP7_75t_R FILLER_219_133 ();
 DECAPx4_ASAP7_75t_R FILLER_219_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_159 ();
 DECAPx10_ASAP7_75t_R FILLER_219_163 ();
 DECAPx10_ASAP7_75t_R FILLER_219_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_207 ();
 DECAPx1_ASAP7_75t_R FILLER_219_242 ();
 DECAPx6_ASAP7_75t_R FILLER_219_266 ();
 DECAPx4_ASAP7_75t_R FILLER_219_286 ();
 DECAPx4_ASAP7_75t_R FILLER_219_308 ();
 FILLER_ASAP7_75t_R FILLER_219_324 ();
 DECAPx4_ASAP7_75t_R FILLER_219_332 ();
 FILLER_ASAP7_75t_R FILLER_219_342 ();
 FILLER_ASAP7_75t_R FILLER_219_358 ();
 DECAPx1_ASAP7_75t_R FILLER_219_368 ();
 DECAPx2_ASAP7_75t_R FILLER_219_382 ();
 FILLER_ASAP7_75t_R FILLER_219_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_402 ();
 DECAPx1_ASAP7_75t_R FILLER_219_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_439 ();
 FILLER_ASAP7_75t_R FILLER_219_446 ();
 DECAPx2_ASAP7_75t_R FILLER_219_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_462 ();
 DECAPx2_ASAP7_75t_R FILLER_219_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_487 ();
 DECAPx4_ASAP7_75t_R FILLER_219_494 ();
 FILLER_ASAP7_75t_R FILLER_219_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_506 ();
 DECAPx2_ASAP7_75t_R FILLER_219_513 ();
 FILLER_ASAP7_75t_R FILLER_219_519 ();
 DECAPx1_ASAP7_75t_R FILLER_219_528 ();
 DECAPx2_ASAP7_75t_R FILLER_219_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_544 ();
 FILLER_ASAP7_75t_R FILLER_219_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_550 ();
 DECAPx4_ASAP7_75t_R FILLER_219_557 ();
 FILLER_ASAP7_75t_R FILLER_219_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_569 ();
 FILLER_ASAP7_75t_R FILLER_219_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_578 ();
 DECAPx10_ASAP7_75t_R FILLER_219_637 ();
 DECAPx10_ASAP7_75t_R FILLER_219_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_681 ();
 DECAPx4_ASAP7_75t_R FILLER_219_688 ();
 FILLER_ASAP7_75t_R FILLER_219_698 ();
 DECAPx1_ASAP7_75t_R FILLER_219_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_753 ();
 FILLER_ASAP7_75t_R FILLER_219_766 ();
 DECAPx2_ASAP7_75t_R FILLER_219_797 ();
 FILLER_ASAP7_75t_R FILLER_219_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_809 ();
 DECAPx2_ASAP7_75t_R FILLER_219_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_819 ();
 DECAPx4_ASAP7_75t_R FILLER_219_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_848 ();
 DECAPx2_ASAP7_75t_R FILLER_219_859 ();
 DECAPx1_ASAP7_75t_R FILLER_219_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_880 ();
 DECAPx1_ASAP7_75t_R FILLER_219_895 ();
 DECAPx1_ASAP7_75t_R FILLER_219_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_923 ();
 FILLER_ASAP7_75t_R FILLER_219_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_928 ();
 FILLER_ASAP7_75t_R FILLER_219_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_951 ();
 DECAPx2_ASAP7_75t_R FILLER_219_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_964 ();
 DECAPx10_ASAP7_75t_R FILLER_219_975 ();
 DECAPx1_ASAP7_75t_R FILLER_219_997 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1014 ();
 FILLER_ASAP7_75t_R FILLER_219_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1036 ();
 FILLER_ASAP7_75t_R FILLER_219_1058 ();
 FILLER_ASAP7_75t_R FILLER_219_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_219_1091 ();
 FILLER_ASAP7_75t_R FILLER_219_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1130 ();
 FILLER_ASAP7_75t_R FILLER_219_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1163 ();
 FILLER_ASAP7_75t_R FILLER_219_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1171 ();
 FILLER_ASAP7_75t_R FILLER_219_1182 ();
 FILLER_ASAP7_75t_R FILLER_219_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1192 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1219 ();
 FILLER_ASAP7_75t_R FILLER_219_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1252 ();
 DECAPx4_ASAP7_75t_R FILLER_219_1285 ();
 FILLER_ASAP7_75t_R FILLER_219_1295 ();
 FILLER_ASAP7_75t_R FILLER_219_1309 ();
 DECAPx6_ASAP7_75t_R FILLER_219_1343 ();
 FILLER_ASAP7_75t_R FILLER_219_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1359 ();
 DECAPx2_ASAP7_75t_R FILLER_220_2 ();
 FILLER_ASAP7_75t_R FILLER_220_8 ();
 DECAPx2_ASAP7_75t_R FILLER_220_42 ();
 FILLER_ASAP7_75t_R FILLER_220_48 ();
 DECAPx6_ASAP7_75t_R FILLER_220_79 ();
 DECAPx2_ASAP7_75t_R FILLER_220_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_99 ();
 DECAPx2_ASAP7_75t_R FILLER_220_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_168 ();
 DECAPx6_ASAP7_75t_R FILLER_220_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_201 ();
 DECAPx2_ASAP7_75t_R FILLER_220_222 ();
 DECAPx4_ASAP7_75t_R FILLER_220_234 ();
 FILLER_ASAP7_75t_R FILLER_220_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_253 ();
 DECAPx2_ASAP7_75t_R FILLER_220_260 ();
 DECAPx4_ASAP7_75t_R FILLER_220_274 ();
 FILLER_ASAP7_75t_R FILLER_220_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_304 ();
 DECAPx1_ASAP7_75t_R FILLER_220_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_355 ();
 FILLER_ASAP7_75t_R FILLER_220_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_364 ();
 DECAPx4_ASAP7_75t_R FILLER_220_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_387 ();
 DECAPx10_ASAP7_75t_R FILLER_220_400 ();
 DECAPx1_ASAP7_75t_R FILLER_220_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_432 ();
 DECAPx2_ASAP7_75t_R FILLER_220_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_461 ();
 FILLER_ASAP7_75t_R FILLER_220_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_466 ();
 DECAPx2_ASAP7_75t_R FILLER_220_473 ();
 FILLER_ASAP7_75t_R FILLER_220_479 ();
 FILLER_ASAP7_75t_R FILLER_220_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_520 ();
 DECAPx1_ASAP7_75t_R FILLER_220_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_531 ();
 DECAPx1_ASAP7_75t_R FILLER_220_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_546 ();
 DECAPx2_ASAP7_75t_R FILLER_220_556 ();
 FILLER_ASAP7_75t_R FILLER_220_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_564 ();
 FILLER_ASAP7_75t_R FILLER_220_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_599 ();
 DECAPx2_ASAP7_75t_R FILLER_220_603 ();
 FILLER_ASAP7_75t_R FILLER_220_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_611 ();
 DECAPx1_ASAP7_75t_R FILLER_220_619 ();
 DECAPx6_ASAP7_75t_R FILLER_220_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_701 ();
 DECAPx2_ASAP7_75t_R FILLER_220_718 ();
 DECAPx1_ASAP7_75t_R FILLER_220_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_750 ();
 DECAPx1_ASAP7_75t_R FILLER_220_761 ();
 FILLER_ASAP7_75t_R FILLER_220_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_777 ();
 DECAPx6_ASAP7_75t_R FILLER_220_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_808 ();
 DECAPx10_ASAP7_75t_R FILLER_220_812 ();
 DECAPx2_ASAP7_75t_R FILLER_220_834 ();
 FILLER_ASAP7_75t_R FILLER_220_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_842 ();
 FILLER_ASAP7_75t_R FILLER_220_875 ();
 DECAPx10_ASAP7_75t_R FILLER_220_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_915 ();
 DECAPx2_ASAP7_75t_R FILLER_220_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_942 ();
 DECAPx6_ASAP7_75t_R FILLER_220_960 ();
 DECAPx1_ASAP7_75t_R FILLER_220_974 ();
 DECAPx4_ASAP7_75t_R FILLER_220_1010 ();
 FILLER_ASAP7_75t_R FILLER_220_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_220_1028 ();
 FILLER_ASAP7_75t_R FILLER_220_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1110 ();
 FILLER_ASAP7_75t_R FILLER_220_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1118 ();
 DECAPx4_ASAP7_75t_R FILLER_220_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1171 ();
 FILLER_ASAP7_75t_R FILLER_220_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1231 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1268 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1277 ();
 FILLER_ASAP7_75t_R FILLER_220_1283 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1295 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1302 ();
 FILLER_ASAP7_75t_R FILLER_220_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1310 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1347 ();
 DECAPx6_ASAP7_75t_R FILLER_220_1354 ();
 FILLER_ASAP7_75t_R FILLER_220_1368 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_221_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_24 ();
 FILLER_ASAP7_75t_R FILLER_221_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_38 ();
 DECAPx2_ASAP7_75t_R FILLER_221_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_54 ();
 DECAPx2_ASAP7_75t_R FILLER_221_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_71 ();
 DECAPx1_ASAP7_75t_R FILLER_221_78 ();
 DECAPx4_ASAP7_75t_R FILLER_221_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_124 ();
 DECAPx2_ASAP7_75t_R FILLER_221_131 ();
 FILLER_ASAP7_75t_R FILLER_221_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_145 ();
 DECAPx4_ASAP7_75t_R FILLER_221_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_159 ();
 DECAPx4_ASAP7_75t_R FILLER_221_170 ();
 FILLER_ASAP7_75t_R FILLER_221_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_202 ();
 DECAPx1_ASAP7_75t_R FILLER_221_213 ();
 FILLER_ASAP7_75t_R FILLER_221_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_225 ();
 DECAPx4_ASAP7_75t_R FILLER_221_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_250 ();
 DECAPx2_ASAP7_75t_R FILLER_221_259 ();
 FILLER_ASAP7_75t_R FILLER_221_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_267 ();
 DECAPx2_ASAP7_75t_R FILLER_221_282 ();
 DECAPx2_ASAP7_75t_R FILLER_221_306 ();
 FILLER_ASAP7_75t_R FILLER_221_312 ();
 DECAPx10_ASAP7_75t_R FILLER_221_323 ();
 DECAPx1_ASAP7_75t_R FILLER_221_345 ();
 DECAPx10_ASAP7_75t_R FILLER_221_355 ();
 DECAPx10_ASAP7_75t_R FILLER_221_390 ();
 DECAPx2_ASAP7_75t_R FILLER_221_412 ();
 FILLER_ASAP7_75t_R FILLER_221_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_420 ();
 FILLER_ASAP7_75t_R FILLER_221_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_455 ();
 DECAPx2_ASAP7_75t_R FILLER_221_478 ();
 FILLER_ASAP7_75t_R FILLER_221_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_549 ();
 DECAPx2_ASAP7_75t_R FILLER_221_576 ();
 FILLER_ASAP7_75t_R FILLER_221_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_584 ();
 FILLER_ASAP7_75t_R FILLER_221_588 ();
 DECAPx2_ASAP7_75t_R FILLER_221_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_600 ();
 FILLER_ASAP7_75t_R FILLER_221_605 ();
 DECAPx4_ASAP7_75t_R FILLER_221_613 ();
 FILLER_ASAP7_75t_R FILLER_221_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_625 ();
 DECAPx4_ASAP7_75t_R FILLER_221_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_643 ();
 DECAPx2_ASAP7_75t_R FILLER_221_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_653 ();
 DECAPx4_ASAP7_75t_R FILLER_221_687 ();
 FILLER_ASAP7_75t_R FILLER_221_697 ();
 DECAPx2_ASAP7_75t_R FILLER_221_709 ();
 FILLER_ASAP7_75t_R FILLER_221_715 ();
 DECAPx4_ASAP7_75t_R FILLER_221_740 ();
 FILLER_ASAP7_75t_R FILLER_221_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_752 ();
 DECAPx2_ASAP7_75t_R FILLER_221_756 ();
 FILLER_ASAP7_75t_R FILLER_221_762 ();
 DECAPx2_ASAP7_75t_R FILLER_221_774 ();
 FILLER_ASAP7_75t_R FILLER_221_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_782 ();
 DECAPx2_ASAP7_75t_R FILLER_221_816 ();
 DECAPx10_ASAP7_75t_R FILLER_221_840 ();
 DECAPx4_ASAP7_75t_R FILLER_221_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_872 ();
 DECAPx6_ASAP7_75t_R FILLER_221_892 ();
 DECAPx4_ASAP7_75t_R FILLER_221_912 ();
 FILLER_ASAP7_75t_R FILLER_221_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_926 ();
 FILLER_ASAP7_75t_R FILLER_221_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_956 ();
 DECAPx2_ASAP7_75t_R FILLER_221_968 ();
 FILLER_ASAP7_75t_R FILLER_221_990 ();
 DECAPx2_ASAP7_75t_R FILLER_221_995 ();
 FILLER_ASAP7_75t_R FILLER_221_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1003 ();
 FILLER_ASAP7_75t_R FILLER_221_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1015 ();
 FILLER_ASAP7_75t_R FILLER_221_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1026 ();
 FILLER_ASAP7_75t_R FILLER_221_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1038 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1065 ();
 FILLER_ASAP7_75t_R FILLER_221_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1086 ();
 FILLER_ASAP7_75t_R FILLER_221_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1097 ();
 DECAPx4_ASAP7_75t_R FILLER_221_1108 ();
 FILLER_ASAP7_75t_R FILLER_221_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1186 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1190 ();
 DECAPx1_ASAP7_75t_R FILLER_221_1204 ();
 DECAPx1_ASAP7_75t_R FILLER_221_1211 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1256 ();
 DECAPx1_ASAP7_75t_R FILLER_221_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1268 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1275 ();
 FILLER_ASAP7_75t_R FILLER_221_1281 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1309 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1328 ();
 DECAPx4_ASAP7_75t_R FILLER_221_1335 ();
 FILLER_ASAP7_75t_R FILLER_221_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_222_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_50 ();
 FILLER_ASAP7_75t_R FILLER_222_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_111 ();
 DECAPx2_ASAP7_75t_R FILLER_222_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_121 ();
 DECAPx6_ASAP7_75t_R FILLER_222_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_149 ();
 DECAPx1_ASAP7_75t_R FILLER_222_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_201 ();
 DECAPx6_ASAP7_75t_R FILLER_222_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_222 ();
 DECAPx2_ASAP7_75t_R FILLER_222_237 ();
 FILLER_ASAP7_75t_R FILLER_222_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_245 ();
 DECAPx1_ASAP7_75t_R FILLER_222_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_260 ();
 DECAPx10_ASAP7_75t_R FILLER_222_267 ();
 DECAPx1_ASAP7_75t_R FILLER_222_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_293 ();
 DECAPx2_ASAP7_75t_R FILLER_222_300 ();
 DECAPx1_ASAP7_75t_R FILLER_222_329 ();
 DECAPx1_ASAP7_75t_R FILLER_222_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_349 ();
 DECAPx2_ASAP7_75t_R FILLER_222_359 ();
 FILLER_ASAP7_75t_R FILLER_222_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_367 ();
 DECAPx1_ASAP7_75t_R FILLER_222_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_389 ();
 DECAPx4_ASAP7_75t_R FILLER_222_426 ();
 DECAPx6_ASAP7_75t_R FILLER_222_442 ();
 DECAPx10_ASAP7_75t_R FILLER_222_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_486 ();
 DECAPx2_ASAP7_75t_R FILLER_222_493 ();
 FILLER_ASAP7_75t_R FILLER_222_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_504 ();
 DECAPx1_ASAP7_75t_R FILLER_222_508 ();
 DECAPx6_ASAP7_75t_R FILLER_222_518 ();
 DECAPx1_ASAP7_75t_R FILLER_222_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_562 ();
 DECAPx2_ASAP7_75t_R FILLER_222_590 ();
 DECAPx4_ASAP7_75t_R FILLER_222_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_641 ();
 DECAPx1_ASAP7_75t_R FILLER_222_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_664 ();
 FILLER_ASAP7_75t_R FILLER_222_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_673 ();
 FILLER_ASAP7_75t_R FILLER_222_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_698 ();
 DECAPx1_ASAP7_75t_R FILLER_222_715 ();
 DECAPx2_ASAP7_75t_R FILLER_222_745 ();
 FILLER_ASAP7_75t_R FILLER_222_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_753 ();
 DECAPx2_ASAP7_75t_R FILLER_222_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_770 ();
 DECAPx1_ASAP7_75t_R FILLER_222_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_785 ();
 DECAPx4_ASAP7_75t_R FILLER_222_792 ();
 FILLER_ASAP7_75t_R FILLER_222_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_804 ();
 DECAPx10_ASAP7_75t_R FILLER_222_808 ();
 DECAPx10_ASAP7_75t_R FILLER_222_830 ();
 DECAPx1_ASAP7_75t_R FILLER_222_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_856 ();
 DECAPx10_ASAP7_75t_R FILLER_222_862 ();
 FILLER_ASAP7_75t_R FILLER_222_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_886 ();
 DECAPx6_ASAP7_75t_R FILLER_222_915 ();
 FILLER_ASAP7_75t_R FILLER_222_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_931 ();
 DECAPx6_ASAP7_75t_R FILLER_222_948 ();
 DECAPx1_ASAP7_75t_R FILLER_222_962 ();
 DECAPx1_ASAP7_75t_R FILLER_222_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_991 ();
 DECAPx4_ASAP7_75t_R FILLER_222_995 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1044 ();
 FILLER_ASAP7_75t_R FILLER_222_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_222_1056 ();
 FILLER_ASAP7_75t_R FILLER_222_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_222_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1115 ();
 FILLER_ASAP7_75t_R FILLER_222_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_222_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1177 ();
 DECAPx4_ASAP7_75t_R FILLER_222_1184 ();
 FILLER_ASAP7_75t_R FILLER_222_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1207 ();
 DECAPx4_ASAP7_75t_R FILLER_222_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_222_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1296 ();
 DECAPx6_ASAP7_75t_R FILLER_222_1300 ();
 FILLER_ASAP7_75t_R FILLER_222_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1322 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1344 ();
 FILLER_ASAP7_75t_R FILLER_222_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1358 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1362 ();
 FILLER_ASAP7_75t_R FILLER_222_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_222_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_223_2 ();
 DECAPx4_ASAP7_75t_R FILLER_223_24 ();
 FILLER_ASAP7_75t_R FILLER_223_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_42 ();
 DECAPx2_ASAP7_75t_R FILLER_223_47 ();
 FILLER_ASAP7_75t_R FILLER_223_59 ();
 DECAPx4_ASAP7_75t_R FILLER_223_70 ();
 FILLER_ASAP7_75t_R FILLER_223_80 ();
 DECAPx2_ASAP7_75t_R FILLER_223_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_94 ();
 DECAPx4_ASAP7_75t_R FILLER_223_104 ();
 FILLER_ASAP7_75t_R FILLER_223_114 ();
 DECAPx10_ASAP7_75t_R FILLER_223_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_164 ();
 FILLER_ASAP7_75t_R FILLER_223_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_193 ();
 FILLER_ASAP7_75t_R FILLER_223_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_221 ();
 DECAPx2_ASAP7_75t_R FILLER_223_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_242 ();
 FILLER_ASAP7_75t_R FILLER_223_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_264 ();
 DECAPx4_ASAP7_75t_R FILLER_223_278 ();
 FILLER_ASAP7_75t_R FILLER_223_294 ();
 DECAPx4_ASAP7_75t_R FILLER_223_322 ();
 FILLER_ASAP7_75t_R FILLER_223_332 ();
 DECAPx2_ASAP7_75t_R FILLER_223_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_366 ();
 FILLER_ASAP7_75t_R FILLER_223_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_380 ();
 DECAPx1_ASAP7_75t_R FILLER_223_388 ();
 DECAPx10_ASAP7_75t_R FILLER_223_410 ();
 FILLER_ASAP7_75t_R FILLER_223_432 ();
 DECAPx10_ASAP7_75t_R FILLER_223_451 ();
 DECAPx1_ASAP7_75t_R FILLER_223_473 ();
 DECAPx6_ASAP7_75t_R FILLER_223_495 ();
 DECAPx2_ASAP7_75t_R FILLER_223_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_518 ();
 DECAPx10_ASAP7_75t_R FILLER_223_527 ();
 DECAPx10_ASAP7_75t_R FILLER_223_549 ();
 DECAPx1_ASAP7_75t_R FILLER_223_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_575 ();
 DECAPx4_ASAP7_75t_R FILLER_223_608 ();
 FILLER_ASAP7_75t_R FILLER_223_618 ();
 DECAPx4_ASAP7_75t_R FILLER_223_623 ();
 FILLER_ASAP7_75t_R FILLER_223_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_635 ();
 DECAPx6_ASAP7_75t_R FILLER_223_654 ();
 DECAPx2_ASAP7_75t_R FILLER_223_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_674 ();
 FILLER_ASAP7_75t_R FILLER_223_681 ();
 DECAPx2_ASAP7_75t_R FILLER_223_715 ();
 DECAPx6_ASAP7_75t_R FILLER_223_733 ();
 DECAPx1_ASAP7_75t_R FILLER_223_747 ();
 DECAPx1_ASAP7_75t_R FILLER_223_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_771 ();
 DECAPx4_ASAP7_75t_R FILLER_223_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_798 ();
 DECAPx10_ASAP7_75t_R FILLER_223_802 ();
 DECAPx6_ASAP7_75t_R FILLER_223_824 ();
 DECAPx1_ASAP7_75t_R FILLER_223_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_842 ();
 DECAPx10_ASAP7_75t_R FILLER_223_869 ();
 DECAPx4_ASAP7_75t_R FILLER_223_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_901 ();
 DECAPx4_ASAP7_75t_R FILLER_223_914 ();
 DECAPx2_ASAP7_75t_R FILLER_223_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_942 ();
 DECAPx6_ASAP7_75t_R FILLER_223_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_992 ();
 DECAPx6_ASAP7_75t_R FILLER_223_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1019 ();
 FILLER_ASAP7_75t_R FILLER_223_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1063 ();
 FILLER_ASAP7_75t_R FILLER_223_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_223_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1189 ();
 FILLER_ASAP7_75t_R FILLER_223_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1240 ();
 FILLER_ASAP7_75t_R FILLER_223_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1284 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1324 ();
 FILLER_ASAP7_75t_R FILLER_223_1330 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1338 ();
 FILLER_ASAP7_75t_R FILLER_223_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_223_1372 ();
 DECAPx6_ASAP7_75t_R FILLER_224_2 ();
 FILLER_ASAP7_75t_R FILLER_224_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_18 ();
 FILLER_ASAP7_75t_R FILLER_224_45 ();
 DECAPx6_ASAP7_75t_R FILLER_224_79 ();
 DECAPx2_ASAP7_75t_R FILLER_224_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_163 ();
 DECAPx2_ASAP7_75t_R FILLER_224_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_179 ();
 DECAPx10_ASAP7_75t_R FILLER_224_195 ();
 DECAPx2_ASAP7_75t_R FILLER_224_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_237 ();
 DECAPx4_ASAP7_75t_R FILLER_224_252 ();
 FILLER_ASAP7_75t_R FILLER_224_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_264 ();
 FILLER_ASAP7_75t_R FILLER_224_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_273 ();
 DECAPx1_ASAP7_75t_R FILLER_224_288 ();
 DECAPx2_ASAP7_75t_R FILLER_224_298 ();
 FILLER_ASAP7_75t_R FILLER_224_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_306 ();
 DECAPx2_ASAP7_75t_R FILLER_224_321 ();
 FILLER_ASAP7_75t_R FILLER_224_327 ();
 DECAPx1_ASAP7_75t_R FILLER_224_345 ();
 DECAPx4_ASAP7_75t_R FILLER_224_358 ();
 DECAPx1_ASAP7_75t_R FILLER_224_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_389 ();
 DECAPx4_ASAP7_75t_R FILLER_224_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_428 ();
 DECAPx2_ASAP7_75t_R FILLER_224_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_461 ();
 DECAPx6_ASAP7_75t_R FILLER_224_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_512 ();
 DECAPx1_ASAP7_75t_R FILLER_224_516 ();
 FILLER_ASAP7_75t_R FILLER_224_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_534 ();
 DECAPx2_ASAP7_75t_R FILLER_224_544 ();
 FILLER_ASAP7_75t_R FILLER_224_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_556 ();
 FILLER_ASAP7_75t_R FILLER_224_593 ();
 DECAPx2_ASAP7_75t_R FILLER_224_601 ();
 DECAPx2_ASAP7_75t_R FILLER_224_610 ();
 FILLER_ASAP7_75t_R FILLER_224_616 ();
 DECAPx6_ASAP7_75t_R FILLER_224_636 ();
 DECAPx2_ASAP7_75t_R FILLER_224_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_656 ();
 DECAPx1_ASAP7_75t_R FILLER_224_694 ();
 DECAPx2_ASAP7_75t_R FILLER_224_711 ();
 FILLER_ASAP7_75t_R FILLER_224_717 ();
 FILLER_ASAP7_75t_R FILLER_224_726 ();
 DECAPx1_ASAP7_75t_R FILLER_224_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_742 ();
 DECAPx4_ASAP7_75t_R FILLER_224_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_779 ();
 DECAPx10_ASAP7_75t_R FILLER_224_806 ();
 DECAPx2_ASAP7_75t_R FILLER_224_828 ();
 FILLER_ASAP7_75t_R FILLER_224_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_836 ();
 DECAPx6_ASAP7_75t_R FILLER_224_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_876 ();
 DECAPx6_ASAP7_75t_R FILLER_224_884 ();
 DECAPx2_ASAP7_75t_R FILLER_224_898 ();
 FILLER_ASAP7_75t_R FILLER_224_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_916 ();
 DECAPx4_ASAP7_75t_R FILLER_224_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_948 ();
 DECAPx6_ASAP7_75t_R FILLER_224_956 ();
 DECAPx2_ASAP7_75t_R FILLER_224_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_976 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_224_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1089 ();
 FILLER_ASAP7_75t_R FILLER_224_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1124 ();
 FILLER_ASAP7_75t_R FILLER_224_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_224_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1159 ();
 FILLER_ASAP7_75t_R FILLER_224_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1175 ();
 FILLER_ASAP7_75t_R FILLER_224_1215 ();
 DECAPx1_ASAP7_75t_R FILLER_224_1224 ();
 FILLER_ASAP7_75t_R FILLER_224_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1233 ();
 FILLER_ASAP7_75t_R FILLER_224_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1243 ();
 FILLER_ASAP7_75t_R FILLER_224_1250 ();
 DECAPx1_ASAP7_75t_R FILLER_224_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1282 ();
 FILLER_ASAP7_75t_R FILLER_224_1315 ();
 DECAPx1_ASAP7_75t_R FILLER_224_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1347 ();
 FILLER_ASAP7_75t_R FILLER_224_1354 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1369 ();
 FILLER_ASAP7_75t_R FILLER_224_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_224_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_225_2 ();
 DECAPx2_ASAP7_75t_R FILLER_225_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_30 ();
 DECAPx10_ASAP7_75t_R FILLER_225_40 ();
 DECAPx4_ASAP7_75t_R FILLER_225_65 ();
 FILLER_ASAP7_75t_R FILLER_225_87 ();
 DECAPx2_ASAP7_75t_R FILLER_225_92 ();
 DECAPx4_ASAP7_75t_R FILLER_225_104 ();
 DECAPx10_ASAP7_75t_R FILLER_225_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_145 ();
 DECAPx1_ASAP7_75t_R FILLER_225_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_160 ();
 DECAPx2_ASAP7_75t_R FILLER_225_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_181 ();
 DECAPx6_ASAP7_75t_R FILLER_225_188 ();
 DECAPx1_ASAP7_75t_R FILLER_225_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_220 ();
 DECAPx6_ASAP7_75t_R FILLER_225_227 ();
 DECAPx4_ASAP7_75t_R FILLER_225_247 ();
 FILLER_ASAP7_75t_R FILLER_225_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_259 ();
 DECAPx6_ASAP7_75t_R FILLER_225_266 ();
 FILLER_ASAP7_75t_R FILLER_225_280 ();
 DECAPx2_ASAP7_75t_R FILLER_225_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_309 ();
 DECAPx10_ASAP7_75t_R FILLER_225_322 ();
 DECAPx2_ASAP7_75t_R FILLER_225_344 ();
 FILLER_ASAP7_75t_R FILLER_225_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_352 ();
 DECAPx1_ASAP7_75t_R FILLER_225_389 ();
 DECAPx6_ASAP7_75t_R FILLER_225_410 ();
 DECAPx1_ASAP7_75t_R FILLER_225_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_442 ();
 DECAPx4_ASAP7_75t_R FILLER_225_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_462 ();
 FILLER_ASAP7_75t_R FILLER_225_481 ();
 DECAPx1_ASAP7_75t_R FILLER_225_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_538 ();
 DECAPx10_ASAP7_75t_R FILLER_225_565 ();
 DECAPx2_ASAP7_75t_R FILLER_225_587 ();
 DECAPx2_ASAP7_75t_R FILLER_225_619 ();
 FILLER_ASAP7_75t_R FILLER_225_625 ();
 DECAPx4_ASAP7_75t_R FILLER_225_688 ();
 FILLER_ASAP7_75t_R FILLER_225_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_753 ();
 DECAPx1_ASAP7_75t_R FILLER_225_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_781 ();
 DECAPx10_ASAP7_75t_R FILLER_225_785 ();
 DECAPx2_ASAP7_75t_R FILLER_225_807 ();
 FILLER_ASAP7_75t_R FILLER_225_813 ();
 DECAPx4_ASAP7_75t_R FILLER_225_825 ();
 DECAPx2_ASAP7_75t_R FILLER_225_849 ();
 FILLER_ASAP7_75t_R FILLER_225_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_857 ();
 FILLER_ASAP7_75t_R FILLER_225_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_870 ();
 DECAPx6_ASAP7_75t_R FILLER_225_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_911 ();
 DECAPx2_ASAP7_75t_R FILLER_225_926 ();
 DECAPx2_ASAP7_75t_R FILLER_225_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_968 ();
 DECAPx2_ASAP7_75t_R FILLER_225_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_981 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1008 ();
 DECAPx6_ASAP7_75t_R FILLER_225_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1030 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1041 ();
 FILLER_ASAP7_75t_R FILLER_225_1047 ();
 FILLER_ASAP7_75t_R FILLER_225_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1075 ();
 FILLER_ASAP7_75t_R FILLER_225_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1109 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1167 ();
 FILLER_ASAP7_75t_R FILLER_225_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1175 ();
 DECAPx6_ASAP7_75t_R FILLER_225_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1208 ();
 DECAPx4_ASAP7_75t_R FILLER_225_1217 ();
 FILLER_ASAP7_75t_R FILLER_225_1227 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1281 ();
 FILLER_ASAP7_75t_R FILLER_225_1297 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1305 ();
 FILLER_ASAP7_75t_R FILLER_225_1348 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1356 ();
 DECAPx6_ASAP7_75t_R FILLER_225_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_226_2 ();
 DECAPx10_ASAP7_75t_R FILLER_226_24 ();
 DECAPx2_ASAP7_75t_R FILLER_226_46 ();
 FILLER_ASAP7_75t_R FILLER_226_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_54 ();
 DECAPx4_ASAP7_75t_R FILLER_226_61 ();
 FILLER_ASAP7_75t_R FILLER_226_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_73 ();
 DECAPx4_ASAP7_75t_R FILLER_226_100 ();
 FILLER_ASAP7_75t_R FILLER_226_110 ();
 DECAPx2_ASAP7_75t_R FILLER_226_115 ();
 FILLER_ASAP7_75t_R FILLER_226_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_123 ();
 DECAPx6_ASAP7_75t_R FILLER_226_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_141 ();
 FILLER_ASAP7_75t_R FILLER_226_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_170 ();
 DECAPx10_ASAP7_75t_R FILLER_226_177 ();
 DECAPx1_ASAP7_75t_R FILLER_226_205 ();
 DECAPx2_ASAP7_75t_R FILLER_226_223 ();
 DECAPx6_ASAP7_75t_R FILLER_226_241 ();
 FILLER_ASAP7_75t_R FILLER_226_255 ();
 DECAPx1_ASAP7_75t_R FILLER_226_277 ();
 FILLER_ASAP7_75t_R FILLER_226_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_290 ();
 DECAPx4_ASAP7_75t_R FILLER_226_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_307 ();
 DECAPx2_ASAP7_75t_R FILLER_226_314 ();
 DECAPx1_ASAP7_75t_R FILLER_226_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_337 ();
 DECAPx10_ASAP7_75t_R FILLER_226_344 ();
 DECAPx2_ASAP7_75t_R FILLER_226_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_372 ();
 DECAPx2_ASAP7_75t_R FILLER_226_386 ();
 FILLER_ASAP7_75t_R FILLER_226_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_394 ();
 DECAPx6_ASAP7_75t_R FILLER_226_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_417 ();
 FILLER_ASAP7_75t_R FILLER_226_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_430 ();
 DECAPx10_ASAP7_75t_R FILLER_226_437 ();
 FILLER_ASAP7_75t_R FILLER_226_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_461 ();
 DECAPx4_ASAP7_75t_R FILLER_226_489 ();
 FILLER_ASAP7_75t_R FILLER_226_499 ();
 DECAPx4_ASAP7_75t_R FILLER_226_515 ();
 DECAPx2_ASAP7_75t_R FILLER_226_531 ();
 FILLER_ASAP7_75t_R FILLER_226_537 ();
 DECAPx2_ASAP7_75t_R FILLER_226_545 ();
 FILLER_ASAP7_75t_R FILLER_226_551 ();
 DECAPx4_ASAP7_75t_R FILLER_226_559 ();
 DECAPx2_ASAP7_75t_R FILLER_226_587 ();
 FILLER_ASAP7_75t_R FILLER_226_593 ();
 DECAPx2_ASAP7_75t_R FILLER_226_601 ();
 DECAPx2_ASAP7_75t_R FILLER_226_639 ();
 FILLER_ASAP7_75t_R FILLER_226_645 ();
 DECAPx10_ASAP7_75t_R FILLER_226_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_672 ();
 DECAPx6_ASAP7_75t_R FILLER_226_683 ();
 FILLER_ASAP7_75t_R FILLER_226_697 ();
 DECAPx4_ASAP7_75t_R FILLER_226_705 ();
 FILLER_ASAP7_75t_R FILLER_226_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_717 ();
 DECAPx6_ASAP7_75t_R FILLER_226_721 ();
 DECAPx2_ASAP7_75t_R FILLER_226_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_741 ();
 DECAPx6_ASAP7_75t_R FILLER_226_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_762 ();
 DECAPx10_ASAP7_75t_R FILLER_226_789 ();
 DECAPx10_ASAP7_75t_R FILLER_226_811 ();
 DECAPx4_ASAP7_75t_R FILLER_226_833 ();
 FILLER_ASAP7_75t_R FILLER_226_843 ();
 DECAPx2_ASAP7_75t_R FILLER_226_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_890 ();
 FILLER_ASAP7_75t_R FILLER_226_901 ();
 DECAPx4_ASAP7_75t_R FILLER_226_929 ();
 FILLER_ASAP7_75t_R FILLER_226_939 ();
 FILLER_ASAP7_75t_R FILLER_226_951 ();
 DECAPx6_ASAP7_75t_R FILLER_226_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_989 ();
 DECAPx2_ASAP7_75t_R FILLER_226_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1052 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1078 ();
 DECAPx4_ASAP7_75t_R FILLER_226_1111 ();
 FILLER_ASAP7_75t_R FILLER_226_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_226_1149 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_226_1172 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1205 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1227 ();
 FILLER_ASAP7_75t_R FILLER_226_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1301 ();
 DECAPx2_ASAP7_75t_R FILLER_226_1323 ();
 FILLER_ASAP7_75t_R FILLER_226_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1331 ();
 DECAPx4_ASAP7_75t_R FILLER_226_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1345 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_227_2 ();
 DECAPx2_ASAP7_75t_R FILLER_227_16 ();
 DECAPx1_ASAP7_75t_R FILLER_227_25 ();
 DECAPx2_ASAP7_75t_R FILLER_227_39 ();
 FILLER_ASAP7_75t_R FILLER_227_75 ();
 FILLER_ASAP7_75t_R FILLER_227_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_123 ();
 DECAPx4_ASAP7_75t_R FILLER_227_137 ();
 FILLER_ASAP7_75t_R FILLER_227_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_149 ();
 FILLER_ASAP7_75t_R FILLER_227_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_196 ();
 DECAPx1_ASAP7_75t_R FILLER_227_205 ();
 DECAPx2_ASAP7_75t_R FILLER_227_223 ();
 DECAPx2_ASAP7_75t_R FILLER_227_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_251 ();
 DECAPx6_ASAP7_75t_R FILLER_227_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_280 ();
 DECAPx6_ASAP7_75t_R FILLER_227_289 ();
 DECAPx1_ASAP7_75t_R FILLER_227_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_333 ();
 DECAPx1_ASAP7_75t_R FILLER_227_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_348 ();
 FILLER_ASAP7_75t_R FILLER_227_373 ();
 DECAPx1_ASAP7_75t_R FILLER_227_386 ();
 DECAPx2_ASAP7_75t_R FILLER_227_401 ();
 FILLER_ASAP7_75t_R FILLER_227_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_433 ();
 DECAPx1_ASAP7_75t_R FILLER_227_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_450 ();
 DECAPx4_ASAP7_75t_R FILLER_227_461 ();
 FILLER_ASAP7_75t_R FILLER_227_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_473 ();
 DECAPx2_ASAP7_75t_R FILLER_227_492 ();
 FILLER_ASAP7_75t_R FILLER_227_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_500 ();
 FILLER_ASAP7_75t_R FILLER_227_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_509 ();
 DECAPx6_ASAP7_75t_R FILLER_227_524 ();
 FILLER_ASAP7_75t_R FILLER_227_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_540 ();
 DECAPx10_ASAP7_75t_R FILLER_227_555 ();
 DECAPx1_ASAP7_75t_R FILLER_227_577 ();
 FILLER_ASAP7_75t_R FILLER_227_599 ();
 DECAPx4_ASAP7_75t_R FILLER_227_638 ();
 FILLER_ASAP7_75t_R FILLER_227_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_650 ();
 FILLER_ASAP7_75t_R FILLER_227_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_656 ();
 DECAPx1_ASAP7_75t_R FILLER_227_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_697 ();
 DECAPx2_ASAP7_75t_R FILLER_227_708 ();
 FILLER_ASAP7_75t_R FILLER_227_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_716 ();
 DECAPx4_ASAP7_75t_R FILLER_227_727 ();
 DECAPx4_ASAP7_75t_R FILLER_227_743 ();
 FILLER_ASAP7_75t_R FILLER_227_753 ();
 DECAPx2_ASAP7_75t_R FILLER_227_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_768 ();
 DECAPx6_ASAP7_75t_R FILLER_227_802 ();
 DECAPx1_ASAP7_75t_R FILLER_227_816 ();
 DECAPx6_ASAP7_75t_R FILLER_227_823 ();
 DECAPx2_ASAP7_75t_R FILLER_227_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_843 ();
 DECAPx2_ASAP7_75t_R FILLER_227_854 ();
 DECAPx6_ASAP7_75t_R FILLER_227_863 ();
 FILLER_ASAP7_75t_R FILLER_227_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_879 ();
 DECAPx1_ASAP7_75t_R FILLER_227_888 ();
 FILLER_ASAP7_75t_R FILLER_227_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_904 ();
 DECAPx1_ASAP7_75t_R FILLER_227_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_916 ();
 DECAPx1_ASAP7_75t_R FILLER_227_920 ();
 DECAPx1_ASAP7_75t_R FILLER_227_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_930 ();
 DECAPx10_ASAP7_75t_R FILLER_227_937 ();
 DECAPx2_ASAP7_75t_R FILLER_227_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_979 ();
 DECAPx1_ASAP7_75t_R FILLER_227_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_997 ();
 FILLER_ASAP7_75t_R FILLER_227_1008 ();
 DECAPx6_ASAP7_75t_R FILLER_227_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_227_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1111 ();
 FILLER_ASAP7_75t_R FILLER_227_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1135 ();
 DECAPx6_ASAP7_75t_R FILLER_227_1146 ();
 FILLER_ASAP7_75t_R FILLER_227_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1188 ();
 FILLER_ASAP7_75t_R FILLER_227_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1196 ();
 DECAPx4_ASAP7_75t_R FILLER_227_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1293 ();
 DECAPx4_ASAP7_75t_R FILLER_227_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1370 ();
 DECAPx2_ASAP7_75t_R FILLER_228_2 ();
 FILLER_ASAP7_75t_R FILLER_228_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_59 ();
 DECAPx2_ASAP7_75t_R FILLER_228_63 ();
 FILLER_ASAP7_75t_R FILLER_228_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_97 ();
 FILLER_ASAP7_75t_R FILLER_228_104 ();
 DECAPx6_ASAP7_75t_R FILLER_228_158 ();
 FILLER_ASAP7_75t_R FILLER_228_172 ();
 DECAPx2_ASAP7_75t_R FILLER_228_180 ();
 DECAPx2_ASAP7_75t_R FILLER_228_206 ();
 FILLER_ASAP7_75t_R FILLER_228_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_214 ();
 FILLER_ASAP7_75t_R FILLER_228_229 ();
 FILLER_ASAP7_75t_R FILLER_228_259 ();
 DECAPx2_ASAP7_75t_R FILLER_228_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_273 ();
 FILLER_ASAP7_75t_R FILLER_228_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_282 ();
 DECAPx2_ASAP7_75t_R FILLER_228_289 ();
 FILLER_ASAP7_75t_R FILLER_228_295 ();
 DECAPx2_ASAP7_75t_R FILLER_228_318 ();
 FILLER_ASAP7_75t_R FILLER_228_324 ();
 DECAPx4_ASAP7_75t_R FILLER_228_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_342 ();
 DECAPx10_ASAP7_75t_R FILLER_228_361 ();
 DECAPx4_ASAP7_75t_R FILLER_228_383 ();
 DECAPx4_ASAP7_75t_R FILLER_228_399 ();
 FILLER_ASAP7_75t_R FILLER_228_409 ();
 DECAPx10_ASAP7_75t_R FILLER_228_429 ();
 FILLER_ASAP7_75t_R FILLER_228_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_453 ();
 FILLER_ASAP7_75t_R FILLER_228_460 ();
 DECAPx1_ASAP7_75t_R FILLER_228_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_479 ();
 FILLER_ASAP7_75t_R FILLER_228_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_488 ();
 DECAPx4_ASAP7_75t_R FILLER_228_500 ();
 DECAPx1_ASAP7_75t_R FILLER_228_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_540 ();
 FILLER_ASAP7_75t_R FILLER_228_547 ();
 DECAPx6_ASAP7_75t_R FILLER_228_558 ();
 DECAPx2_ASAP7_75t_R FILLER_228_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_581 ();
 DECAPx2_ASAP7_75t_R FILLER_228_594 ();
 FILLER_ASAP7_75t_R FILLER_228_600 ();
 DECAPx2_ASAP7_75t_R FILLER_228_605 ();
 FILLER_ASAP7_75t_R FILLER_228_611 ();
 DECAPx2_ASAP7_75t_R FILLER_228_620 ();
 FILLER_ASAP7_75t_R FILLER_228_626 ();
 DECAPx2_ASAP7_75t_R FILLER_228_663 ();
 FILLER_ASAP7_75t_R FILLER_228_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_671 ();
 FILLER_ASAP7_75t_R FILLER_228_675 ();
 DECAPx1_ASAP7_75t_R FILLER_228_709 ();
 DECAPx4_ASAP7_75t_R FILLER_228_781 ();
 DECAPx4_ASAP7_75t_R FILLER_228_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_804 ();
 DECAPx4_ASAP7_75t_R FILLER_228_831 ();
 FILLER_ASAP7_75t_R FILLER_228_841 ();
 DECAPx10_ASAP7_75t_R FILLER_228_850 ();
 DECAPx4_ASAP7_75t_R FILLER_228_872 ();
 DECAPx6_ASAP7_75t_R FILLER_228_888 ();
 DECAPx1_ASAP7_75t_R FILLER_228_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_906 ();
 DECAPx4_ASAP7_75t_R FILLER_228_915 ();
 FILLER_ASAP7_75t_R FILLER_228_925 ();
 DECAPx4_ASAP7_75t_R FILLER_228_942 ();
 FILLER_ASAP7_75t_R FILLER_228_952 ();
 DECAPx6_ASAP7_75t_R FILLER_228_964 ();
 FILLER_ASAP7_75t_R FILLER_228_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_980 ();
 DECAPx4_ASAP7_75t_R FILLER_228_995 ();
 FILLER_ASAP7_75t_R FILLER_228_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_228_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1044 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1061 ();
 DECAPx4_ASAP7_75t_R FILLER_228_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1078 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_228_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_228_1151 ();
 FILLER_ASAP7_75t_R FILLER_228_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1159 ();
 FILLER_ASAP7_75t_R FILLER_228_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1175 ();
 FILLER_ASAP7_75t_R FILLER_228_1179 ();
 FILLER_ASAP7_75t_R FILLER_228_1193 ();
 FILLER_ASAP7_75t_R FILLER_228_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_228_1273 ();
 FILLER_ASAP7_75t_R FILLER_228_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1321 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1328 ();
 FILLER_ASAP7_75t_R FILLER_228_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1357 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_229_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_24 ();
 DECAPx10_ASAP7_75t_R FILLER_229_51 ();
 FILLER_ASAP7_75t_R FILLER_229_73 ();
 DECAPx1_ASAP7_75t_R FILLER_229_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_85 ();
 DECAPx10_ASAP7_75t_R FILLER_229_98 ();
 FILLER_ASAP7_75t_R FILLER_229_120 ();
 FILLER_ASAP7_75t_R FILLER_229_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_141 ();
 DECAPx2_ASAP7_75t_R FILLER_229_152 ();
 FILLER_ASAP7_75t_R FILLER_229_158 ();
 DECAPx6_ASAP7_75t_R FILLER_229_166 ();
 FILLER_ASAP7_75t_R FILLER_229_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_182 ();
 DECAPx4_ASAP7_75t_R FILLER_229_197 ();
 FILLER_ASAP7_75t_R FILLER_229_207 ();
 DECAPx6_ASAP7_75t_R FILLER_229_223 ();
 FILLER_ASAP7_75t_R FILLER_229_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_239 ();
 FILLER_ASAP7_75t_R FILLER_229_246 ();
 DECAPx1_ASAP7_75t_R FILLER_229_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_260 ();
 DECAPx1_ASAP7_75t_R FILLER_229_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_285 ();
 DECAPx10_ASAP7_75t_R FILLER_229_307 ();
 DECAPx4_ASAP7_75t_R FILLER_229_329 ();
 FILLER_ASAP7_75t_R FILLER_229_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_358 ();
 FILLER_ASAP7_75t_R FILLER_229_372 ();
 DECAPx4_ASAP7_75t_R FILLER_229_380 ();
 FILLER_ASAP7_75t_R FILLER_229_390 ();
 DECAPx2_ASAP7_75t_R FILLER_229_395 ();
 FILLER_ASAP7_75t_R FILLER_229_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_403 ();
 DECAPx1_ASAP7_75t_R FILLER_229_407 ();
 DECAPx6_ASAP7_75t_R FILLER_229_419 ();
 DECAPx2_ASAP7_75t_R FILLER_229_439 ();
 DECAPx6_ASAP7_75t_R FILLER_229_464 ();
 DECAPx2_ASAP7_75t_R FILLER_229_478 ();
 DECAPx4_ASAP7_75t_R FILLER_229_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_506 ();
 DECAPx6_ASAP7_75t_R FILLER_229_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_551 ();
 DECAPx1_ASAP7_75t_R FILLER_229_584 ();
 DECAPx6_ASAP7_75t_R FILLER_229_614 ();
 DECAPx2_ASAP7_75t_R FILLER_229_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_634 ();
 DECAPx10_ASAP7_75t_R FILLER_229_642 ();
 DECAPx4_ASAP7_75t_R FILLER_229_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_674 ();
 DECAPx6_ASAP7_75t_R FILLER_229_682 ();
 FILLER_ASAP7_75t_R FILLER_229_696 ();
 DECAPx2_ASAP7_75t_R FILLER_229_701 ();
 FILLER_ASAP7_75t_R FILLER_229_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_719 ();
 FILLER_ASAP7_75t_R FILLER_229_732 ();
 DECAPx2_ASAP7_75t_R FILLER_229_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_766 ();
 DECAPx10_ASAP7_75t_R FILLER_229_779 ();
 DECAPx6_ASAP7_75t_R FILLER_229_801 ();
 FILLER_ASAP7_75t_R FILLER_229_832 ();
 FILLER_ASAP7_75t_R FILLER_229_840 ();
 FILLER_ASAP7_75t_R FILLER_229_848 ();
 DECAPx6_ASAP7_75t_R FILLER_229_886 ();
 FILLER_ASAP7_75t_R FILLER_229_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_902 ();
 FILLER_ASAP7_75t_R FILLER_229_922 ();
 DECAPx4_ASAP7_75t_R FILLER_229_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_962 ();
 DECAPx4_ASAP7_75t_R FILLER_229_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_979 ();
 DECAPx4_ASAP7_75t_R FILLER_229_995 ();
 FILLER_ASAP7_75t_R FILLER_229_1005 ();
 FILLER_ASAP7_75t_R FILLER_229_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1019 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1090 ();
 DECAPx4_ASAP7_75t_R FILLER_229_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1143 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1213 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1220 ();
 FILLER_ASAP7_75t_R FILLER_229_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1228 ();
 FILLER_ASAP7_75t_R FILLER_229_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1234 ();
 FILLER_ASAP7_75t_R FILLER_229_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1250 ();
 FILLER_ASAP7_75t_R FILLER_229_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1278 ();
 FILLER_ASAP7_75t_R FILLER_229_1308 ();
 FILLER_ASAP7_75t_R FILLER_229_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1315 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1322 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1329 ();
 FILLER_ASAP7_75t_R FILLER_229_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1351 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1373 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1387 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_230_2 ();
 DECAPx1_ASAP7_75t_R FILLER_230_24 ();
 FILLER_ASAP7_75t_R FILLER_230_34 ();
 DECAPx2_ASAP7_75t_R FILLER_230_45 ();
 FILLER_ASAP7_75t_R FILLER_230_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_68 ();
 FILLER_ASAP7_75t_R FILLER_230_79 ();
 DECAPx1_ASAP7_75t_R FILLER_230_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_137 ();
 FILLER_ASAP7_75t_R FILLER_230_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_166 ();
 FILLER_ASAP7_75t_R FILLER_230_173 ();
 DECAPx1_ASAP7_75t_R FILLER_230_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_182 ();
 DECAPx2_ASAP7_75t_R FILLER_230_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_198 ();
 DECAPx2_ASAP7_75t_R FILLER_230_205 ();
 DECAPx2_ASAP7_75t_R FILLER_230_217 ();
 FILLER_ASAP7_75t_R FILLER_230_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_225 ();
 DECAPx1_ASAP7_75t_R FILLER_230_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_257 ();
 DECAPx6_ASAP7_75t_R FILLER_230_278 ();
 DECAPx2_ASAP7_75t_R FILLER_230_304 ();
 FILLER_ASAP7_75t_R FILLER_230_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_312 ();
 DECAPx1_ASAP7_75t_R FILLER_230_319 ();
 DECAPx6_ASAP7_75t_R FILLER_230_332 ();
 DECAPx1_ASAP7_75t_R FILLER_230_346 ();
 DECAPx1_ASAP7_75t_R FILLER_230_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_416 ();
 DECAPx1_ASAP7_75t_R FILLER_230_423 ();
 DECAPx1_ASAP7_75t_R FILLER_230_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_447 ();
 DECAPx2_ASAP7_75t_R FILLER_230_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_470 ();
 FILLER_ASAP7_75t_R FILLER_230_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_489 ();
 DECAPx1_ASAP7_75t_R FILLER_230_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_504 ();
 DECAPx1_ASAP7_75t_R FILLER_230_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_517 ();
 DECAPx1_ASAP7_75t_R FILLER_230_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_539 ();
 DECAPx2_ASAP7_75t_R FILLER_230_548 ();
 FILLER_ASAP7_75t_R FILLER_230_554 ();
 FILLER_ASAP7_75t_R FILLER_230_588 ();
 FILLER_ASAP7_75t_R FILLER_230_593 ();
 DECAPx1_ASAP7_75t_R FILLER_230_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_602 ();
 FILLER_ASAP7_75t_R FILLER_230_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_631 ();
 DECAPx1_ASAP7_75t_R FILLER_230_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_649 ();
 DECAPx1_ASAP7_75t_R FILLER_230_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_657 ();
 DECAPx6_ASAP7_75t_R FILLER_230_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_698 ();
 DECAPx6_ASAP7_75t_R FILLER_230_706 ();
 FILLER_ASAP7_75t_R FILLER_230_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_722 ();
 DECAPx6_ASAP7_75t_R FILLER_230_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_747 ();
 DECAPx6_ASAP7_75t_R FILLER_230_751 ();
 FILLER_ASAP7_75t_R FILLER_230_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_767 ();
 DECAPx10_ASAP7_75t_R FILLER_230_774 ();
 DECAPx2_ASAP7_75t_R FILLER_230_796 ();
 FILLER_ASAP7_75t_R FILLER_230_802 ();
 DECAPx2_ASAP7_75t_R FILLER_230_807 ();
 FILLER_ASAP7_75t_R FILLER_230_813 ();
 FILLER_ASAP7_75t_R FILLER_230_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_829 ();
 FILLER_ASAP7_75t_R FILLER_230_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_843 ();
 DECAPx1_ASAP7_75t_R FILLER_230_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_861 ();
 DECAPx1_ASAP7_75t_R FILLER_230_873 ();
 DECAPx6_ASAP7_75t_R FILLER_230_916 ();
 DECAPx1_ASAP7_75t_R FILLER_230_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_934 ();
 FILLER_ASAP7_75t_R FILLER_230_941 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1008 ();
 FILLER_ASAP7_75t_R FILLER_230_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_230_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1065 ();
 FILLER_ASAP7_75t_R FILLER_230_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1109 ();
 FILLER_ASAP7_75t_R FILLER_230_1115 ();
 DECAPx6_ASAP7_75t_R FILLER_230_1120 ();
 FILLER_ASAP7_75t_R FILLER_230_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_230_1152 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1173 ();
 FILLER_ASAP7_75t_R FILLER_230_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_230_1188 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1206 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_230_1246 ();
 FILLER_ASAP7_75t_R FILLER_230_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1269 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1299 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1321 ();
 FILLER_ASAP7_75t_R FILLER_230_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1378 ();
 FILLER_ASAP7_75t_R FILLER_230_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_231_2 ();
 DECAPx4_ASAP7_75t_R FILLER_231_24 ();
 FILLER_ASAP7_75t_R FILLER_231_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_43 ();
 FILLER_ASAP7_75t_R FILLER_231_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_50 ();
 FILLER_ASAP7_75t_R FILLER_231_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_79 ();
 DECAPx4_ASAP7_75t_R FILLER_231_86 ();
 DECAPx2_ASAP7_75t_R FILLER_231_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_111 ();
 DECAPx1_ASAP7_75t_R FILLER_231_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_120 ();
 DECAPx10_ASAP7_75t_R FILLER_231_124 ();
 DECAPx2_ASAP7_75t_R FILLER_231_146 ();
 DECAPx1_ASAP7_75t_R FILLER_231_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_186 ();
 FILLER_ASAP7_75t_R FILLER_231_213 ();
 FILLER_ASAP7_75t_R FILLER_231_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_220 ();
 DECAPx1_ASAP7_75t_R FILLER_231_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_232 ();
 DECAPx1_ASAP7_75t_R FILLER_231_241 ();
 DECAPx4_ASAP7_75t_R FILLER_231_251 ();
 DECAPx2_ASAP7_75t_R FILLER_231_267 ();
 FILLER_ASAP7_75t_R FILLER_231_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_275 ();
 DECAPx10_ASAP7_75t_R FILLER_231_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_304 ();
 DECAPx2_ASAP7_75t_R FILLER_231_334 ();
 FILLER_ASAP7_75t_R FILLER_231_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_342 ();
 DECAPx2_ASAP7_75t_R FILLER_231_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_357 ();
 DECAPx1_ASAP7_75t_R FILLER_231_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_368 ();
 DECAPx4_ASAP7_75t_R FILLER_231_375 ();
 FILLER_ASAP7_75t_R FILLER_231_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_387 ();
 FILLER_ASAP7_75t_R FILLER_231_394 ();
 DECAPx1_ASAP7_75t_R FILLER_231_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_406 ();
 FILLER_ASAP7_75t_R FILLER_231_413 ();
 DECAPx4_ASAP7_75t_R FILLER_231_421 ();
 DECAPx2_ASAP7_75t_R FILLER_231_437 ();
 FILLER_ASAP7_75t_R FILLER_231_443 ();
 DECAPx6_ASAP7_75t_R FILLER_231_457 ();
 FILLER_ASAP7_75t_R FILLER_231_471 ();
 DECAPx1_ASAP7_75t_R FILLER_231_479 ();
 FILLER_ASAP7_75t_R FILLER_231_503 ();
 FILLER_ASAP7_75t_R FILLER_231_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_519 ();
 DECAPx4_ASAP7_75t_R FILLER_231_528 ();
 DECAPx2_ASAP7_75t_R FILLER_231_561 ();
 FILLER_ASAP7_75t_R FILLER_231_567 ();
 DECAPx1_ASAP7_75t_R FILLER_231_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_605 ();
 DECAPx1_ASAP7_75t_R FILLER_231_632 ();
 DECAPx4_ASAP7_75t_R FILLER_231_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_672 ();
 FILLER_ASAP7_75t_R FILLER_231_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_747 ();
 FILLER_ASAP7_75t_R FILLER_231_761 ();
 FILLER_ASAP7_75t_R FILLER_231_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_775 ();
 DECAPx4_ASAP7_75t_R FILLER_231_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_789 ();
 FILLER_ASAP7_75t_R FILLER_231_833 ();
 DECAPx1_ASAP7_75t_R FILLER_231_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_863 ();
 DECAPx2_ASAP7_75t_R FILLER_231_867 ();
 FILLER_ASAP7_75t_R FILLER_231_873 ();
 DECAPx2_ASAP7_75t_R FILLER_231_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_907 ();
 DECAPx4_ASAP7_75t_R FILLER_231_914 ();
 DECAPx2_ASAP7_75t_R FILLER_231_935 ();
 FILLER_ASAP7_75t_R FILLER_231_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_943 ();
 DECAPx4_ASAP7_75t_R FILLER_231_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_963 ();
 DECAPx2_ASAP7_75t_R FILLER_231_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_976 ();
 DECAPx4_ASAP7_75t_R FILLER_231_986 ();
 FILLER_ASAP7_75t_R FILLER_231_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1001 ();
 DECAPx6_ASAP7_75t_R FILLER_231_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_231_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1034 ();
 FILLER_ASAP7_75t_R FILLER_231_1051 ();
 FILLER_ASAP7_75t_R FILLER_231_1063 ();
 DECAPx4_ASAP7_75t_R FILLER_231_1071 ();
 FILLER_ASAP7_75t_R FILLER_231_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1083 ();
 FILLER_ASAP7_75t_R FILLER_231_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_231_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1159 ();
 FILLER_ASAP7_75t_R FILLER_231_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1167 ();
 DECAPx4_ASAP7_75t_R FILLER_231_1171 ();
 FILLER_ASAP7_75t_R FILLER_231_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_231_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1204 ();
 DECAPx1_ASAP7_75t_R FILLER_231_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1221 ();
 DECAPx4_ASAP7_75t_R FILLER_231_1225 ();
 FILLER_ASAP7_75t_R FILLER_231_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1237 ();
 FILLER_ASAP7_75t_R FILLER_231_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1250 ();
 FILLER_ASAP7_75t_R FILLER_231_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1256 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1283 ();
 DECAPx1_ASAP7_75t_R FILLER_231_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1312 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1349 ();
 DECAPx6_ASAP7_75t_R FILLER_231_1371 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1385 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1391 ();
 DECAPx6_ASAP7_75t_R FILLER_232_2 ();
 DECAPx1_ASAP7_75t_R FILLER_232_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_20 ();
 DECAPx6_ASAP7_75t_R FILLER_232_47 ();
 FILLER_ASAP7_75t_R FILLER_232_61 ();
 FILLER_ASAP7_75t_R FILLER_232_115 ();
 DECAPx6_ASAP7_75t_R FILLER_232_129 ();
 DECAPx2_ASAP7_75t_R FILLER_232_143 ();
 FILLER_ASAP7_75t_R FILLER_232_156 ();
 DECAPx6_ASAP7_75t_R FILLER_232_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_184 ();
 DECAPx4_ASAP7_75t_R FILLER_232_191 ();
 DECAPx1_ASAP7_75t_R FILLER_232_204 ();
 DECAPx6_ASAP7_75t_R FILLER_232_240 ();
 FILLER_ASAP7_75t_R FILLER_232_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_256 ();
 FILLER_ASAP7_75t_R FILLER_232_265 ();
 FILLER_ASAP7_75t_R FILLER_232_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_275 ();
 DECAPx1_ASAP7_75t_R FILLER_232_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_292 ();
 DECAPx1_ASAP7_75t_R FILLER_232_299 ();
 DECAPx1_ASAP7_75t_R FILLER_232_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_332 ();
 DECAPx4_ASAP7_75t_R FILLER_232_359 ();
 FILLER_ASAP7_75t_R FILLER_232_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_389 ();
 FILLER_ASAP7_75t_R FILLER_232_411 ();
 DECAPx1_ASAP7_75t_R FILLER_232_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_431 ();
 DECAPx2_ASAP7_75t_R FILLER_232_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_450 ();
 DECAPx1_ASAP7_75t_R FILLER_232_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_461 ();
 FILLER_ASAP7_75t_R FILLER_232_464 ();
 DECAPx6_ASAP7_75t_R FILLER_232_480 ();
 DECAPx2_ASAP7_75t_R FILLER_232_502 ();
 FILLER_ASAP7_75t_R FILLER_232_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_510 ();
 DECAPx10_ASAP7_75t_R FILLER_232_525 ();
 DECAPx10_ASAP7_75t_R FILLER_232_547 ();
 FILLER_ASAP7_75t_R FILLER_232_569 ();
 DECAPx4_ASAP7_75t_R FILLER_232_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_584 ();
 DECAPx10_ASAP7_75t_R FILLER_232_591 ();
 DECAPx1_ASAP7_75t_R FILLER_232_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_617 ();
 DECAPx1_ASAP7_75t_R FILLER_232_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_625 ();
 DECAPx10_ASAP7_75t_R FILLER_232_652 ();
 DECAPx4_ASAP7_75t_R FILLER_232_674 ();
 FILLER_ASAP7_75t_R FILLER_232_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_686 ();
 DECAPx6_ASAP7_75t_R FILLER_232_791 ();
 DECAPx2_ASAP7_75t_R FILLER_232_805 ();
 DECAPx2_ASAP7_75t_R FILLER_232_827 ();
 DECAPx6_ASAP7_75t_R FILLER_232_848 ();
 DECAPx1_ASAP7_75t_R FILLER_232_862 ();
 DECAPx1_ASAP7_75t_R FILLER_232_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_876 ();
 DECAPx6_ASAP7_75t_R FILLER_232_892 ();
 FILLER_ASAP7_75t_R FILLER_232_906 ();
 FILLER_ASAP7_75t_R FILLER_232_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_924 ();
 DECAPx4_ASAP7_75t_R FILLER_232_934 ();
 DECAPx4_ASAP7_75t_R FILLER_232_950 ();
 FILLER_ASAP7_75t_R FILLER_232_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_962 ();
 DECAPx10_ASAP7_75t_R FILLER_232_977 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1030 ();
 FILLER_ASAP7_75t_R FILLER_232_1062 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1080 ();
 FILLER_ASAP7_75t_R FILLER_232_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1092 ();
 FILLER_ASAP7_75t_R FILLER_232_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_232_1103 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1130 ();
 FILLER_ASAP7_75t_R FILLER_232_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1205 ();
 DECAPx6_ASAP7_75t_R FILLER_232_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1263 ();
 FILLER_ASAP7_75t_R FILLER_232_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_232_1275 ();
 FILLER_ASAP7_75t_R FILLER_232_1325 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1332 ();
 FILLER_ASAP7_75t_R FILLER_232_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1378 ();
 FILLER_ASAP7_75t_R FILLER_232_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_233_2 ();
 DECAPx4_ASAP7_75t_R FILLER_233_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_34 ();
 DECAPx4_ASAP7_75t_R FILLER_233_68 ();
 DECAPx10_ASAP7_75t_R FILLER_233_81 ();
 FILLER_ASAP7_75t_R FILLER_233_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_138 ();
 DECAPx4_ASAP7_75t_R FILLER_233_165 ();
 FILLER_ASAP7_75t_R FILLER_233_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_177 ();
 DECAPx4_ASAP7_75t_R FILLER_233_186 ();
 FILLER_ASAP7_75t_R FILLER_233_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_198 ();
 DECAPx6_ASAP7_75t_R FILLER_233_205 ();
 FILLER_ASAP7_75t_R FILLER_233_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_221 ();
 FILLER_ASAP7_75t_R FILLER_233_225 ();
 DECAPx2_ASAP7_75t_R FILLER_233_241 ();
 FILLER_ASAP7_75t_R FILLER_233_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_266 ();
 DECAPx2_ASAP7_75t_R FILLER_233_281 ();
 DECAPx2_ASAP7_75t_R FILLER_233_313 ();
 DECAPx2_ASAP7_75t_R FILLER_233_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_331 ();
 DECAPx10_ASAP7_75t_R FILLER_233_338 ();
 DECAPx4_ASAP7_75t_R FILLER_233_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_370 ();
 DECAPx1_ASAP7_75t_R FILLER_233_389 ();
 DECAPx4_ASAP7_75t_R FILLER_233_401 ();
 DECAPx2_ASAP7_75t_R FILLER_233_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_432 ();
 DECAPx4_ASAP7_75t_R FILLER_233_455 ();
 FILLER_ASAP7_75t_R FILLER_233_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_467 ();
 DECAPx1_ASAP7_75t_R FILLER_233_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_480 ();
 DECAPx2_ASAP7_75t_R FILLER_233_489 ();
 DECAPx2_ASAP7_75t_R FILLER_233_501 ();
 FILLER_ASAP7_75t_R FILLER_233_516 ();
 DECAPx1_ASAP7_75t_R FILLER_233_524 ();
 DECAPx4_ASAP7_75t_R FILLER_233_531 ();
 DECAPx2_ASAP7_75t_R FILLER_233_549 ();
 FILLER_ASAP7_75t_R FILLER_233_555 ();
 DECAPx1_ASAP7_75t_R FILLER_233_581 ();
 DECAPx10_ASAP7_75t_R FILLER_233_617 ();
 FILLER_ASAP7_75t_R FILLER_233_639 ();
 DECAPx10_ASAP7_75t_R FILLER_233_644 ();
 DECAPx10_ASAP7_75t_R FILLER_233_666 ();
 DECAPx6_ASAP7_75t_R FILLER_233_688 ();
 FILLER_ASAP7_75t_R FILLER_233_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_704 ();
 DECAPx2_ASAP7_75t_R FILLER_233_708 ();
 FILLER_ASAP7_75t_R FILLER_233_714 ();
 DECAPx1_ASAP7_75t_R FILLER_233_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_727 ();
 DECAPx1_ASAP7_75t_R FILLER_233_731 ();
 DECAPx4_ASAP7_75t_R FILLER_233_741 ();
 FILLER_ASAP7_75t_R FILLER_233_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_753 ();
 DECAPx10_ASAP7_75t_R FILLER_233_757 ();
 DECAPx2_ASAP7_75t_R FILLER_233_779 ();
 FILLER_ASAP7_75t_R FILLER_233_785 ();
 DECAPx1_ASAP7_75t_R FILLER_233_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_817 ();
 FILLER_ASAP7_75t_R FILLER_233_824 ();
 DECAPx1_ASAP7_75t_R FILLER_233_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_833 ();
 DECAPx4_ASAP7_75t_R FILLER_233_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_861 ();
 DECAPx6_ASAP7_75t_R FILLER_233_878 ();
 DECAPx1_ASAP7_75t_R FILLER_233_892 ();
 FILLER_ASAP7_75t_R FILLER_233_922 ();
 DECAPx1_ASAP7_75t_R FILLER_233_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_940 ();
 FILLER_ASAP7_75t_R FILLER_233_965 ();
 FILLER_ASAP7_75t_R FILLER_233_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_995 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1023 ();
 DECAPx6_ASAP7_75t_R FILLER_233_1033 ();
 FILLER_ASAP7_75t_R FILLER_233_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1049 ();
 FILLER_ASAP7_75t_R FILLER_233_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1055 ();
 FILLER_ASAP7_75t_R FILLER_233_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_233_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1186 ();
 FILLER_ASAP7_75t_R FILLER_233_1193 ();
 FILLER_ASAP7_75t_R FILLER_233_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1239 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1250 ();
 FILLER_ASAP7_75t_R FILLER_233_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_233_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1309 ();
 FILLER_ASAP7_75t_R FILLER_233_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1317 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1324 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1386 ();
 DECAPx10_ASAP7_75t_R FILLER_234_2 ();
 DECAPx6_ASAP7_75t_R FILLER_234_24 ();
 FILLER_ASAP7_75t_R FILLER_234_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_82 ();
 DECAPx1_ASAP7_75t_R FILLER_234_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_93 ();
 FILLER_ASAP7_75t_R FILLER_234_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_102 ();
 FILLER_ASAP7_75t_R FILLER_234_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_146 ();
 FILLER_ASAP7_75t_R FILLER_234_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_152 ();
 DECAPx6_ASAP7_75t_R FILLER_234_156 ();
 FILLER_ASAP7_75t_R FILLER_234_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_172 ();
 DECAPx1_ASAP7_75t_R FILLER_234_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_242 ();
 DECAPx6_ASAP7_75t_R FILLER_234_257 ();
 FILLER_ASAP7_75t_R FILLER_234_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_273 ();
 DECAPx2_ASAP7_75t_R FILLER_234_282 ();
 FILLER_ASAP7_75t_R FILLER_234_288 ();
 DECAPx1_ASAP7_75t_R FILLER_234_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_300 ();
 DECAPx10_ASAP7_75t_R FILLER_234_310 ();
 DECAPx4_ASAP7_75t_R FILLER_234_332 ();
 DECAPx1_ASAP7_75t_R FILLER_234_352 ();
 DECAPx2_ASAP7_75t_R FILLER_234_374 ();
 FILLER_ASAP7_75t_R FILLER_234_380 ();
 DECAPx6_ASAP7_75t_R FILLER_234_396 ();
 DECAPx4_ASAP7_75t_R FILLER_234_426 ();
 FILLER_ASAP7_75t_R FILLER_234_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_438 ();
 DECAPx1_ASAP7_75t_R FILLER_234_442 ();
 DECAPx1_ASAP7_75t_R FILLER_234_458 ();
 FILLER_ASAP7_75t_R FILLER_234_480 ();
 DECAPx2_ASAP7_75t_R FILLER_234_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_497 ();
 DECAPx4_ASAP7_75t_R FILLER_234_501 ();
 FILLER_ASAP7_75t_R FILLER_234_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_513 ();
 FILLER_ASAP7_75t_R FILLER_234_540 ();
 DECAPx1_ASAP7_75t_R FILLER_234_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_554 ();
 DECAPx1_ASAP7_75t_R FILLER_234_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_609 ();
 DECAPx10_ASAP7_75t_R FILLER_234_636 ();
 DECAPx10_ASAP7_75t_R FILLER_234_658 ();
 DECAPx10_ASAP7_75t_R FILLER_234_680 ();
 DECAPx10_ASAP7_75t_R FILLER_234_702 ();
 DECAPx10_ASAP7_75t_R FILLER_234_724 ();
 DECAPx10_ASAP7_75t_R FILLER_234_746 ();
 DECAPx10_ASAP7_75t_R FILLER_234_768 ();
 DECAPx4_ASAP7_75t_R FILLER_234_790 ();
 FILLER_ASAP7_75t_R FILLER_234_800 ();
 DECAPx1_ASAP7_75t_R FILLER_234_805 ();
 FILLER_ASAP7_75t_R FILLER_234_819 ();
 DECAPx4_ASAP7_75t_R FILLER_234_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_892 ();
 FILLER_ASAP7_75t_R FILLER_234_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_905 ();
 DECAPx6_ASAP7_75t_R FILLER_234_931 ();
 DECAPx2_ASAP7_75t_R FILLER_234_955 ();
 FILLER_ASAP7_75t_R FILLER_234_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_963 ();
 DECAPx1_ASAP7_75t_R FILLER_234_972 ();
 FILLER_ASAP7_75t_R FILLER_234_979 ();
 DECAPx2_ASAP7_75t_R FILLER_234_984 ();
 FILLER_ASAP7_75t_R FILLER_234_990 ();
 DECAPx2_ASAP7_75t_R FILLER_234_1032 ();
 FILLER_ASAP7_75t_R FILLER_234_1038 ();
 DECAPx4_ASAP7_75t_R FILLER_234_1043 ();
 FILLER_ASAP7_75t_R FILLER_234_1053 ();
 DECAPx4_ASAP7_75t_R FILLER_234_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1091 ();
 DECAPx4_ASAP7_75t_R FILLER_234_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_234_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_234_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_234_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1163 ();
 FILLER_ASAP7_75t_R FILLER_234_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1192 ();
 DECAPx2_ASAP7_75t_R FILLER_234_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_234_1213 ();
 FILLER_ASAP7_75t_R FILLER_234_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1247 ();
 DECAPx6_ASAP7_75t_R FILLER_234_1280 ();
 DECAPx6_ASAP7_75t_R FILLER_234_1297 ();
 FILLER_ASAP7_75t_R FILLER_234_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_235_2 ();
 DECAPx10_ASAP7_75t_R FILLER_235_24 ();
 DECAPx2_ASAP7_75t_R FILLER_235_46 ();
 FILLER_ASAP7_75t_R FILLER_235_52 ();
 DECAPx2_ASAP7_75t_R FILLER_235_66 ();
 DECAPx2_ASAP7_75t_R FILLER_235_106 ();
 FILLER_ASAP7_75t_R FILLER_235_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_141 ();
 DECAPx1_ASAP7_75t_R FILLER_235_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_149 ();
 FILLER_ASAP7_75t_R FILLER_235_156 ();
 DECAPx1_ASAP7_75t_R FILLER_235_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_174 ();
 DECAPx6_ASAP7_75t_R FILLER_235_196 ();
 FILLER_ASAP7_75t_R FILLER_235_210 ();
 DECAPx10_ASAP7_75t_R FILLER_235_215 ();
 DECAPx2_ASAP7_75t_R FILLER_235_237 ();
 FILLER_ASAP7_75t_R FILLER_235_243 ();
 DECAPx1_ASAP7_75t_R FILLER_235_251 ();
 DECAPx4_ASAP7_75t_R FILLER_235_261 ();
 DECAPx4_ASAP7_75t_R FILLER_235_280 ();
 FILLER_ASAP7_75t_R FILLER_235_290 ();
 DECAPx1_ASAP7_75t_R FILLER_235_300 ();
 DECAPx1_ASAP7_75t_R FILLER_235_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_314 ();
 FILLER_ASAP7_75t_R FILLER_235_329 ();
 DECAPx6_ASAP7_75t_R FILLER_235_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_377 ();
 DECAPx2_ASAP7_75t_R FILLER_235_428 ();
 DECAPx2_ASAP7_75t_R FILLER_235_440 ();
 DECAPx6_ASAP7_75t_R FILLER_235_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_466 ();
 FILLER_ASAP7_75t_R FILLER_235_473 ();
 FILLER_ASAP7_75t_R FILLER_235_481 ();
 DECAPx1_ASAP7_75t_R FILLER_235_509 ();
 DECAPx2_ASAP7_75t_R FILLER_235_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_536 ();
 DECAPx2_ASAP7_75t_R FILLER_235_550 ();
 FILLER_ASAP7_75t_R FILLER_235_556 ();
 DECAPx10_ASAP7_75t_R FILLER_235_566 ();
 DECAPx1_ASAP7_75t_R FILLER_235_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_592 ();
 FILLER_ASAP7_75t_R FILLER_235_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_598 ();
 DECAPx2_ASAP7_75t_R FILLER_235_602 ();
 FILLER_ASAP7_75t_R FILLER_235_608 ();
 DECAPx2_ASAP7_75t_R FILLER_235_616 ();
 FILLER_ASAP7_75t_R FILLER_235_622 ();
 DECAPx1_ASAP7_75t_R FILLER_235_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_631 ();
 DECAPx10_ASAP7_75t_R FILLER_235_650 ();
 DECAPx10_ASAP7_75t_R FILLER_235_672 ();
 DECAPx10_ASAP7_75t_R FILLER_235_694 ();
 DECAPx10_ASAP7_75t_R FILLER_235_716 ();
 DECAPx10_ASAP7_75t_R FILLER_235_738 ();
 DECAPx10_ASAP7_75t_R FILLER_235_760 ();
 DECAPx2_ASAP7_75t_R FILLER_235_782 ();
 DECAPx4_ASAP7_75t_R FILLER_235_814 ();
 DECAPx2_ASAP7_75t_R FILLER_235_833 ();
 FILLER_ASAP7_75t_R FILLER_235_839 ();
 DECAPx4_ASAP7_75t_R FILLER_235_849 ();
 FILLER_ASAP7_75t_R FILLER_235_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_861 ();
 DECAPx6_ASAP7_75t_R FILLER_235_874 ();
 DECAPx2_ASAP7_75t_R FILLER_235_888 ();
 DECAPx6_ASAP7_75t_R FILLER_235_904 ();
 DECAPx2_ASAP7_75t_R FILLER_235_918 ();
 DECAPx6_ASAP7_75t_R FILLER_235_926 ();
 FILLER_ASAP7_75t_R FILLER_235_940 ();
 DECAPx4_ASAP7_75t_R FILLER_235_978 ();
 DECAPx1_ASAP7_75t_R FILLER_235_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_235_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_235_1069 ();
 FILLER_ASAP7_75t_R FILLER_235_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_235_1100 ();
 FILLER_ASAP7_75t_R FILLER_235_1106 ();
 DECAPx4_ASAP7_75t_R FILLER_235_1114 ();
 DECAPx4_ASAP7_75t_R FILLER_235_1129 ();
 FILLER_ASAP7_75t_R FILLER_235_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1141 ();
 FILLER_ASAP7_75t_R FILLER_235_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1154 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1182 ();
 FILLER_ASAP7_75t_R FILLER_235_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1233 ();
 DECAPx6_ASAP7_75t_R FILLER_235_1237 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1251 ();
 DECAPx2_ASAP7_75t_R FILLER_235_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1268 ();
 DECAPx4_ASAP7_75t_R FILLER_235_1285 ();
 DECAPx2_ASAP7_75t_R FILLER_235_1301 ();
 FILLER_ASAP7_75t_R FILLER_235_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1357 ();
 DECAPx4_ASAP7_75t_R FILLER_235_1379 ();
 FILLER_ASAP7_75t_R FILLER_235_1389 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_236_2 ();
 DECAPx10_ASAP7_75t_R FILLER_236_24 ();
 DECAPx10_ASAP7_75t_R FILLER_236_46 ();
 FILLER_ASAP7_75t_R FILLER_236_68 ();
 DECAPx2_ASAP7_75t_R FILLER_236_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_79 ();
 DECAPx1_ASAP7_75t_R FILLER_236_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_90 ();
 FILLER_ASAP7_75t_R FILLER_236_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_96 ();
 FILLER_ASAP7_75t_R FILLER_236_103 ();
 DECAPx1_ASAP7_75t_R FILLER_236_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_112 ();
 DECAPx4_ASAP7_75t_R FILLER_236_117 ();
 FILLER_ASAP7_75t_R FILLER_236_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_129 ();
 DECAPx4_ASAP7_75t_R FILLER_236_133 ();
 FILLER_ASAP7_75t_R FILLER_236_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_153 ();
 DECAPx2_ASAP7_75t_R FILLER_236_180 ();
 DECAPx2_ASAP7_75t_R FILLER_236_195 ();
 DECAPx6_ASAP7_75t_R FILLER_236_204 ();
 DECAPx2_ASAP7_75t_R FILLER_236_218 ();
 DECAPx6_ASAP7_75t_R FILLER_236_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_254 ();
 DECAPx1_ASAP7_75t_R FILLER_236_281 ();
 FILLER_ASAP7_75t_R FILLER_236_311 ();
 DECAPx1_ASAP7_75t_R FILLER_236_339 ();
 DECAPx6_ASAP7_75t_R FILLER_236_369 ();
 FILLER_ASAP7_75t_R FILLER_236_383 ();
 FILLER_ASAP7_75t_R FILLER_236_391 ();
 DECAPx10_ASAP7_75t_R FILLER_236_396 ();
 DECAPx4_ASAP7_75t_R FILLER_236_418 ();
 DECAPx2_ASAP7_75t_R FILLER_236_454 ();
 FILLER_ASAP7_75t_R FILLER_236_460 ();
 DECAPx2_ASAP7_75t_R FILLER_236_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_483 ();
 DECAPx1_ASAP7_75t_R FILLER_236_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_494 ();
 DECAPx6_ASAP7_75t_R FILLER_236_527 ();
 FILLER_ASAP7_75t_R FILLER_236_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_549 ();
 DECAPx6_ASAP7_75t_R FILLER_236_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_585 ();
 DECAPx2_ASAP7_75t_R FILLER_236_589 ();
 FILLER_ASAP7_75t_R FILLER_236_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_597 ();
 DECAPx10_ASAP7_75t_R FILLER_236_616 ();
 DECAPx10_ASAP7_75t_R FILLER_236_638 ();
 DECAPx10_ASAP7_75t_R FILLER_236_660 ();
 DECAPx10_ASAP7_75t_R FILLER_236_682 ();
 DECAPx10_ASAP7_75t_R FILLER_236_704 ();
 DECAPx10_ASAP7_75t_R FILLER_236_726 ();
 DECAPx10_ASAP7_75t_R FILLER_236_748 ();
 DECAPx10_ASAP7_75t_R FILLER_236_770 ();
 DECAPx4_ASAP7_75t_R FILLER_236_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_802 ();
 DECAPx4_ASAP7_75t_R FILLER_236_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_816 ();
 DECAPx10_ASAP7_75t_R FILLER_236_823 ();
 DECAPx6_ASAP7_75t_R FILLER_236_845 ();
 DECAPx2_ASAP7_75t_R FILLER_236_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_865 ();
 DECAPx2_ASAP7_75t_R FILLER_236_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_878 ();
 DECAPx2_ASAP7_75t_R FILLER_236_887 ();
 FILLER_ASAP7_75t_R FILLER_236_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_905 ();
 DECAPx10_ASAP7_75t_R FILLER_236_938 ();
 DECAPx6_ASAP7_75t_R FILLER_236_960 ();
 DECAPx2_ASAP7_75t_R FILLER_236_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_980 ();
 DECAPx2_ASAP7_75t_R FILLER_236_989 ();
 FILLER_ASAP7_75t_R FILLER_236_995 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1039 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1043 ();
 FILLER_ASAP7_75t_R FILLER_236_1057 ();
 FILLER_ASAP7_75t_R FILLER_236_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1179 ();
 FILLER_ASAP7_75t_R FILLER_236_1196 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1224 ();
 FILLER_ASAP7_75t_R FILLER_236_1238 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1250 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1268 ();
 FILLER_ASAP7_75t_R FILLER_236_1276 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1349 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_237_2 ();
 DECAPx10_ASAP7_75t_R FILLER_237_24 ();
 DECAPx10_ASAP7_75t_R FILLER_237_46 ();
 DECAPx10_ASAP7_75t_R FILLER_237_68 ();
 FILLER_ASAP7_75t_R FILLER_237_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_118 ();
 FILLER_ASAP7_75t_R FILLER_237_125 ();
 DECAPx2_ASAP7_75t_R FILLER_237_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_139 ();
 FILLER_ASAP7_75t_R FILLER_237_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_168 ();
 DECAPx6_ASAP7_75t_R FILLER_237_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_186 ();
 DECAPx2_ASAP7_75t_R FILLER_237_245 ();
 FILLER_ASAP7_75t_R FILLER_237_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_253 ();
 DECAPx2_ASAP7_75t_R FILLER_237_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_269 ();
 DECAPx6_ASAP7_75t_R FILLER_237_279 ();
 DECAPx2_ASAP7_75t_R FILLER_237_293 ();
 DECAPx4_ASAP7_75t_R FILLER_237_302 ();
 FILLER_ASAP7_75t_R FILLER_237_312 ();
 DECAPx6_ASAP7_75t_R FILLER_237_335 ();
 DECAPx1_ASAP7_75t_R FILLER_237_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_353 ();
 DECAPx1_ASAP7_75t_R FILLER_237_363 ();
 FILLER_ASAP7_75t_R FILLER_237_393 ();
 FILLER_ASAP7_75t_R FILLER_237_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_409 ();
 FILLER_ASAP7_75t_R FILLER_237_413 ();
 DECAPx1_ASAP7_75t_R FILLER_237_422 ();
 DECAPx1_ASAP7_75t_R FILLER_237_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_442 ();
 FILLER_ASAP7_75t_R FILLER_237_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_448 ();
 DECAPx1_ASAP7_75t_R FILLER_237_452 ();
 DECAPx1_ASAP7_75t_R FILLER_237_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_486 ();
 DECAPx4_ASAP7_75t_R FILLER_237_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_503 ();
 DECAPx2_ASAP7_75t_R FILLER_237_510 ();
 DECAPx1_ASAP7_75t_R FILLER_237_519 ();
 DECAPx2_ASAP7_75t_R FILLER_237_529 ();
 DECAPx6_ASAP7_75t_R FILLER_237_541 ();
 DECAPx1_ASAP7_75t_R FILLER_237_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_627 ();
 DECAPx10_ASAP7_75t_R FILLER_237_646 ();
 DECAPx10_ASAP7_75t_R FILLER_237_668 ();
 DECAPx10_ASAP7_75t_R FILLER_237_690 ();
 DECAPx10_ASAP7_75t_R FILLER_237_712 ();
 DECAPx10_ASAP7_75t_R FILLER_237_734 ();
 DECAPx10_ASAP7_75t_R FILLER_237_756 ();
 DECAPx2_ASAP7_75t_R FILLER_237_778 ();
 DECAPx1_ASAP7_75t_R FILLER_237_810 ();
 FILLER_ASAP7_75t_R FILLER_237_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_830 ();
 DECAPx6_ASAP7_75t_R FILLER_237_840 ();
 DECAPx1_ASAP7_75t_R FILLER_237_854 ();
 DECAPx2_ASAP7_75t_R FILLER_237_867 ();
 FILLER_ASAP7_75t_R FILLER_237_873 ();
 DECAPx1_ASAP7_75t_R FILLER_237_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_889 ();
 DECAPx6_ASAP7_75t_R FILLER_237_893 ();
 FILLER_ASAP7_75t_R FILLER_237_907 ();
 DECAPx4_ASAP7_75t_R FILLER_237_965 ();
 DECAPx6_ASAP7_75t_R FILLER_237_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1011 ();
 FILLER_ASAP7_75t_R FILLER_237_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1035 ();
 FILLER_ASAP7_75t_R FILLER_237_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1093 ();
 FILLER_ASAP7_75t_R FILLER_237_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1101 ();
 FILLER_ASAP7_75t_R FILLER_237_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1119 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1155 ();
 FILLER_ASAP7_75t_R FILLER_237_1165 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1170 ();
 FILLER_ASAP7_75t_R FILLER_237_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1219 ();
 DECAPx1_ASAP7_75t_R FILLER_237_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1239 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1386 ();
 DECAPx10_ASAP7_75t_R FILLER_238_2 ();
 DECAPx10_ASAP7_75t_R FILLER_238_24 ();
 DECAPx10_ASAP7_75t_R FILLER_238_46 ();
 DECAPx10_ASAP7_75t_R FILLER_238_68 ();
 FILLER_ASAP7_75t_R FILLER_238_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_92 ();
 DECAPx6_ASAP7_75t_R FILLER_238_99 ();
 DECAPx1_ASAP7_75t_R FILLER_238_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_154 ();
 DECAPx4_ASAP7_75t_R FILLER_238_158 ();
 FILLER_ASAP7_75t_R FILLER_238_168 ();
 FILLER_ASAP7_75t_R FILLER_238_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_184 ();
 DECAPx6_ASAP7_75t_R FILLER_238_188 ();
 DECAPx1_ASAP7_75t_R FILLER_238_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_206 ();
 FILLER_ASAP7_75t_R FILLER_238_237 ();
 FILLER_ASAP7_75t_R FILLER_238_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_247 ();
 FILLER_ASAP7_75t_R FILLER_238_283 ();
 DECAPx4_ASAP7_75t_R FILLER_238_300 ();
 DECAPx10_ASAP7_75t_R FILLER_238_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_335 ();
 DECAPx1_ASAP7_75t_R FILLER_238_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_358 ();
 DECAPx1_ASAP7_75t_R FILLER_238_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_387 ();
 FILLER_ASAP7_75t_R FILLER_238_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_416 ();
 DECAPx1_ASAP7_75t_R FILLER_238_424 ();
 DECAPx2_ASAP7_75t_R FILLER_238_434 ();
 FILLER_ASAP7_75t_R FILLER_238_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_442 ();
 DECAPx4_ASAP7_75t_R FILLER_238_446 ();
 FILLER_ASAP7_75t_R FILLER_238_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_478 ();
 FILLER_ASAP7_75t_R FILLER_238_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_487 ();
 DECAPx1_ASAP7_75t_R FILLER_238_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_501 ();
 DECAPx6_ASAP7_75t_R FILLER_238_508 ();
 FILLER_ASAP7_75t_R FILLER_238_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_524 ();
 DECAPx1_ASAP7_75t_R FILLER_238_528 ();
 DECAPx2_ASAP7_75t_R FILLER_238_588 ();
 FILLER_ASAP7_75t_R FILLER_238_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_603 ();
 DECAPx10_ASAP7_75t_R FILLER_238_636 ();
 DECAPx10_ASAP7_75t_R FILLER_238_658 ();
 DECAPx10_ASAP7_75t_R FILLER_238_680 ();
 DECAPx10_ASAP7_75t_R FILLER_238_702 ();
 DECAPx10_ASAP7_75t_R FILLER_238_724 ();
 DECAPx10_ASAP7_75t_R FILLER_238_746 ();
 DECAPx10_ASAP7_75t_R FILLER_238_768 ();
 DECAPx2_ASAP7_75t_R FILLER_238_790 ();
 FILLER_ASAP7_75t_R FILLER_238_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_798 ();
 DECAPx2_ASAP7_75t_R FILLER_238_802 ();
 FILLER_ASAP7_75t_R FILLER_238_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_824 ();
 FILLER_ASAP7_75t_R FILLER_238_839 ();
 FILLER_ASAP7_75t_R FILLER_238_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_853 ();
 FILLER_ASAP7_75t_R FILLER_238_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_869 ();
 FILLER_ASAP7_75t_R FILLER_238_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_921 ();
 DECAPx1_ASAP7_75t_R FILLER_238_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_932 ();
 DECAPx4_ASAP7_75t_R FILLER_238_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_959 ();
 DECAPx1_ASAP7_75t_R FILLER_238_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_974 ();
 FILLER_ASAP7_75t_R FILLER_238_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1003 ();
 FILLER_ASAP7_75t_R FILLER_238_1030 ();
 DECAPx6_ASAP7_75t_R FILLER_238_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1093 ();
 FILLER_ASAP7_75t_R FILLER_238_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1136 ();
 FILLER_ASAP7_75t_R FILLER_238_1142 ();
 FILLER_ASAP7_75t_R FILLER_238_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_238_1157 ();
 FILLER_ASAP7_75t_R FILLER_238_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1244 ();
 DECAPx4_ASAP7_75t_R FILLER_238_1266 ();
 FILLER_ASAP7_75t_R FILLER_238_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_238_1370 ();
 FILLER_ASAP7_75t_R FILLER_238_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_239_2 ();
 DECAPx10_ASAP7_75t_R FILLER_239_24 ();
 DECAPx10_ASAP7_75t_R FILLER_239_46 ();
 DECAPx10_ASAP7_75t_R FILLER_239_68 ();
 DECAPx10_ASAP7_75t_R FILLER_239_90 ();
 DECAPx6_ASAP7_75t_R FILLER_239_112 ();
 FILLER_ASAP7_75t_R FILLER_239_126 ();
 DECAPx4_ASAP7_75t_R FILLER_239_131 ();
 FILLER_ASAP7_75t_R FILLER_239_141 ();
 FILLER_ASAP7_75t_R FILLER_239_169 ();
 DECAPx4_ASAP7_75t_R FILLER_239_200 ();
 DECAPx2_ASAP7_75t_R FILLER_239_216 ();
 DECAPx4_ASAP7_75t_R FILLER_239_225 ();
 DECAPx4_ASAP7_75t_R FILLER_239_261 ();
 DECAPx2_ASAP7_75t_R FILLER_239_297 ();
 DECAPx4_ASAP7_75t_R FILLER_239_315 ();
 FILLER_ASAP7_75t_R FILLER_239_325 ();
 FILLER_ASAP7_75t_R FILLER_239_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_332 ();
 FILLER_ASAP7_75t_R FILLER_239_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_361 ();
 DECAPx4_ASAP7_75t_R FILLER_239_388 ();
 DECAPx1_ASAP7_75t_R FILLER_239_425 ();
 DECAPx6_ASAP7_75t_R FILLER_239_455 ();
 DECAPx1_ASAP7_75t_R FILLER_239_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_473 ();
 FILLER_ASAP7_75t_R FILLER_239_503 ();
 DECAPx1_ASAP7_75t_R FILLER_239_513 ();
 DECAPx2_ASAP7_75t_R FILLER_239_537 ();
 DECAPx6_ASAP7_75t_R FILLER_239_559 ();
 DECAPx1_ASAP7_75t_R FILLER_239_573 ();
 DECAPx2_ASAP7_75t_R FILLER_239_580 ();
 DECAPx2_ASAP7_75t_R FILLER_239_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_610 ();
 DECAPx10_ASAP7_75t_R FILLER_239_614 ();
 DECAPx10_ASAP7_75t_R FILLER_239_636 ();
 DECAPx10_ASAP7_75t_R FILLER_239_658 ();
 DECAPx10_ASAP7_75t_R FILLER_239_680 ();
 DECAPx10_ASAP7_75t_R FILLER_239_702 ();
 DECAPx10_ASAP7_75t_R FILLER_239_724 ();
 DECAPx10_ASAP7_75t_R FILLER_239_746 ();
 DECAPx6_ASAP7_75t_R FILLER_239_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_782 ();
 DECAPx2_ASAP7_75t_R FILLER_239_823 ();
 FILLER_ASAP7_75t_R FILLER_239_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_872 ();
 DECAPx4_ASAP7_75t_R FILLER_239_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_897 ();
 FILLER_ASAP7_75t_R FILLER_239_912 ();
 DECAPx1_ASAP7_75t_R FILLER_239_920 ();
 FILLER_ASAP7_75t_R FILLER_239_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_928 ();
 DECAPx6_ASAP7_75t_R FILLER_239_942 ();
 DECAPx2_ASAP7_75t_R FILLER_239_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_995 ();
 FILLER_ASAP7_75t_R FILLER_239_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_239_1054 ();
 DECAPx1_ASAP7_75t_R FILLER_239_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_239_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_239_1101 ();
 FILLER_ASAP7_75t_R FILLER_239_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1125 ();
 FILLER_ASAP7_75t_R FILLER_239_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1355 ();
 DECAPx6_ASAP7_75t_R FILLER_239_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_240_2 ();
 DECAPx10_ASAP7_75t_R FILLER_240_24 ();
 DECAPx10_ASAP7_75t_R FILLER_240_46 ();
 DECAPx10_ASAP7_75t_R FILLER_240_68 ();
 FILLER_ASAP7_75t_R FILLER_240_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_92 ();
 DECAPx1_ASAP7_75t_R FILLER_240_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_133 ();
 DECAPx1_ASAP7_75t_R FILLER_240_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_144 ();
 DECAPx2_ASAP7_75t_R FILLER_240_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_157 ();
 DECAPx2_ASAP7_75t_R FILLER_240_161 ();
 DECAPx6_ASAP7_75t_R FILLER_240_171 ();
 FILLER_ASAP7_75t_R FILLER_240_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_191 ();
 DECAPx2_ASAP7_75t_R FILLER_240_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_210 ();
 DECAPx6_ASAP7_75t_R FILLER_240_217 ();
 DECAPx2_ASAP7_75t_R FILLER_240_231 ();
 DECAPx2_ASAP7_75t_R FILLER_240_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_252 ();
 DECAPx2_ASAP7_75t_R FILLER_240_259 ();
 FILLER_ASAP7_75t_R FILLER_240_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_267 ();
 FILLER_ASAP7_75t_R FILLER_240_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_273 ();
 DECAPx2_ASAP7_75t_R FILLER_240_280 ();
 DECAPx4_ASAP7_75t_R FILLER_240_289 ();
 FILLER_ASAP7_75t_R FILLER_240_299 ();
 DECAPx4_ASAP7_75t_R FILLER_240_335 ();
 FILLER_ASAP7_75t_R FILLER_240_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_351 ();
 DECAPx6_ASAP7_75t_R FILLER_240_358 ();
 DECAPx1_ASAP7_75t_R FILLER_240_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_380 ();
 DECAPx4_ASAP7_75t_R FILLER_240_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_420 ();
 DECAPx10_ASAP7_75t_R FILLER_240_427 ();
 DECAPx2_ASAP7_75t_R FILLER_240_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_461 ();
 DECAPx1_ASAP7_75t_R FILLER_240_464 ();
 DECAPx4_ASAP7_75t_R FILLER_240_471 ();
 FILLER_ASAP7_75t_R FILLER_240_481 ();
 FILLER_ASAP7_75t_R FILLER_240_489 ();
 DECAPx2_ASAP7_75t_R FILLER_240_494 ();
 DECAPx6_ASAP7_75t_R FILLER_240_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_546 ();
 DECAPx1_ASAP7_75t_R FILLER_240_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_554 ();
 DECAPx6_ASAP7_75t_R FILLER_240_564 ();
 DECAPx1_ASAP7_75t_R FILLER_240_578 ();
 DECAPx6_ASAP7_75t_R FILLER_240_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_606 ();
 DECAPx10_ASAP7_75t_R FILLER_240_617 ();
 DECAPx10_ASAP7_75t_R FILLER_240_639 ();
 DECAPx10_ASAP7_75t_R FILLER_240_661 ();
 DECAPx10_ASAP7_75t_R FILLER_240_683 ();
 DECAPx10_ASAP7_75t_R FILLER_240_705 ();
 DECAPx10_ASAP7_75t_R FILLER_240_727 ();
 DECAPx10_ASAP7_75t_R FILLER_240_749 ();
 DECAPx10_ASAP7_75t_R FILLER_240_771 ();
 DECAPx1_ASAP7_75t_R FILLER_240_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_800 ();
 DECAPx2_ASAP7_75t_R FILLER_240_825 ();
 FILLER_ASAP7_75t_R FILLER_240_831 ();
 DECAPx1_ASAP7_75t_R FILLER_240_839 ();
 DECAPx2_ASAP7_75t_R FILLER_240_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_855 ();
 FILLER_ASAP7_75t_R FILLER_240_874 ();
 DECAPx6_ASAP7_75t_R FILLER_240_882 ();
 DECAPx6_ASAP7_75t_R FILLER_240_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_923 ();
 DECAPx1_ASAP7_75t_R FILLER_240_931 ();
 DECAPx2_ASAP7_75t_R FILLER_240_948 ();
 DECAPx6_ASAP7_75t_R FILLER_240_957 ();
 DECAPx2_ASAP7_75t_R FILLER_240_971 ();
 DECAPx6_ASAP7_75t_R FILLER_240_987 ();
 DECAPx2_ASAP7_75t_R FILLER_240_1011 ();
 FILLER_ASAP7_75t_R FILLER_240_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1019 ();
 DECAPx4_ASAP7_75t_R FILLER_240_1023 ();
 FILLER_ASAP7_75t_R FILLER_240_1033 ();
 FILLER_ASAP7_75t_R FILLER_240_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_240_1074 ();
 FILLER_ASAP7_75t_R FILLER_240_1080 ();
 FILLER_ASAP7_75t_R FILLER_240_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1110 ();
 DECAPx4_ASAP7_75t_R FILLER_240_1137 ();
 FILLER_ASAP7_75t_R FILLER_240_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_240_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1349 ();
 DECAPx6_ASAP7_75t_R FILLER_240_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_241_2 ();
 DECAPx10_ASAP7_75t_R FILLER_241_24 ();
 DECAPx10_ASAP7_75t_R FILLER_241_46 ();
 DECAPx10_ASAP7_75t_R FILLER_241_68 ();
 DECAPx10_ASAP7_75t_R FILLER_241_90 ();
 FILLER_ASAP7_75t_R FILLER_241_112 ();
 FILLER_ASAP7_75t_R FILLER_241_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_152 ();
 DECAPx1_ASAP7_75t_R FILLER_241_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_160 ();
 DECAPx2_ASAP7_75t_R FILLER_241_167 ();
 DECAPx1_ASAP7_75t_R FILLER_241_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_203 ();
 DECAPx1_ASAP7_75t_R FILLER_241_239 ();
 DECAPx1_ASAP7_75t_R FILLER_241_251 ();
 DECAPx2_ASAP7_75t_R FILLER_241_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_292 ();
 DECAPx1_ASAP7_75t_R FILLER_241_319 ();
 DECAPx1_ASAP7_75t_R FILLER_241_326 ();
 FILLER_ASAP7_75t_R FILLER_241_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_358 ();
 DECAPx10_ASAP7_75t_R FILLER_241_365 ();
 DECAPx10_ASAP7_75t_R FILLER_241_387 ();
 DECAPx6_ASAP7_75t_R FILLER_241_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_426 ();
 FILLER_ASAP7_75t_R FILLER_241_440 ();
 FILLER_ASAP7_75t_R FILLER_241_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_447 ();
 DECAPx6_ASAP7_75t_R FILLER_241_480 ();
 DECAPx2_ASAP7_75t_R FILLER_241_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_500 ();
 FILLER_ASAP7_75t_R FILLER_241_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_506 ();
 DECAPx2_ASAP7_75t_R FILLER_241_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_519 ();
 DECAPx6_ASAP7_75t_R FILLER_241_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_537 ();
 FILLER_ASAP7_75t_R FILLER_241_556 ();
 DECAPx1_ASAP7_75t_R FILLER_241_584 ();
 DECAPx1_ASAP7_75t_R FILLER_241_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_602 ();
 DECAPx10_ASAP7_75t_R FILLER_241_613 ();
 DECAPx10_ASAP7_75t_R FILLER_241_635 ();
 DECAPx10_ASAP7_75t_R FILLER_241_657 ();
 DECAPx10_ASAP7_75t_R FILLER_241_679 ();
 DECAPx10_ASAP7_75t_R FILLER_241_701 ();
 DECAPx10_ASAP7_75t_R FILLER_241_723 ();
 DECAPx10_ASAP7_75t_R FILLER_241_745 ();
 DECAPx10_ASAP7_75t_R FILLER_241_767 ();
 DECAPx2_ASAP7_75t_R FILLER_241_789 ();
 FILLER_ASAP7_75t_R FILLER_241_795 ();
 DECAPx4_ASAP7_75t_R FILLER_241_800 ();
 DECAPx10_ASAP7_75t_R FILLER_241_819 ();
 DECAPx10_ASAP7_75t_R FILLER_241_841 ();
 DECAPx10_ASAP7_75t_R FILLER_241_863 ();
 DECAPx1_ASAP7_75t_R FILLER_241_885 ();
 DECAPx2_ASAP7_75t_R FILLER_241_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_916 ();
 FILLER_ASAP7_75t_R FILLER_241_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_928 ();
 FILLER_ASAP7_75t_R FILLER_241_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_939 ();
 DECAPx10_ASAP7_75t_R FILLER_241_966 ();
 DECAPx10_ASAP7_75t_R FILLER_241_988 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_241_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1058 ();
 DECAPx6_ASAP7_75t_R FILLER_241_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_241_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_241_1087 ();
 FILLER_ASAP7_75t_R FILLER_241_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_241_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_241_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1348 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1370 ();
 DECAPx10_ASAP7_75t_R FILLER_242_2 ();
 DECAPx10_ASAP7_75t_R FILLER_242_24 ();
 DECAPx10_ASAP7_75t_R FILLER_242_46 ();
 DECAPx10_ASAP7_75t_R FILLER_242_68 ();
 DECAPx10_ASAP7_75t_R FILLER_242_90 ();
 DECAPx4_ASAP7_75t_R FILLER_242_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_155 ();
 DECAPx4_ASAP7_75t_R FILLER_242_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_196 ();
 DECAPx1_ASAP7_75t_R FILLER_242_204 ();
 DECAPx1_ASAP7_75t_R FILLER_242_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_222 ();
 DECAPx1_ASAP7_75t_R FILLER_242_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_262 ();
 FILLER_ASAP7_75t_R FILLER_242_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_268 ();
 FILLER_ASAP7_75t_R FILLER_242_281 ();
 DECAPx4_ASAP7_75t_R FILLER_242_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_383 ();
 DECAPx2_ASAP7_75t_R FILLER_242_393 ();
 FILLER_ASAP7_75t_R FILLER_242_399 ();
 FILLER_ASAP7_75t_R FILLER_242_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_410 ();
 DECAPx1_ASAP7_75t_R FILLER_242_414 ();
 FILLER_ASAP7_75t_R FILLER_242_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_426 ();
 FILLER_ASAP7_75t_R FILLER_242_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_455 ();
 FILLER_ASAP7_75t_R FILLER_242_464 ();
 FILLER_ASAP7_75t_R FILLER_242_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_483 ();
 DECAPx4_ASAP7_75t_R FILLER_242_508 ();
 FILLER_ASAP7_75t_R FILLER_242_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_520 ();
 DECAPx6_ASAP7_75t_R FILLER_242_530 ();
 FILLER_ASAP7_75t_R FILLER_242_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_553 ();
 DECAPx4_ASAP7_75t_R FILLER_242_560 ();
 FILLER_ASAP7_75t_R FILLER_242_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_572 ();
 DECAPx10_ASAP7_75t_R FILLER_242_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_598 ();
 DECAPx2_ASAP7_75t_R FILLER_242_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_625 ();
 DECAPx10_ASAP7_75t_R FILLER_242_644 ();
 DECAPx10_ASAP7_75t_R FILLER_242_666 ();
 DECAPx10_ASAP7_75t_R FILLER_242_688 ();
 DECAPx10_ASAP7_75t_R FILLER_242_710 ();
 DECAPx10_ASAP7_75t_R FILLER_242_732 ();
 DECAPx10_ASAP7_75t_R FILLER_242_754 ();
 DECAPx2_ASAP7_75t_R FILLER_242_776 ();
 FILLER_ASAP7_75t_R FILLER_242_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_810 ();
 DECAPx1_ASAP7_75t_R FILLER_242_829 ();
 DECAPx4_ASAP7_75t_R FILLER_242_842 ();
 DECAPx6_ASAP7_75t_R FILLER_242_861 ();
 DECAPx1_ASAP7_75t_R FILLER_242_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_879 ();
 DECAPx1_ASAP7_75t_R FILLER_242_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_920 ();
 DECAPx6_ASAP7_75t_R FILLER_242_927 ();
 DECAPx1_ASAP7_75t_R FILLER_242_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_945 ();
 FILLER_ASAP7_75t_R FILLER_242_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_958 ();
 DECAPx2_ASAP7_75t_R FILLER_242_969 ();
 DECAPx1_ASAP7_75t_R FILLER_242_993 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_242_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1045 ();
 FILLER_ASAP7_75t_R FILLER_242_1051 ();
 FILLER_ASAP7_75t_R FILLER_242_1069 ();
 FILLER_ASAP7_75t_R FILLER_242_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1081 ();
 FILLER_ASAP7_75t_R FILLER_242_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1123 ();
 DECAPx4_ASAP7_75t_R FILLER_242_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1347 ();
 DECAPx6_ASAP7_75t_R FILLER_242_1369 ();
 FILLER_ASAP7_75t_R FILLER_242_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_242_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_243_2 ();
 DECAPx10_ASAP7_75t_R FILLER_243_24 ();
 DECAPx10_ASAP7_75t_R FILLER_243_46 ();
 DECAPx10_ASAP7_75t_R FILLER_243_68 ();
 DECAPx10_ASAP7_75t_R FILLER_243_90 ();
 DECAPx6_ASAP7_75t_R FILLER_243_112 ();
 DECAPx1_ASAP7_75t_R FILLER_243_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_130 ();
 DECAPx1_ASAP7_75t_R FILLER_243_140 ();
 DECAPx4_ASAP7_75t_R FILLER_243_147 ();
 DECAPx6_ASAP7_75t_R FILLER_243_179 ();
 FILLER_ASAP7_75t_R FILLER_243_193 ();
 DECAPx2_ASAP7_75t_R FILLER_243_221 ();
 FILLER_ASAP7_75t_R FILLER_243_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_237 ();
 FILLER_ASAP7_75t_R FILLER_243_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_305 ();
 FILLER_ASAP7_75t_R FILLER_243_312 ();
 DECAPx6_ASAP7_75t_R FILLER_243_327 ();
 DECAPx1_ASAP7_75t_R FILLER_243_341 ();
 DECAPx2_ASAP7_75t_R FILLER_243_348 ();
 DECAPx1_ASAP7_75t_R FILLER_243_361 ();
 FILLER_ASAP7_75t_R FILLER_243_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_370 ();
 DECAPx1_ASAP7_75t_R FILLER_243_423 ();
 FILLER_ASAP7_75t_R FILLER_243_440 ();
 DECAPx2_ASAP7_75t_R FILLER_243_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_451 ();
 DECAPx1_ASAP7_75t_R FILLER_243_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_482 ();
 DECAPx1_ASAP7_75t_R FILLER_243_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_519 ();
 DECAPx1_ASAP7_75t_R FILLER_243_546 ();
 DECAPx6_ASAP7_75t_R FILLER_243_576 ();
 FILLER_ASAP7_75t_R FILLER_243_590 ();
 DECAPx6_ASAP7_75t_R FILLER_243_602 ();
 DECAPx1_ASAP7_75t_R FILLER_243_616 ();
 DECAPx10_ASAP7_75t_R FILLER_243_638 ();
 DECAPx10_ASAP7_75t_R FILLER_243_660 ();
 DECAPx10_ASAP7_75t_R FILLER_243_682 ();
 DECAPx10_ASAP7_75t_R FILLER_243_704 ();
 DECAPx10_ASAP7_75t_R FILLER_243_726 ();
 DECAPx10_ASAP7_75t_R FILLER_243_748 ();
 DECAPx10_ASAP7_75t_R FILLER_243_770 ();
 DECAPx2_ASAP7_75t_R FILLER_243_792 ();
 DECAPx2_ASAP7_75t_R FILLER_243_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_807 ();
 DECAPx2_ASAP7_75t_R FILLER_243_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_832 ();
 DECAPx1_ASAP7_75t_R FILLER_243_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_863 ();
 DECAPx2_ASAP7_75t_R FILLER_243_890 ();
 FILLER_ASAP7_75t_R FILLER_243_896 ();
 DECAPx1_ASAP7_75t_R FILLER_243_904 ();
 DECAPx4_ASAP7_75t_R FILLER_243_911 ();
 DECAPx2_ASAP7_75t_R FILLER_243_926 ();
 FILLER_ASAP7_75t_R FILLER_243_932 ();
 DECAPx6_ASAP7_75t_R FILLER_243_944 ();
 DECAPx2_ASAP7_75t_R FILLER_243_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_243_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1036 ();
 DECAPx6_ASAP7_75t_R FILLER_243_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_243_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1085 ();
 DECAPx1_ASAP7_75t_R FILLER_243_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_243_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1110 ();
 DECAPx4_ASAP7_75t_R FILLER_243_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1125 ();
 FILLER_ASAP7_75t_R FILLER_243_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_243_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1353 ();
 DECAPx6_ASAP7_75t_R FILLER_243_1375 ();
 FILLER_ASAP7_75t_R FILLER_243_1389 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_244_2 ();
 DECAPx10_ASAP7_75t_R FILLER_244_24 ();
 DECAPx10_ASAP7_75t_R FILLER_244_46 ();
 DECAPx10_ASAP7_75t_R FILLER_244_68 ();
 DECAPx10_ASAP7_75t_R FILLER_244_90 ();
 DECAPx10_ASAP7_75t_R FILLER_244_112 ();
 DECAPx10_ASAP7_75t_R FILLER_244_134 ();
 DECAPx1_ASAP7_75t_R FILLER_244_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_160 ();
 DECAPx2_ASAP7_75t_R FILLER_244_193 ();
 FILLER_ASAP7_75t_R FILLER_244_199 ();
 FILLER_ASAP7_75t_R FILLER_244_207 ();
 DECAPx10_ASAP7_75t_R FILLER_244_212 ();
 DECAPx10_ASAP7_75t_R FILLER_244_234 ();
 DECAPx6_ASAP7_75t_R FILLER_244_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_270 ();
 DECAPx1_ASAP7_75t_R FILLER_244_277 ();
 DECAPx1_ASAP7_75t_R FILLER_244_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_288 ();
 DECAPx2_ASAP7_75t_R FILLER_244_292 ();
 FILLER_ASAP7_75t_R FILLER_244_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_300 ();
 DECAPx1_ASAP7_75t_R FILLER_244_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_348 ();
 DECAPx6_ASAP7_75t_R FILLER_244_355 ();
 DECAPx2_ASAP7_75t_R FILLER_244_369 ();
 DECAPx2_ASAP7_75t_R FILLER_244_399 ();
 FILLER_ASAP7_75t_R FILLER_244_405 ();
 DECAPx6_ASAP7_75t_R FILLER_244_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_427 ();
 DECAPx2_ASAP7_75t_R FILLER_244_454 ();
 FILLER_ASAP7_75t_R FILLER_244_460 ();
 FILLER_ASAP7_75t_R FILLER_244_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_466 ();
 FILLER_ASAP7_75t_R FILLER_244_470 ();
 DECAPx4_ASAP7_75t_R FILLER_244_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_498 ();
 DECAPx1_ASAP7_75t_R FILLER_244_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_538 ();
 FILLER_ASAP7_75t_R FILLER_244_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_559 ();
 DECAPx10_ASAP7_75t_R FILLER_244_599 ();
 DECAPx10_ASAP7_75t_R FILLER_244_621 ();
 DECAPx10_ASAP7_75t_R FILLER_244_643 ();
 DECAPx10_ASAP7_75t_R FILLER_244_665 ();
 DECAPx10_ASAP7_75t_R FILLER_244_687 ();
 DECAPx10_ASAP7_75t_R FILLER_244_709 ();
 DECAPx10_ASAP7_75t_R FILLER_244_731 ();
 DECAPx10_ASAP7_75t_R FILLER_244_753 ();
 DECAPx2_ASAP7_75t_R FILLER_244_775 ();
 FILLER_ASAP7_75t_R FILLER_244_781 ();
 DECAPx2_ASAP7_75t_R FILLER_244_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_815 ();
 DECAPx6_ASAP7_75t_R FILLER_244_822 ();
 FILLER_ASAP7_75t_R FILLER_244_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_864 ();
 DECAPx10_ASAP7_75t_R FILLER_244_890 ();
 FILLER_ASAP7_75t_R FILLER_244_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_914 ();
 DECAPx4_ASAP7_75t_R FILLER_244_926 ();
 FILLER_ASAP7_75t_R FILLER_244_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_938 ();
 DECAPx4_ASAP7_75t_R FILLER_244_947 ();
 FILLER_ASAP7_75t_R FILLER_244_957 ();
 DECAPx4_ASAP7_75t_R FILLER_244_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1025 ();
 DECAPx4_ASAP7_75t_R FILLER_244_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1047 ();
 FILLER_ASAP7_75t_R FILLER_244_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_244_1075 ();
 FILLER_ASAP7_75t_R FILLER_244_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1091 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_244_1120 ();
 FILLER_ASAP7_75t_R FILLER_244_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1128 ();
 DECAPx4_ASAP7_75t_R FILLER_244_1135 ();
 FILLER_ASAP7_75t_R FILLER_244_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1147 ();
 DECAPx4_ASAP7_75t_R FILLER_244_1151 ();
 FILLER_ASAP7_75t_R FILLER_244_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_244_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_245_2 ();
 DECAPx10_ASAP7_75t_R FILLER_245_24 ();
 DECAPx10_ASAP7_75t_R FILLER_245_46 ();
 DECAPx10_ASAP7_75t_R FILLER_245_68 ();
 DECAPx10_ASAP7_75t_R FILLER_245_90 ();
 DECAPx10_ASAP7_75t_R FILLER_245_112 ();
 DECAPx6_ASAP7_75t_R FILLER_245_134 ();
 FILLER_ASAP7_75t_R FILLER_245_148 ();
 DECAPx2_ASAP7_75t_R FILLER_245_161 ();
 FILLER_ASAP7_75t_R FILLER_245_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_169 ();
 FILLER_ASAP7_75t_R FILLER_245_174 ();
 FILLER_ASAP7_75t_R FILLER_245_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_211 ();
 FILLER_ASAP7_75t_R FILLER_245_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_221 ();
 FILLER_ASAP7_75t_R FILLER_245_225 ();
 DECAPx6_ASAP7_75t_R FILLER_245_233 ();
 DECAPx4_ASAP7_75t_R FILLER_245_260 ();
 FILLER_ASAP7_75t_R FILLER_245_270 ();
 DECAPx6_ASAP7_75t_R FILLER_245_275 ();
 DECAPx2_ASAP7_75t_R FILLER_245_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_295 ();
 DECAPx1_ASAP7_75t_R FILLER_245_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_326 ();
 DECAPx2_ASAP7_75t_R FILLER_245_330 ();
 DECAPx6_ASAP7_75t_R FILLER_245_362 ();
 DECAPx1_ASAP7_75t_R FILLER_245_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_380 ();
 FILLER_ASAP7_75t_R FILLER_245_413 ();
 DECAPx2_ASAP7_75t_R FILLER_245_418 ();
 FILLER_ASAP7_75t_R FILLER_245_424 ();
 FILLER_ASAP7_75t_R FILLER_245_432 ();
 DECAPx6_ASAP7_75t_R FILLER_245_446 ();
 FILLER_ASAP7_75t_R FILLER_245_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_462 ();
 DECAPx4_ASAP7_75t_R FILLER_245_469 ();
 DECAPx6_ASAP7_75t_R FILLER_245_489 ();
 DECAPx2_ASAP7_75t_R FILLER_245_506 ();
 FILLER_ASAP7_75t_R FILLER_245_512 ();
 DECAPx10_ASAP7_75t_R FILLER_245_517 ();
 DECAPx4_ASAP7_75t_R FILLER_245_539 ();
 DECAPx10_ASAP7_75t_R FILLER_245_555 ();
 DECAPx4_ASAP7_75t_R FILLER_245_577 ();
 FILLER_ASAP7_75t_R FILLER_245_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_589 ();
 DECAPx6_ASAP7_75t_R FILLER_245_600 ();
 DECAPx1_ASAP7_75t_R FILLER_245_614 ();
 DECAPx10_ASAP7_75t_R FILLER_245_628 ();
 DECAPx10_ASAP7_75t_R FILLER_245_650 ();
 DECAPx10_ASAP7_75t_R FILLER_245_672 ();
 DECAPx10_ASAP7_75t_R FILLER_245_694 ();
 DECAPx10_ASAP7_75t_R FILLER_245_716 ();
 DECAPx10_ASAP7_75t_R FILLER_245_738 ();
 DECAPx10_ASAP7_75t_R FILLER_245_760 ();
 DECAPx10_ASAP7_75t_R FILLER_245_782 ();
 DECAPx2_ASAP7_75t_R FILLER_245_804 ();
 FILLER_ASAP7_75t_R FILLER_245_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_812 ();
 DECAPx2_ASAP7_75t_R FILLER_245_819 ();
 FILLER_ASAP7_75t_R FILLER_245_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_827 ();
 DECAPx6_ASAP7_75t_R FILLER_245_841 ();
 DECAPx1_ASAP7_75t_R FILLER_245_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_870 ();
 DECAPx10_ASAP7_75t_R FILLER_245_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_901 ();
 FILLER_ASAP7_75t_R FILLER_245_919 ();
 FILLER_ASAP7_75t_R FILLER_245_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_928 ();
 DECAPx2_ASAP7_75t_R FILLER_245_947 ();
 DECAPx2_ASAP7_75t_R FILLER_245_956 ();
 FILLER_ASAP7_75t_R FILLER_245_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_964 ();
 DECAPx4_ASAP7_75t_R FILLER_245_975 ();
 FILLER_ASAP7_75t_R FILLER_245_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_987 ();
 DECAPx1_ASAP7_75t_R FILLER_245_998 ();
 DECAPx1_ASAP7_75t_R FILLER_245_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_245_1031 ();
 FILLER_ASAP7_75t_R FILLER_245_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1039 ();
 DECAPx6_ASAP7_75t_R FILLER_245_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1068 ();
 DECAPx4_ASAP7_75t_R FILLER_245_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_245_1097 ();
 FILLER_ASAP7_75t_R FILLER_245_1124 ();
 DECAPx6_ASAP7_75t_R FILLER_245_1148 ();
 FILLER_ASAP7_75t_R FILLER_245_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1346 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1368 ();
 FILLER_ASAP7_75t_R FILLER_245_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_246_2 ();
 DECAPx10_ASAP7_75t_R FILLER_246_24 ();
 DECAPx10_ASAP7_75t_R FILLER_246_46 ();
 DECAPx10_ASAP7_75t_R FILLER_246_68 ();
 DECAPx10_ASAP7_75t_R FILLER_246_90 ();
 DECAPx10_ASAP7_75t_R FILLER_246_112 ();
 DECAPx2_ASAP7_75t_R FILLER_246_134 ();
 FILLER_ASAP7_75t_R FILLER_246_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_142 ();
 DECAPx6_ASAP7_75t_R FILLER_246_169 ();
 FILLER_ASAP7_75t_R FILLER_246_183 ();
 DECAPx1_ASAP7_75t_R FILLER_246_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_195 ();
 DECAPx2_ASAP7_75t_R FILLER_246_199 ();
 FILLER_ASAP7_75t_R FILLER_246_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_239 ();
 DECAPx1_ASAP7_75t_R FILLER_246_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_283 ();
 DECAPx6_ASAP7_75t_R FILLER_246_297 ();
 DECAPx10_ASAP7_75t_R FILLER_246_314 ();
 DECAPx2_ASAP7_75t_R FILLER_246_336 ();
 FILLER_ASAP7_75t_R FILLER_246_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_350 ();
 FILLER_ASAP7_75t_R FILLER_246_354 ();
 DECAPx1_ASAP7_75t_R FILLER_246_368 ();
 DECAPx2_ASAP7_75t_R FILLER_246_378 ();
 FILLER_ASAP7_75t_R FILLER_246_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_386 ();
 FILLER_ASAP7_75t_R FILLER_246_393 ();
 FILLER_ASAP7_75t_R FILLER_246_398 ();
 DECAPx1_ASAP7_75t_R FILLER_246_432 ();
 DECAPx1_ASAP7_75t_R FILLER_246_470 ();
 DECAPx6_ASAP7_75t_R FILLER_246_506 ();
 FILLER_ASAP7_75t_R FILLER_246_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_522 ();
 DECAPx4_ASAP7_75t_R FILLER_246_529 ();
 DECAPx6_ASAP7_75t_R FILLER_246_545 ();
 FILLER_ASAP7_75t_R FILLER_246_559 ();
 DECAPx4_ASAP7_75t_R FILLER_246_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_577 ();
 FILLER_ASAP7_75t_R FILLER_246_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_584 ();
 DECAPx10_ASAP7_75t_R FILLER_246_595 ();
 DECAPx10_ASAP7_75t_R FILLER_246_617 ();
 DECAPx10_ASAP7_75t_R FILLER_246_639 ();
 DECAPx10_ASAP7_75t_R FILLER_246_661 ();
 DECAPx10_ASAP7_75t_R FILLER_246_683 ();
 DECAPx10_ASAP7_75t_R FILLER_246_705 ();
 DECAPx10_ASAP7_75t_R FILLER_246_727 ();
 DECAPx10_ASAP7_75t_R FILLER_246_749 ();
 DECAPx6_ASAP7_75t_R FILLER_246_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_812 ();
 DECAPx6_ASAP7_75t_R FILLER_246_843 ();
 FILLER_ASAP7_75t_R FILLER_246_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_859 ();
 DECAPx6_ASAP7_75t_R FILLER_246_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_891 ();
 DECAPx4_ASAP7_75t_R FILLER_246_964 ();
 DECAPx2_ASAP7_75t_R FILLER_246_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_998 ();
 DECAPx2_ASAP7_75t_R FILLER_246_1013 ();
 FILLER_ASAP7_75t_R FILLER_246_1019 ();
 DECAPx4_ASAP7_75t_R FILLER_246_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1040 ();
 FILLER_ASAP7_75t_R FILLER_246_1047 ();
 FILLER_ASAP7_75t_R FILLER_246_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_246_1078 ();
 FILLER_ASAP7_75t_R FILLER_246_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_246_1097 ();
 FILLER_ASAP7_75t_R FILLER_246_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1117 ();
 FILLER_ASAP7_75t_R FILLER_246_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1252 ();
 DECAPx2_ASAP7_75t_R FILLER_246_1274 ();
 FILLER_ASAP7_75t_R FILLER_246_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1354 ();
 DECAPx4_ASAP7_75t_R FILLER_246_1376 ();
 DECAPx1_ASAP7_75t_R FILLER_246_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_247_2 ();
 DECAPx10_ASAP7_75t_R FILLER_247_24 ();
 DECAPx10_ASAP7_75t_R FILLER_247_46 ();
 DECAPx10_ASAP7_75t_R FILLER_247_68 ();
 DECAPx10_ASAP7_75t_R FILLER_247_90 ();
 DECAPx10_ASAP7_75t_R FILLER_247_112 ();
 DECAPx6_ASAP7_75t_R FILLER_247_134 ();
 DECAPx1_ASAP7_75t_R FILLER_247_148 ();
 DECAPx10_ASAP7_75t_R FILLER_247_158 ();
 FILLER_ASAP7_75t_R FILLER_247_180 ();
 DECAPx6_ASAP7_75t_R FILLER_247_196 ();
 DECAPx2_ASAP7_75t_R FILLER_247_210 ();
 DECAPx4_ASAP7_75t_R FILLER_247_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_252 ();
 FILLER_ASAP7_75t_R FILLER_247_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_310 ();
 DECAPx4_ASAP7_75t_R FILLER_247_321 ();
 FILLER_ASAP7_75t_R FILLER_247_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_333 ();
 DECAPx2_ASAP7_75t_R FILLER_247_343 ();
 FILLER_ASAP7_75t_R FILLER_247_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_351 ();
 DECAPx6_ASAP7_75t_R FILLER_247_384 ();
 DECAPx2_ASAP7_75t_R FILLER_247_398 ();
 DECAPx1_ASAP7_75t_R FILLER_247_410 ();
 FILLER_ASAP7_75t_R FILLER_247_417 ();
 FILLER_ASAP7_75t_R FILLER_247_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_451 ();
 FILLER_ASAP7_75t_R FILLER_247_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_490 ();
 FILLER_ASAP7_75t_R FILLER_247_553 ();
 DECAPx10_ASAP7_75t_R FILLER_247_585 ();
 DECAPx10_ASAP7_75t_R FILLER_247_607 ();
 DECAPx10_ASAP7_75t_R FILLER_247_629 ();
 DECAPx10_ASAP7_75t_R FILLER_247_651 ();
 DECAPx10_ASAP7_75t_R FILLER_247_673 ();
 DECAPx10_ASAP7_75t_R FILLER_247_695 ();
 DECAPx10_ASAP7_75t_R FILLER_247_717 ();
 DECAPx10_ASAP7_75t_R FILLER_247_739 ();
 DECAPx10_ASAP7_75t_R FILLER_247_761 ();
 DECAPx6_ASAP7_75t_R FILLER_247_783 ();
 FILLER_ASAP7_75t_R FILLER_247_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_799 ();
 FILLER_ASAP7_75t_R FILLER_247_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_805 ();
 FILLER_ASAP7_75t_R FILLER_247_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_834 ();
 FILLER_ASAP7_75t_R FILLER_247_847 ();
 FILLER_ASAP7_75t_R FILLER_247_853 ();
 DECAPx4_ASAP7_75t_R FILLER_247_873 ();
 DECAPx1_ASAP7_75t_R FILLER_247_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_897 ();
 FILLER_ASAP7_75t_R FILLER_247_904 ();
 FILLER_ASAP7_75t_R FILLER_247_909 ();
 DECAPx2_ASAP7_75t_R FILLER_247_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_923 ();
 FILLER_ASAP7_75t_R FILLER_247_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_928 ();
 DECAPx6_ASAP7_75t_R FILLER_247_943 ();
 FILLER_ASAP7_75t_R FILLER_247_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_959 ();
 DECAPx1_ASAP7_75t_R FILLER_247_970 ();
 DECAPx4_ASAP7_75t_R FILLER_247_984 ();
 FILLER_ASAP7_75t_R FILLER_247_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_247_1013 ();
 FILLER_ASAP7_75t_R FILLER_247_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_247_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1105 ();
 DECAPx6_ASAP7_75t_R FILLER_247_1112 ();
 FILLER_ASAP7_75t_R FILLER_247_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1128 ();
 DECAPx4_ASAP7_75t_R FILLER_247_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1354 ();
 DECAPx6_ASAP7_75t_R FILLER_247_1376 ();
 FILLER_ASAP7_75t_R FILLER_247_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_248_2 ();
 DECAPx10_ASAP7_75t_R FILLER_248_24 ();
 DECAPx10_ASAP7_75t_R FILLER_248_46 ();
 DECAPx10_ASAP7_75t_R FILLER_248_68 ();
 DECAPx10_ASAP7_75t_R FILLER_248_90 ();
 DECAPx10_ASAP7_75t_R FILLER_248_112 ();
 DECAPx10_ASAP7_75t_R FILLER_248_134 ();
 DECAPx1_ASAP7_75t_R FILLER_248_156 ();
 FILLER_ASAP7_75t_R FILLER_248_172 ();
 DECAPx4_ASAP7_75t_R FILLER_248_214 ();
 DECAPx10_ASAP7_75t_R FILLER_248_234 ();
 DECAPx4_ASAP7_75t_R FILLER_248_256 ();
 FILLER_ASAP7_75t_R FILLER_248_279 ();
 DECAPx4_ASAP7_75t_R FILLER_248_284 ();
 FILLER_ASAP7_75t_R FILLER_248_294 ();
 FILLER_ASAP7_75t_R FILLER_248_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_339 ();
 FILLER_ASAP7_75t_R FILLER_248_346 ();
 DECAPx4_ASAP7_75t_R FILLER_248_374 ();
 FILLER_ASAP7_75t_R FILLER_248_399 ();
 DECAPx6_ASAP7_75t_R FILLER_248_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_418 ();
 DECAPx6_ASAP7_75t_R FILLER_248_445 ();
 FILLER_ASAP7_75t_R FILLER_248_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_461 ();
 DECAPx1_ASAP7_75t_R FILLER_248_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_468 ();
 DECAPx6_ASAP7_75t_R FILLER_248_475 ();
 DECAPx2_ASAP7_75t_R FILLER_248_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_498 ();
 DECAPx4_ASAP7_75t_R FILLER_248_505 ();
 FILLER_ASAP7_75t_R FILLER_248_518 ();
 DECAPx1_ASAP7_75t_R FILLER_248_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_534 ();
 FILLER_ASAP7_75t_R FILLER_248_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_572 ();
 DECAPx10_ASAP7_75t_R FILLER_248_576 ();
 DECAPx10_ASAP7_75t_R FILLER_248_598 ();
 DECAPx10_ASAP7_75t_R FILLER_248_620 ();
 DECAPx10_ASAP7_75t_R FILLER_248_642 ();
 DECAPx10_ASAP7_75t_R FILLER_248_664 ();
 DECAPx10_ASAP7_75t_R FILLER_248_686 ();
 DECAPx10_ASAP7_75t_R FILLER_248_708 ();
 DECAPx10_ASAP7_75t_R FILLER_248_730 ();
 DECAPx10_ASAP7_75t_R FILLER_248_752 ();
 DECAPx4_ASAP7_75t_R FILLER_248_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_868 ();
 FILLER_ASAP7_75t_R FILLER_248_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_879 ();
 DECAPx2_ASAP7_75t_R FILLER_248_901 ();
 FILLER_ASAP7_75t_R FILLER_248_917 ();
 DECAPx2_ASAP7_75t_R FILLER_248_926 ();
 FILLER_ASAP7_75t_R FILLER_248_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_934 ();
 DECAPx6_ASAP7_75t_R FILLER_248_946 ();
 FILLER_ASAP7_75t_R FILLER_248_960 ();
 DECAPx2_ASAP7_75t_R FILLER_248_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_986 ();
 DECAPx2_ASAP7_75t_R FILLER_248_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_248_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_248_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_248_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_248_1116 ();
 DECAPx2_ASAP7_75t_R FILLER_248_1123 ();
 FILLER_ASAP7_75t_R FILLER_248_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_248_1377 ();
 FILLER_ASAP7_75t_R FILLER_248_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_248_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_249_2 ();
 DECAPx10_ASAP7_75t_R FILLER_249_24 ();
 DECAPx10_ASAP7_75t_R FILLER_249_46 ();
 DECAPx10_ASAP7_75t_R FILLER_249_68 ();
 DECAPx10_ASAP7_75t_R FILLER_249_90 ();
 DECAPx10_ASAP7_75t_R FILLER_249_112 ();
 DECAPx10_ASAP7_75t_R FILLER_249_134 ();
 FILLER_ASAP7_75t_R FILLER_249_156 ();
 DECAPx1_ASAP7_75t_R FILLER_249_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_215 ();
 DECAPx6_ASAP7_75t_R FILLER_249_223 ();
 FILLER_ASAP7_75t_R FILLER_249_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_249 ();
 DECAPx2_ASAP7_75t_R FILLER_249_260 ();
 DECAPx1_ASAP7_75t_R FILLER_249_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_322 ();
 DECAPx2_ASAP7_75t_R FILLER_249_349 ();
 FILLER_ASAP7_75t_R FILLER_249_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_357 ();
 DECAPx6_ASAP7_75t_R FILLER_249_367 ();
 DECAPx6_ASAP7_75t_R FILLER_249_407 ();
 DECAPx1_ASAP7_75t_R FILLER_249_421 ();
 DECAPx1_ASAP7_75t_R FILLER_249_477 ();
 FILLER_ASAP7_75t_R FILLER_249_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_487 ();
 DECAPx10_ASAP7_75t_R FILLER_249_494 ();
 DECAPx6_ASAP7_75t_R FILLER_249_520 ();
 DECAPx1_ASAP7_75t_R FILLER_249_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_538 ();
 DECAPx2_ASAP7_75t_R FILLER_249_545 ();
 FILLER_ASAP7_75t_R FILLER_249_551 ();
 DECAPx10_ASAP7_75t_R FILLER_249_556 ();
 DECAPx10_ASAP7_75t_R FILLER_249_578 ();
 DECAPx10_ASAP7_75t_R FILLER_249_600 ();
 DECAPx10_ASAP7_75t_R FILLER_249_622 ();
 DECAPx10_ASAP7_75t_R FILLER_249_644 ();
 DECAPx10_ASAP7_75t_R FILLER_249_666 ();
 DECAPx10_ASAP7_75t_R FILLER_249_688 ();
 DECAPx10_ASAP7_75t_R FILLER_249_710 ();
 DECAPx10_ASAP7_75t_R FILLER_249_732 ();
 DECAPx10_ASAP7_75t_R FILLER_249_754 ();
 DECAPx10_ASAP7_75t_R FILLER_249_776 ();
 FILLER_ASAP7_75t_R FILLER_249_798 ();
 FILLER_ASAP7_75t_R FILLER_249_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_836 ();
 FILLER_ASAP7_75t_R FILLER_249_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_854 ();
 DECAPx1_ASAP7_75t_R FILLER_249_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_936 ();
 DECAPx4_ASAP7_75t_R FILLER_249_953 ();
 DECAPx2_ASAP7_75t_R FILLER_249_973 ();
 FILLER_ASAP7_75t_R FILLER_249_979 ();
 DECAPx10_ASAP7_75t_R FILLER_249_989 ();
 DECAPx2_ASAP7_75t_R FILLER_249_1011 ();
 FILLER_ASAP7_75t_R FILLER_249_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1019 ();
 DECAPx6_ASAP7_75t_R FILLER_249_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1058 ();
 FILLER_ASAP7_75t_R FILLER_249_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1071 ();
 FILLER_ASAP7_75t_R FILLER_249_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_249_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1346 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1368 ();
 FILLER_ASAP7_75t_R FILLER_249_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_250_2 ();
 DECAPx10_ASAP7_75t_R FILLER_250_24 ();
 DECAPx10_ASAP7_75t_R FILLER_250_46 ();
 DECAPx10_ASAP7_75t_R FILLER_250_68 ();
 DECAPx10_ASAP7_75t_R FILLER_250_90 ();
 DECAPx10_ASAP7_75t_R FILLER_250_112 ();
 DECAPx10_ASAP7_75t_R FILLER_250_134 ();
 DECAPx6_ASAP7_75t_R FILLER_250_156 ();
 FILLER_ASAP7_75t_R FILLER_250_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_172 ();
 DECAPx6_ASAP7_75t_R FILLER_250_176 ();
 FILLER_ASAP7_75t_R FILLER_250_196 ();
 FILLER_ASAP7_75t_R FILLER_250_201 ();
 DECAPx4_ASAP7_75t_R FILLER_250_258 ();
 DECAPx6_ASAP7_75t_R FILLER_250_281 ();
 DECAPx2_ASAP7_75t_R FILLER_250_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_301 ();
 FILLER_ASAP7_75t_R FILLER_250_308 ();
 DECAPx2_ASAP7_75t_R FILLER_250_313 ();
 DECAPx1_ASAP7_75t_R FILLER_250_323 ();
 DECAPx2_ASAP7_75t_R FILLER_250_330 ();
 FILLER_ASAP7_75t_R FILLER_250_336 ();
 DECAPx2_ASAP7_75t_R FILLER_250_341 ();
 DECAPx6_ASAP7_75t_R FILLER_250_353 ();
 DECAPx2_ASAP7_75t_R FILLER_250_367 ();
 DECAPx2_ASAP7_75t_R FILLER_250_385 ();
 FILLER_ASAP7_75t_R FILLER_250_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_393 ();
 DECAPx2_ASAP7_75t_R FILLER_250_398 ();
 DECAPx1_ASAP7_75t_R FILLER_250_437 ();
 DECAPx4_ASAP7_75t_R FILLER_250_444 ();
 FILLER_ASAP7_75t_R FILLER_250_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_464 ();
 DECAPx2_ASAP7_75t_R FILLER_250_468 ();
 FILLER_ASAP7_75t_R FILLER_250_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_484 ();
 DECAPx10_ASAP7_75t_R FILLER_250_520 ();
 DECAPx10_ASAP7_75t_R FILLER_250_542 ();
 DECAPx10_ASAP7_75t_R FILLER_250_564 ();
 DECAPx10_ASAP7_75t_R FILLER_250_586 ();
 DECAPx10_ASAP7_75t_R FILLER_250_608 ();
 DECAPx10_ASAP7_75t_R FILLER_250_630 ();
 DECAPx10_ASAP7_75t_R FILLER_250_652 ();
 DECAPx10_ASAP7_75t_R FILLER_250_674 ();
 DECAPx10_ASAP7_75t_R FILLER_250_696 ();
 DECAPx10_ASAP7_75t_R FILLER_250_718 ();
 DECAPx10_ASAP7_75t_R FILLER_250_740 ();
 DECAPx10_ASAP7_75t_R FILLER_250_762 ();
 DECAPx10_ASAP7_75t_R FILLER_250_784 ();
 DECAPx2_ASAP7_75t_R FILLER_250_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_868 ();
 DECAPx6_ASAP7_75t_R FILLER_250_872 ();
 DECAPx2_ASAP7_75t_R FILLER_250_886 ();
 DECAPx10_ASAP7_75t_R FILLER_250_954 ();
 DECAPx2_ASAP7_75t_R FILLER_250_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_982 ();
 DECAPx4_ASAP7_75t_R FILLER_250_991 ();
 FILLER_ASAP7_75t_R FILLER_250_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_250_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_250_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_250_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1083 ();
 DECAPx6_ASAP7_75t_R FILLER_250_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1347 ();
 DECAPx6_ASAP7_75t_R FILLER_250_1369 ();
 FILLER_ASAP7_75t_R FILLER_250_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_250_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_251_2 ();
 DECAPx10_ASAP7_75t_R FILLER_251_24 ();
 DECAPx10_ASAP7_75t_R FILLER_251_46 ();
 DECAPx10_ASAP7_75t_R FILLER_251_68 ();
 DECAPx10_ASAP7_75t_R FILLER_251_90 ();
 DECAPx10_ASAP7_75t_R FILLER_251_112 ();
 DECAPx10_ASAP7_75t_R FILLER_251_134 ();
 DECAPx10_ASAP7_75t_R FILLER_251_156 ();
 DECAPx10_ASAP7_75t_R FILLER_251_178 ();
 DECAPx10_ASAP7_75t_R FILLER_251_200 ();
 DECAPx2_ASAP7_75t_R FILLER_251_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_237 ();
 DECAPx2_ASAP7_75t_R FILLER_251_244 ();
 FILLER_ASAP7_75t_R FILLER_251_250 ();
 DECAPx2_ASAP7_75t_R FILLER_251_261 ();
 FILLER_ASAP7_75t_R FILLER_251_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_269 ();
 DECAPx6_ASAP7_75t_R FILLER_251_296 ();
 DECAPx10_ASAP7_75t_R FILLER_251_316 ();
 DECAPx2_ASAP7_75t_R FILLER_251_338 ();
 FILLER_ASAP7_75t_R FILLER_251_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_346 ();
 DECAPx2_ASAP7_75t_R FILLER_251_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_359 ();
 DECAPx1_ASAP7_75t_R FILLER_251_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_374 ();
 FILLER_ASAP7_75t_R FILLER_251_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_403 ();
 DECAPx1_ASAP7_75t_R FILLER_251_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_434 ();
 DECAPx6_ASAP7_75t_R FILLER_251_441 ();
 DECAPx4_ASAP7_75t_R FILLER_251_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_529 ();
 DECAPx10_ASAP7_75t_R FILLER_251_533 ();
 DECAPx10_ASAP7_75t_R FILLER_251_555 ();
 DECAPx10_ASAP7_75t_R FILLER_251_577 ();
 DECAPx10_ASAP7_75t_R FILLER_251_599 ();
 DECAPx10_ASAP7_75t_R FILLER_251_621 ();
 DECAPx10_ASAP7_75t_R FILLER_251_643 ();
 DECAPx10_ASAP7_75t_R FILLER_251_665 ();
 DECAPx10_ASAP7_75t_R FILLER_251_687 ();
 DECAPx10_ASAP7_75t_R FILLER_251_709 ();
 DECAPx10_ASAP7_75t_R FILLER_251_731 ();
 DECAPx10_ASAP7_75t_R FILLER_251_753 ();
 DECAPx10_ASAP7_75t_R FILLER_251_775 ();
 DECAPx6_ASAP7_75t_R FILLER_251_797 ();
 DECAPx6_ASAP7_75t_R FILLER_251_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_828 ();
 DECAPx6_ASAP7_75t_R FILLER_251_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_849 ();
 DECAPx10_ASAP7_75t_R FILLER_251_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_875 ();
 DECAPx2_ASAP7_75t_R FILLER_251_905 ();
 DECAPx2_ASAP7_75t_R FILLER_251_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_923 ();
 DECAPx2_ASAP7_75t_R FILLER_251_926 ();
 FILLER_ASAP7_75t_R FILLER_251_932 ();
 DECAPx1_ASAP7_75t_R FILLER_251_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_974 ();
 DECAPx2_ASAP7_75t_R FILLER_251_978 ();
 FILLER_ASAP7_75t_R FILLER_251_984 ();
 DECAPx2_ASAP7_75t_R FILLER_251_1051 ();
 FILLER_ASAP7_75t_R FILLER_251_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1085 ();
 FILLER_ASAP7_75t_R FILLER_251_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_251_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1289 ();
 DECAPx6_ASAP7_75t_R FILLER_251_1311 ();
 DECAPx1_ASAP7_75t_R FILLER_251_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1357 ();
 DECAPx4_ASAP7_75t_R FILLER_251_1379 ();
 FILLER_ASAP7_75t_R FILLER_251_1389 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_252_2 ();
 DECAPx10_ASAP7_75t_R FILLER_252_24 ();
 DECAPx10_ASAP7_75t_R FILLER_252_46 ();
 DECAPx10_ASAP7_75t_R FILLER_252_68 ();
 DECAPx10_ASAP7_75t_R FILLER_252_90 ();
 DECAPx10_ASAP7_75t_R FILLER_252_112 ();
 DECAPx10_ASAP7_75t_R FILLER_252_134 ();
 DECAPx10_ASAP7_75t_R FILLER_252_156 ();
 DECAPx10_ASAP7_75t_R FILLER_252_178 ();
 DECAPx10_ASAP7_75t_R FILLER_252_200 ();
 DECAPx4_ASAP7_75t_R FILLER_252_222 ();
 FILLER_ASAP7_75t_R FILLER_252_232 ();
 DECAPx10_ASAP7_75t_R FILLER_252_260 ();
 FILLER_ASAP7_75t_R FILLER_252_282 ();
 FILLER_ASAP7_75t_R FILLER_252_287 ();
 FILLER_ASAP7_75t_R FILLER_252_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_321 ();
 DECAPx2_ASAP7_75t_R FILLER_252_326 ();
 FILLER_ASAP7_75t_R FILLER_252_332 ();
 DECAPx6_ASAP7_75t_R FILLER_252_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_399 ();
 DECAPx6_ASAP7_75t_R FILLER_252_403 ();
 DECAPx1_ASAP7_75t_R FILLER_252_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_421 ();
 FILLER_ASAP7_75t_R FILLER_252_448 ();
 FILLER_ASAP7_75t_R FILLER_252_453 ();
 FILLER_ASAP7_75t_R FILLER_252_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_461 ();
 DECAPx1_ASAP7_75t_R FILLER_252_464 ();
 DECAPx1_ASAP7_75t_R FILLER_252_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_485 ();
 DECAPx4_ASAP7_75t_R FILLER_252_489 ();
 DECAPx10_ASAP7_75t_R FILLER_252_542 ();
 DECAPx10_ASAP7_75t_R FILLER_252_564 ();
 DECAPx10_ASAP7_75t_R FILLER_252_586 ();
 DECAPx10_ASAP7_75t_R FILLER_252_608 ();
 DECAPx10_ASAP7_75t_R FILLER_252_630 ();
 DECAPx10_ASAP7_75t_R FILLER_252_652 ();
 DECAPx10_ASAP7_75t_R FILLER_252_674 ();
 DECAPx10_ASAP7_75t_R FILLER_252_696 ();
 DECAPx10_ASAP7_75t_R FILLER_252_718 ();
 DECAPx10_ASAP7_75t_R FILLER_252_740 ();
 DECAPx10_ASAP7_75t_R FILLER_252_762 ();
 DECAPx4_ASAP7_75t_R FILLER_252_784 ();
 FILLER_ASAP7_75t_R FILLER_252_794 ();
 FILLER_ASAP7_75t_R FILLER_252_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_839 ();
 DECAPx4_ASAP7_75t_R FILLER_252_849 ();
 FILLER_ASAP7_75t_R FILLER_252_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_861 ();
 DECAPx6_ASAP7_75t_R FILLER_252_871 ();
 DECAPx1_ASAP7_75t_R FILLER_252_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_889 ();
 DECAPx10_ASAP7_75t_R FILLER_252_893 ();
 DECAPx2_ASAP7_75t_R FILLER_252_915 ();
 FILLER_ASAP7_75t_R FILLER_252_924 ();
 DECAPx1_ASAP7_75t_R FILLER_252_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_947 ();
 DECAPx6_ASAP7_75t_R FILLER_252_951 ();
 FILLER_ASAP7_75t_R FILLER_252_965 ();
 FILLER_ASAP7_75t_R FILLER_252_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_252_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_252_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1073 ();
 FILLER_ASAP7_75t_R FILLER_252_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_252_1097 ();
 FILLER_ASAP7_75t_R FILLER_252_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_252_1378 ();
 FILLER_ASAP7_75t_R FILLER_252_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_252_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_253_2 ();
 DECAPx10_ASAP7_75t_R FILLER_253_24 ();
 DECAPx10_ASAP7_75t_R FILLER_253_46 ();
 DECAPx10_ASAP7_75t_R FILLER_253_68 ();
 DECAPx10_ASAP7_75t_R FILLER_253_90 ();
 DECAPx10_ASAP7_75t_R FILLER_253_112 ();
 DECAPx10_ASAP7_75t_R FILLER_253_134 ();
 DECAPx10_ASAP7_75t_R FILLER_253_156 ();
 DECAPx10_ASAP7_75t_R FILLER_253_178 ();
 DECAPx10_ASAP7_75t_R FILLER_253_200 ();
 DECAPx10_ASAP7_75t_R FILLER_253_222 ();
 DECAPx1_ASAP7_75t_R FILLER_253_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_263 ();
 DECAPx1_ASAP7_75t_R FILLER_253_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_272 ();
 DECAPx1_ASAP7_75t_R FILLER_253_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_291 ();
 FILLER_ASAP7_75t_R FILLER_253_303 ();
 FILLER_ASAP7_75t_R FILLER_253_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_333 ();
 FILLER_ASAP7_75t_R FILLER_253_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_342 ();
 DECAPx4_ASAP7_75t_R FILLER_253_369 ();
 FILLER_ASAP7_75t_R FILLER_253_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_381 ();
 DECAPx6_ASAP7_75t_R FILLER_253_408 ();
 FILLER_ASAP7_75t_R FILLER_253_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_424 ();
 DECAPx1_ASAP7_75t_R FILLER_253_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_461 ();
 DECAPx10_ASAP7_75t_R FILLER_253_474 ();
 DECAPx6_ASAP7_75t_R FILLER_253_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_510 ();
 DECAPx1_ASAP7_75t_R FILLER_253_514 ();
 DECAPx10_ASAP7_75t_R FILLER_253_524 ();
 DECAPx10_ASAP7_75t_R FILLER_253_546 ();
 DECAPx10_ASAP7_75t_R FILLER_253_568 ();
 DECAPx10_ASAP7_75t_R FILLER_253_590 ();
 DECAPx10_ASAP7_75t_R FILLER_253_612 ();
 DECAPx10_ASAP7_75t_R FILLER_253_634 ();
 DECAPx10_ASAP7_75t_R FILLER_253_656 ();
 DECAPx10_ASAP7_75t_R FILLER_253_678 ();
 DECAPx10_ASAP7_75t_R FILLER_253_700 ();
 DECAPx10_ASAP7_75t_R FILLER_253_722 ();
 DECAPx10_ASAP7_75t_R FILLER_253_744 ();
 DECAPx10_ASAP7_75t_R FILLER_253_766 ();
 FILLER_ASAP7_75t_R FILLER_253_788 ();
 DECAPx4_ASAP7_75t_R FILLER_253_816 ();
 DECAPx1_ASAP7_75t_R FILLER_253_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_836 ();
 DECAPx2_ASAP7_75t_R FILLER_253_852 ();
 DECAPx10_ASAP7_75t_R FILLER_253_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_898 ();
 DECAPx4_ASAP7_75t_R FILLER_253_911 ();
 FILLER_ASAP7_75t_R FILLER_253_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_926 ();
 FILLER_ASAP7_75t_R FILLER_253_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_932 ();
 DECAPx4_ASAP7_75t_R FILLER_253_945 ();
 FILLER_ASAP7_75t_R FILLER_253_955 ();
 DECAPx4_ASAP7_75t_R FILLER_253_996 ();
 FILLER_ASAP7_75t_R FILLER_253_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_253_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_253_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1053 ();
 DECAPx4_ASAP7_75t_R FILLER_253_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1085 ();
 DECAPx1_ASAP7_75t_R FILLER_253_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1101 ();
 FILLER_ASAP7_75t_R FILLER_253_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1346 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1368 ();
 FILLER_ASAP7_75t_R FILLER_253_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_254_2 ();
 DECAPx10_ASAP7_75t_R FILLER_254_24 ();
 DECAPx10_ASAP7_75t_R FILLER_254_46 ();
 DECAPx10_ASAP7_75t_R FILLER_254_68 ();
 DECAPx10_ASAP7_75t_R FILLER_254_90 ();
 DECAPx10_ASAP7_75t_R FILLER_254_112 ();
 DECAPx10_ASAP7_75t_R FILLER_254_134 ();
 DECAPx10_ASAP7_75t_R FILLER_254_156 ();
 DECAPx10_ASAP7_75t_R FILLER_254_178 ();
 DECAPx10_ASAP7_75t_R FILLER_254_200 ();
 DECAPx6_ASAP7_75t_R FILLER_254_222 ();
 DECAPx2_ASAP7_75t_R FILLER_254_236 ();
 DECAPx2_ASAP7_75t_R FILLER_254_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_345 ();
 DECAPx2_ASAP7_75t_R FILLER_254_352 ();
 DECAPx10_ASAP7_75t_R FILLER_254_361 ();
 FILLER_ASAP7_75t_R FILLER_254_383 ();
 DECAPx6_ASAP7_75t_R FILLER_254_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_416 ();
 DECAPx2_ASAP7_75t_R FILLER_254_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_441 ();
 DECAPx6_ASAP7_75t_R FILLER_254_446 ();
 FILLER_ASAP7_75t_R FILLER_254_460 ();
 DECAPx10_ASAP7_75t_R FILLER_254_496 ();
 DECAPx10_ASAP7_75t_R FILLER_254_518 ();
 DECAPx10_ASAP7_75t_R FILLER_254_540 ();
 DECAPx10_ASAP7_75t_R FILLER_254_562 ();
 DECAPx10_ASAP7_75t_R FILLER_254_584 ();
 DECAPx10_ASAP7_75t_R FILLER_254_606 ();
 DECAPx10_ASAP7_75t_R FILLER_254_628 ();
 DECAPx10_ASAP7_75t_R FILLER_254_650 ();
 DECAPx10_ASAP7_75t_R FILLER_254_672 ();
 DECAPx10_ASAP7_75t_R FILLER_254_694 ();
 DECAPx10_ASAP7_75t_R FILLER_254_716 ();
 DECAPx10_ASAP7_75t_R FILLER_254_738 ();
 DECAPx10_ASAP7_75t_R FILLER_254_760 ();
 DECAPx4_ASAP7_75t_R FILLER_254_782 ();
 DECAPx2_ASAP7_75t_R FILLER_254_835 ();
 FILLER_ASAP7_75t_R FILLER_254_841 ();
 DECAPx2_ASAP7_75t_R FILLER_254_857 ();
 FILLER_ASAP7_75t_R FILLER_254_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_865 ();
 FILLER_ASAP7_75t_R FILLER_254_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_894 ();
 FILLER_ASAP7_75t_R FILLER_254_967 ();
 FILLER_ASAP7_75t_R FILLER_254_983 ();
 DECAPx2_ASAP7_75t_R FILLER_254_1001 ();
 FILLER_ASAP7_75t_R FILLER_254_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_254_1024 ();
 DECAPx6_ASAP7_75t_R FILLER_254_1044 ();
 FILLER_ASAP7_75t_R FILLER_254_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_254_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1094 ();
 FILLER_ASAP7_75t_R FILLER_254_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_254_1370 ();
 FILLER_ASAP7_75t_R FILLER_254_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_254_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_255_2 ();
 DECAPx10_ASAP7_75t_R FILLER_255_24 ();
 DECAPx10_ASAP7_75t_R FILLER_255_46 ();
 DECAPx10_ASAP7_75t_R FILLER_255_68 ();
 DECAPx10_ASAP7_75t_R FILLER_255_90 ();
 DECAPx10_ASAP7_75t_R FILLER_255_112 ();
 DECAPx10_ASAP7_75t_R FILLER_255_134 ();
 DECAPx10_ASAP7_75t_R FILLER_255_156 ();
 DECAPx10_ASAP7_75t_R FILLER_255_178 ();
 DECAPx10_ASAP7_75t_R FILLER_255_200 ();
 DECAPx10_ASAP7_75t_R FILLER_255_222 ();
 DECAPx4_ASAP7_75t_R FILLER_255_244 ();
 FILLER_ASAP7_75t_R FILLER_255_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_256 ();
 DECAPx10_ASAP7_75t_R FILLER_255_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_282 ();
 DECAPx10_ASAP7_75t_R FILLER_255_286 ();
 DECAPx4_ASAP7_75t_R FILLER_255_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_318 ();
 DECAPx2_ASAP7_75t_R FILLER_255_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_328 ();
 DECAPx4_ASAP7_75t_R FILLER_255_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_342 ();
 DECAPx2_ASAP7_75t_R FILLER_255_359 ();
 FILLER_ASAP7_75t_R FILLER_255_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_385 ();
 DECAPx4_ASAP7_75t_R FILLER_255_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_433 ();
 DECAPx2_ASAP7_75t_R FILLER_255_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_446 ();
 DECAPx4_ASAP7_75t_R FILLER_255_451 ();
 FILLER_ASAP7_75t_R FILLER_255_461 ();
 DECAPx10_ASAP7_75t_R FILLER_255_489 ();
 DECAPx10_ASAP7_75t_R FILLER_255_511 ();
 DECAPx10_ASAP7_75t_R FILLER_255_533 ();
 DECAPx10_ASAP7_75t_R FILLER_255_555 ();
 DECAPx10_ASAP7_75t_R FILLER_255_577 ();
 DECAPx10_ASAP7_75t_R FILLER_255_599 ();
 DECAPx10_ASAP7_75t_R FILLER_255_621 ();
 DECAPx10_ASAP7_75t_R FILLER_255_643 ();
 DECAPx10_ASAP7_75t_R FILLER_255_665 ();
 DECAPx10_ASAP7_75t_R FILLER_255_687 ();
 DECAPx10_ASAP7_75t_R FILLER_255_709 ();
 DECAPx10_ASAP7_75t_R FILLER_255_731 ();
 DECAPx10_ASAP7_75t_R FILLER_255_753 ();
 DECAPx10_ASAP7_75t_R FILLER_255_775 ();
 DECAPx2_ASAP7_75t_R FILLER_255_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_803 ();
 DECAPx1_ASAP7_75t_R FILLER_255_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_814 ();
 DECAPx1_ASAP7_75t_R FILLER_255_840 ();
 DECAPx2_ASAP7_75t_R FILLER_255_850 ();
 FILLER_ASAP7_75t_R FILLER_255_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_858 ();
 FILLER_ASAP7_75t_R FILLER_255_875 ();
 DECAPx2_ASAP7_75t_R FILLER_255_911 ();
 DECAPx1_ASAP7_75t_R FILLER_255_920 ();
 DECAPx4_ASAP7_75t_R FILLER_255_926 ();
 DECAPx6_ASAP7_75t_R FILLER_255_946 ();
 DECAPx1_ASAP7_75t_R FILLER_255_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_964 ();
 DECAPx6_ASAP7_75t_R FILLER_255_972 ();
 DECAPx2_ASAP7_75t_R FILLER_255_986 ();
 DECAPx4_ASAP7_75t_R FILLER_255_1018 ();
 DECAPx1_ASAP7_75t_R FILLER_255_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1046 ();
 DECAPx6_ASAP7_75t_R FILLER_255_1056 ();
 FILLER_ASAP7_75t_R FILLER_255_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_255_1077 ();
 FILLER_ASAP7_75t_R FILLER_255_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1085 ();
 FILLER_ASAP7_75t_R FILLER_255_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_255_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1111 ();
 FILLER_ASAP7_75t_R FILLER_255_1118 ();
 DECAPx4_ASAP7_75t_R FILLER_255_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_255_1383 ();
 FILLER_ASAP7_75t_R FILLER_255_1389 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_256_2 ();
 DECAPx10_ASAP7_75t_R FILLER_256_24 ();
 DECAPx10_ASAP7_75t_R FILLER_256_46 ();
 DECAPx10_ASAP7_75t_R FILLER_256_68 ();
 DECAPx10_ASAP7_75t_R FILLER_256_90 ();
 DECAPx10_ASAP7_75t_R FILLER_256_112 ();
 DECAPx10_ASAP7_75t_R FILLER_256_134 ();
 DECAPx10_ASAP7_75t_R FILLER_256_156 ();
 DECAPx10_ASAP7_75t_R FILLER_256_178 ();
 DECAPx10_ASAP7_75t_R FILLER_256_200 ();
 DECAPx10_ASAP7_75t_R FILLER_256_222 ();
 DECAPx10_ASAP7_75t_R FILLER_256_244 ();
 DECAPx10_ASAP7_75t_R FILLER_256_266 ();
 DECAPx10_ASAP7_75t_R FILLER_256_288 ();
 DECAPx6_ASAP7_75t_R FILLER_256_310 ();
 FILLER_ASAP7_75t_R FILLER_256_350 ();
 FILLER_ASAP7_75t_R FILLER_256_358 ();
 FILLER_ASAP7_75t_R FILLER_256_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_396 ();
 FILLER_ASAP7_75t_R FILLER_256_411 ();
 FILLER_ASAP7_75t_R FILLER_256_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_453 ();
 DECAPx1_ASAP7_75t_R FILLER_256_458 ();
 DECAPx4_ASAP7_75t_R FILLER_256_464 ();
 FILLER_ASAP7_75t_R FILLER_256_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_476 ();
 DECAPx1_ASAP7_75t_R FILLER_256_480 ();
 DECAPx10_ASAP7_75t_R FILLER_256_487 ();
 DECAPx10_ASAP7_75t_R FILLER_256_509 ();
 DECAPx10_ASAP7_75t_R FILLER_256_531 ();
 DECAPx10_ASAP7_75t_R FILLER_256_553 ();
 DECAPx10_ASAP7_75t_R FILLER_256_575 ();
 DECAPx10_ASAP7_75t_R FILLER_256_597 ();
 DECAPx10_ASAP7_75t_R FILLER_256_619 ();
 DECAPx10_ASAP7_75t_R FILLER_256_641 ();
 DECAPx10_ASAP7_75t_R FILLER_256_663 ();
 DECAPx10_ASAP7_75t_R FILLER_256_685 ();
 DECAPx10_ASAP7_75t_R FILLER_256_707 ();
 DECAPx10_ASAP7_75t_R FILLER_256_729 ();
 DECAPx10_ASAP7_75t_R FILLER_256_751 ();
 FILLER_ASAP7_75t_R FILLER_256_773 ();
 FILLER_ASAP7_75t_R FILLER_256_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_821 ();
 DECAPx6_ASAP7_75t_R FILLER_256_840 ();
 DECAPx1_ASAP7_75t_R FILLER_256_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_882 ();
 FILLER_ASAP7_75t_R FILLER_256_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_891 ();
 DECAPx1_ASAP7_75t_R FILLER_256_895 ();
 DECAPx10_ASAP7_75t_R FILLER_256_906 ();
 DECAPx2_ASAP7_75t_R FILLER_256_928 ();
 DECAPx2_ASAP7_75t_R FILLER_256_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_947 ();
 DECAPx2_ASAP7_75t_R FILLER_256_961 ();
 DECAPx2_ASAP7_75t_R FILLER_256_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_983 ();
 DECAPx1_ASAP7_75t_R FILLER_256_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_992 ();
 DECAPx4_ASAP7_75t_R FILLER_256_999 ();
 FILLER_ASAP7_75t_R FILLER_256_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_256_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_256_1060 ();
 FILLER_ASAP7_75t_R FILLER_256_1083 ();
 DECAPx6_ASAP7_75t_R FILLER_256_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_256_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_256_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_256_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_256_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_257_2 ();
 DECAPx10_ASAP7_75t_R FILLER_257_24 ();
 DECAPx10_ASAP7_75t_R FILLER_257_46 ();
 DECAPx10_ASAP7_75t_R FILLER_257_68 ();
 DECAPx10_ASAP7_75t_R FILLER_257_90 ();
 DECAPx10_ASAP7_75t_R FILLER_257_112 ();
 DECAPx10_ASAP7_75t_R FILLER_257_134 ();
 DECAPx10_ASAP7_75t_R FILLER_257_156 ();
 DECAPx10_ASAP7_75t_R FILLER_257_178 ();
 DECAPx10_ASAP7_75t_R FILLER_257_200 ();
 DECAPx10_ASAP7_75t_R FILLER_257_222 ();
 DECAPx10_ASAP7_75t_R FILLER_257_244 ();
 DECAPx10_ASAP7_75t_R FILLER_257_266 ();
 DECAPx10_ASAP7_75t_R FILLER_257_288 ();
 DECAPx10_ASAP7_75t_R FILLER_257_310 ();
 DECAPx2_ASAP7_75t_R FILLER_257_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_338 ();
 FILLER_ASAP7_75t_R FILLER_257_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_344 ();
 DECAPx1_ASAP7_75t_R FILLER_257_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_384 ();
 FILLER_ASAP7_75t_R FILLER_257_388 ();
 DECAPx4_ASAP7_75t_R FILLER_257_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_429 ();
 DECAPx10_ASAP7_75t_R FILLER_257_462 ();
 DECAPx10_ASAP7_75t_R FILLER_257_484 ();
 DECAPx10_ASAP7_75t_R FILLER_257_506 ();
 DECAPx10_ASAP7_75t_R FILLER_257_528 ();
 DECAPx10_ASAP7_75t_R FILLER_257_550 ();
 DECAPx10_ASAP7_75t_R FILLER_257_572 ();
 DECAPx10_ASAP7_75t_R FILLER_257_594 ();
 DECAPx10_ASAP7_75t_R FILLER_257_616 ();
 DECAPx10_ASAP7_75t_R FILLER_257_638 ();
 DECAPx10_ASAP7_75t_R FILLER_257_660 ();
 DECAPx10_ASAP7_75t_R FILLER_257_682 ();
 DECAPx10_ASAP7_75t_R FILLER_257_704 ();
 DECAPx10_ASAP7_75t_R FILLER_257_726 ();
 DECAPx10_ASAP7_75t_R FILLER_257_748 ();
 DECAPx10_ASAP7_75t_R FILLER_257_770 ();
 DECAPx6_ASAP7_75t_R FILLER_257_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_806 ();
 DECAPx6_ASAP7_75t_R FILLER_257_810 ();
 DECAPx1_ASAP7_75t_R FILLER_257_824 ();
 DECAPx6_ASAP7_75t_R FILLER_257_834 ();
 DECAPx4_ASAP7_75t_R FILLER_257_854 ();
 FILLER_ASAP7_75t_R FILLER_257_864 ();
 FILLER_ASAP7_75t_R FILLER_257_875 ();
 DECAPx10_ASAP7_75t_R FILLER_257_880 ();
 DECAPx1_ASAP7_75t_R FILLER_257_914 ();
 FILLER_ASAP7_75t_R FILLER_257_926 ();
 DECAPx2_ASAP7_75t_R FILLER_257_934 ();
 FILLER_ASAP7_75t_R FILLER_257_940 ();
 DECAPx1_ASAP7_75t_R FILLER_257_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_981 ();
 FILLER_ASAP7_75t_R FILLER_257_989 ();
 DECAPx4_ASAP7_75t_R FILLER_257_997 ();
 FILLER_ASAP7_75t_R FILLER_257_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_257_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1088 ();
 FILLER_ASAP7_75t_R FILLER_257_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1346 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1368 ();
 FILLER_ASAP7_75t_R FILLER_257_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_258_2 ();
 DECAPx10_ASAP7_75t_R FILLER_258_24 ();
 DECAPx10_ASAP7_75t_R FILLER_258_46 ();
 DECAPx10_ASAP7_75t_R FILLER_258_68 ();
 DECAPx10_ASAP7_75t_R FILLER_258_90 ();
 DECAPx10_ASAP7_75t_R FILLER_258_112 ();
 DECAPx10_ASAP7_75t_R FILLER_258_134 ();
 DECAPx10_ASAP7_75t_R FILLER_258_156 ();
 DECAPx10_ASAP7_75t_R FILLER_258_178 ();
 DECAPx10_ASAP7_75t_R FILLER_258_200 ();
 DECAPx10_ASAP7_75t_R FILLER_258_222 ();
 DECAPx10_ASAP7_75t_R FILLER_258_244 ();
 DECAPx10_ASAP7_75t_R FILLER_258_266 ();
 DECAPx10_ASAP7_75t_R FILLER_258_288 ();
 DECAPx10_ASAP7_75t_R FILLER_258_310 ();
 DECAPx4_ASAP7_75t_R FILLER_258_332 ();
 FILLER_ASAP7_75t_R FILLER_258_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_344 ();
 DECAPx2_ASAP7_75t_R FILLER_258_351 ();
 FILLER_ASAP7_75t_R FILLER_258_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_359 ();
 DECAPx2_ASAP7_75t_R FILLER_258_363 ();
 FILLER_ASAP7_75t_R FILLER_258_369 ();
 DECAPx2_ASAP7_75t_R FILLER_258_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_403 ();
 DECAPx10_ASAP7_75t_R FILLER_258_407 ();
 DECAPx4_ASAP7_75t_R FILLER_258_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_439 ();
 DECAPx2_ASAP7_75t_R FILLER_258_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_449 ();
 DECAPx2_ASAP7_75t_R FILLER_258_453 ();
 FILLER_ASAP7_75t_R FILLER_258_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_461 ();
 DECAPx10_ASAP7_75t_R FILLER_258_464 ();
 DECAPx10_ASAP7_75t_R FILLER_258_486 ();
 DECAPx10_ASAP7_75t_R FILLER_258_508 ();
 DECAPx10_ASAP7_75t_R FILLER_258_530 ();
 DECAPx10_ASAP7_75t_R FILLER_258_552 ();
 DECAPx10_ASAP7_75t_R FILLER_258_574 ();
 DECAPx10_ASAP7_75t_R FILLER_258_596 ();
 DECAPx10_ASAP7_75t_R FILLER_258_618 ();
 DECAPx10_ASAP7_75t_R FILLER_258_640 ();
 DECAPx10_ASAP7_75t_R FILLER_258_662 ();
 DECAPx10_ASAP7_75t_R FILLER_258_684 ();
 DECAPx10_ASAP7_75t_R FILLER_258_706 ();
 DECAPx10_ASAP7_75t_R FILLER_258_728 ();
 DECAPx10_ASAP7_75t_R FILLER_258_750 ();
 DECAPx6_ASAP7_75t_R FILLER_258_772 ();
 DECAPx1_ASAP7_75t_R FILLER_258_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_790 ();
 FILLER_ASAP7_75t_R FILLER_258_817 ();
 FILLER_ASAP7_75t_R FILLER_258_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_828 ();
 FILLER_ASAP7_75t_R FILLER_258_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_840 ();
 FILLER_ASAP7_75t_R FILLER_258_847 ();
 DECAPx2_ASAP7_75t_R FILLER_258_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_867 ();
 DECAPx6_ASAP7_75t_R FILLER_258_876 ();
 FILLER_ASAP7_75t_R FILLER_258_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_954 ();
 FILLER_ASAP7_75t_R FILLER_258_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_977 ();
 FILLER_ASAP7_75t_R FILLER_258_997 ();
 DECAPx2_ASAP7_75t_R FILLER_258_1020 ();
 FILLER_ASAP7_75t_R FILLER_258_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_1028 ();
 DECAPx4_ASAP7_75t_R FILLER_258_1039 ();
 FILLER_ASAP7_75t_R FILLER_258_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_258_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_1068 ();
 FILLER_ASAP7_75t_R FILLER_258_1080 ();
 FILLER_ASAP7_75t_R FILLER_258_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_258_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_258_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_258_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_259_2 ();
 DECAPx10_ASAP7_75t_R FILLER_259_24 ();
 DECAPx10_ASAP7_75t_R FILLER_259_46 ();
 DECAPx10_ASAP7_75t_R FILLER_259_68 ();
 DECAPx10_ASAP7_75t_R FILLER_259_90 ();
 DECAPx10_ASAP7_75t_R FILLER_259_112 ();
 DECAPx10_ASAP7_75t_R FILLER_259_134 ();
 DECAPx10_ASAP7_75t_R FILLER_259_156 ();
 DECAPx10_ASAP7_75t_R FILLER_259_178 ();
 DECAPx10_ASAP7_75t_R FILLER_259_200 ();
 DECAPx10_ASAP7_75t_R FILLER_259_222 ();
 DECAPx10_ASAP7_75t_R FILLER_259_244 ();
 DECAPx10_ASAP7_75t_R FILLER_259_266 ();
 DECAPx10_ASAP7_75t_R FILLER_259_288 ();
 DECAPx10_ASAP7_75t_R FILLER_259_310 ();
 DECAPx10_ASAP7_75t_R FILLER_259_332 ();
 DECAPx10_ASAP7_75t_R FILLER_259_354 ();
 DECAPx10_ASAP7_75t_R FILLER_259_376 ();
 DECAPx10_ASAP7_75t_R FILLER_259_398 ();
 DECAPx10_ASAP7_75t_R FILLER_259_420 ();
 DECAPx10_ASAP7_75t_R FILLER_259_442 ();
 DECAPx10_ASAP7_75t_R FILLER_259_464 ();
 DECAPx10_ASAP7_75t_R FILLER_259_486 ();
 DECAPx10_ASAP7_75t_R FILLER_259_508 ();
 DECAPx10_ASAP7_75t_R FILLER_259_530 ();
 DECAPx10_ASAP7_75t_R FILLER_259_552 ();
 DECAPx10_ASAP7_75t_R FILLER_259_574 ();
 DECAPx10_ASAP7_75t_R FILLER_259_596 ();
 DECAPx10_ASAP7_75t_R FILLER_259_618 ();
 DECAPx10_ASAP7_75t_R FILLER_259_640 ();
 DECAPx10_ASAP7_75t_R FILLER_259_662 ();
 DECAPx10_ASAP7_75t_R FILLER_259_684 ();
 DECAPx10_ASAP7_75t_R FILLER_259_706 ();
 DECAPx10_ASAP7_75t_R FILLER_259_728 ();
 DECAPx10_ASAP7_75t_R FILLER_259_750 ();
 DECAPx4_ASAP7_75t_R FILLER_259_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_830 ();
 DECAPx1_ASAP7_75t_R FILLER_259_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_859 ();
 DECAPx4_ASAP7_75t_R FILLER_259_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_926 ();
 DECAPx2_ASAP7_75t_R FILLER_259_931 ();
 DECAPx6_ASAP7_75t_R FILLER_259_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_968 ();
 DECAPx2_ASAP7_75t_R FILLER_259_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_978 ();
 DECAPx1_ASAP7_75t_R FILLER_259_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_996 ();
 DECAPx6_ASAP7_75t_R FILLER_259_1014 ();
 FILLER_ASAP7_75t_R FILLER_259_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1030 ();
 FILLER_ASAP7_75t_R FILLER_259_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1040 ();
 FILLER_ASAP7_75t_R FILLER_259_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_259_1069 ();
 FILLER_ASAP7_75t_R FILLER_259_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1085 ();
 DECAPx1_ASAP7_75t_R FILLER_259_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1102 ();
 FILLER_ASAP7_75t_R FILLER_259_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1351 ();
 DECAPx6_ASAP7_75t_R FILLER_259_1373 ();
 DECAPx1_ASAP7_75t_R FILLER_259_1387 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_260_2 ();
 DECAPx10_ASAP7_75t_R FILLER_260_24 ();
 DECAPx10_ASAP7_75t_R FILLER_260_46 ();
 DECAPx10_ASAP7_75t_R FILLER_260_68 ();
 DECAPx10_ASAP7_75t_R FILLER_260_90 ();
 DECAPx10_ASAP7_75t_R FILLER_260_112 ();
 DECAPx10_ASAP7_75t_R FILLER_260_134 ();
 DECAPx10_ASAP7_75t_R FILLER_260_156 ();
 DECAPx10_ASAP7_75t_R FILLER_260_178 ();
 DECAPx10_ASAP7_75t_R FILLER_260_200 ();
 DECAPx10_ASAP7_75t_R FILLER_260_222 ();
 DECAPx10_ASAP7_75t_R FILLER_260_244 ();
 DECAPx10_ASAP7_75t_R FILLER_260_266 ();
 DECAPx10_ASAP7_75t_R FILLER_260_288 ();
 DECAPx10_ASAP7_75t_R FILLER_260_310 ();
 DECAPx10_ASAP7_75t_R FILLER_260_332 ();
 DECAPx10_ASAP7_75t_R FILLER_260_354 ();
 DECAPx10_ASAP7_75t_R FILLER_260_376 ();
 DECAPx10_ASAP7_75t_R FILLER_260_398 ();
 DECAPx10_ASAP7_75t_R FILLER_260_420 ();
 DECAPx6_ASAP7_75t_R FILLER_260_442 ();
 DECAPx2_ASAP7_75t_R FILLER_260_456 ();
 DECAPx10_ASAP7_75t_R FILLER_260_464 ();
 DECAPx10_ASAP7_75t_R FILLER_260_486 ();
 DECAPx10_ASAP7_75t_R FILLER_260_508 ();
 DECAPx10_ASAP7_75t_R FILLER_260_530 ();
 DECAPx10_ASAP7_75t_R FILLER_260_552 ();
 DECAPx10_ASAP7_75t_R FILLER_260_574 ();
 DECAPx10_ASAP7_75t_R FILLER_260_596 ();
 DECAPx10_ASAP7_75t_R FILLER_260_618 ();
 DECAPx10_ASAP7_75t_R FILLER_260_640 ();
 DECAPx10_ASAP7_75t_R FILLER_260_662 ();
 DECAPx10_ASAP7_75t_R FILLER_260_684 ();
 DECAPx10_ASAP7_75t_R FILLER_260_706 ();
 DECAPx10_ASAP7_75t_R FILLER_260_728 ();
 DECAPx10_ASAP7_75t_R FILLER_260_750 ();
 DECAPx10_ASAP7_75t_R FILLER_260_772 ();
 FILLER_ASAP7_75t_R FILLER_260_794 ();
 DECAPx2_ASAP7_75t_R FILLER_260_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_805 ();
 DECAPx4_ASAP7_75t_R FILLER_260_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_819 ();
 DECAPx2_ASAP7_75t_R FILLER_260_823 ();
 FILLER_ASAP7_75t_R FILLER_260_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_842 ();
 FILLER_ASAP7_75t_R FILLER_260_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_857 ();
 DECAPx4_ASAP7_75t_R FILLER_260_884 ();
 DECAPx2_ASAP7_75t_R FILLER_260_910 ();
 DECAPx10_ASAP7_75t_R FILLER_260_919 ();
 DECAPx2_ASAP7_75t_R FILLER_260_947 ();
 FILLER_ASAP7_75t_R FILLER_260_953 ();
 FILLER_ASAP7_75t_R FILLER_260_981 ();
 FILLER_ASAP7_75t_R FILLER_260_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_994 ();
 DECAPx2_ASAP7_75t_R FILLER_260_1021 ();
 FILLER_ASAP7_75t_R FILLER_260_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1029 ();
 DECAPx1_ASAP7_75t_R FILLER_260_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1043 ();
 DECAPx4_ASAP7_75t_R FILLER_260_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1087 ();
 DECAPx4_ASAP7_75t_R FILLER_260_1103 ();
 FILLER_ASAP7_75t_R FILLER_260_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_260_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1361 ();
 FILLER_ASAP7_75t_R FILLER_260_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_260_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_261_2 ();
 DECAPx10_ASAP7_75t_R FILLER_261_24 ();
 DECAPx10_ASAP7_75t_R FILLER_261_46 ();
 DECAPx10_ASAP7_75t_R FILLER_261_68 ();
 DECAPx10_ASAP7_75t_R FILLER_261_90 ();
 DECAPx10_ASAP7_75t_R FILLER_261_112 ();
 DECAPx10_ASAP7_75t_R FILLER_261_134 ();
 DECAPx10_ASAP7_75t_R FILLER_261_156 ();
 DECAPx10_ASAP7_75t_R FILLER_261_178 ();
 DECAPx10_ASAP7_75t_R FILLER_261_200 ();
 DECAPx10_ASAP7_75t_R FILLER_261_222 ();
 DECAPx10_ASAP7_75t_R FILLER_261_244 ();
 DECAPx10_ASAP7_75t_R FILLER_261_266 ();
 DECAPx10_ASAP7_75t_R FILLER_261_288 ();
 DECAPx10_ASAP7_75t_R FILLER_261_310 ();
 DECAPx10_ASAP7_75t_R FILLER_261_332 ();
 DECAPx10_ASAP7_75t_R FILLER_261_354 ();
 DECAPx10_ASAP7_75t_R FILLER_261_376 ();
 DECAPx10_ASAP7_75t_R FILLER_261_398 ();
 DECAPx10_ASAP7_75t_R FILLER_261_420 ();
 DECAPx10_ASAP7_75t_R FILLER_261_442 ();
 DECAPx10_ASAP7_75t_R FILLER_261_464 ();
 DECAPx10_ASAP7_75t_R FILLER_261_486 ();
 DECAPx10_ASAP7_75t_R FILLER_261_508 ();
 DECAPx10_ASAP7_75t_R FILLER_261_530 ();
 DECAPx10_ASAP7_75t_R FILLER_261_552 ();
 DECAPx10_ASAP7_75t_R FILLER_261_574 ();
 DECAPx10_ASAP7_75t_R FILLER_261_596 ();
 DECAPx10_ASAP7_75t_R FILLER_261_618 ();
 DECAPx10_ASAP7_75t_R FILLER_261_640 ();
 DECAPx10_ASAP7_75t_R FILLER_261_662 ();
 DECAPx10_ASAP7_75t_R FILLER_261_684 ();
 DECAPx10_ASAP7_75t_R FILLER_261_706 ();
 DECAPx10_ASAP7_75t_R FILLER_261_728 ();
 DECAPx10_ASAP7_75t_R FILLER_261_750 ();
 DECAPx10_ASAP7_75t_R FILLER_261_772 ();
 DECAPx6_ASAP7_75t_R FILLER_261_794 ();
 DECAPx2_ASAP7_75t_R FILLER_261_808 ();
 DECAPx10_ASAP7_75t_R FILLER_261_829 ();
 DECAPx6_ASAP7_75t_R FILLER_261_851 ();
 DECAPx1_ASAP7_75t_R FILLER_261_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_869 ();
 DECAPx2_ASAP7_75t_R FILLER_261_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_889 ();
 DECAPx10_ASAP7_75t_R FILLER_261_900 ();
 FILLER_ASAP7_75t_R FILLER_261_922 ();
 FILLER_ASAP7_75t_R FILLER_261_926 ();
 FILLER_ASAP7_75t_R FILLER_261_934 ();
 DECAPx2_ASAP7_75t_R FILLER_261_953 ();
 FILLER_ASAP7_75t_R FILLER_261_959 ();
 DECAPx10_ASAP7_75t_R FILLER_261_964 ();
 DECAPx6_ASAP7_75t_R FILLER_261_994 ();
 FILLER_ASAP7_75t_R FILLER_261_1008 ();
 FILLER_ASAP7_75t_R FILLER_261_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_261_1070 ();
 DECAPx4_ASAP7_75t_R FILLER_261_1103 ();
 DECAPx2_ASAP7_75t_R FILLER_261_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1347 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_262_2 ();
 DECAPx10_ASAP7_75t_R FILLER_262_24 ();
 DECAPx10_ASAP7_75t_R FILLER_262_46 ();
 DECAPx10_ASAP7_75t_R FILLER_262_68 ();
 DECAPx10_ASAP7_75t_R FILLER_262_90 ();
 DECAPx10_ASAP7_75t_R FILLER_262_112 ();
 DECAPx10_ASAP7_75t_R FILLER_262_134 ();
 DECAPx10_ASAP7_75t_R FILLER_262_156 ();
 DECAPx10_ASAP7_75t_R FILLER_262_178 ();
 DECAPx10_ASAP7_75t_R FILLER_262_200 ();
 DECAPx10_ASAP7_75t_R FILLER_262_222 ();
 DECAPx10_ASAP7_75t_R FILLER_262_244 ();
 DECAPx10_ASAP7_75t_R FILLER_262_266 ();
 DECAPx10_ASAP7_75t_R FILLER_262_288 ();
 DECAPx10_ASAP7_75t_R FILLER_262_310 ();
 DECAPx10_ASAP7_75t_R FILLER_262_332 ();
 DECAPx10_ASAP7_75t_R FILLER_262_354 ();
 DECAPx10_ASAP7_75t_R FILLER_262_376 ();
 DECAPx10_ASAP7_75t_R FILLER_262_398 ();
 DECAPx10_ASAP7_75t_R FILLER_262_420 ();
 DECAPx6_ASAP7_75t_R FILLER_262_442 ();
 DECAPx2_ASAP7_75t_R FILLER_262_456 ();
 DECAPx10_ASAP7_75t_R FILLER_262_464 ();
 DECAPx10_ASAP7_75t_R FILLER_262_486 ();
 DECAPx10_ASAP7_75t_R FILLER_262_508 ();
 DECAPx10_ASAP7_75t_R FILLER_262_530 ();
 DECAPx10_ASAP7_75t_R FILLER_262_552 ();
 DECAPx10_ASAP7_75t_R FILLER_262_574 ();
 DECAPx10_ASAP7_75t_R FILLER_262_596 ();
 DECAPx10_ASAP7_75t_R FILLER_262_618 ();
 DECAPx10_ASAP7_75t_R FILLER_262_640 ();
 DECAPx10_ASAP7_75t_R FILLER_262_662 ();
 DECAPx10_ASAP7_75t_R FILLER_262_684 ();
 DECAPx10_ASAP7_75t_R FILLER_262_706 ();
 DECAPx10_ASAP7_75t_R FILLER_262_728 ();
 DECAPx10_ASAP7_75t_R FILLER_262_750 ();
 DECAPx10_ASAP7_75t_R FILLER_262_772 ();
 DECAPx2_ASAP7_75t_R FILLER_262_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_800 ();
 DECAPx6_ASAP7_75t_R FILLER_262_804 ();
 FILLER_ASAP7_75t_R FILLER_262_818 ();
 DECAPx2_ASAP7_75t_R FILLER_262_832 ();
 DECAPx2_ASAP7_75t_R FILLER_262_844 ();
 DECAPx2_ASAP7_75t_R FILLER_262_876 ();
 FILLER_ASAP7_75t_R FILLER_262_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_945 ();
 DECAPx4_ASAP7_75t_R FILLER_262_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_982 ();
 DECAPx6_ASAP7_75t_R FILLER_262_992 ();
 FILLER_ASAP7_75t_R FILLER_262_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1066 ();
 DECAPx1_ASAP7_75t_R FILLER_262_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_262_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_262_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_262_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_263_2 ();
 DECAPx10_ASAP7_75t_R FILLER_263_24 ();
 DECAPx10_ASAP7_75t_R FILLER_263_46 ();
 DECAPx10_ASAP7_75t_R FILLER_263_68 ();
 DECAPx10_ASAP7_75t_R FILLER_263_90 ();
 DECAPx10_ASAP7_75t_R FILLER_263_112 ();
 DECAPx10_ASAP7_75t_R FILLER_263_134 ();
 DECAPx10_ASAP7_75t_R FILLER_263_156 ();
 DECAPx10_ASAP7_75t_R FILLER_263_178 ();
 DECAPx10_ASAP7_75t_R FILLER_263_200 ();
 DECAPx10_ASAP7_75t_R FILLER_263_222 ();
 DECAPx10_ASAP7_75t_R FILLER_263_244 ();
 DECAPx10_ASAP7_75t_R FILLER_263_266 ();
 DECAPx10_ASAP7_75t_R FILLER_263_288 ();
 DECAPx10_ASAP7_75t_R FILLER_263_310 ();
 DECAPx10_ASAP7_75t_R FILLER_263_332 ();
 DECAPx10_ASAP7_75t_R FILLER_263_354 ();
 DECAPx10_ASAP7_75t_R FILLER_263_376 ();
 DECAPx10_ASAP7_75t_R FILLER_263_398 ();
 DECAPx10_ASAP7_75t_R FILLER_263_420 ();
 DECAPx10_ASAP7_75t_R FILLER_263_442 ();
 DECAPx10_ASAP7_75t_R FILLER_263_464 ();
 DECAPx10_ASAP7_75t_R FILLER_263_486 ();
 DECAPx10_ASAP7_75t_R FILLER_263_508 ();
 DECAPx10_ASAP7_75t_R FILLER_263_530 ();
 DECAPx10_ASAP7_75t_R FILLER_263_552 ();
 DECAPx10_ASAP7_75t_R FILLER_263_574 ();
 DECAPx10_ASAP7_75t_R FILLER_263_596 ();
 DECAPx10_ASAP7_75t_R FILLER_263_618 ();
 DECAPx10_ASAP7_75t_R FILLER_263_640 ();
 DECAPx10_ASAP7_75t_R FILLER_263_662 ();
 DECAPx10_ASAP7_75t_R FILLER_263_684 ();
 DECAPx10_ASAP7_75t_R FILLER_263_706 ();
 DECAPx10_ASAP7_75t_R FILLER_263_728 ();
 DECAPx10_ASAP7_75t_R FILLER_263_750 ();
 DECAPx6_ASAP7_75t_R FILLER_263_772 ();
 FILLER_ASAP7_75t_R FILLER_263_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_814 ();
 DECAPx2_ASAP7_75t_R FILLER_263_827 ();
 FILLER_ASAP7_75t_R FILLER_263_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_835 ();
 DECAPx10_ASAP7_75t_R FILLER_263_868 ();
 DECAPx4_ASAP7_75t_R FILLER_263_890 ();
 FILLER_ASAP7_75t_R FILLER_263_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_902 ();
 FILLER_ASAP7_75t_R FILLER_263_926 ();
 FILLER_ASAP7_75t_R FILLER_263_942 ();
 DECAPx10_ASAP7_75t_R FILLER_263_950 ();
 DECAPx1_ASAP7_75t_R FILLER_263_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_976 ();
 DECAPx4_ASAP7_75t_R FILLER_263_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1013 ();
 FILLER_ASAP7_75t_R FILLER_263_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_263_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_263_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_263_1078 ();
 DECAPx1_ASAP7_75t_R FILLER_263_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_263_1386 ();
 DECAPx10_ASAP7_75t_R FILLER_264_2 ();
 DECAPx10_ASAP7_75t_R FILLER_264_24 ();
 DECAPx10_ASAP7_75t_R FILLER_264_46 ();
 DECAPx10_ASAP7_75t_R FILLER_264_68 ();
 DECAPx10_ASAP7_75t_R FILLER_264_90 ();
 DECAPx10_ASAP7_75t_R FILLER_264_112 ();
 DECAPx10_ASAP7_75t_R FILLER_264_134 ();
 DECAPx10_ASAP7_75t_R FILLER_264_156 ();
 DECAPx10_ASAP7_75t_R FILLER_264_178 ();
 DECAPx10_ASAP7_75t_R FILLER_264_200 ();
 DECAPx10_ASAP7_75t_R FILLER_264_222 ();
 DECAPx10_ASAP7_75t_R FILLER_264_244 ();
 DECAPx10_ASAP7_75t_R FILLER_264_266 ();
 DECAPx10_ASAP7_75t_R FILLER_264_288 ();
 DECAPx10_ASAP7_75t_R FILLER_264_310 ();
 DECAPx10_ASAP7_75t_R FILLER_264_332 ();
 DECAPx10_ASAP7_75t_R FILLER_264_354 ();
 DECAPx10_ASAP7_75t_R FILLER_264_376 ();
 DECAPx10_ASAP7_75t_R FILLER_264_398 ();
 DECAPx10_ASAP7_75t_R FILLER_264_420 ();
 DECAPx6_ASAP7_75t_R FILLER_264_442 ();
 DECAPx2_ASAP7_75t_R FILLER_264_456 ();
 DECAPx10_ASAP7_75t_R FILLER_264_464 ();
 DECAPx10_ASAP7_75t_R FILLER_264_486 ();
 DECAPx10_ASAP7_75t_R FILLER_264_508 ();
 DECAPx10_ASAP7_75t_R FILLER_264_530 ();
 DECAPx10_ASAP7_75t_R FILLER_264_552 ();
 DECAPx10_ASAP7_75t_R FILLER_264_574 ();
 DECAPx10_ASAP7_75t_R FILLER_264_596 ();
 DECAPx10_ASAP7_75t_R FILLER_264_618 ();
 DECAPx10_ASAP7_75t_R FILLER_264_640 ();
 DECAPx10_ASAP7_75t_R FILLER_264_662 ();
 DECAPx10_ASAP7_75t_R FILLER_264_684 ();
 DECAPx10_ASAP7_75t_R FILLER_264_706 ();
 DECAPx10_ASAP7_75t_R FILLER_264_728 ();
 DECAPx10_ASAP7_75t_R FILLER_264_750 ();
 DECAPx6_ASAP7_75t_R FILLER_264_772 ();
 FILLER_ASAP7_75t_R FILLER_264_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_814 ();
 FILLER_ASAP7_75t_R FILLER_264_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_838 ();
 DECAPx2_ASAP7_75t_R FILLER_264_845 ();
 DECAPx1_ASAP7_75t_R FILLER_264_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_858 ();
 DECAPx4_ASAP7_75t_R FILLER_264_868 ();
 FILLER_ASAP7_75t_R FILLER_264_878 ();
 DECAPx6_ASAP7_75t_R FILLER_264_886 ();
 FILLER_ASAP7_75t_R FILLER_264_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_902 ();
 DECAPx4_ASAP7_75t_R FILLER_264_913 ();
 FILLER_ASAP7_75t_R FILLER_264_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_925 ();
 FILLER_ASAP7_75t_R FILLER_264_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_939 ();
 DECAPx2_ASAP7_75t_R FILLER_264_948 ();
 FILLER_ASAP7_75t_R FILLER_264_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_956 ();
 DECAPx4_ASAP7_75t_R FILLER_264_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_973 ();
 DECAPx2_ASAP7_75t_R FILLER_264_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_990 ();
 DECAPx1_ASAP7_75t_R FILLER_264_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_998 ();
 DECAPx4_ASAP7_75t_R FILLER_264_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_264_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_1031 ();
 DECAPx1_ASAP7_75t_R FILLER_264_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_264_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_264_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_264_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_265_2 ();
 DECAPx10_ASAP7_75t_R FILLER_265_24 ();
 DECAPx10_ASAP7_75t_R FILLER_265_46 ();
 DECAPx10_ASAP7_75t_R FILLER_265_68 ();
 DECAPx10_ASAP7_75t_R FILLER_265_90 ();
 DECAPx10_ASAP7_75t_R FILLER_265_112 ();
 DECAPx10_ASAP7_75t_R FILLER_265_134 ();
 DECAPx10_ASAP7_75t_R FILLER_265_156 ();
 DECAPx10_ASAP7_75t_R FILLER_265_178 ();
 DECAPx10_ASAP7_75t_R FILLER_265_200 ();
 DECAPx10_ASAP7_75t_R FILLER_265_222 ();
 DECAPx10_ASAP7_75t_R FILLER_265_244 ();
 DECAPx10_ASAP7_75t_R FILLER_265_266 ();
 DECAPx10_ASAP7_75t_R FILLER_265_288 ();
 DECAPx10_ASAP7_75t_R FILLER_265_310 ();
 DECAPx10_ASAP7_75t_R FILLER_265_332 ();
 DECAPx10_ASAP7_75t_R FILLER_265_354 ();
 DECAPx10_ASAP7_75t_R FILLER_265_376 ();
 DECAPx10_ASAP7_75t_R FILLER_265_398 ();
 DECAPx10_ASAP7_75t_R FILLER_265_420 ();
 DECAPx10_ASAP7_75t_R FILLER_265_442 ();
 DECAPx10_ASAP7_75t_R FILLER_265_464 ();
 DECAPx10_ASAP7_75t_R FILLER_265_486 ();
 DECAPx10_ASAP7_75t_R FILLER_265_508 ();
 DECAPx10_ASAP7_75t_R FILLER_265_530 ();
 DECAPx10_ASAP7_75t_R FILLER_265_552 ();
 DECAPx10_ASAP7_75t_R FILLER_265_574 ();
 DECAPx10_ASAP7_75t_R FILLER_265_596 ();
 DECAPx10_ASAP7_75t_R FILLER_265_618 ();
 DECAPx10_ASAP7_75t_R FILLER_265_640 ();
 DECAPx10_ASAP7_75t_R FILLER_265_662 ();
 DECAPx10_ASAP7_75t_R FILLER_265_684 ();
 DECAPx10_ASAP7_75t_R FILLER_265_706 ();
 DECAPx10_ASAP7_75t_R FILLER_265_728 ();
 DECAPx10_ASAP7_75t_R FILLER_265_750 ();
 DECAPx10_ASAP7_75t_R FILLER_265_772 ();
 DECAPx2_ASAP7_75t_R FILLER_265_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_800 ();
 DECAPx2_ASAP7_75t_R FILLER_265_804 ();
 FILLER_ASAP7_75t_R FILLER_265_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_829 ();
 DECAPx6_ASAP7_75t_R FILLER_265_844 ();
 DECAPx4_ASAP7_75t_R FILLER_265_864 ();
 FILLER_ASAP7_75t_R FILLER_265_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_879 ();
 DECAPx2_ASAP7_75t_R FILLER_265_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_892 ();
 DECAPx4_ASAP7_75t_R FILLER_265_896 ();
 DECAPx2_ASAP7_75t_R FILLER_265_912 ();
 FILLER_ASAP7_75t_R FILLER_265_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_926 ();
 FILLER_ASAP7_75t_R FILLER_265_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_938 ();
 DECAPx1_ASAP7_75t_R FILLER_265_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_957 ();
 DECAPx2_ASAP7_75t_R FILLER_265_984 ();
 FILLER_ASAP7_75t_R FILLER_265_990 ();
 FILLER_ASAP7_75t_R FILLER_265_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_997 ();
 DECAPx2_ASAP7_75t_R FILLER_265_1009 ();
 FILLER_ASAP7_75t_R FILLER_265_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_265_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_265_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_265_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_265_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_266_2 ();
 DECAPx10_ASAP7_75t_R FILLER_266_24 ();
 DECAPx10_ASAP7_75t_R FILLER_266_46 ();
 DECAPx10_ASAP7_75t_R FILLER_266_68 ();
 DECAPx10_ASAP7_75t_R FILLER_266_90 ();
 DECAPx10_ASAP7_75t_R FILLER_266_112 ();
 DECAPx10_ASAP7_75t_R FILLER_266_134 ();
 DECAPx10_ASAP7_75t_R FILLER_266_156 ();
 DECAPx10_ASAP7_75t_R FILLER_266_178 ();
 DECAPx10_ASAP7_75t_R FILLER_266_200 ();
 DECAPx10_ASAP7_75t_R FILLER_266_222 ();
 DECAPx10_ASAP7_75t_R FILLER_266_244 ();
 DECAPx10_ASAP7_75t_R FILLER_266_266 ();
 DECAPx10_ASAP7_75t_R FILLER_266_288 ();
 DECAPx10_ASAP7_75t_R FILLER_266_310 ();
 DECAPx10_ASAP7_75t_R FILLER_266_332 ();
 DECAPx10_ASAP7_75t_R FILLER_266_354 ();
 DECAPx10_ASAP7_75t_R FILLER_266_376 ();
 DECAPx10_ASAP7_75t_R FILLER_266_398 ();
 DECAPx10_ASAP7_75t_R FILLER_266_420 ();
 DECAPx6_ASAP7_75t_R FILLER_266_442 ();
 DECAPx2_ASAP7_75t_R FILLER_266_456 ();
 DECAPx10_ASAP7_75t_R FILLER_266_464 ();
 DECAPx10_ASAP7_75t_R FILLER_266_486 ();
 DECAPx10_ASAP7_75t_R FILLER_266_508 ();
 DECAPx10_ASAP7_75t_R FILLER_266_530 ();
 DECAPx10_ASAP7_75t_R FILLER_266_552 ();
 DECAPx10_ASAP7_75t_R FILLER_266_574 ();
 DECAPx10_ASAP7_75t_R FILLER_266_596 ();
 DECAPx10_ASAP7_75t_R FILLER_266_618 ();
 DECAPx10_ASAP7_75t_R FILLER_266_640 ();
 DECAPx10_ASAP7_75t_R FILLER_266_662 ();
 DECAPx10_ASAP7_75t_R FILLER_266_684 ();
 DECAPx10_ASAP7_75t_R FILLER_266_706 ();
 DECAPx10_ASAP7_75t_R FILLER_266_728 ();
 DECAPx10_ASAP7_75t_R FILLER_266_750 ();
 DECAPx10_ASAP7_75t_R FILLER_266_772 ();
 DECAPx6_ASAP7_75t_R FILLER_266_794 ();
 DECAPx1_ASAP7_75t_R FILLER_266_808 ();
 DECAPx2_ASAP7_75t_R FILLER_266_822 ();
 FILLER_ASAP7_75t_R FILLER_266_828 ();
 FILLER_ASAP7_75t_R FILLER_266_834 ();
 FILLER_ASAP7_75t_R FILLER_266_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_844 ();
 DECAPx2_ASAP7_75t_R FILLER_266_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_867 ();
 FILLER_ASAP7_75t_R FILLER_266_876 ();
 FILLER_ASAP7_75t_R FILLER_266_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_906 ();
 DECAPx1_ASAP7_75t_R FILLER_266_919 ();
 FILLER_ASAP7_75t_R FILLER_266_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_937 ();
 DECAPx2_ASAP7_75t_R FILLER_266_950 ();
 DECAPx4_ASAP7_75t_R FILLER_266_962 ();
 FILLER_ASAP7_75t_R FILLER_266_975 ();
 DECAPx2_ASAP7_75t_R FILLER_266_1009 ();
 FILLER_ASAP7_75t_R FILLER_266_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1017 ();
 DECAPx6_ASAP7_75t_R FILLER_266_1032 ();
 FILLER_ASAP7_75t_R FILLER_266_1046 ();
 FILLER_ASAP7_75t_R FILLER_266_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1064 ();
 FILLER_ASAP7_75t_R FILLER_266_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1076 ();
 FILLER_ASAP7_75t_R FILLER_266_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1345 ();
 DECAPx6_ASAP7_75t_R FILLER_266_1367 ();
 DECAPx1_ASAP7_75t_R FILLER_266_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_266_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_267_2 ();
 DECAPx10_ASAP7_75t_R FILLER_267_24 ();
 DECAPx10_ASAP7_75t_R FILLER_267_46 ();
 DECAPx10_ASAP7_75t_R FILLER_267_68 ();
 DECAPx10_ASAP7_75t_R FILLER_267_90 ();
 DECAPx10_ASAP7_75t_R FILLER_267_112 ();
 DECAPx10_ASAP7_75t_R FILLER_267_134 ();
 DECAPx10_ASAP7_75t_R FILLER_267_156 ();
 DECAPx10_ASAP7_75t_R FILLER_267_178 ();
 DECAPx10_ASAP7_75t_R FILLER_267_200 ();
 DECAPx10_ASAP7_75t_R FILLER_267_222 ();
 DECAPx10_ASAP7_75t_R FILLER_267_244 ();
 DECAPx10_ASAP7_75t_R FILLER_267_266 ();
 DECAPx10_ASAP7_75t_R FILLER_267_288 ();
 DECAPx10_ASAP7_75t_R FILLER_267_310 ();
 DECAPx10_ASAP7_75t_R FILLER_267_332 ();
 DECAPx10_ASAP7_75t_R FILLER_267_354 ();
 DECAPx10_ASAP7_75t_R FILLER_267_376 ();
 DECAPx10_ASAP7_75t_R FILLER_267_398 ();
 DECAPx10_ASAP7_75t_R FILLER_267_420 ();
 DECAPx10_ASAP7_75t_R FILLER_267_442 ();
 DECAPx10_ASAP7_75t_R FILLER_267_464 ();
 DECAPx10_ASAP7_75t_R FILLER_267_486 ();
 DECAPx10_ASAP7_75t_R FILLER_267_508 ();
 DECAPx10_ASAP7_75t_R FILLER_267_530 ();
 DECAPx10_ASAP7_75t_R FILLER_267_552 ();
 DECAPx10_ASAP7_75t_R FILLER_267_574 ();
 DECAPx10_ASAP7_75t_R FILLER_267_596 ();
 DECAPx10_ASAP7_75t_R FILLER_267_618 ();
 DECAPx10_ASAP7_75t_R FILLER_267_640 ();
 DECAPx10_ASAP7_75t_R FILLER_267_662 ();
 DECAPx10_ASAP7_75t_R FILLER_267_684 ();
 DECAPx10_ASAP7_75t_R FILLER_267_706 ();
 DECAPx10_ASAP7_75t_R FILLER_267_728 ();
 DECAPx10_ASAP7_75t_R FILLER_267_750 ();
 DECAPx10_ASAP7_75t_R FILLER_267_772 ();
 DECAPx6_ASAP7_75t_R FILLER_267_794 ();
 DECAPx1_ASAP7_75t_R FILLER_267_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_812 ();
 FILLER_ASAP7_75t_R FILLER_267_839 ();
 FILLER_ASAP7_75t_R FILLER_267_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_859 ();
 FILLER_ASAP7_75t_R FILLER_267_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_874 ();
 DECAPx1_ASAP7_75t_R FILLER_267_881 ();
 FILLER_ASAP7_75t_R FILLER_267_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_897 ();
 DECAPx6_ASAP7_75t_R FILLER_267_926 ();
 FILLER_ASAP7_75t_R FILLER_267_940 ();
 FILLER_ASAP7_75t_R FILLER_267_954 ();
 DECAPx2_ASAP7_75t_R FILLER_267_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_978 ();
 DECAPx2_ASAP7_75t_R FILLER_267_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_995 ();
 FILLER_ASAP7_75t_R FILLER_267_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_267_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1035 ();
 DECAPx4_ASAP7_75t_R FILLER_267_1039 ();
 FILLER_ASAP7_75t_R FILLER_267_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_267_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1352 ();
 DECAPx6_ASAP7_75t_R FILLER_267_1374 ();
 DECAPx1_ASAP7_75t_R FILLER_267_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_268_2 ();
 DECAPx10_ASAP7_75t_R FILLER_268_24 ();
 DECAPx10_ASAP7_75t_R FILLER_268_46 ();
 DECAPx10_ASAP7_75t_R FILLER_268_68 ();
 DECAPx10_ASAP7_75t_R FILLER_268_90 ();
 DECAPx10_ASAP7_75t_R FILLER_268_112 ();
 DECAPx10_ASAP7_75t_R FILLER_268_134 ();
 DECAPx10_ASAP7_75t_R FILLER_268_156 ();
 DECAPx10_ASAP7_75t_R FILLER_268_178 ();
 DECAPx10_ASAP7_75t_R FILLER_268_200 ();
 DECAPx10_ASAP7_75t_R FILLER_268_222 ();
 DECAPx10_ASAP7_75t_R FILLER_268_244 ();
 DECAPx10_ASAP7_75t_R FILLER_268_266 ();
 DECAPx10_ASAP7_75t_R FILLER_268_288 ();
 DECAPx10_ASAP7_75t_R FILLER_268_310 ();
 DECAPx10_ASAP7_75t_R FILLER_268_332 ();
 DECAPx10_ASAP7_75t_R FILLER_268_354 ();
 DECAPx10_ASAP7_75t_R FILLER_268_376 ();
 DECAPx10_ASAP7_75t_R FILLER_268_398 ();
 DECAPx10_ASAP7_75t_R FILLER_268_420 ();
 DECAPx6_ASAP7_75t_R FILLER_268_442 ();
 DECAPx2_ASAP7_75t_R FILLER_268_456 ();
 DECAPx10_ASAP7_75t_R FILLER_268_464 ();
 DECAPx10_ASAP7_75t_R FILLER_268_486 ();
 DECAPx10_ASAP7_75t_R FILLER_268_508 ();
 DECAPx10_ASAP7_75t_R FILLER_268_530 ();
 DECAPx10_ASAP7_75t_R FILLER_268_552 ();
 DECAPx10_ASAP7_75t_R FILLER_268_574 ();
 DECAPx10_ASAP7_75t_R FILLER_268_596 ();
 DECAPx10_ASAP7_75t_R FILLER_268_618 ();
 DECAPx10_ASAP7_75t_R FILLER_268_640 ();
 DECAPx10_ASAP7_75t_R FILLER_268_662 ();
 DECAPx10_ASAP7_75t_R FILLER_268_684 ();
 DECAPx10_ASAP7_75t_R FILLER_268_706 ();
 DECAPx10_ASAP7_75t_R FILLER_268_728 ();
 DECAPx10_ASAP7_75t_R FILLER_268_750 ();
 DECAPx10_ASAP7_75t_R FILLER_268_772 ();
 DECAPx6_ASAP7_75t_R FILLER_268_794 ();
 DECAPx1_ASAP7_75t_R FILLER_268_808 ();
 DECAPx6_ASAP7_75t_R FILLER_268_824 ();
 DECAPx1_ASAP7_75t_R FILLER_268_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_859 ();
 DECAPx4_ASAP7_75t_R FILLER_268_867 ();
 FILLER_ASAP7_75t_R FILLER_268_877 ();
 DECAPx6_ASAP7_75t_R FILLER_268_885 ();
 FILLER_ASAP7_75t_R FILLER_268_899 ();
 DECAPx2_ASAP7_75t_R FILLER_268_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_913 ();
 DECAPx4_ASAP7_75t_R FILLER_268_917 ();
 DECAPx2_ASAP7_75t_R FILLER_268_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_945 ();
 DECAPx6_ASAP7_75t_R FILLER_268_984 ();
 DECAPx1_ASAP7_75t_R FILLER_268_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1010 ();
 FILLER_ASAP7_75t_R FILLER_268_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1021 ();
 FILLER_ASAP7_75t_R FILLER_268_1033 ();
 DECAPx6_ASAP7_75t_R FILLER_268_1046 ();
 FILLER_ASAP7_75t_R FILLER_268_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1062 ();
 DECAPx4_ASAP7_75t_R FILLER_268_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_268_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_268_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_268_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_269_2 ();
 DECAPx10_ASAP7_75t_R FILLER_269_24 ();
 DECAPx10_ASAP7_75t_R FILLER_269_46 ();
 DECAPx10_ASAP7_75t_R FILLER_269_68 ();
 DECAPx10_ASAP7_75t_R FILLER_269_90 ();
 DECAPx10_ASAP7_75t_R FILLER_269_112 ();
 DECAPx10_ASAP7_75t_R FILLER_269_134 ();
 DECAPx10_ASAP7_75t_R FILLER_269_156 ();
 DECAPx10_ASAP7_75t_R FILLER_269_178 ();
 DECAPx10_ASAP7_75t_R FILLER_269_200 ();
 DECAPx10_ASAP7_75t_R FILLER_269_222 ();
 DECAPx10_ASAP7_75t_R FILLER_269_244 ();
 DECAPx10_ASAP7_75t_R FILLER_269_266 ();
 DECAPx10_ASAP7_75t_R FILLER_269_288 ();
 DECAPx10_ASAP7_75t_R FILLER_269_310 ();
 DECAPx10_ASAP7_75t_R FILLER_269_332 ();
 DECAPx10_ASAP7_75t_R FILLER_269_354 ();
 DECAPx10_ASAP7_75t_R FILLER_269_376 ();
 DECAPx10_ASAP7_75t_R FILLER_269_398 ();
 DECAPx10_ASAP7_75t_R FILLER_269_420 ();
 DECAPx10_ASAP7_75t_R FILLER_269_442 ();
 DECAPx10_ASAP7_75t_R FILLER_269_464 ();
 DECAPx10_ASAP7_75t_R FILLER_269_486 ();
 DECAPx10_ASAP7_75t_R FILLER_269_508 ();
 DECAPx10_ASAP7_75t_R FILLER_269_530 ();
 DECAPx10_ASAP7_75t_R FILLER_269_552 ();
 DECAPx10_ASAP7_75t_R FILLER_269_574 ();
 DECAPx10_ASAP7_75t_R FILLER_269_596 ();
 DECAPx10_ASAP7_75t_R FILLER_269_618 ();
 DECAPx10_ASAP7_75t_R FILLER_269_640 ();
 DECAPx10_ASAP7_75t_R FILLER_269_662 ();
 DECAPx10_ASAP7_75t_R FILLER_269_684 ();
 DECAPx10_ASAP7_75t_R FILLER_269_706 ();
 DECAPx10_ASAP7_75t_R FILLER_269_728 ();
 DECAPx10_ASAP7_75t_R FILLER_269_750 ();
 DECAPx10_ASAP7_75t_R FILLER_269_772 ();
 DECAPx10_ASAP7_75t_R FILLER_269_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_816 ();
 DECAPx2_ASAP7_75t_R FILLER_269_829 ();
 FILLER_ASAP7_75t_R FILLER_269_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_837 ();
 DECAPx4_ASAP7_75t_R FILLER_269_844 ();
 FILLER_ASAP7_75t_R FILLER_269_854 ();
 FILLER_ASAP7_75t_R FILLER_269_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_864 ();
 DECAPx2_ASAP7_75t_R FILLER_269_871 ();
 DECAPx4_ASAP7_75t_R FILLER_269_889 ();
 FILLER_ASAP7_75t_R FILLER_269_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_901 ();
 DECAPx6_ASAP7_75t_R FILLER_269_908 ();
 FILLER_ASAP7_75t_R FILLER_269_922 ();
 FILLER_ASAP7_75t_R FILLER_269_932 ();
 DECAPx4_ASAP7_75t_R FILLER_269_943 ();
 FILLER_ASAP7_75t_R FILLER_269_953 ();
 DECAPx4_ASAP7_75t_R FILLER_269_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_971 ();
 DECAPx4_ASAP7_75t_R FILLER_269_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_985 ();
 DECAPx1_ASAP7_75t_R FILLER_269_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1048 ();
 FILLER_ASAP7_75t_R FILLER_269_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_269_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_270_2 ();
 DECAPx10_ASAP7_75t_R FILLER_270_24 ();
 DECAPx10_ASAP7_75t_R FILLER_270_46 ();
 DECAPx10_ASAP7_75t_R FILLER_270_68 ();
 DECAPx10_ASAP7_75t_R FILLER_270_90 ();
 DECAPx10_ASAP7_75t_R FILLER_270_112 ();
 DECAPx10_ASAP7_75t_R FILLER_270_134 ();
 DECAPx10_ASAP7_75t_R FILLER_270_156 ();
 DECAPx10_ASAP7_75t_R FILLER_270_178 ();
 DECAPx10_ASAP7_75t_R FILLER_270_200 ();
 DECAPx10_ASAP7_75t_R FILLER_270_222 ();
 DECAPx10_ASAP7_75t_R FILLER_270_244 ();
 DECAPx10_ASAP7_75t_R FILLER_270_266 ();
 DECAPx10_ASAP7_75t_R FILLER_270_288 ();
 DECAPx10_ASAP7_75t_R FILLER_270_310 ();
 DECAPx10_ASAP7_75t_R FILLER_270_332 ();
 DECAPx10_ASAP7_75t_R FILLER_270_354 ();
 DECAPx10_ASAP7_75t_R FILLER_270_376 ();
 DECAPx10_ASAP7_75t_R FILLER_270_398 ();
 DECAPx10_ASAP7_75t_R FILLER_270_420 ();
 DECAPx6_ASAP7_75t_R FILLER_270_442 ();
 DECAPx2_ASAP7_75t_R FILLER_270_456 ();
 DECAPx10_ASAP7_75t_R FILLER_270_464 ();
 DECAPx10_ASAP7_75t_R FILLER_270_486 ();
 DECAPx10_ASAP7_75t_R FILLER_270_508 ();
 DECAPx10_ASAP7_75t_R FILLER_270_530 ();
 DECAPx10_ASAP7_75t_R FILLER_270_552 ();
 DECAPx10_ASAP7_75t_R FILLER_270_574 ();
 DECAPx10_ASAP7_75t_R FILLER_270_596 ();
 DECAPx10_ASAP7_75t_R FILLER_270_618 ();
 DECAPx10_ASAP7_75t_R FILLER_270_640 ();
 DECAPx10_ASAP7_75t_R FILLER_270_662 ();
 DECAPx10_ASAP7_75t_R FILLER_270_684 ();
 DECAPx10_ASAP7_75t_R FILLER_270_706 ();
 DECAPx10_ASAP7_75t_R FILLER_270_728 ();
 DECAPx10_ASAP7_75t_R FILLER_270_750 ();
 DECAPx10_ASAP7_75t_R FILLER_270_772 ();
 DECAPx6_ASAP7_75t_R FILLER_270_794 ();
 FILLER_ASAP7_75t_R FILLER_270_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_810 ();
 FILLER_ASAP7_75t_R FILLER_270_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_837 ();
 FILLER_ASAP7_75t_R FILLER_270_850 ();
 DECAPx2_ASAP7_75t_R FILLER_270_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_885 ();
 DECAPx6_ASAP7_75t_R FILLER_270_906 ();
 FILLER_ASAP7_75t_R FILLER_270_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_922 ();
 FILLER_ASAP7_75t_R FILLER_270_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_937 ();
 DECAPx4_ASAP7_75t_R FILLER_270_947 ();
 DECAPx10_ASAP7_75t_R FILLER_270_963 ();
 DECAPx2_ASAP7_75t_R FILLER_270_985 ();
 FILLER_ASAP7_75t_R FILLER_270_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_993 ();
 FILLER_ASAP7_75t_R FILLER_270_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1002 ();
 FILLER_ASAP7_75t_R FILLER_270_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_270_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1023 ();
 FILLER_ASAP7_75t_R FILLER_270_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1353 ();
 DECAPx4_ASAP7_75t_R FILLER_270_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_270_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_271_2 ();
 DECAPx10_ASAP7_75t_R FILLER_271_24 ();
 DECAPx10_ASAP7_75t_R FILLER_271_46 ();
 DECAPx10_ASAP7_75t_R FILLER_271_68 ();
 DECAPx10_ASAP7_75t_R FILLER_271_90 ();
 DECAPx10_ASAP7_75t_R FILLER_271_112 ();
 DECAPx10_ASAP7_75t_R FILLER_271_134 ();
 DECAPx10_ASAP7_75t_R FILLER_271_156 ();
 DECAPx10_ASAP7_75t_R FILLER_271_178 ();
 DECAPx10_ASAP7_75t_R FILLER_271_200 ();
 DECAPx10_ASAP7_75t_R FILLER_271_222 ();
 DECAPx10_ASAP7_75t_R FILLER_271_244 ();
 DECAPx10_ASAP7_75t_R FILLER_271_266 ();
 DECAPx10_ASAP7_75t_R FILLER_271_288 ();
 DECAPx10_ASAP7_75t_R FILLER_271_310 ();
 DECAPx10_ASAP7_75t_R FILLER_271_332 ();
 DECAPx10_ASAP7_75t_R FILLER_271_354 ();
 DECAPx10_ASAP7_75t_R FILLER_271_376 ();
 DECAPx10_ASAP7_75t_R FILLER_271_398 ();
 DECAPx10_ASAP7_75t_R FILLER_271_420 ();
 DECAPx10_ASAP7_75t_R FILLER_271_442 ();
 DECAPx10_ASAP7_75t_R FILLER_271_464 ();
 DECAPx10_ASAP7_75t_R FILLER_271_486 ();
 DECAPx10_ASAP7_75t_R FILLER_271_508 ();
 DECAPx10_ASAP7_75t_R FILLER_271_530 ();
 DECAPx10_ASAP7_75t_R FILLER_271_552 ();
 DECAPx10_ASAP7_75t_R FILLER_271_574 ();
 DECAPx10_ASAP7_75t_R FILLER_271_596 ();
 DECAPx10_ASAP7_75t_R FILLER_271_618 ();
 DECAPx10_ASAP7_75t_R FILLER_271_640 ();
 DECAPx10_ASAP7_75t_R FILLER_271_662 ();
 DECAPx10_ASAP7_75t_R FILLER_271_684 ();
 DECAPx10_ASAP7_75t_R FILLER_271_706 ();
 DECAPx10_ASAP7_75t_R FILLER_271_728 ();
 DECAPx10_ASAP7_75t_R FILLER_271_750 ();
 DECAPx10_ASAP7_75t_R FILLER_271_772 ();
 DECAPx6_ASAP7_75t_R FILLER_271_794 ();
 DECAPx4_ASAP7_75t_R FILLER_271_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_844 ();
 DECAPx1_ASAP7_75t_R FILLER_271_848 ();
 DECAPx6_ASAP7_75t_R FILLER_271_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_909 ();
 DECAPx4_ASAP7_75t_R FILLER_271_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_942 ();
 DECAPx2_ASAP7_75t_R FILLER_271_949 ();
 FILLER_ASAP7_75t_R FILLER_271_955 ();
 DECAPx2_ASAP7_75t_R FILLER_271_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_975 ();
 DECAPx4_ASAP7_75t_R FILLER_271_979 ();
 DECAPx4_ASAP7_75t_R FILLER_271_1015 ();
 FILLER_ASAP7_75t_R FILLER_271_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_271_1385 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_272_2 ();
 DECAPx10_ASAP7_75t_R FILLER_272_24 ();
 DECAPx10_ASAP7_75t_R FILLER_272_46 ();
 DECAPx10_ASAP7_75t_R FILLER_272_68 ();
 DECAPx10_ASAP7_75t_R FILLER_272_90 ();
 DECAPx10_ASAP7_75t_R FILLER_272_112 ();
 DECAPx10_ASAP7_75t_R FILLER_272_134 ();
 DECAPx10_ASAP7_75t_R FILLER_272_156 ();
 DECAPx10_ASAP7_75t_R FILLER_272_178 ();
 DECAPx10_ASAP7_75t_R FILLER_272_200 ();
 DECAPx10_ASAP7_75t_R FILLER_272_222 ();
 DECAPx10_ASAP7_75t_R FILLER_272_244 ();
 DECAPx10_ASAP7_75t_R FILLER_272_266 ();
 DECAPx10_ASAP7_75t_R FILLER_272_288 ();
 DECAPx10_ASAP7_75t_R FILLER_272_310 ();
 DECAPx10_ASAP7_75t_R FILLER_272_332 ();
 DECAPx10_ASAP7_75t_R FILLER_272_354 ();
 DECAPx10_ASAP7_75t_R FILLER_272_376 ();
 DECAPx10_ASAP7_75t_R FILLER_272_398 ();
 DECAPx10_ASAP7_75t_R FILLER_272_420 ();
 DECAPx6_ASAP7_75t_R FILLER_272_442 ();
 DECAPx2_ASAP7_75t_R FILLER_272_456 ();
 DECAPx10_ASAP7_75t_R FILLER_272_464 ();
 DECAPx10_ASAP7_75t_R FILLER_272_486 ();
 DECAPx10_ASAP7_75t_R FILLER_272_508 ();
 DECAPx10_ASAP7_75t_R FILLER_272_530 ();
 DECAPx10_ASAP7_75t_R FILLER_272_552 ();
 DECAPx10_ASAP7_75t_R FILLER_272_574 ();
 DECAPx10_ASAP7_75t_R FILLER_272_596 ();
 DECAPx10_ASAP7_75t_R FILLER_272_618 ();
 DECAPx10_ASAP7_75t_R FILLER_272_640 ();
 DECAPx10_ASAP7_75t_R FILLER_272_662 ();
 DECAPx10_ASAP7_75t_R FILLER_272_684 ();
 DECAPx10_ASAP7_75t_R FILLER_272_706 ();
 DECAPx10_ASAP7_75t_R FILLER_272_728 ();
 DECAPx10_ASAP7_75t_R FILLER_272_750 ();
 DECAPx10_ASAP7_75t_R FILLER_272_772 ();
 DECAPx10_ASAP7_75t_R FILLER_272_794 ();
 FILLER_ASAP7_75t_R FILLER_272_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_818 ();
 FILLER_ASAP7_75t_R FILLER_272_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_830 ();
 DECAPx6_ASAP7_75t_R FILLER_272_857 ();
 DECAPx2_ASAP7_75t_R FILLER_272_884 ();
 FILLER_ASAP7_75t_R FILLER_272_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_903 ();
 DECAPx1_ASAP7_75t_R FILLER_272_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_920 ();
 FILLER_ASAP7_75t_R FILLER_272_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_961 ();
 DECAPx2_ASAP7_75t_R FILLER_272_1014 ();
 FILLER_ASAP7_75t_R FILLER_272_1020 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_272_1378 ();
 FILLER_ASAP7_75t_R FILLER_272_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_272_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_273_2 ();
 DECAPx10_ASAP7_75t_R FILLER_273_24 ();
 DECAPx10_ASAP7_75t_R FILLER_273_46 ();
 DECAPx10_ASAP7_75t_R FILLER_273_68 ();
 DECAPx10_ASAP7_75t_R FILLER_273_90 ();
 DECAPx10_ASAP7_75t_R FILLER_273_112 ();
 DECAPx10_ASAP7_75t_R FILLER_273_134 ();
 DECAPx10_ASAP7_75t_R FILLER_273_156 ();
 DECAPx10_ASAP7_75t_R FILLER_273_178 ();
 DECAPx10_ASAP7_75t_R FILLER_273_200 ();
 DECAPx10_ASAP7_75t_R FILLER_273_222 ();
 DECAPx10_ASAP7_75t_R FILLER_273_244 ();
 DECAPx10_ASAP7_75t_R FILLER_273_266 ();
 DECAPx10_ASAP7_75t_R FILLER_273_288 ();
 DECAPx10_ASAP7_75t_R FILLER_273_310 ();
 DECAPx10_ASAP7_75t_R FILLER_273_332 ();
 DECAPx10_ASAP7_75t_R FILLER_273_354 ();
 DECAPx10_ASAP7_75t_R FILLER_273_376 ();
 DECAPx10_ASAP7_75t_R FILLER_273_398 ();
 DECAPx10_ASAP7_75t_R FILLER_273_420 ();
 DECAPx10_ASAP7_75t_R FILLER_273_442 ();
 DECAPx10_ASAP7_75t_R FILLER_273_464 ();
 DECAPx10_ASAP7_75t_R FILLER_273_486 ();
 DECAPx10_ASAP7_75t_R FILLER_273_508 ();
 DECAPx10_ASAP7_75t_R FILLER_273_530 ();
 DECAPx10_ASAP7_75t_R FILLER_273_552 ();
 DECAPx10_ASAP7_75t_R FILLER_273_574 ();
 DECAPx10_ASAP7_75t_R FILLER_273_596 ();
 DECAPx10_ASAP7_75t_R FILLER_273_618 ();
 DECAPx10_ASAP7_75t_R FILLER_273_640 ();
 DECAPx10_ASAP7_75t_R FILLER_273_662 ();
 DECAPx10_ASAP7_75t_R FILLER_273_684 ();
 DECAPx10_ASAP7_75t_R FILLER_273_706 ();
 DECAPx10_ASAP7_75t_R FILLER_273_728 ();
 DECAPx10_ASAP7_75t_R FILLER_273_750 ();
 DECAPx10_ASAP7_75t_R FILLER_273_772 ();
 DECAPx10_ASAP7_75t_R FILLER_273_794 ();
 DECAPx4_ASAP7_75t_R FILLER_273_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_826 ();
 DECAPx2_ASAP7_75t_R FILLER_273_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_836 ();
 DECAPx2_ASAP7_75t_R FILLER_273_847 ();
 FILLER_ASAP7_75t_R FILLER_273_853 ();
 DECAPx2_ASAP7_75t_R FILLER_273_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_887 ();
 DECAPx1_ASAP7_75t_R FILLER_273_904 ();
 DECAPx1_ASAP7_75t_R FILLER_273_920 ();
 FILLER_ASAP7_75t_R FILLER_273_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_940 ();
 DECAPx10_ASAP7_75t_R FILLER_273_962 ();
 DECAPx6_ASAP7_75t_R FILLER_273_984 ();
 DECAPx1_ASAP7_75t_R FILLER_273_998 ();
 DECAPx4_ASAP7_75t_R FILLER_273_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1352 ();
 DECAPx6_ASAP7_75t_R FILLER_273_1374 ();
 DECAPx1_ASAP7_75t_R FILLER_273_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_274_2 ();
 DECAPx10_ASAP7_75t_R FILLER_274_24 ();
 DECAPx10_ASAP7_75t_R FILLER_274_46 ();
 DECAPx10_ASAP7_75t_R FILLER_274_68 ();
 DECAPx10_ASAP7_75t_R FILLER_274_90 ();
 DECAPx10_ASAP7_75t_R FILLER_274_112 ();
 DECAPx10_ASAP7_75t_R FILLER_274_134 ();
 DECAPx10_ASAP7_75t_R FILLER_274_156 ();
 DECAPx10_ASAP7_75t_R FILLER_274_178 ();
 DECAPx10_ASAP7_75t_R FILLER_274_200 ();
 DECAPx10_ASAP7_75t_R FILLER_274_222 ();
 DECAPx10_ASAP7_75t_R FILLER_274_244 ();
 DECAPx10_ASAP7_75t_R FILLER_274_266 ();
 DECAPx10_ASAP7_75t_R FILLER_274_288 ();
 DECAPx10_ASAP7_75t_R FILLER_274_310 ();
 DECAPx10_ASAP7_75t_R FILLER_274_332 ();
 DECAPx10_ASAP7_75t_R FILLER_274_354 ();
 DECAPx10_ASAP7_75t_R FILLER_274_376 ();
 DECAPx10_ASAP7_75t_R FILLER_274_398 ();
 DECAPx10_ASAP7_75t_R FILLER_274_420 ();
 DECAPx6_ASAP7_75t_R FILLER_274_442 ();
 DECAPx2_ASAP7_75t_R FILLER_274_456 ();
 DECAPx10_ASAP7_75t_R FILLER_274_464 ();
 DECAPx10_ASAP7_75t_R FILLER_274_486 ();
 DECAPx10_ASAP7_75t_R FILLER_274_508 ();
 DECAPx10_ASAP7_75t_R FILLER_274_530 ();
 DECAPx10_ASAP7_75t_R FILLER_274_552 ();
 DECAPx10_ASAP7_75t_R FILLER_274_574 ();
 DECAPx10_ASAP7_75t_R FILLER_274_596 ();
 DECAPx10_ASAP7_75t_R FILLER_274_618 ();
 DECAPx10_ASAP7_75t_R FILLER_274_640 ();
 DECAPx10_ASAP7_75t_R FILLER_274_662 ();
 DECAPx10_ASAP7_75t_R FILLER_274_684 ();
 DECAPx10_ASAP7_75t_R FILLER_274_706 ();
 DECAPx10_ASAP7_75t_R FILLER_274_728 ();
 DECAPx10_ASAP7_75t_R FILLER_274_750 ();
 DECAPx10_ASAP7_75t_R FILLER_274_772 ();
 DECAPx6_ASAP7_75t_R FILLER_274_794 ();
 DECAPx1_ASAP7_75t_R FILLER_274_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_812 ();
 FILLER_ASAP7_75t_R FILLER_274_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_868 ();
 DECAPx10_ASAP7_75t_R FILLER_274_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_894 ();
 DECAPx4_ASAP7_75t_R FILLER_274_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_929 ();
 DECAPx4_ASAP7_75t_R FILLER_274_933 ();
 FILLER_ASAP7_75t_R FILLER_274_943 ();
 DECAPx2_ASAP7_75t_R FILLER_274_948 ();
 DECAPx2_ASAP7_75t_R FILLER_274_960 ();
 FILLER_ASAP7_75t_R FILLER_274_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_968 ();
 DECAPx1_ASAP7_75t_R FILLER_274_972 ();
 DECAPx10_ASAP7_75t_R FILLER_274_986 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1008 ();
 FILLER_ASAP7_75t_R FILLER_274_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_274_1370 ();
 FILLER_ASAP7_75t_R FILLER_274_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_274_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_275_2 ();
 DECAPx10_ASAP7_75t_R FILLER_275_24 ();
 DECAPx10_ASAP7_75t_R FILLER_275_46 ();
 DECAPx10_ASAP7_75t_R FILLER_275_68 ();
 DECAPx10_ASAP7_75t_R FILLER_275_90 ();
 DECAPx10_ASAP7_75t_R FILLER_275_112 ();
 DECAPx10_ASAP7_75t_R FILLER_275_134 ();
 DECAPx10_ASAP7_75t_R FILLER_275_156 ();
 DECAPx10_ASAP7_75t_R FILLER_275_178 ();
 DECAPx10_ASAP7_75t_R FILLER_275_200 ();
 DECAPx10_ASAP7_75t_R FILLER_275_222 ();
 DECAPx10_ASAP7_75t_R FILLER_275_244 ();
 DECAPx10_ASAP7_75t_R FILLER_275_266 ();
 DECAPx10_ASAP7_75t_R FILLER_275_288 ();
 DECAPx10_ASAP7_75t_R FILLER_275_310 ();
 DECAPx10_ASAP7_75t_R FILLER_275_332 ();
 DECAPx10_ASAP7_75t_R FILLER_275_354 ();
 DECAPx10_ASAP7_75t_R FILLER_275_376 ();
 DECAPx10_ASAP7_75t_R FILLER_275_398 ();
 DECAPx10_ASAP7_75t_R FILLER_275_420 ();
 DECAPx10_ASAP7_75t_R FILLER_275_442 ();
 DECAPx10_ASAP7_75t_R FILLER_275_464 ();
 DECAPx10_ASAP7_75t_R FILLER_275_486 ();
 DECAPx10_ASAP7_75t_R FILLER_275_508 ();
 DECAPx10_ASAP7_75t_R FILLER_275_530 ();
 DECAPx10_ASAP7_75t_R FILLER_275_552 ();
 DECAPx10_ASAP7_75t_R FILLER_275_574 ();
 DECAPx10_ASAP7_75t_R FILLER_275_596 ();
 DECAPx10_ASAP7_75t_R FILLER_275_618 ();
 DECAPx4_ASAP7_75t_R FILLER_275_640 ();
 DECAPx2_ASAP7_75t_R FILLER_275_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_662 ();
 DECAPx10_ASAP7_75t_R FILLER_275_681 ();
 DECAPx10_ASAP7_75t_R FILLER_275_703 ();
 DECAPx10_ASAP7_75t_R FILLER_275_725 ();
 DECAPx10_ASAP7_75t_R FILLER_275_747 ();
 DECAPx10_ASAP7_75t_R FILLER_275_769 ();
 DECAPx10_ASAP7_75t_R FILLER_275_791 ();
 DECAPx10_ASAP7_75t_R FILLER_275_813 ();
 DECAPx10_ASAP7_75t_R FILLER_275_835 ();
 DECAPx2_ASAP7_75t_R FILLER_275_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_866 ();
 DECAPx6_ASAP7_75t_R FILLER_275_893 ();
 DECAPx2_ASAP7_75t_R FILLER_275_907 ();
 DECAPx2_ASAP7_75t_R FILLER_275_916 ();
 FILLER_ASAP7_75t_R FILLER_275_922 ();
 DECAPx2_ASAP7_75t_R FILLER_275_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_935 ();
 DECAPx6_ASAP7_75t_R FILLER_275_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_953 ();
 DECAPx10_ASAP7_75t_R FILLER_275_980 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1354 ();
 DECAPx6_ASAP7_75t_R FILLER_275_1376 ();
 FILLER_ASAP7_75t_R FILLER_275_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_276_2 ();
 DECAPx10_ASAP7_75t_R FILLER_276_24 ();
 DECAPx10_ASAP7_75t_R FILLER_276_46 ();
 DECAPx10_ASAP7_75t_R FILLER_276_68 ();
 DECAPx10_ASAP7_75t_R FILLER_276_90 ();
 DECAPx10_ASAP7_75t_R FILLER_276_112 ();
 DECAPx10_ASAP7_75t_R FILLER_276_134 ();
 DECAPx10_ASAP7_75t_R FILLER_276_156 ();
 DECAPx10_ASAP7_75t_R FILLER_276_178 ();
 DECAPx10_ASAP7_75t_R FILLER_276_200 ();
 DECAPx10_ASAP7_75t_R FILLER_276_222 ();
 DECAPx10_ASAP7_75t_R FILLER_276_244 ();
 DECAPx10_ASAP7_75t_R FILLER_276_266 ();
 DECAPx10_ASAP7_75t_R FILLER_276_288 ();
 DECAPx10_ASAP7_75t_R FILLER_276_310 ();
 DECAPx10_ASAP7_75t_R FILLER_276_332 ();
 DECAPx10_ASAP7_75t_R FILLER_276_354 ();
 DECAPx10_ASAP7_75t_R FILLER_276_376 ();
 DECAPx10_ASAP7_75t_R FILLER_276_398 ();
 DECAPx10_ASAP7_75t_R FILLER_276_420 ();
 DECAPx6_ASAP7_75t_R FILLER_276_442 ();
 DECAPx2_ASAP7_75t_R FILLER_276_456 ();
 DECAPx10_ASAP7_75t_R FILLER_276_464 ();
 DECAPx10_ASAP7_75t_R FILLER_276_486 ();
 DECAPx10_ASAP7_75t_R FILLER_276_508 ();
 DECAPx10_ASAP7_75t_R FILLER_276_530 ();
 DECAPx10_ASAP7_75t_R FILLER_276_552 ();
 DECAPx10_ASAP7_75t_R FILLER_276_574 ();
 DECAPx10_ASAP7_75t_R FILLER_276_596 ();
 DECAPx10_ASAP7_75t_R FILLER_276_618 ();
 DECAPx2_ASAP7_75t_R FILLER_276_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_646 ();
 DECAPx1_ASAP7_75t_R FILLER_276_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_703 ();
 DECAPx4_ASAP7_75t_R FILLER_276_710 ();
 DECAPx6_ASAP7_75t_R FILLER_276_726 ();
 DECAPx1_ASAP7_75t_R FILLER_276_740 ();
 DECAPx2_ASAP7_75t_R FILLER_276_750 ();
 FILLER_ASAP7_75t_R FILLER_276_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_758 ();
 DECAPx2_ASAP7_75t_R FILLER_276_765 ();
 DECAPx10_ASAP7_75t_R FILLER_276_777 ();
 DECAPx10_ASAP7_75t_R FILLER_276_799 ();
 DECAPx10_ASAP7_75t_R FILLER_276_821 ();
 DECAPx10_ASAP7_75t_R FILLER_276_843 ();
 DECAPx2_ASAP7_75t_R FILLER_276_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_871 ();
 DECAPx10_ASAP7_75t_R FILLER_276_950 ();
 DECAPx10_ASAP7_75t_R FILLER_276_972 ();
 DECAPx10_ASAP7_75t_R FILLER_276_994 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_276_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_276_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_276_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_277_2 ();
 DECAPx10_ASAP7_75t_R FILLER_277_24 ();
 DECAPx10_ASAP7_75t_R FILLER_277_46 ();
 DECAPx10_ASAP7_75t_R FILLER_277_68 ();
 DECAPx10_ASAP7_75t_R FILLER_277_90 ();
 DECAPx10_ASAP7_75t_R FILLER_277_112 ();
 DECAPx10_ASAP7_75t_R FILLER_277_134 ();
 DECAPx10_ASAP7_75t_R FILLER_277_156 ();
 DECAPx10_ASAP7_75t_R FILLER_277_178 ();
 DECAPx10_ASAP7_75t_R FILLER_277_200 ();
 DECAPx10_ASAP7_75t_R FILLER_277_222 ();
 DECAPx10_ASAP7_75t_R FILLER_277_244 ();
 DECAPx10_ASAP7_75t_R FILLER_277_266 ();
 DECAPx10_ASAP7_75t_R FILLER_277_288 ();
 DECAPx10_ASAP7_75t_R FILLER_277_310 ();
 DECAPx10_ASAP7_75t_R FILLER_277_332 ();
 DECAPx10_ASAP7_75t_R FILLER_277_354 ();
 DECAPx10_ASAP7_75t_R FILLER_277_376 ();
 DECAPx10_ASAP7_75t_R FILLER_277_398 ();
 DECAPx10_ASAP7_75t_R FILLER_277_420 ();
 DECAPx6_ASAP7_75t_R FILLER_277_442 ();
 DECAPx2_ASAP7_75t_R FILLER_277_456 ();
 DECAPx10_ASAP7_75t_R FILLER_277_464 ();
 DECAPx10_ASAP7_75t_R FILLER_277_486 ();
 DECAPx10_ASAP7_75t_R FILLER_277_508 ();
 DECAPx10_ASAP7_75t_R FILLER_277_530 ();
 DECAPx10_ASAP7_75t_R FILLER_277_552 ();
 DECAPx10_ASAP7_75t_R FILLER_277_574 ();
 DECAPx10_ASAP7_75t_R FILLER_277_596 ();
 DECAPx10_ASAP7_75t_R FILLER_277_618 ();
 FILLER_ASAP7_75t_R FILLER_277_640 ();
 DECAPx1_ASAP7_75t_R FILLER_277_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_662 ();
 DECAPx4_ASAP7_75t_R FILLER_277_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_727 ();
 DECAPx2_ASAP7_75t_R FILLER_277_734 ();
 FILLER_ASAP7_75t_R FILLER_277_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_742 ();
 DECAPx2_ASAP7_75t_R FILLER_277_749 ();
 DECAPx10_ASAP7_75t_R FILLER_277_785 ();
 DECAPx10_ASAP7_75t_R FILLER_277_807 ();
 DECAPx10_ASAP7_75t_R FILLER_277_829 ();
 DECAPx10_ASAP7_75t_R FILLER_277_851 ();
 DECAPx2_ASAP7_75t_R FILLER_277_873 ();
 FILLER_ASAP7_75t_R FILLER_277_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_885 ();
 DECAPx10_ASAP7_75t_R FILLER_277_889 ();
 DECAPx4_ASAP7_75t_R FILLER_277_911 ();
 FILLER_ASAP7_75t_R FILLER_277_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_923 ();
 DECAPx10_ASAP7_75t_R FILLER_277_952 ();
 DECAPx10_ASAP7_75t_R FILLER_277_974 ();
 DECAPx10_ASAP7_75t_R FILLER_277_996 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_277_1370 ();
 FILLER_ASAP7_75t_R FILLER_277_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_277_1388 ();
endmodule
