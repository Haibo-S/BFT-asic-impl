module t_switch (ce,
    clk,
    done,
    rst,
    l_i,
    l_o,
    r_i,
    r_o,
    u0_i,
    u0_o);
 input ce;
 input clk;
 output done;
 input rst;
 input [36:0] l_i;
 output [36:0] l_o;
 input [36:0] r_i;
 output [36:0] r_o;
 input [36:0] u0_i;
 output [36:0] u0_o;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire _486_;
 wire _487_;
 wire _488_;
 wire _489_;
 wire _490_;
 wire _491_;
 wire _492_;
 wire _493_;
 wire clknet_0_clk;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net219;
 wire net220;
 wire net221;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 BUFx12f_ASAP7_75t_R _495_ (.A(net102),
    .Y(_218_));
 BUFx6f_ASAP7_75t_R _496_ (.A(_218_),
    .Y(_219_));
 OR3x1_ASAP7_75t_R _497_ (.A(_219_),
    .B(net65),
    .C(net29),
    .Y(_220_));
 INVx1_ASAP7_75t_R _498_ (.A(_220_),
    .Y(_000_));
 INVx1_ASAP7_75t_R _499_ (.A(_001_),
    .Y(net218));
 INVx1_ASAP7_75t_R _500_ (.A(_002_),
    .Y(net217));
 INVx1_ASAP7_75t_R _501_ (.A(_003_),
    .Y(net216));
 INVx1_ASAP7_75t_R _502_ (.A(_004_),
    .Y(net215));
 INVx1_ASAP7_75t_R _503_ (.A(_005_),
    .Y(net214));
 INVx1_ASAP7_75t_R _504_ (.A(_006_),
    .Y(net213));
 INVx1_ASAP7_75t_R _505_ (.A(_007_),
    .Y(net212));
 INVx1_ASAP7_75t_R _506_ (.A(_008_),
    .Y(net211));
 INVx1_ASAP7_75t_R _507_ (.A(_009_),
    .Y(net210));
 INVx1_ASAP7_75t_R _508_ (.A(_010_),
    .Y(net209));
 INVx1_ASAP7_75t_R _509_ (.A(_011_),
    .Y(net208));
 INVx1_ASAP7_75t_R _510_ (.A(_012_),
    .Y(net207));
 INVx1_ASAP7_75t_R _511_ (.A(_013_),
    .Y(net206));
 INVx1_ASAP7_75t_R _512_ (.A(_014_),
    .Y(net205));
 INVx1_ASAP7_75t_R _513_ (.A(_015_),
    .Y(net204));
 INVx1_ASAP7_75t_R _514_ (.A(_016_),
    .Y(net203));
 INVx1_ASAP7_75t_R _515_ (.A(_017_),
    .Y(net202));
 INVx1_ASAP7_75t_R _516_ (.A(_018_),
    .Y(net201));
 INVx1_ASAP7_75t_R _517_ (.A(_019_),
    .Y(net200));
 INVx1_ASAP7_75t_R _518_ (.A(_020_),
    .Y(net199));
 INVx1_ASAP7_75t_R _519_ (.A(_021_),
    .Y(net198));
 INVx1_ASAP7_75t_R _520_ (.A(_022_),
    .Y(net197));
 INVx1_ASAP7_75t_R _521_ (.A(_023_),
    .Y(net196));
 INVx1_ASAP7_75t_R _522_ (.A(_024_),
    .Y(net195));
 INVx1_ASAP7_75t_R _523_ (.A(_025_),
    .Y(net194));
 INVx1_ASAP7_75t_R _524_ (.A(_026_),
    .Y(net193));
 INVx1_ASAP7_75t_R _525_ (.A(_027_),
    .Y(net192));
 INVx1_ASAP7_75t_R _526_ (.A(_028_),
    .Y(net191));
 INVx1_ASAP7_75t_R _527_ (.A(_029_),
    .Y(net190));
 INVx1_ASAP7_75t_R _528_ (.A(_030_),
    .Y(net189));
 INVx1_ASAP7_75t_R _529_ (.A(_031_),
    .Y(net188));
 INVx1_ASAP7_75t_R _530_ (.A(_032_),
    .Y(net187));
 INVx1_ASAP7_75t_R _531_ (.A(_033_),
    .Y(net186));
 INVx1_ASAP7_75t_R _532_ (.A(_034_),
    .Y(net185));
 INVx1_ASAP7_75t_R _533_ (.A(_035_),
    .Y(net184));
 INVx1_ASAP7_75t_R _534_ (.A(_036_),
    .Y(net183));
 INVx1_ASAP7_75t_R _535_ (.A(_037_),
    .Y(net182));
 INVx1_ASAP7_75t_R _536_ (.A(_038_),
    .Y(net181));
 INVx1_ASAP7_75t_R _537_ (.A(_039_),
    .Y(net180));
 INVx1_ASAP7_75t_R _538_ (.A(_040_),
    .Y(net179));
 INVx1_ASAP7_75t_R _539_ (.A(_041_),
    .Y(net178));
 INVx1_ASAP7_75t_R _540_ (.A(_042_),
    .Y(net177));
 INVx1_ASAP7_75t_R _541_ (.A(_043_),
    .Y(net176));
 INVx1_ASAP7_75t_R _542_ (.A(_044_),
    .Y(net175));
 INVx1_ASAP7_75t_R _543_ (.A(_045_),
    .Y(net174));
 INVx1_ASAP7_75t_R _544_ (.A(_046_),
    .Y(net173));
 INVx1_ASAP7_75t_R _545_ (.A(_047_),
    .Y(net172));
 INVx1_ASAP7_75t_R _546_ (.A(_048_),
    .Y(net171));
 INVx1_ASAP7_75t_R _547_ (.A(_049_),
    .Y(net170));
 INVx1_ASAP7_75t_R _548_ (.A(_050_),
    .Y(net169));
 INVx1_ASAP7_75t_R _549_ (.A(_051_),
    .Y(net168));
 INVx1_ASAP7_75t_R _550_ (.A(_052_),
    .Y(net167));
 INVx1_ASAP7_75t_R _551_ (.A(_053_),
    .Y(net166));
 INVx1_ASAP7_75t_R _552_ (.A(_054_),
    .Y(net165));
 INVx1_ASAP7_75t_R _553_ (.A(_055_),
    .Y(net164));
 INVx1_ASAP7_75t_R _554_ (.A(_056_),
    .Y(net163));
 INVx1_ASAP7_75t_R _555_ (.A(_057_),
    .Y(net162));
 INVx1_ASAP7_75t_R _556_ (.A(_058_),
    .Y(net161));
 INVx1_ASAP7_75t_R _557_ (.A(_059_),
    .Y(net160));
 INVx1_ASAP7_75t_R _558_ (.A(_060_),
    .Y(net159));
 INVx1_ASAP7_75t_R _559_ (.A(_061_),
    .Y(net158));
 INVx1_ASAP7_75t_R _560_ (.A(_062_),
    .Y(net157));
 INVx1_ASAP7_75t_R _561_ (.A(_063_),
    .Y(net156));
 INVx1_ASAP7_75t_R _562_ (.A(_064_),
    .Y(net155));
 INVx1_ASAP7_75t_R _563_ (.A(_065_),
    .Y(net154));
 INVx1_ASAP7_75t_R _564_ (.A(_066_),
    .Y(net153));
 INVx1_ASAP7_75t_R _565_ (.A(_067_),
    .Y(net152));
 INVx1_ASAP7_75t_R _566_ (.A(_068_),
    .Y(net151));
 INVx1_ASAP7_75t_R _567_ (.A(_069_),
    .Y(net150));
 INVx1_ASAP7_75t_R _568_ (.A(_070_),
    .Y(net149));
 INVx1_ASAP7_75t_R _569_ (.A(_071_),
    .Y(net148));
 INVx1_ASAP7_75t_R _570_ (.A(_072_),
    .Y(net147));
 INVx1_ASAP7_75t_R _571_ (.A(_073_),
    .Y(net146));
 INVx1_ASAP7_75t_R _572_ (.A(_074_),
    .Y(net145));
 INVx1_ASAP7_75t_R _573_ (.A(_075_),
    .Y(net144));
 INVx1_ASAP7_75t_R _574_ (.A(_076_),
    .Y(net143));
 INVx1_ASAP7_75t_R _575_ (.A(_077_),
    .Y(net142));
 INVx1_ASAP7_75t_R _576_ (.A(_078_),
    .Y(net141));
 INVx1_ASAP7_75t_R _577_ (.A(_079_),
    .Y(net140));
 INVx1_ASAP7_75t_R _578_ (.A(_080_),
    .Y(net139));
 INVx1_ASAP7_75t_R _579_ (.A(_081_),
    .Y(net138));
 INVx1_ASAP7_75t_R _580_ (.A(_082_),
    .Y(net137));
 INVx1_ASAP7_75t_R _581_ (.A(_083_),
    .Y(net136));
 INVx1_ASAP7_75t_R _582_ (.A(_084_),
    .Y(net135));
 INVx1_ASAP7_75t_R _583_ (.A(_085_),
    .Y(net134));
 INVx1_ASAP7_75t_R _584_ (.A(_086_),
    .Y(net133));
 INVx1_ASAP7_75t_R _585_ (.A(_087_),
    .Y(net132));
 INVx1_ASAP7_75t_R _586_ (.A(_088_),
    .Y(net131));
 INVx1_ASAP7_75t_R _587_ (.A(_089_),
    .Y(net130));
 INVx1_ASAP7_75t_R _588_ (.A(_090_),
    .Y(net129));
 INVx1_ASAP7_75t_R _589_ (.A(_091_),
    .Y(net128));
 INVx1_ASAP7_75t_R _590_ (.A(_092_),
    .Y(net127));
 INVx1_ASAP7_75t_R _591_ (.A(_093_),
    .Y(net126));
 INVx1_ASAP7_75t_R _592_ (.A(_094_),
    .Y(net125));
 INVx1_ASAP7_75t_R _593_ (.A(_095_),
    .Y(net124));
 INVx1_ASAP7_75t_R _594_ (.A(_096_),
    .Y(net123));
 INVx1_ASAP7_75t_R _595_ (.A(_097_),
    .Y(net122));
 INVx1_ASAP7_75t_R _596_ (.A(_098_),
    .Y(net121));
 INVx1_ASAP7_75t_R _597_ (.A(_099_),
    .Y(net120));
 INVx1_ASAP7_75t_R _598_ (.A(_100_),
    .Y(net119));
 INVx1_ASAP7_75t_R _599_ (.A(_101_),
    .Y(net118));
 INVx1_ASAP7_75t_R _600_ (.A(_102_),
    .Y(net117));
 INVx1_ASAP7_75t_R _601_ (.A(_103_),
    .Y(net116));
 INVx1_ASAP7_75t_R _602_ (.A(_104_),
    .Y(net115));
 INVx1_ASAP7_75t_R _603_ (.A(_105_),
    .Y(net114));
 INVx1_ASAP7_75t_R _604_ (.A(_106_),
    .Y(net113));
 INVx1_ASAP7_75t_R _605_ (.A(_107_),
    .Y(net112));
 INVx1_ASAP7_75t_R _606_ (.A(_108_),
    .Y(net111));
 INVx1_ASAP7_75t_R _607_ (.A(_109_),
    .Y(net110));
 INVx3_ASAP7_75t_R _608_ (.A(net73),
    .Y(_221_));
 BUFx6f_ASAP7_75t_R _609_ (.A(_221_),
    .Y(_222_));
 BUFx6f_ASAP7_75t_R _610_ (.A(_222_),
    .Y(_223_));
 INVx5_ASAP7_75t_R _611_ (.A(net99),
    .Y(_224_));
 NAND2x2_ASAP7_75t_R _612_ (.A(_218_),
    .B(_224_),
    .Y(_225_));
 BUFx6f_ASAP7_75t_R _613_ (.A(_225_),
    .Y(_226_));
 BUFx6f_ASAP7_75t_R _614_ (.A(_224_),
    .Y(_227_));
 AND3x1_ASAP7_75t_R _615_ (.A(_219_),
    .B(_227_),
    .C(net74),
    .Y(_228_));
 AO21x1_ASAP7_75t_R _616_ (.A1(net37),
    .A2(_226_),
    .B(_228_),
    .Y(_229_));
 AND2x2_ASAP7_75t_R _617_ (.A(_223_),
    .B(_229_),
    .Y(_110_));
 AND3x1_ASAP7_75t_R _618_ (.A(_219_),
    .B(_227_),
    .C(net75),
    .Y(_230_));
 AO21x1_ASAP7_75t_R _619_ (.A1(net38),
    .A2(_226_),
    .B(_230_),
    .Y(_231_));
 AND2x2_ASAP7_75t_R _620_ (.A(_223_),
    .B(_231_),
    .Y(_111_));
 AND3x1_ASAP7_75t_R _621_ (.A(_219_),
    .B(_227_),
    .C(net76),
    .Y(_232_));
 AO21x1_ASAP7_75t_R _622_ (.A1(net39),
    .A2(_226_),
    .B(_232_),
    .Y(_233_));
 AND2x2_ASAP7_75t_R _623_ (.A(_223_),
    .B(_233_),
    .Y(_112_));
 AND3x1_ASAP7_75t_R _624_ (.A(_219_),
    .B(_227_),
    .C(net77),
    .Y(_234_));
 AO21x1_ASAP7_75t_R _625_ (.A1(net40),
    .A2(_226_),
    .B(_234_),
    .Y(_235_));
 AND2x2_ASAP7_75t_R _626_ (.A(_223_),
    .B(_235_),
    .Y(_113_));
 AND3x1_ASAP7_75t_R _627_ (.A(_219_),
    .B(_227_),
    .C(net78),
    .Y(_236_));
 AO21x1_ASAP7_75t_R _628_ (.A1(net41),
    .A2(_226_),
    .B(_236_),
    .Y(_237_));
 AND2x2_ASAP7_75t_R _629_ (.A(_223_),
    .B(_237_),
    .Y(_114_));
 AND3x1_ASAP7_75t_R _630_ (.A(_219_),
    .B(_227_),
    .C(net79),
    .Y(_238_));
 AO21x1_ASAP7_75t_R _631_ (.A1(net42),
    .A2(_226_),
    .B(_238_),
    .Y(_239_));
 AND2x2_ASAP7_75t_R _632_ (.A(_223_),
    .B(_239_),
    .Y(_115_));
 AND3x1_ASAP7_75t_R _633_ (.A(_219_),
    .B(_227_),
    .C(net80),
    .Y(_240_));
 AO21x1_ASAP7_75t_R _634_ (.A1(net43),
    .A2(_226_),
    .B(_240_),
    .Y(_241_));
 AND2x2_ASAP7_75t_R _635_ (.A(_223_),
    .B(_241_),
    .Y(_116_));
 AND3x1_ASAP7_75t_R _636_ (.A(_219_),
    .B(_227_),
    .C(net81),
    .Y(_242_));
 AO21x1_ASAP7_75t_R _637_ (.A1(net44),
    .A2(_226_),
    .B(_242_),
    .Y(_243_));
 AND2x2_ASAP7_75t_R _638_ (.A(_223_),
    .B(_243_),
    .Y(_117_));
 BUFx6f_ASAP7_75t_R _639_ (.A(_218_),
    .Y(_244_));
 AND3x1_ASAP7_75t_R _640_ (.A(_244_),
    .B(_227_),
    .C(net82),
    .Y(_245_));
 AO21x1_ASAP7_75t_R _641_ (.A1(net45),
    .A2(_226_),
    .B(_245_),
    .Y(_246_));
 AND2x2_ASAP7_75t_R _642_ (.A(_223_),
    .B(_246_),
    .Y(_118_));
 BUFx6f_ASAP7_75t_R _643_ (.A(_225_),
    .Y(_247_));
 AND3x1_ASAP7_75t_R _644_ (.A(_244_),
    .B(_227_),
    .C(net83),
    .Y(_248_));
 AO21x1_ASAP7_75t_R _645_ (.A1(net46),
    .A2(_247_),
    .B(_248_),
    .Y(_249_));
 AND2x2_ASAP7_75t_R _646_ (.A(_223_),
    .B(_249_),
    .Y(_119_));
 BUFx6f_ASAP7_75t_R _647_ (.A(_222_),
    .Y(_250_));
 BUFx6f_ASAP7_75t_R _648_ (.A(_224_),
    .Y(_251_));
 AND3x1_ASAP7_75t_R _649_ (.A(_244_),
    .B(_251_),
    .C(net84),
    .Y(_252_));
 AO21x1_ASAP7_75t_R _650_ (.A1(net47),
    .A2(_247_),
    .B(_252_),
    .Y(_253_));
 AND2x2_ASAP7_75t_R _651_ (.A(_250_),
    .B(_253_),
    .Y(_120_));
 AND3x1_ASAP7_75t_R _652_ (.A(_244_),
    .B(_251_),
    .C(net85),
    .Y(_254_));
 AO21x1_ASAP7_75t_R _653_ (.A1(net48),
    .A2(_247_),
    .B(_254_),
    .Y(_255_));
 AND2x2_ASAP7_75t_R _654_ (.A(_250_),
    .B(_255_),
    .Y(_121_));
 AND3x1_ASAP7_75t_R _655_ (.A(_244_),
    .B(_251_),
    .C(net86),
    .Y(_256_));
 AO21x1_ASAP7_75t_R _656_ (.A1(net49),
    .A2(_247_),
    .B(_256_),
    .Y(_257_));
 AND2x2_ASAP7_75t_R _657_ (.A(_250_),
    .B(_257_),
    .Y(_122_));
 AND3x1_ASAP7_75t_R _658_ (.A(_244_),
    .B(_251_),
    .C(net87),
    .Y(_258_));
 AO21x1_ASAP7_75t_R _659_ (.A1(net50),
    .A2(_247_),
    .B(_258_),
    .Y(_259_));
 AND2x2_ASAP7_75t_R _660_ (.A(_250_),
    .B(_259_),
    .Y(_123_));
 AND3x1_ASAP7_75t_R _661_ (.A(_244_),
    .B(_251_),
    .C(net88),
    .Y(_260_));
 AO21x1_ASAP7_75t_R _662_ (.A1(net51),
    .A2(_247_),
    .B(_260_),
    .Y(_261_));
 AND2x2_ASAP7_75t_R _663_ (.A(_250_),
    .B(_261_),
    .Y(_124_));
 AND3x1_ASAP7_75t_R _664_ (.A(_244_),
    .B(_251_),
    .C(net89),
    .Y(_262_));
 AO21x1_ASAP7_75t_R _665_ (.A1(net52),
    .A2(_247_),
    .B(_262_),
    .Y(_263_));
 AND2x2_ASAP7_75t_R _666_ (.A(_250_),
    .B(_263_),
    .Y(_125_));
 AND3x1_ASAP7_75t_R _667_ (.A(_244_),
    .B(_251_),
    .C(net90),
    .Y(_264_));
 AO21x1_ASAP7_75t_R _668_ (.A1(net53),
    .A2(_247_),
    .B(_264_),
    .Y(_265_));
 AND2x2_ASAP7_75t_R _669_ (.A(_250_),
    .B(_265_),
    .Y(_126_));
 AND3x1_ASAP7_75t_R _670_ (.A(_244_),
    .B(_251_),
    .C(net91),
    .Y(_266_));
 AO21x1_ASAP7_75t_R _671_ (.A1(net54),
    .A2(_247_),
    .B(_266_),
    .Y(_267_));
 AND2x2_ASAP7_75t_R _672_ (.A(_250_),
    .B(_267_),
    .Y(_127_));
 BUFx6f_ASAP7_75t_R _673_ (.A(_218_),
    .Y(_268_));
 AND3x1_ASAP7_75t_R _674_ (.A(_268_),
    .B(_251_),
    .C(net92),
    .Y(_269_));
 AO21x1_ASAP7_75t_R _675_ (.A1(net55),
    .A2(_247_),
    .B(_269_),
    .Y(_270_));
 AND2x2_ASAP7_75t_R _676_ (.A(_250_),
    .B(_270_),
    .Y(_128_));
 BUFx6f_ASAP7_75t_R _677_ (.A(_225_),
    .Y(_271_));
 AND3x1_ASAP7_75t_R _678_ (.A(_268_),
    .B(_251_),
    .C(net93),
    .Y(_272_));
 AO21x1_ASAP7_75t_R _679_ (.A1(net56),
    .A2(_271_),
    .B(_272_),
    .Y(_273_));
 AND2x2_ASAP7_75t_R _680_ (.A(_250_),
    .B(_273_),
    .Y(_129_));
 BUFx6f_ASAP7_75t_R _681_ (.A(_222_),
    .Y(_274_));
 BUFx6f_ASAP7_75t_R _682_ (.A(_224_),
    .Y(_275_));
 AND3x1_ASAP7_75t_R _683_ (.A(_268_),
    .B(_275_),
    .C(net94),
    .Y(_276_));
 AO21x1_ASAP7_75t_R _684_ (.A1(net57),
    .A2(_271_),
    .B(_276_),
    .Y(_277_));
 AND2x2_ASAP7_75t_R _685_ (.A(_274_),
    .B(_277_),
    .Y(_130_));
 AND3x1_ASAP7_75t_R _686_ (.A(_268_),
    .B(_275_),
    .C(net95),
    .Y(_278_));
 AO21x1_ASAP7_75t_R _687_ (.A1(net58),
    .A2(_271_),
    .B(_278_),
    .Y(_279_));
 AND2x2_ASAP7_75t_R _688_ (.A(_274_),
    .B(_279_),
    .Y(_131_));
 AND3x1_ASAP7_75t_R _689_ (.A(_268_),
    .B(_275_),
    .C(net96),
    .Y(_280_));
 AO21x1_ASAP7_75t_R _690_ (.A1(net59),
    .A2(_271_),
    .B(_280_),
    .Y(_281_));
 AND2x2_ASAP7_75t_R _691_ (.A(_274_),
    .B(_281_),
    .Y(_132_));
 AND3x1_ASAP7_75t_R _692_ (.A(_268_),
    .B(_275_),
    .C(net97),
    .Y(_282_));
 AO21x1_ASAP7_75t_R _693_ (.A1(net60),
    .A2(_271_),
    .B(_282_),
    .Y(_283_));
 AND2x2_ASAP7_75t_R _694_ (.A(_274_),
    .B(_283_),
    .Y(_133_));
 AND3x1_ASAP7_75t_R _695_ (.A(_268_),
    .B(_275_),
    .C(net98),
    .Y(_284_));
 AO21x1_ASAP7_75t_R _696_ (.A1(net61),
    .A2(_271_),
    .B(_284_),
    .Y(_285_));
 AND2x2_ASAP7_75t_R _697_ (.A(_274_),
    .B(_285_),
    .Y(_134_));
 BUFx6f_ASAP7_75t_R _698_ (.A(_221_),
    .Y(_286_));
 BUFx6f_ASAP7_75t_R _699_ (.A(_286_),
    .Y(_287_));
 AND3x1_ASAP7_75t_R _700_ (.A(net62),
    .B(_287_),
    .C(_226_),
    .Y(_135_));
 AND3x1_ASAP7_75t_R _701_ (.A(_268_),
    .B(_275_),
    .C(net100),
    .Y(_288_));
 AO21x1_ASAP7_75t_R _702_ (.A1(net63),
    .A2(_271_),
    .B(_288_),
    .Y(_289_));
 AND2x2_ASAP7_75t_R _703_ (.A(_274_),
    .B(_289_),
    .Y(_136_));
 AND3x1_ASAP7_75t_R _704_ (.A(_268_),
    .B(_275_),
    .C(net101),
    .Y(_290_));
 AO21x1_ASAP7_75t_R _705_ (.A1(net64),
    .A2(_271_),
    .B(_290_),
    .Y(_291_));
 AND2x2_ASAP7_75t_R _706_ (.A(_274_),
    .B(_291_),
    .Y(_137_));
 OR2x6_ASAP7_75t_R _707_ (.A(net64),
    .B(net63),
    .Y(_292_));
 OAI21x1_ASAP7_75t_R _708_ (.A1(net28),
    .A2(net27),
    .B(net29),
    .Y(_293_));
 INVx1_ASAP7_75t_R _709_ (.A(net65),
    .Y(_294_));
 AO21x1_ASAP7_75t_R _710_ (.A1(_292_),
    .A2(_293_),
    .B(_294_),
    .Y(_295_));
 BUFx6f_ASAP7_75t_R _711_ (.A(net99),
    .Y(_296_));
 INVx2_ASAP7_75t_R _712_ (.A(net102),
    .Y(_297_));
 AO21x1_ASAP7_75t_R _713_ (.A1(_296_),
    .A2(_294_),
    .B(_297_),
    .Y(_298_));
 AOI21x1_ASAP7_75t_R _714_ (.A1(_295_),
    .A2(_298_),
    .B(net73),
    .Y(_138_));
 AND3x1_ASAP7_75t_R _715_ (.A(_268_),
    .B(_275_),
    .C(net103),
    .Y(_299_));
 AO21x1_ASAP7_75t_R _716_ (.A1(net66),
    .A2(_271_),
    .B(_299_),
    .Y(_300_));
 AND2x2_ASAP7_75t_R _717_ (.A(_274_),
    .B(_300_),
    .Y(_139_));
 BUFx6f_ASAP7_75t_R _718_ (.A(_218_),
    .Y(_301_));
 AND3x1_ASAP7_75t_R _719_ (.A(_301_),
    .B(_275_),
    .C(net104),
    .Y(_302_));
 AO21x1_ASAP7_75t_R _720_ (.A1(net67),
    .A2(_271_),
    .B(_302_),
    .Y(_303_));
 AND2x2_ASAP7_75t_R _721_ (.A(_274_),
    .B(_303_),
    .Y(_140_));
 AND3x1_ASAP7_75t_R _722_ (.A(_301_),
    .B(_275_),
    .C(net105),
    .Y(_304_));
 AO21x1_ASAP7_75t_R _723_ (.A1(net68),
    .A2(_225_),
    .B(_304_),
    .Y(_305_));
 AND2x2_ASAP7_75t_R _724_ (.A(_274_),
    .B(_305_),
    .Y(_141_));
 BUFx6f_ASAP7_75t_R _725_ (.A(_222_),
    .Y(_306_));
 AND3x1_ASAP7_75t_R _726_ (.A(_301_),
    .B(_224_),
    .C(net106),
    .Y(_307_));
 AO21x1_ASAP7_75t_R _727_ (.A1(net69),
    .A2(_225_),
    .B(_307_),
    .Y(_308_));
 AND2x2_ASAP7_75t_R _728_ (.A(_306_),
    .B(_308_),
    .Y(_142_));
 AND3x1_ASAP7_75t_R _729_ (.A(_301_),
    .B(_224_),
    .C(net107),
    .Y(_309_));
 AO21x1_ASAP7_75t_R _730_ (.A1(net70),
    .A2(_225_),
    .B(_309_),
    .Y(_310_));
 AND2x2_ASAP7_75t_R _731_ (.A(_306_),
    .B(_310_),
    .Y(_143_));
 AND3x1_ASAP7_75t_R _732_ (.A(_301_),
    .B(_224_),
    .C(net108),
    .Y(_311_));
 AO21x1_ASAP7_75t_R _733_ (.A1(net71),
    .A2(_225_),
    .B(_311_),
    .Y(_312_));
 AND2x2_ASAP7_75t_R _734_ (.A(_306_),
    .B(_312_),
    .Y(_144_));
 AND3x1_ASAP7_75t_R _735_ (.A(_301_),
    .B(_224_),
    .C(net109),
    .Y(_313_));
 AO21x1_ASAP7_75t_R _736_ (.A1(net72),
    .A2(_225_),
    .B(_313_),
    .Y(_314_));
 AND2x2_ASAP7_75t_R _737_ (.A(_306_),
    .B(_314_),
    .Y(_145_));
 NAND2x2_ASAP7_75t_R _738_ (.A(_218_),
    .B(net99),
    .Y(_315_));
 BUFx6f_ASAP7_75t_R _739_ (.A(_315_),
    .Y(_316_));
 AND3x1_ASAP7_75t_R _740_ (.A(_301_),
    .B(_296_),
    .C(net74),
    .Y(_317_));
 AO21x1_ASAP7_75t_R _741_ (.A1(net1),
    .A2(_316_),
    .B(_317_),
    .Y(_318_));
 AND2x2_ASAP7_75t_R _742_ (.A(_306_),
    .B(_318_),
    .Y(_146_));
 AND3x1_ASAP7_75t_R _743_ (.A(_301_),
    .B(_296_),
    .C(net75),
    .Y(_319_));
 AO21x1_ASAP7_75t_R _744_ (.A1(net2),
    .A2(_316_),
    .B(_319_),
    .Y(_320_));
 AND2x2_ASAP7_75t_R _745_ (.A(_306_),
    .B(_320_),
    .Y(_147_));
 AND3x1_ASAP7_75t_R _746_ (.A(_301_),
    .B(_296_),
    .C(net76),
    .Y(_321_));
 AO21x1_ASAP7_75t_R _747_ (.A1(net3),
    .A2(_316_),
    .B(_321_),
    .Y(_322_));
 AND2x2_ASAP7_75t_R _748_ (.A(_306_),
    .B(_322_),
    .Y(_148_));
 AND3x1_ASAP7_75t_R _749_ (.A(_301_),
    .B(_296_),
    .C(net77),
    .Y(_323_));
 AO21x1_ASAP7_75t_R _750_ (.A1(net4),
    .A2(_316_),
    .B(_323_),
    .Y(_324_));
 AND2x2_ASAP7_75t_R _751_ (.A(_306_),
    .B(_324_),
    .Y(_149_));
 BUFx6f_ASAP7_75t_R _752_ (.A(_218_),
    .Y(_325_));
 AND3x1_ASAP7_75t_R _753_ (.A(_325_),
    .B(_296_),
    .C(net78),
    .Y(_326_));
 AO21x1_ASAP7_75t_R _754_ (.A1(net5),
    .A2(_316_),
    .B(_326_),
    .Y(_327_));
 AND2x2_ASAP7_75t_R _755_ (.A(_306_),
    .B(_327_),
    .Y(_150_));
 AND3x1_ASAP7_75t_R _756_ (.A(_325_),
    .B(_296_),
    .C(net79),
    .Y(_328_));
 AO21x1_ASAP7_75t_R _757_ (.A1(net6),
    .A2(_316_),
    .B(_328_),
    .Y(_329_));
 AND2x2_ASAP7_75t_R _758_ (.A(_306_),
    .B(_329_),
    .Y(_151_));
 BUFx6f_ASAP7_75t_R _759_ (.A(_222_),
    .Y(_330_));
 AND3x1_ASAP7_75t_R _760_ (.A(_325_),
    .B(_296_),
    .C(net80),
    .Y(_331_));
 AO21x1_ASAP7_75t_R _761_ (.A1(net7),
    .A2(_316_),
    .B(_331_),
    .Y(_332_));
 AND2x2_ASAP7_75t_R _762_ (.A(_330_),
    .B(_332_),
    .Y(_152_));
 AND3x1_ASAP7_75t_R _763_ (.A(_325_),
    .B(_296_),
    .C(net81),
    .Y(_333_));
 AO21x1_ASAP7_75t_R _764_ (.A1(net8),
    .A2(_316_),
    .B(_333_),
    .Y(_334_));
 AND2x2_ASAP7_75t_R _765_ (.A(_330_),
    .B(_334_),
    .Y(_153_));
 AND3x1_ASAP7_75t_R _766_ (.A(_325_),
    .B(_296_),
    .C(net82),
    .Y(_335_));
 AO21x1_ASAP7_75t_R _767_ (.A1(net9),
    .A2(_316_),
    .B(_335_),
    .Y(_336_));
 AND2x2_ASAP7_75t_R _768_ (.A(_330_),
    .B(_336_),
    .Y(_154_));
 BUFx6f_ASAP7_75t_R _769_ (.A(_315_),
    .Y(_337_));
 BUFx6f_ASAP7_75t_R _770_ (.A(net99),
    .Y(_338_));
 BUFx6f_ASAP7_75t_R _771_ (.A(_338_),
    .Y(_339_));
 AND3x1_ASAP7_75t_R _772_ (.A(_325_),
    .B(_339_),
    .C(net83),
    .Y(_340_));
 AO21x1_ASAP7_75t_R _773_ (.A1(net10),
    .A2(_337_),
    .B(_340_),
    .Y(_341_));
 AND2x2_ASAP7_75t_R _774_ (.A(_330_),
    .B(_341_),
    .Y(_155_));
 AND3x1_ASAP7_75t_R _775_ (.A(_325_),
    .B(_339_),
    .C(net84),
    .Y(_342_));
 AO21x1_ASAP7_75t_R _776_ (.A1(net11),
    .A2(_337_),
    .B(_342_),
    .Y(_343_));
 AND2x2_ASAP7_75t_R _777_ (.A(_330_),
    .B(_343_),
    .Y(_156_));
 AND3x1_ASAP7_75t_R _778_ (.A(_325_),
    .B(_339_),
    .C(net85),
    .Y(_344_));
 AO21x1_ASAP7_75t_R _779_ (.A1(net12),
    .A2(_337_),
    .B(_344_),
    .Y(_345_));
 AND2x2_ASAP7_75t_R _780_ (.A(_330_),
    .B(_345_),
    .Y(_157_));
 AND3x1_ASAP7_75t_R _781_ (.A(_325_),
    .B(_339_),
    .C(net86),
    .Y(_346_));
 AO21x1_ASAP7_75t_R _782_ (.A1(net13),
    .A2(_337_),
    .B(_346_),
    .Y(_347_));
 AND2x2_ASAP7_75t_R _783_ (.A(_330_),
    .B(_347_),
    .Y(_158_));
 AND3x1_ASAP7_75t_R _784_ (.A(_325_),
    .B(_339_),
    .C(net87),
    .Y(_348_));
 AO21x1_ASAP7_75t_R _785_ (.A1(net14),
    .A2(_337_),
    .B(_348_),
    .Y(_349_));
 AND2x2_ASAP7_75t_R _786_ (.A(_330_),
    .B(_349_),
    .Y(_159_));
 BUFx6f_ASAP7_75t_R _787_ (.A(_218_),
    .Y(_350_));
 AND3x1_ASAP7_75t_R _788_ (.A(_350_),
    .B(_339_),
    .C(net88),
    .Y(_351_));
 AO21x1_ASAP7_75t_R _789_ (.A1(net15),
    .A2(_337_),
    .B(_351_),
    .Y(_352_));
 AND2x2_ASAP7_75t_R _790_ (.A(_330_),
    .B(_352_),
    .Y(_160_));
 AND3x1_ASAP7_75t_R _791_ (.A(_350_),
    .B(_339_),
    .C(net89),
    .Y(_353_));
 AO21x1_ASAP7_75t_R _792_ (.A1(net16),
    .A2(_337_),
    .B(_353_),
    .Y(_354_));
 AND2x2_ASAP7_75t_R _793_ (.A(_330_),
    .B(_354_),
    .Y(_161_));
 BUFx6f_ASAP7_75t_R _794_ (.A(_221_),
    .Y(_355_));
 BUFx6f_ASAP7_75t_R _795_ (.A(_355_),
    .Y(_356_));
 AND3x1_ASAP7_75t_R _796_ (.A(_350_),
    .B(_339_),
    .C(net90),
    .Y(_357_));
 AO21x1_ASAP7_75t_R _797_ (.A1(net17),
    .A2(_337_),
    .B(_357_),
    .Y(_358_));
 AND2x2_ASAP7_75t_R _798_ (.A(_356_),
    .B(_358_),
    .Y(_162_));
 AND3x1_ASAP7_75t_R _799_ (.A(_350_),
    .B(_339_),
    .C(net91),
    .Y(_359_));
 AO21x1_ASAP7_75t_R _800_ (.A1(net18),
    .A2(_337_),
    .B(_359_),
    .Y(_360_));
 AND2x2_ASAP7_75t_R _801_ (.A(_356_),
    .B(_360_),
    .Y(_163_));
 AND3x1_ASAP7_75t_R _802_ (.A(_350_),
    .B(_339_),
    .C(net92),
    .Y(_361_));
 AO21x1_ASAP7_75t_R _803_ (.A1(net19),
    .A2(_337_),
    .B(_361_),
    .Y(_362_));
 AND2x2_ASAP7_75t_R _804_ (.A(_356_),
    .B(_362_),
    .Y(_164_));
 BUFx6f_ASAP7_75t_R _805_ (.A(_315_),
    .Y(_363_));
 BUFx6f_ASAP7_75t_R _806_ (.A(_338_),
    .Y(_364_));
 AND3x1_ASAP7_75t_R _807_ (.A(_350_),
    .B(_364_),
    .C(net93),
    .Y(_365_));
 AO21x1_ASAP7_75t_R _808_ (.A1(net20),
    .A2(_363_),
    .B(_365_),
    .Y(_366_));
 AND2x2_ASAP7_75t_R _809_ (.A(_356_),
    .B(_366_),
    .Y(_165_));
 AND3x1_ASAP7_75t_R _810_ (.A(_350_),
    .B(_364_),
    .C(net94),
    .Y(_367_));
 AO21x1_ASAP7_75t_R _811_ (.A1(net21),
    .A2(_363_),
    .B(_367_),
    .Y(_368_));
 AND2x2_ASAP7_75t_R _812_ (.A(_356_),
    .B(_368_),
    .Y(_166_));
 AND3x1_ASAP7_75t_R _813_ (.A(_350_),
    .B(_364_),
    .C(net95),
    .Y(_369_));
 AO21x1_ASAP7_75t_R _814_ (.A1(net22),
    .A2(_363_),
    .B(_369_),
    .Y(_370_));
 AND2x2_ASAP7_75t_R _815_ (.A(_356_),
    .B(_370_),
    .Y(_167_));
 AND3x1_ASAP7_75t_R _816_ (.A(_350_),
    .B(_364_),
    .C(net96),
    .Y(_371_));
 AO21x1_ASAP7_75t_R _817_ (.A1(net23),
    .A2(_363_),
    .B(_371_),
    .Y(_372_));
 AND2x2_ASAP7_75t_R _818_ (.A(_356_),
    .B(_372_),
    .Y(_168_));
 AND3x1_ASAP7_75t_R _819_ (.A(_350_),
    .B(_364_),
    .C(net97),
    .Y(_373_));
 AO21x1_ASAP7_75t_R _820_ (.A1(net24),
    .A2(_363_),
    .B(_373_),
    .Y(_374_));
 AND2x2_ASAP7_75t_R _821_ (.A(_356_),
    .B(_374_),
    .Y(_169_));
 BUFx6f_ASAP7_75t_R _822_ (.A(_218_),
    .Y(_375_));
 AND3x1_ASAP7_75t_R _823_ (.A(_375_),
    .B(_364_),
    .C(net98),
    .Y(_376_));
 AO21x1_ASAP7_75t_R _824_ (.A1(net25),
    .A2(_363_),
    .B(_376_),
    .Y(_377_));
 AND2x2_ASAP7_75t_R _825_ (.A(_356_),
    .B(_377_),
    .Y(_170_));
 INVx1_ASAP7_75t_R _826_ (.A(net26),
    .Y(_378_));
 AOI21x1_ASAP7_75t_R _827_ (.A1(_378_),
    .A2(_316_),
    .B(net73),
    .Y(_171_));
 AND3x1_ASAP7_75t_R _828_ (.A(_375_),
    .B(_364_),
    .C(net100),
    .Y(_379_));
 AO21x1_ASAP7_75t_R _829_ (.A1(net27),
    .A2(_363_),
    .B(_379_),
    .Y(_380_));
 AND2x2_ASAP7_75t_R _830_ (.A(_356_),
    .B(_380_),
    .Y(_172_));
 AND3x1_ASAP7_75t_R _831_ (.A(_375_),
    .B(_364_),
    .C(net101),
    .Y(_381_));
 AO21x1_ASAP7_75t_R _832_ (.A1(net28),
    .A2(_363_),
    .B(_381_),
    .Y(_382_));
 AND2x2_ASAP7_75t_R _833_ (.A(_287_),
    .B(_382_),
    .Y(_173_));
 INVx1_ASAP7_75t_R _834_ (.A(net28),
    .Y(_383_));
 INVx1_ASAP7_75t_R _835_ (.A(net27),
    .Y(_384_));
 AO21x1_ASAP7_75t_R _836_ (.A1(net65),
    .A2(net29),
    .B(_338_),
    .Y(_385_));
 AO32x1_ASAP7_75t_R _837_ (.A1(net29),
    .A2(_383_),
    .A3(_384_),
    .B1(_385_),
    .B2(_219_),
    .Y(_386_));
 AND2x2_ASAP7_75t_R _838_ (.A(_287_),
    .B(_386_),
    .Y(_174_));
 AND3x1_ASAP7_75t_R _839_ (.A(_375_),
    .B(_364_),
    .C(net103),
    .Y(_387_));
 AO21x1_ASAP7_75t_R _840_ (.A1(net30),
    .A2(_363_),
    .B(_387_),
    .Y(_388_));
 AND2x2_ASAP7_75t_R _841_ (.A(_287_),
    .B(_388_),
    .Y(_175_));
 AND3x1_ASAP7_75t_R _842_ (.A(_375_),
    .B(_364_),
    .C(net104),
    .Y(_389_));
 AO21x1_ASAP7_75t_R _843_ (.A1(net31),
    .A2(_363_),
    .B(_389_),
    .Y(_390_));
 AND2x2_ASAP7_75t_R _844_ (.A(_287_),
    .B(_390_),
    .Y(_176_));
 AND3x1_ASAP7_75t_R _845_ (.A(_375_),
    .B(_338_),
    .C(net105),
    .Y(_391_));
 AO21x1_ASAP7_75t_R _846_ (.A1(net32),
    .A2(_315_),
    .B(_391_),
    .Y(_392_));
 AND2x2_ASAP7_75t_R _847_ (.A(_287_),
    .B(_392_),
    .Y(_177_));
 AND3x1_ASAP7_75t_R _848_ (.A(_375_),
    .B(_338_),
    .C(net106),
    .Y(_393_));
 AO21x1_ASAP7_75t_R _849_ (.A1(net33),
    .A2(_315_),
    .B(_393_),
    .Y(_394_));
 AND2x2_ASAP7_75t_R _850_ (.A(_287_),
    .B(_394_),
    .Y(_178_));
 AND3x1_ASAP7_75t_R _851_ (.A(_375_),
    .B(_338_),
    .C(net107),
    .Y(_395_));
 AO21x1_ASAP7_75t_R _852_ (.A1(net34),
    .A2(_315_),
    .B(_395_),
    .Y(_396_));
 AND2x2_ASAP7_75t_R _853_ (.A(_287_),
    .B(_396_),
    .Y(_179_));
 AND3x1_ASAP7_75t_R _854_ (.A(_375_),
    .B(_338_),
    .C(net108),
    .Y(_397_));
 AO21x1_ASAP7_75t_R _855_ (.A1(net35),
    .A2(_315_),
    .B(_397_),
    .Y(_398_));
 AND2x2_ASAP7_75t_R _856_ (.A(_287_),
    .B(_398_),
    .Y(_180_));
 AND3x1_ASAP7_75t_R _857_ (.A(_375_),
    .B(_338_),
    .C(net109),
    .Y(_399_));
 AO21x1_ASAP7_75t_R _858_ (.A1(net36),
    .A2(_315_),
    .B(_399_),
    .Y(_400_));
 AND2x2_ASAP7_75t_R _859_ (.A(_287_),
    .B(_400_),
    .Y(_181_));
 AND4x1_ASAP7_75t_R _860_ (.A(_297_),
    .B(net65),
    .C(_292_),
    .D(_293_),
    .Y(_401_));
 BUFx6f_ASAP7_75t_R _861_ (.A(_401_),
    .Y(_402_));
 AND3x1_ASAP7_75t_R _862_ (.A(_218_),
    .B(_224_),
    .C(net65),
    .Y(_403_));
 BUFx6f_ASAP7_75t_R _863_ (.A(_403_),
    .Y(_404_));
 NOR2x2_ASAP7_75t_R _864_ (.A(_402_),
    .B(_404_),
    .Y(_405_));
 BUFx6f_ASAP7_75t_R _865_ (.A(_405_),
    .Y(_406_));
 BUFx6f_ASAP7_75t_R _866_ (.A(_286_),
    .Y(_407_));
 AND2x2_ASAP7_75t_R _867_ (.A(_407_),
    .B(net1),
    .Y(_408_));
 BUFx6f_ASAP7_75t_R _868_ (.A(_402_),
    .Y(_409_));
 BUFx6f_ASAP7_75t_R _869_ (.A(_404_),
    .Y(_410_));
 OA211x2_ASAP7_75t_R _870_ (.A1(_409_),
    .A2(_410_),
    .B(_355_),
    .C(net37),
    .Y(_411_));
 AO21x1_ASAP7_75t_R _871_ (.A1(_406_),
    .A2(_408_),
    .B(_411_),
    .Y(_182_));
 AND2x2_ASAP7_75t_R _872_ (.A(_407_),
    .B(net2),
    .Y(_412_));
 OA211x2_ASAP7_75t_R _873_ (.A1(_409_),
    .A2(_410_),
    .B(_355_),
    .C(net38),
    .Y(_413_));
 AO21x1_ASAP7_75t_R _874_ (.A1(_406_),
    .A2(_412_),
    .B(_413_),
    .Y(_183_));
 AND2x2_ASAP7_75t_R _875_ (.A(_407_),
    .B(net3),
    .Y(_414_));
 OA211x2_ASAP7_75t_R _876_ (.A1(_409_),
    .A2(_410_),
    .B(_355_),
    .C(net39),
    .Y(_415_));
 AO21x1_ASAP7_75t_R _877_ (.A1(_406_),
    .A2(_414_),
    .B(_415_),
    .Y(_184_));
 AND2x2_ASAP7_75t_R _878_ (.A(_407_),
    .B(net4),
    .Y(_416_));
 OA211x2_ASAP7_75t_R _879_ (.A1(_409_),
    .A2(_410_),
    .B(_355_),
    .C(net40),
    .Y(_417_));
 AO21x1_ASAP7_75t_R _880_ (.A1(_406_),
    .A2(_416_),
    .B(_417_),
    .Y(_185_));
 AND2x2_ASAP7_75t_R _881_ (.A(_407_),
    .B(net5),
    .Y(_418_));
 OA211x2_ASAP7_75t_R _882_ (.A1(_409_),
    .A2(_410_),
    .B(_355_),
    .C(net41),
    .Y(_419_));
 AO21x1_ASAP7_75t_R _883_ (.A1(_406_),
    .A2(_418_),
    .B(_419_),
    .Y(_186_));
 AND2x2_ASAP7_75t_R _884_ (.A(_407_),
    .B(net6),
    .Y(_420_));
 OA211x2_ASAP7_75t_R _885_ (.A1(_409_),
    .A2(_410_),
    .B(_355_),
    .C(net42),
    .Y(_421_));
 AO21x1_ASAP7_75t_R _886_ (.A1(_406_),
    .A2(_420_),
    .B(_421_),
    .Y(_187_));
 AND2x2_ASAP7_75t_R _887_ (.A(_407_),
    .B(net7),
    .Y(_422_));
 OA211x2_ASAP7_75t_R _888_ (.A1(_409_),
    .A2(_410_),
    .B(_355_),
    .C(net43),
    .Y(_423_));
 AO21x1_ASAP7_75t_R _889_ (.A1(_406_),
    .A2(_422_),
    .B(_423_),
    .Y(_188_));
 AND2x2_ASAP7_75t_R _890_ (.A(_407_),
    .B(net8),
    .Y(_424_));
 OA211x2_ASAP7_75t_R _891_ (.A1(_409_),
    .A2(_410_),
    .B(_355_),
    .C(net44),
    .Y(_425_));
 AO21x1_ASAP7_75t_R _892_ (.A1(_406_),
    .A2(_424_),
    .B(_425_),
    .Y(_189_));
 AND2x2_ASAP7_75t_R _893_ (.A(_407_),
    .B(net9),
    .Y(_426_));
 OA211x2_ASAP7_75t_R _894_ (.A1(_409_),
    .A2(_410_),
    .B(_355_),
    .C(net45),
    .Y(_427_));
 AO21x1_ASAP7_75t_R _895_ (.A1(_406_),
    .A2(_426_),
    .B(_427_),
    .Y(_190_));
 AND2x2_ASAP7_75t_R _896_ (.A(_407_),
    .B(net10),
    .Y(_428_));
 BUFx3_ASAP7_75t_R _897_ (.A(_221_),
    .Y(_429_));
 OA211x2_ASAP7_75t_R _898_ (.A1(_409_),
    .A2(_410_),
    .B(_429_),
    .C(net46),
    .Y(_430_));
 AO21x1_ASAP7_75t_R _899_ (.A1(_406_),
    .A2(_428_),
    .B(_430_),
    .Y(_191_));
 BUFx6f_ASAP7_75t_R _900_ (.A(_405_),
    .Y(_431_));
 BUFx6f_ASAP7_75t_R _901_ (.A(_286_),
    .Y(_432_));
 AND2x2_ASAP7_75t_R _902_ (.A(_432_),
    .B(net11),
    .Y(_433_));
 BUFx6f_ASAP7_75t_R _903_ (.A(_402_),
    .Y(_434_));
 BUFx6f_ASAP7_75t_R _904_ (.A(_404_),
    .Y(_435_));
 OA211x2_ASAP7_75t_R _905_ (.A1(_434_),
    .A2(_435_),
    .B(_429_),
    .C(net47),
    .Y(_436_));
 AO21x1_ASAP7_75t_R _906_ (.A1(_431_),
    .A2(_433_),
    .B(_436_),
    .Y(_192_));
 AND2x2_ASAP7_75t_R _907_ (.A(_432_),
    .B(net12),
    .Y(_437_));
 OA211x2_ASAP7_75t_R _908_ (.A1(_434_),
    .A2(_435_),
    .B(_429_),
    .C(net48),
    .Y(_438_));
 AO21x1_ASAP7_75t_R _909_ (.A1(_431_),
    .A2(_437_),
    .B(_438_),
    .Y(_193_));
 AND2x2_ASAP7_75t_R _910_ (.A(_432_),
    .B(net13),
    .Y(_439_));
 OA211x2_ASAP7_75t_R _911_ (.A1(_434_),
    .A2(_435_),
    .B(_429_),
    .C(net49),
    .Y(_440_));
 AO21x1_ASAP7_75t_R _912_ (.A1(_431_),
    .A2(_439_),
    .B(_440_),
    .Y(_194_));
 AND2x2_ASAP7_75t_R _913_ (.A(_432_),
    .B(net14),
    .Y(_441_));
 OA211x2_ASAP7_75t_R _914_ (.A1(_434_),
    .A2(_435_),
    .B(_429_),
    .C(net50),
    .Y(_442_));
 AO21x1_ASAP7_75t_R _915_ (.A1(_431_),
    .A2(_441_),
    .B(_442_),
    .Y(_195_));
 AND2x2_ASAP7_75t_R _916_ (.A(_432_),
    .B(net15),
    .Y(_443_));
 OA211x2_ASAP7_75t_R _917_ (.A1(_434_),
    .A2(_435_),
    .B(_429_),
    .C(net51),
    .Y(_444_));
 AO21x1_ASAP7_75t_R _918_ (.A1(_431_),
    .A2(_443_),
    .B(_444_),
    .Y(_196_));
 AND2x2_ASAP7_75t_R _919_ (.A(_432_),
    .B(net16),
    .Y(_445_));
 OA211x2_ASAP7_75t_R _920_ (.A1(_434_),
    .A2(_435_),
    .B(_429_),
    .C(net52),
    .Y(_446_));
 AO21x1_ASAP7_75t_R _921_ (.A1(_431_),
    .A2(_445_),
    .B(_446_),
    .Y(_197_));
 AND2x2_ASAP7_75t_R _922_ (.A(_432_),
    .B(net17),
    .Y(_447_));
 OA211x2_ASAP7_75t_R _923_ (.A1(_434_),
    .A2(_435_),
    .B(_429_),
    .C(net53),
    .Y(_448_));
 AO21x1_ASAP7_75t_R _924_ (.A1(_431_),
    .A2(_447_),
    .B(_448_),
    .Y(_198_));
 AND2x2_ASAP7_75t_R _925_ (.A(_432_),
    .B(net18),
    .Y(_449_));
 OA211x2_ASAP7_75t_R _926_ (.A1(_434_),
    .A2(_435_),
    .B(_429_),
    .C(net54),
    .Y(_450_));
 AO21x1_ASAP7_75t_R _927_ (.A1(_431_),
    .A2(_449_),
    .B(_450_),
    .Y(_199_));
 AND2x2_ASAP7_75t_R _928_ (.A(_432_),
    .B(net19),
    .Y(_451_));
 OA211x2_ASAP7_75t_R _929_ (.A1(_434_),
    .A2(_435_),
    .B(_429_),
    .C(net55),
    .Y(_452_));
 AO21x1_ASAP7_75t_R _930_ (.A1(_431_),
    .A2(_451_),
    .B(_452_),
    .Y(_200_));
 AND2x2_ASAP7_75t_R _931_ (.A(_432_),
    .B(net20),
    .Y(_453_));
 BUFx6f_ASAP7_75t_R _932_ (.A(_221_),
    .Y(_454_));
 OA211x2_ASAP7_75t_R _933_ (.A1(_434_),
    .A2(_435_),
    .B(_454_),
    .C(net56),
    .Y(_455_));
 AO21x1_ASAP7_75t_R _934_ (.A1(_431_),
    .A2(_453_),
    .B(_455_),
    .Y(_201_));
 BUFx6f_ASAP7_75t_R _935_ (.A(_405_),
    .Y(_456_));
 BUFx6f_ASAP7_75t_R _936_ (.A(_286_),
    .Y(_457_));
 AND2x2_ASAP7_75t_R _937_ (.A(_457_),
    .B(net21),
    .Y(_458_));
 BUFx6f_ASAP7_75t_R _938_ (.A(_402_),
    .Y(_459_));
 BUFx6f_ASAP7_75t_R _939_ (.A(_404_),
    .Y(_460_));
 OA211x2_ASAP7_75t_R _940_ (.A1(_459_),
    .A2(_460_),
    .B(_454_),
    .C(net57),
    .Y(_461_));
 AO21x1_ASAP7_75t_R _941_ (.A1(_456_),
    .A2(_458_),
    .B(_461_),
    .Y(_202_));
 AND2x2_ASAP7_75t_R _942_ (.A(_457_),
    .B(net22),
    .Y(_462_));
 OA211x2_ASAP7_75t_R _943_ (.A1(_459_),
    .A2(_460_),
    .B(_454_),
    .C(net58),
    .Y(_463_));
 AO21x1_ASAP7_75t_R _944_ (.A1(_456_),
    .A2(_462_),
    .B(_463_),
    .Y(_203_));
 AND2x2_ASAP7_75t_R _945_ (.A(_457_),
    .B(net23),
    .Y(_464_));
 OA211x2_ASAP7_75t_R _946_ (.A1(_459_),
    .A2(_460_),
    .B(_454_),
    .C(net59),
    .Y(_465_));
 AO21x1_ASAP7_75t_R _947_ (.A1(_456_),
    .A2(_464_),
    .B(_465_),
    .Y(_204_));
 AND2x2_ASAP7_75t_R _948_ (.A(_457_),
    .B(net24),
    .Y(_466_));
 OA211x2_ASAP7_75t_R _949_ (.A1(_459_),
    .A2(_460_),
    .B(_454_),
    .C(net60),
    .Y(_467_));
 AO21x1_ASAP7_75t_R _950_ (.A1(_456_),
    .A2(_466_),
    .B(_467_),
    .Y(_205_));
 AND2x2_ASAP7_75t_R _951_ (.A(_457_),
    .B(net25),
    .Y(_468_));
 OA211x2_ASAP7_75t_R _952_ (.A1(_459_),
    .A2(_460_),
    .B(_454_),
    .C(net61),
    .Y(_469_));
 AO21x1_ASAP7_75t_R _953_ (.A1(_456_),
    .A2(_468_),
    .B(_469_),
    .Y(_206_));
 AND2x2_ASAP7_75t_R _954_ (.A(net26),
    .B(_222_),
    .Y(_470_));
 OA211x2_ASAP7_75t_R _955_ (.A1(_459_),
    .A2(_460_),
    .B(net62),
    .C(_286_),
    .Y(_471_));
 AO21x1_ASAP7_75t_R _956_ (.A1(_456_),
    .A2(_470_),
    .B(_471_),
    .Y(_207_));
 AND2x2_ASAP7_75t_R _957_ (.A(net27),
    .B(_222_),
    .Y(_472_));
 OA211x2_ASAP7_75t_R _958_ (.A1(_459_),
    .A2(_460_),
    .B(net63),
    .C(_286_),
    .Y(_473_));
 AO21x1_ASAP7_75t_R _959_ (.A1(_456_),
    .A2(_472_),
    .B(_473_),
    .Y(_208_));
 AND2x2_ASAP7_75t_R _960_ (.A(net28),
    .B(_222_),
    .Y(_474_));
 OA211x2_ASAP7_75t_R _961_ (.A1(_459_),
    .A2(_460_),
    .B(net64),
    .C(_286_),
    .Y(_475_));
 AO21x1_ASAP7_75t_R _962_ (.A1(_456_),
    .A2(_474_),
    .B(_475_),
    .Y(_209_));
 NAND2x1_ASAP7_75t_R _963_ (.A(_338_),
    .B(net29),
    .Y(_476_));
 OA21x2_ASAP7_75t_R _964_ (.A1(_338_),
    .A2(_294_),
    .B(_476_),
    .Y(_477_));
 NAND3x1_ASAP7_75t_R _965_ (.A(_297_),
    .B(net65),
    .C(_292_),
    .Y(_478_));
 OA211x2_ASAP7_75t_R _966_ (.A1(_297_),
    .A2(_477_),
    .B(_478_),
    .C(_293_),
    .Y(_479_));
 NOR2x1_ASAP7_75t_R _967_ (.A(net73),
    .B(_479_),
    .Y(_210_));
 AND2x2_ASAP7_75t_R _968_ (.A(_457_),
    .B(net30),
    .Y(_480_));
 OA211x2_ASAP7_75t_R _969_ (.A1(_459_),
    .A2(_460_),
    .B(_454_),
    .C(net66),
    .Y(_481_));
 AO21x1_ASAP7_75t_R _970_ (.A1(_456_),
    .A2(_480_),
    .B(_481_),
    .Y(_211_));
 AND2x2_ASAP7_75t_R _971_ (.A(_457_),
    .B(net31),
    .Y(_482_));
 OA211x2_ASAP7_75t_R _972_ (.A1(_459_),
    .A2(_460_),
    .B(_454_),
    .C(net67),
    .Y(_483_));
 AO21x1_ASAP7_75t_R _973_ (.A1(_456_),
    .A2(_482_),
    .B(_483_),
    .Y(_212_));
 AND2x2_ASAP7_75t_R _974_ (.A(_457_),
    .B(net32),
    .Y(_484_));
 OA211x2_ASAP7_75t_R _975_ (.A1(_402_),
    .A2(_404_),
    .B(_454_),
    .C(net68),
    .Y(_485_));
 AO21x1_ASAP7_75t_R _976_ (.A1(_405_),
    .A2(_484_),
    .B(_485_),
    .Y(_213_));
 AND2x2_ASAP7_75t_R _977_ (.A(_457_),
    .B(net33),
    .Y(_486_));
 OA211x2_ASAP7_75t_R _978_ (.A1(_402_),
    .A2(_404_),
    .B(_454_),
    .C(net69),
    .Y(_487_));
 AO21x1_ASAP7_75t_R _979_ (.A1(_405_),
    .A2(_486_),
    .B(_487_),
    .Y(_214_));
 AND2x2_ASAP7_75t_R _980_ (.A(_457_),
    .B(net34),
    .Y(_488_));
 OA211x2_ASAP7_75t_R _981_ (.A1(_402_),
    .A2(_404_),
    .B(_286_),
    .C(net70),
    .Y(_489_));
 AO21x1_ASAP7_75t_R _982_ (.A1(_405_),
    .A2(_488_),
    .B(_489_),
    .Y(_215_));
 AND2x2_ASAP7_75t_R _983_ (.A(_222_),
    .B(net35),
    .Y(_490_));
 OA211x2_ASAP7_75t_R _984_ (.A1(_402_),
    .A2(_404_),
    .B(_286_),
    .C(net71),
    .Y(_491_));
 AO21x1_ASAP7_75t_R _985_ (.A1(_405_),
    .A2(_490_),
    .B(_491_),
    .Y(_216_));
 AND2x2_ASAP7_75t_R _986_ (.A(_222_),
    .B(net36),
    .Y(_492_));
 OA211x2_ASAP7_75t_R _987_ (.A1(_402_),
    .A2(_404_),
    .B(_286_),
    .C(net72),
    .Y(_493_));
 AO21x1_ASAP7_75t_R _988_ (.A1(_405_),
    .A2(_492_),
    .B(_493_),
    .Y(_217_));
 BUFx2_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx2_ASAP7_75t_R _990_ (.A(net219),
    .Y(l_o[35]));
 BUFx2_ASAP7_75t_R _991_ (.A(net220),
    .Y(r_o[35]));
 BUFx2_ASAP7_75t_R _992_ (.A(net221),
    .Y(u0_o[35]));
 DFFHQNx1_ASAP7_75t_R \done_sig$_DFF_P_  (.CLK(clknet_3_0__leaf_clk),
    .D(_000_),
    .QN(_109_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_110_),
    .QN(_108_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[10]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_111_),
    .QN(_107_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[11]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_112_),
    .QN(_106_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[12]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_113_),
    .QN(_105_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[13]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_114_),
    .QN(_104_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[14]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_115_),
    .QN(_103_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[15]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_116_),
    .QN(_102_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[16]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_117_),
    .QN(_101_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[17]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_118_),
    .QN(_100_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[18]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_119_),
    .QN(_099_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[19]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_120_),
    .QN(_098_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_121_),
    .QN(_097_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[20]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_122_),
    .QN(_096_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[21]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_123_),
    .QN(_095_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[22]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_124_),
    .QN(_094_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[23]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_125_),
    .QN(_093_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[24]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_126_),
    .QN(_092_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[25]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_127_),
    .QN(_091_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[26]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_128_),
    .QN(_090_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[27]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_129_),
    .QN(_089_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[28]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_130_),
    .QN(_088_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[29]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_131_),
    .QN(_087_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_132_),
    .QN(_086_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[30]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_133_),
    .QN(_085_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_134_),
    .QN(_084_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_3_1__leaf_clk),
    .D(_135_),
    .QN(_083_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_136_),
    .QN(_082_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_137_),
    .QN(_081_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_3_1__leaf_clk),
    .D(_138_),
    .QN(_080_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_139_),
    .QN(_079_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_140_),
    .QN(_078_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[5]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_141_),
    .QN(_077_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[6]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_142_),
    .QN(_076_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[7]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_143_),
    .QN(_075_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[8]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_144_),
    .QN(_074_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[9]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_145_),
    .QN(_073_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_146_),
    .QN(_072_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[10]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_147_),
    .QN(_071_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[11]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_148_),
    .QN(_070_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[12]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_149_),
    .QN(_069_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[13]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_150_),
    .QN(_068_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[14]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_151_),
    .QN(_067_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[15]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_152_),
    .QN(_066_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[16]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_153_),
    .QN(_065_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[17]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_154_),
    .QN(_064_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[18]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_155_),
    .QN(_063_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[19]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_156_),
    .QN(_062_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_157_),
    .QN(_061_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[20]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_158_),
    .QN(_060_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[21]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_159_),
    .QN(_059_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[22]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_160_),
    .QN(_058_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[23]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_161_),
    .QN(_057_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[24]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_162_),
    .QN(_056_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[25]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_163_),
    .QN(_055_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[26]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_164_),
    .QN(_054_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[27]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_165_),
    .QN(_053_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[28]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_166_),
    .QN(_052_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[29]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_167_),
    .QN(_051_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_168_),
    .QN(_050_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[30]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_169_),
    .QN(_049_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_170_),
    .QN(_048_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_171_),
    .QN(_047_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_172_),
    .QN(_046_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_3_1__leaf_clk),
    .D(_173_),
    .QN(_045_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_3_1__leaf_clk),
    .D(_174_),
    .QN(_044_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_3_1__leaf_clk),
    .D(_175_),
    .QN(_043_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_3_1__leaf_clk),
    .D(_176_),
    .QN(_042_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[5]$_SDFF_PP0_  (.CLK(clknet_3_1__leaf_clk),
    .D(_177_),
    .QN(_041_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[6]$_SDFF_PP0_  (.CLK(clknet_3_1__leaf_clk),
    .D(_178_),
    .QN(_040_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[7]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_179_),
    .QN(_039_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[8]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_180_),
    .QN(_038_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[9]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_181_),
    .QN(_037_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_182_),
    .QN(_036_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[10]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_183_),
    .QN(_035_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[11]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_184_),
    .QN(_034_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[12]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_185_),
    .QN(_033_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[13]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_186_),
    .QN(_032_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[14]$_SDFF_PP0_  (.CLK(clknet_3_2__leaf_clk),
    .D(_187_),
    .QN(_031_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[15]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_188_),
    .QN(_030_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[16]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_189_),
    .QN(_029_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[17]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_190_),
    .QN(_028_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[18]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_191_),
    .QN(_027_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[19]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_192_),
    .QN(_026_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_193_),
    .QN(_025_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[20]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_194_),
    .QN(_024_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[21]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_195_),
    .QN(_023_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[22]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_196_),
    .QN(_022_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[23]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_197_),
    .QN(_021_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[24]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_198_),
    .QN(_020_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[25]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_199_),
    .QN(_019_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[26]$_SDFF_PP0_  (.CLK(clknet_3_7__leaf_clk),
    .D(_200_),
    .QN(_018_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[27]$_SDFF_PP0_  (.CLK(clknet_3_6__leaf_clk),
    .D(_201_),
    .QN(_017_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[28]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_202_),
    .QN(_016_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[29]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_203_),
    .QN(_015_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_204_),
    .QN(_014_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[30]$_SDFF_PP0_  (.CLK(clknet_3_5__leaf_clk),
    .D(_205_),
    .QN(_013_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_206_),
    .QN(_012_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_207_),
    .QN(_011_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_208_),
    .QN(_010_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_209_),
    .QN(_009_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_3_3__leaf_clk),
    .D(_210_),
    .QN(_008_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_211_),
    .QN(_007_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .D(_212_),
    .QN(_006_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[5]$_SDFF_PP0_  (.CLK(clknet_3_1__leaf_clk),
    .D(_213_),
    .QN(_005_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[6]$_SDFF_PP0_  (.CLK(clknet_3_1__leaf_clk),
    .D(_214_),
    .QN(_004_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[7]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_215_),
    .QN(_003_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[8]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_216_),
    .QN(_002_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[9]$_SDFF_PP0_  (.CLK(clknet_3_0__leaf_clk),
    .D(_217_),
    .QN(_001_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_95 ();
 BUFx3_ASAP7_75t_R input1 (.A(l_i[0]),
    .Y(net1));
 BUFx3_ASAP7_75t_R input2 (.A(l_i[10]),
    .Y(net2));
 BUFx3_ASAP7_75t_R input3 (.A(l_i[11]),
    .Y(net3));
 BUFx3_ASAP7_75t_R input4 (.A(l_i[12]),
    .Y(net4));
 BUFx3_ASAP7_75t_R input5 (.A(l_i[13]),
    .Y(net5));
 BUFx3_ASAP7_75t_R input6 (.A(l_i[14]),
    .Y(net6));
 BUFx3_ASAP7_75t_R input7 (.A(l_i[15]),
    .Y(net7));
 BUFx3_ASAP7_75t_R input8 (.A(l_i[16]),
    .Y(net8));
 BUFx3_ASAP7_75t_R input9 (.A(l_i[17]),
    .Y(net9));
 BUFx3_ASAP7_75t_R input10 (.A(l_i[18]),
    .Y(net10));
 BUFx3_ASAP7_75t_R input11 (.A(l_i[19]),
    .Y(net11));
 BUFx3_ASAP7_75t_R input12 (.A(l_i[1]),
    .Y(net12));
 BUFx3_ASAP7_75t_R input13 (.A(l_i[20]),
    .Y(net13));
 BUFx3_ASAP7_75t_R input14 (.A(l_i[21]),
    .Y(net14));
 BUFx3_ASAP7_75t_R input15 (.A(l_i[22]),
    .Y(net15));
 BUFx3_ASAP7_75t_R input16 (.A(l_i[23]),
    .Y(net16));
 BUFx3_ASAP7_75t_R input17 (.A(l_i[24]),
    .Y(net17));
 BUFx3_ASAP7_75t_R input18 (.A(l_i[25]),
    .Y(net18));
 BUFx3_ASAP7_75t_R input19 (.A(l_i[26]),
    .Y(net19));
 BUFx3_ASAP7_75t_R input20 (.A(l_i[27]),
    .Y(net20));
 BUFx3_ASAP7_75t_R input21 (.A(l_i[28]),
    .Y(net21));
 BUFx3_ASAP7_75t_R input22 (.A(l_i[29]),
    .Y(net22));
 BUFx3_ASAP7_75t_R input23 (.A(l_i[2]),
    .Y(net23));
 BUFx3_ASAP7_75t_R input24 (.A(l_i[30]),
    .Y(net24));
 BUFx3_ASAP7_75t_R input25 (.A(l_i[31]),
    .Y(net25));
 BUFx3_ASAP7_75t_R input26 (.A(l_i[32]),
    .Y(net26));
 BUFx3_ASAP7_75t_R input27 (.A(l_i[33]),
    .Y(net27));
 BUFx3_ASAP7_75t_R input28 (.A(l_i[34]),
    .Y(net28));
 BUFx3_ASAP7_75t_R input29 (.A(l_i[36]),
    .Y(net29));
 BUFx3_ASAP7_75t_R input30 (.A(l_i[3]),
    .Y(net30));
 BUFx3_ASAP7_75t_R input31 (.A(l_i[4]),
    .Y(net31));
 BUFx3_ASAP7_75t_R input32 (.A(l_i[5]),
    .Y(net32));
 BUFx3_ASAP7_75t_R input33 (.A(l_i[6]),
    .Y(net33));
 BUFx3_ASAP7_75t_R input34 (.A(l_i[7]),
    .Y(net34));
 BUFx3_ASAP7_75t_R input35 (.A(l_i[8]),
    .Y(net35));
 BUFx3_ASAP7_75t_R input36 (.A(l_i[9]),
    .Y(net36));
 BUFx3_ASAP7_75t_R input37 (.A(r_i[0]),
    .Y(net37));
 BUFx3_ASAP7_75t_R input38 (.A(r_i[10]),
    .Y(net38));
 BUFx3_ASAP7_75t_R input39 (.A(r_i[11]),
    .Y(net39));
 BUFx3_ASAP7_75t_R input40 (.A(r_i[12]),
    .Y(net40));
 BUFx3_ASAP7_75t_R input41 (.A(r_i[13]),
    .Y(net41));
 BUFx3_ASAP7_75t_R input42 (.A(r_i[14]),
    .Y(net42));
 BUFx3_ASAP7_75t_R input43 (.A(r_i[15]),
    .Y(net43));
 BUFx3_ASAP7_75t_R input44 (.A(r_i[16]),
    .Y(net44));
 BUFx3_ASAP7_75t_R input45 (.A(r_i[17]),
    .Y(net45));
 BUFx3_ASAP7_75t_R input46 (.A(r_i[18]),
    .Y(net46));
 BUFx3_ASAP7_75t_R input47 (.A(r_i[19]),
    .Y(net47));
 BUFx3_ASAP7_75t_R input48 (.A(r_i[1]),
    .Y(net48));
 BUFx3_ASAP7_75t_R input49 (.A(r_i[20]),
    .Y(net49));
 BUFx3_ASAP7_75t_R input50 (.A(r_i[21]),
    .Y(net50));
 BUFx3_ASAP7_75t_R input51 (.A(r_i[22]),
    .Y(net51));
 BUFx3_ASAP7_75t_R input52 (.A(r_i[23]),
    .Y(net52));
 BUFx3_ASAP7_75t_R input53 (.A(r_i[24]),
    .Y(net53));
 BUFx3_ASAP7_75t_R input54 (.A(r_i[25]),
    .Y(net54));
 BUFx3_ASAP7_75t_R input55 (.A(r_i[26]),
    .Y(net55));
 BUFx3_ASAP7_75t_R input56 (.A(r_i[27]),
    .Y(net56));
 BUFx3_ASAP7_75t_R input57 (.A(r_i[28]),
    .Y(net57));
 BUFx3_ASAP7_75t_R input58 (.A(r_i[29]),
    .Y(net58));
 BUFx3_ASAP7_75t_R input59 (.A(r_i[2]),
    .Y(net59));
 BUFx3_ASAP7_75t_R input60 (.A(r_i[30]),
    .Y(net60));
 BUFx3_ASAP7_75t_R input61 (.A(r_i[31]),
    .Y(net61));
 BUFx3_ASAP7_75t_R input62 (.A(r_i[32]),
    .Y(net62));
 BUFx3_ASAP7_75t_R input63 (.A(r_i[33]),
    .Y(net63));
 BUFx3_ASAP7_75t_R input64 (.A(r_i[34]),
    .Y(net64));
 BUFx3_ASAP7_75t_R input65 (.A(r_i[36]),
    .Y(net65));
 BUFx3_ASAP7_75t_R input66 (.A(r_i[3]),
    .Y(net66));
 BUFx3_ASAP7_75t_R input67 (.A(r_i[4]),
    .Y(net67));
 BUFx3_ASAP7_75t_R input68 (.A(r_i[5]),
    .Y(net68));
 BUFx3_ASAP7_75t_R input69 (.A(r_i[6]),
    .Y(net69));
 BUFx3_ASAP7_75t_R input70 (.A(r_i[7]),
    .Y(net70));
 BUFx3_ASAP7_75t_R input71 (.A(r_i[8]),
    .Y(net71));
 BUFx3_ASAP7_75t_R input72 (.A(r_i[9]),
    .Y(net72));
 BUFx6f_ASAP7_75t_R input73 (.A(rst),
    .Y(net73));
 BUFx3_ASAP7_75t_R input74 (.A(u0_i[0]),
    .Y(net74));
 BUFx3_ASAP7_75t_R input75 (.A(u0_i[10]),
    .Y(net75));
 BUFx3_ASAP7_75t_R input76 (.A(u0_i[11]),
    .Y(net76));
 BUFx3_ASAP7_75t_R input77 (.A(u0_i[12]),
    .Y(net77));
 BUFx3_ASAP7_75t_R input78 (.A(u0_i[13]),
    .Y(net78));
 BUFx3_ASAP7_75t_R input79 (.A(u0_i[14]),
    .Y(net79));
 BUFx3_ASAP7_75t_R input80 (.A(u0_i[15]),
    .Y(net80));
 BUFx3_ASAP7_75t_R input81 (.A(u0_i[16]),
    .Y(net81));
 BUFx3_ASAP7_75t_R input82 (.A(u0_i[17]),
    .Y(net82));
 BUFx3_ASAP7_75t_R input83 (.A(u0_i[18]),
    .Y(net83));
 BUFx3_ASAP7_75t_R input84 (.A(u0_i[19]),
    .Y(net84));
 BUFx3_ASAP7_75t_R input85 (.A(u0_i[1]),
    .Y(net85));
 BUFx3_ASAP7_75t_R input86 (.A(u0_i[20]),
    .Y(net86));
 BUFx3_ASAP7_75t_R input87 (.A(u0_i[21]),
    .Y(net87));
 BUFx3_ASAP7_75t_R input88 (.A(u0_i[22]),
    .Y(net88));
 BUFx3_ASAP7_75t_R input89 (.A(u0_i[23]),
    .Y(net89));
 BUFx3_ASAP7_75t_R input90 (.A(u0_i[24]),
    .Y(net90));
 BUFx3_ASAP7_75t_R input91 (.A(u0_i[25]),
    .Y(net91));
 BUFx3_ASAP7_75t_R input92 (.A(u0_i[26]),
    .Y(net92));
 BUFx3_ASAP7_75t_R input93 (.A(u0_i[27]),
    .Y(net93));
 BUFx3_ASAP7_75t_R input94 (.A(u0_i[28]),
    .Y(net94));
 BUFx3_ASAP7_75t_R input95 (.A(u0_i[29]),
    .Y(net95));
 BUFx3_ASAP7_75t_R input96 (.A(u0_i[2]),
    .Y(net96));
 BUFx3_ASAP7_75t_R input97 (.A(u0_i[30]),
    .Y(net97));
 BUFx3_ASAP7_75t_R input98 (.A(u0_i[31]),
    .Y(net98));
 BUFx6f_ASAP7_75t_R input99 (.A(u0_i[32]),
    .Y(net99));
 BUFx3_ASAP7_75t_R input100 (.A(u0_i[33]),
    .Y(net100));
 BUFx3_ASAP7_75t_R input101 (.A(u0_i[34]),
    .Y(net101));
 BUFx3_ASAP7_75t_R input102 (.A(u0_i[36]),
    .Y(net102));
 BUFx3_ASAP7_75t_R input103 (.A(u0_i[3]),
    .Y(net103));
 BUFx3_ASAP7_75t_R input104 (.A(u0_i[4]),
    .Y(net104));
 BUFx3_ASAP7_75t_R input105 (.A(u0_i[5]),
    .Y(net105));
 BUFx3_ASAP7_75t_R input106 (.A(u0_i[6]),
    .Y(net106));
 BUFx3_ASAP7_75t_R input107 (.A(u0_i[7]),
    .Y(net107));
 BUFx3_ASAP7_75t_R input108 (.A(u0_i[8]),
    .Y(net108));
 BUFx3_ASAP7_75t_R input109 (.A(u0_i[9]),
    .Y(net109));
 BUFx3_ASAP7_75t_R output110 (.A(net110),
    .Y(done));
 BUFx3_ASAP7_75t_R output111 (.A(net111),
    .Y(l_o[0]));
 BUFx3_ASAP7_75t_R output112 (.A(net112),
    .Y(l_o[10]));
 BUFx3_ASAP7_75t_R output113 (.A(net113),
    .Y(l_o[11]));
 BUFx3_ASAP7_75t_R output114 (.A(net114),
    .Y(l_o[12]));
 BUFx3_ASAP7_75t_R output115 (.A(net115),
    .Y(l_o[13]));
 BUFx3_ASAP7_75t_R output116 (.A(net116),
    .Y(l_o[14]));
 BUFx3_ASAP7_75t_R output117 (.A(net117),
    .Y(l_o[15]));
 BUFx3_ASAP7_75t_R output118 (.A(net118),
    .Y(l_o[16]));
 BUFx3_ASAP7_75t_R output119 (.A(net119),
    .Y(l_o[17]));
 BUFx3_ASAP7_75t_R output120 (.A(net120),
    .Y(l_o[18]));
 BUFx3_ASAP7_75t_R output121 (.A(net121),
    .Y(l_o[19]));
 BUFx3_ASAP7_75t_R output122 (.A(net122),
    .Y(l_o[1]));
 BUFx3_ASAP7_75t_R output123 (.A(net123),
    .Y(l_o[20]));
 BUFx3_ASAP7_75t_R output124 (.A(net124),
    .Y(l_o[21]));
 BUFx3_ASAP7_75t_R output125 (.A(net125),
    .Y(l_o[22]));
 BUFx3_ASAP7_75t_R output126 (.A(net126),
    .Y(l_o[23]));
 BUFx3_ASAP7_75t_R output127 (.A(net127),
    .Y(l_o[24]));
 BUFx3_ASAP7_75t_R output128 (.A(net128),
    .Y(l_o[25]));
 BUFx3_ASAP7_75t_R output129 (.A(net129),
    .Y(l_o[26]));
 BUFx3_ASAP7_75t_R output130 (.A(net130),
    .Y(l_o[27]));
 BUFx3_ASAP7_75t_R output131 (.A(net131),
    .Y(l_o[28]));
 BUFx3_ASAP7_75t_R output132 (.A(net132),
    .Y(l_o[29]));
 BUFx3_ASAP7_75t_R output133 (.A(net133),
    .Y(l_o[2]));
 BUFx3_ASAP7_75t_R output134 (.A(net134),
    .Y(l_o[30]));
 BUFx3_ASAP7_75t_R output135 (.A(net135),
    .Y(l_o[31]));
 BUFx3_ASAP7_75t_R output136 (.A(net136),
    .Y(l_o[32]));
 BUFx3_ASAP7_75t_R output137 (.A(net137),
    .Y(l_o[33]));
 BUFx3_ASAP7_75t_R output138 (.A(net138),
    .Y(l_o[34]));
 BUFx3_ASAP7_75t_R output139 (.A(net139),
    .Y(l_o[36]));
 BUFx3_ASAP7_75t_R output140 (.A(net140),
    .Y(l_o[3]));
 BUFx3_ASAP7_75t_R output141 (.A(net141),
    .Y(l_o[4]));
 BUFx3_ASAP7_75t_R output142 (.A(net142),
    .Y(l_o[5]));
 BUFx3_ASAP7_75t_R output143 (.A(net143),
    .Y(l_o[6]));
 BUFx3_ASAP7_75t_R output144 (.A(net144),
    .Y(l_o[7]));
 BUFx3_ASAP7_75t_R output145 (.A(net145),
    .Y(l_o[8]));
 BUFx3_ASAP7_75t_R output146 (.A(net146),
    .Y(l_o[9]));
 BUFx3_ASAP7_75t_R output147 (.A(net147),
    .Y(r_o[0]));
 BUFx3_ASAP7_75t_R output148 (.A(net148),
    .Y(r_o[10]));
 BUFx3_ASAP7_75t_R output149 (.A(net149),
    .Y(r_o[11]));
 BUFx3_ASAP7_75t_R output150 (.A(net150),
    .Y(r_o[12]));
 BUFx3_ASAP7_75t_R output151 (.A(net151),
    .Y(r_o[13]));
 BUFx3_ASAP7_75t_R output152 (.A(net152),
    .Y(r_o[14]));
 BUFx3_ASAP7_75t_R output153 (.A(net153),
    .Y(r_o[15]));
 BUFx3_ASAP7_75t_R output154 (.A(net154),
    .Y(r_o[16]));
 BUFx3_ASAP7_75t_R output155 (.A(net155),
    .Y(r_o[17]));
 BUFx3_ASAP7_75t_R output156 (.A(net156),
    .Y(r_o[18]));
 BUFx3_ASAP7_75t_R output157 (.A(net157),
    .Y(r_o[19]));
 BUFx3_ASAP7_75t_R output158 (.A(net158),
    .Y(r_o[1]));
 BUFx3_ASAP7_75t_R output159 (.A(net159),
    .Y(r_o[20]));
 BUFx3_ASAP7_75t_R output160 (.A(net160),
    .Y(r_o[21]));
 BUFx3_ASAP7_75t_R output161 (.A(net161),
    .Y(r_o[22]));
 BUFx3_ASAP7_75t_R output162 (.A(net162),
    .Y(r_o[23]));
 BUFx3_ASAP7_75t_R output163 (.A(net163),
    .Y(r_o[24]));
 BUFx3_ASAP7_75t_R output164 (.A(net164),
    .Y(r_o[25]));
 BUFx3_ASAP7_75t_R output165 (.A(net165),
    .Y(r_o[26]));
 BUFx3_ASAP7_75t_R output166 (.A(net166),
    .Y(r_o[27]));
 BUFx3_ASAP7_75t_R output167 (.A(net167),
    .Y(r_o[28]));
 BUFx3_ASAP7_75t_R output168 (.A(net168),
    .Y(r_o[29]));
 BUFx3_ASAP7_75t_R output169 (.A(net169),
    .Y(r_o[2]));
 BUFx3_ASAP7_75t_R output170 (.A(net170),
    .Y(r_o[30]));
 BUFx3_ASAP7_75t_R output171 (.A(net171),
    .Y(r_o[31]));
 BUFx3_ASAP7_75t_R output172 (.A(net172),
    .Y(r_o[32]));
 BUFx3_ASAP7_75t_R output173 (.A(net173),
    .Y(r_o[33]));
 BUFx3_ASAP7_75t_R output174 (.A(net174),
    .Y(r_o[34]));
 BUFx3_ASAP7_75t_R output175 (.A(net175),
    .Y(r_o[36]));
 BUFx3_ASAP7_75t_R output176 (.A(net176),
    .Y(r_o[3]));
 BUFx3_ASAP7_75t_R output177 (.A(net177),
    .Y(r_o[4]));
 BUFx3_ASAP7_75t_R output178 (.A(net178),
    .Y(r_o[5]));
 BUFx3_ASAP7_75t_R output179 (.A(net179),
    .Y(r_o[6]));
 BUFx3_ASAP7_75t_R output180 (.A(net180),
    .Y(r_o[7]));
 BUFx3_ASAP7_75t_R output181 (.A(net181),
    .Y(r_o[8]));
 BUFx3_ASAP7_75t_R output182 (.A(net182),
    .Y(r_o[9]));
 BUFx3_ASAP7_75t_R output183 (.A(net183),
    .Y(u0_o[0]));
 BUFx3_ASAP7_75t_R output184 (.A(net184),
    .Y(u0_o[10]));
 BUFx3_ASAP7_75t_R output185 (.A(net185),
    .Y(u0_o[11]));
 BUFx3_ASAP7_75t_R output186 (.A(net186),
    .Y(u0_o[12]));
 BUFx3_ASAP7_75t_R output187 (.A(net187),
    .Y(u0_o[13]));
 BUFx3_ASAP7_75t_R output188 (.A(net188),
    .Y(u0_o[14]));
 BUFx3_ASAP7_75t_R output189 (.A(net189),
    .Y(u0_o[15]));
 BUFx3_ASAP7_75t_R output190 (.A(net190),
    .Y(u0_o[16]));
 BUFx3_ASAP7_75t_R output191 (.A(net191),
    .Y(u0_o[17]));
 BUFx3_ASAP7_75t_R output192 (.A(net192),
    .Y(u0_o[18]));
 BUFx3_ASAP7_75t_R output193 (.A(net193),
    .Y(u0_o[19]));
 BUFx3_ASAP7_75t_R output194 (.A(net194),
    .Y(u0_o[1]));
 BUFx3_ASAP7_75t_R output195 (.A(net195),
    .Y(u0_o[20]));
 BUFx3_ASAP7_75t_R output196 (.A(net196),
    .Y(u0_o[21]));
 BUFx3_ASAP7_75t_R output197 (.A(net197),
    .Y(u0_o[22]));
 BUFx3_ASAP7_75t_R output198 (.A(net198),
    .Y(u0_o[23]));
 BUFx3_ASAP7_75t_R output199 (.A(net199),
    .Y(u0_o[24]));
 BUFx3_ASAP7_75t_R output200 (.A(net200),
    .Y(u0_o[25]));
 BUFx3_ASAP7_75t_R output201 (.A(net201),
    .Y(u0_o[26]));
 BUFx3_ASAP7_75t_R output202 (.A(net202),
    .Y(u0_o[27]));
 BUFx3_ASAP7_75t_R output203 (.A(net203),
    .Y(u0_o[28]));
 BUFx3_ASAP7_75t_R output204 (.A(net204),
    .Y(u0_o[29]));
 BUFx3_ASAP7_75t_R output205 (.A(net205),
    .Y(u0_o[2]));
 BUFx3_ASAP7_75t_R output206 (.A(net206),
    .Y(u0_o[30]));
 BUFx3_ASAP7_75t_R output207 (.A(net207),
    .Y(u0_o[31]));
 BUFx3_ASAP7_75t_R output208 (.A(net208),
    .Y(u0_o[32]));
 BUFx3_ASAP7_75t_R output209 (.A(net209),
    .Y(u0_o[33]));
 BUFx3_ASAP7_75t_R output210 (.A(net210),
    .Y(u0_o[34]));
 BUFx3_ASAP7_75t_R output211 (.A(net211),
    .Y(u0_o[36]));
 BUFx3_ASAP7_75t_R output212 (.A(net212),
    .Y(u0_o[3]));
 BUFx3_ASAP7_75t_R output213 (.A(net213),
    .Y(u0_o[4]));
 BUFx3_ASAP7_75t_R output214 (.A(net214),
    .Y(u0_o[5]));
 BUFx3_ASAP7_75t_R output215 (.A(net215),
    .Y(u0_o[6]));
 BUFx3_ASAP7_75t_R output216 (.A(net216),
    .Y(u0_o[7]));
 BUFx3_ASAP7_75t_R output217 (.A(net217),
    .Y(u0_o[8]));
 BUFx3_ASAP7_75t_R output218 (.A(net218),
    .Y(u0_o[9]));
 TIELOx1_ASAP7_75t_R _990__219 (.L(net219));
 TIELOx1_ASAP7_75t_R _991__220 (.L(net220));
 TIELOx1_ASAP7_75t_R _992__221 (.L(net221));
 BUFx2_ASAP7_75t_R clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_0__leaf_clk));
 BUFx2_ASAP7_75t_R clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_1__leaf_clk));
 BUFx2_ASAP7_75t_R clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_2__leaf_clk));
 BUFx2_ASAP7_75t_R clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_3__leaf_clk));
 BUFx2_ASAP7_75t_R clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_4__leaf_clk));
 BUFx2_ASAP7_75t_R clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_5__leaf_clk));
 BUFx2_ASAP7_75t_R clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_6__leaf_clk));
 BUFx2_ASAP7_75t_R clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_7__leaf_clk));
 BUFx12_ASAP7_75t_R clkload0 (.A(clknet_3_0__leaf_clk));
 INVx5_ASAP7_75t_R clkload1 (.A(clknet_3_1__leaf_clk));
 BUFx4f_ASAP7_75t_R clkload2 (.A(clknet_3_3__leaf_clk));
 INVxp67_ASAP7_75t_R clkload3 (.A(clknet_3_4__leaf_clk));
 BUFx4f_ASAP7_75t_R clkload4 (.A(clknet_3_5__leaf_clk));
 INVx3_ASAP7_75t_R clkload5 (.A(clknet_3_6__leaf_clk));
 INVxp67_ASAP7_75t_R clkload6 (.A(clknet_3_7__leaf_clk));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30 ();
 DECAPx4_ASAP7_75t_R FILLER_0_36 ();
 FILLER_ASAP7_75t_R FILLER_0_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48 ();
 FILLER_ASAP7_75t_R FILLER_0_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 FILLER_ASAP7_75t_R FILLER_1_24 ();
 DECAPx6_ASAP7_75t_R FILLER_1_37 ();
 DECAPx2_ASAP7_75t_R FILLER_1_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_57 ();
 FILLER_ASAP7_75t_R FILLER_1_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_155 ();
 DECAPx10_ASAP7_75t_R FILLER_1_214 ();
 DECAPx2_ASAP7_75t_R FILLER_1_236 ();
 FILLER_ASAP7_75t_R FILLER_1_242 ();
 DECAPx6_ASAP7_75t_R FILLER_2_2 ();
 DECAPx2_ASAP7_75t_R FILLER_2_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_22 ();
 DECAPx6_ASAP7_75t_R FILLER_2_31 ();
 DECAPx2_ASAP7_75t_R FILLER_2_45 ();
 FILLER_ASAP7_75t_R FILLER_2_132 ();
 FILLER_ASAP7_75t_R FILLER_2_206 ();
 DECAPx10_ASAP7_75t_R FILLER_2_211 ();
 DECAPx4_ASAP7_75t_R FILLER_2_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_243 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx1_ASAP7_75t_R FILLER_3_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_73 ();
 DECAPx2_ASAP7_75t_R FILLER_3_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_89 ();
 FILLER_ASAP7_75t_R FILLER_3_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_124 ();
 DECAPx4_ASAP7_75t_R FILLER_3_169 ();
 DECAPx10_ASAP7_75t_R FILLER_3_211 ();
 DECAPx4_ASAP7_75t_R FILLER_3_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_243 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx6_ASAP7_75t_R FILLER_4_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_96 ();
 FILLER_ASAP7_75t_R FILLER_4_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_148 ();
 DECAPx1_ASAP7_75t_R FILLER_4_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_171 ();
 DECAPx6_ASAP7_75t_R FILLER_4_187 ();
 DECAPx10_ASAP7_75t_R FILLER_4_207 ();
 DECAPx6_ASAP7_75t_R FILLER_4_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_243 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx6_ASAP7_75t_R FILLER_5_24 ();
 DECAPx2_ASAP7_75t_R FILLER_5_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_44 ();
 DECAPx10_ASAP7_75t_R FILLER_5_51 ();
 DECAPx10_ASAP7_75t_R FILLER_5_73 ();
 DECAPx1_ASAP7_75t_R FILLER_5_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_99 ();
 FILLER_ASAP7_75t_R FILLER_5_155 ();
 DECAPx1_ASAP7_75t_R FILLER_5_169 ();
 DECAPx10_ASAP7_75t_R FILLER_5_185 ();
 DECAPx10_ASAP7_75t_R FILLER_5_207 ();
 DECAPx6_ASAP7_75t_R FILLER_5_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_243 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_76 ();
 DECAPx10_ASAP7_75t_R FILLER_6_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_102 ();
 DECAPx2_ASAP7_75t_R FILLER_6_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_168 ();
 DECAPx4_ASAP7_75t_R FILLER_6_187 ();
 FILLER_ASAP7_75t_R FILLER_6_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_199 ();
 DECAPx2_ASAP7_75t_R FILLER_6_220 ();
 FILLER_ASAP7_75t_R FILLER_6_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_231 ();
 DECAPx2_ASAP7_75t_R FILLER_6_238 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 FILLER_ASAP7_75t_R FILLER_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_7_29 ();
 DECAPx2_ASAP7_75t_R FILLER_7_51 ();
 DECAPx1_ASAP7_75t_R FILLER_7_63 ();
 DECAPx2_ASAP7_75t_R FILLER_7_102 ();
 FILLER_ASAP7_75t_R FILLER_7_108 ();
 DECAPx2_ASAP7_75t_R FILLER_7_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_130 ();
 DECAPx10_ASAP7_75t_R FILLER_7_139 ();
 FILLER_ASAP7_75t_R FILLER_7_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_171 ();
 DECAPx2_ASAP7_75t_R FILLER_7_209 ();
 FILLER_ASAP7_75t_R FILLER_7_215 ();
 FILLER_ASAP7_75t_R FILLER_7_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_222 ();
 DECAPx1_ASAP7_75t_R FILLER_7_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_243 ();
 DECAPx4_ASAP7_75t_R FILLER_8_2 ();
 FILLER_ASAP7_75t_R FILLER_8_12 ();
 DECAPx6_ASAP7_75t_R FILLER_8_103 ();
 DECAPx1_ASAP7_75t_R FILLER_8_117 ();
 FILLER_ASAP7_75t_R FILLER_8_135 ();
 DECAPx1_ASAP7_75t_R FILLER_8_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_171 ();
 FILLER_ASAP7_75t_R FILLER_8_180 ();
 DECAPx10_ASAP7_75t_R FILLER_8_208 ();
 DECAPx6_ASAP7_75t_R FILLER_8_230 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_24 ();
 FILLER_ASAP7_75t_R FILLER_9_45 ();
 DECAPx6_ASAP7_75t_R FILLER_9_87 ();
 DECAPx2_ASAP7_75t_R FILLER_9_101 ();
 FILLER_ASAP7_75t_R FILLER_9_123 ();
 FILLER_ASAP7_75t_R FILLER_9_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_139 ();
 DECAPx4_ASAP7_75t_R FILLER_9_146 ();
 FILLER_ASAP7_75t_R FILLER_9_156 ();
 DECAPx10_ASAP7_75t_R FILLER_9_200 ();
 DECAPx10_ASAP7_75t_R FILLER_9_222 ();
 DECAPx6_ASAP7_75t_R FILLER_10_8 ();
 FILLER_ASAP7_75t_R FILLER_10_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_51 ();
 DECAPx1_ASAP7_75t_R FILLER_10_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_64 ();
 DECAPx10_ASAP7_75t_R FILLER_10_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_107 ();
 DECAPx4_ASAP7_75t_R FILLER_10_118 ();
 FILLER_ASAP7_75t_R FILLER_10_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_130 ();
 DECAPx1_ASAP7_75t_R FILLER_10_137 ();
 DECAPx10_ASAP7_75t_R FILLER_10_164 ();
 DECAPx6_ASAP7_75t_R FILLER_10_186 ();
 FILLER_ASAP7_75t_R FILLER_10_200 ();
 DECAPx4_ASAP7_75t_R FILLER_10_222 ();
 FILLER_ASAP7_75t_R FILLER_10_232 ();
 DECAPx1_ASAP7_75t_R FILLER_10_240 ();
 DECAPx2_ASAP7_75t_R FILLER_11_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_26 ();
 FILLER_ASAP7_75t_R FILLER_11_33 ();
 FILLER_ASAP7_75t_R FILLER_11_41 ();
 FILLER_ASAP7_75t_R FILLER_11_49 ();
 DECAPx1_ASAP7_75t_R FILLER_11_69 ();
 DECAPx2_ASAP7_75t_R FILLER_11_79 ();
 FILLER_ASAP7_75t_R FILLER_11_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_110 ();
 DECAPx2_ASAP7_75t_R FILLER_11_131 ();
 FILLER_ASAP7_75t_R FILLER_11_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_139 ();
 DECAPx2_ASAP7_75t_R FILLER_11_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_175 ();
 DECAPx4_ASAP7_75t_R FILLER_11_182 ();
 FILLER_ASAP7_75t_R FILLER_11_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_194 ();
 DECAPx6_ASAP7_75t_R FILLER_11_218 ();
 DECAPx1_ASAP7_75t_R FILLER_11_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_243 ();
 DECAPx2_ASAP7_75t_R FILLER_12_2 ();
 FILLER_ASAP7_75t_R FILLER_12_8 ();
 DECAPx10_ASAP7_75t_R FILLER_12_46 ();
 DECAPx6_ASAP7_75t_R FILLER_12_68 ();
 DECAPx2_ASAP7_75t_R FILLER_12_82 ();
 DECAPx6_ASAP7_75t_R FILLER_12_97 ();
 DECAPx1_ASAP7_75t_R FILLER_12_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_115 ();
 DECAPx10_ASAP7_75t_R FILLER_12_126 ();
 DECAPx4_ASAP7_75t_R FILLER_12_148 ();
 FILLER_ASAP7_75t_R FILLER_12_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_160 ();
 FILLER_ASAP7_75t_R FILLER_12_167 ();
 FILLER_ASAP7_75t_R FILLER_12_175 ();
 DECAPx2_ASAP7_75t_R FILLER_12_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_189 ();
 DECAPx2_ASAP7_75t_R FILLER_12_196 ();
 FILLER_ASAP7_75t_R FILLER_12_202 ();
 FILLER_ASAP7_75t_R FILLER_12_224 ();
 FILLER_ASAP7_75t_R FILLER_12_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_42 ();
 DECAPx4_ASAP7_75t_R FILLER_13_59 ();
 FILLER_ASAP7_75t_R FILLER_13_69 ();
 DECAPx2_ASAP7_75t_R FILLER_13_77 ();
 FILLER_ASAP7_75t_R FILLER_13_83 ();
 FILLER_ASAP7_75t_R FILLER_13_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_93 ();
 FILLER_ASAP7_75t_R FILLER_13_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_114 ();
 DECAPx10_ASAP7_75t_R FILLER_13_125 ();
 DECAPx6_ASAP7_75t_R FILLER_13_147 ();
 FILLER_ASAP7_75t_R FILLER_13_161 ();
 DECAPx1_ASAP7_75t_R FILLER_13_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_193 ();
 DECAPx1_ASAP7_75t_R FILLER_13_220 ();
 DECAPx6_ASAP7_75t_R FILLER_13_227 ();
 FILLER_ASAP7_75t_R FILLER_13_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_243 ();
 FILLER_ASAP7_75t_R FILLER_14_8 ();
 DECAPx2_ASAP7_75t_R FILLER_14_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_42 ();
 DECAPx2_ASAP7_75t_R FILLER_14_49 ();
 FILLER_ASAP7_75t_R FILLER_14_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_78 ();
 FILLER_ASAP7_75t_R FILLER_14_98 ();
 DECAPx1_ASAP7_75t_R FILLER_14_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_114 ();
 FILLER_ASAP7_75t_R FILLER_14_128 ();
 FILLER_ASAP7_75t_R FILLER_14_140 ();
 DECAPx4_ASAP7_75t_R FILLER_14_152 ();
 FILLER_ASAP7_75t_R FILLER_14_188 ();
 DECAPx2_ASAP7_75t_R FILLER_14_196 ();
 FILLER_ASAP7_75t_R FILLER_14_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_224 ();
 DECAPx4_ASAP7_75t_R FILLER_14_228 ();
 DECAPx2_ASAP7_75t_R FILLER_15_14 ();
 FILLER_ASAP7_75t_R FILLER_15_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_22 ();
 DECAPx1_ASAP7_75t_R FILLER_15_29 ();
 FILLER_ASAP7_75t_R FILLER_15_45 ();
 DECAPx1_ASAP7_75t_R FILLER_15_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_59 ();
 FILLER_ASAP7_75t_R FILLER_15_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_74 ();
 DECAPx4_ASAP7_75t_R FILLER_15_96 ();
 DECAPx4_ASAP7_75t_R FILLER_15_126 ();
 DECAPx10_ASAP7_75t_R FILLER_15_139 ();
 DECAPx1_ASAP7_75t_R FILLER_15_161 ();
 DECAPx1_ASAP7_75t_R FILLER_15_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_182 ();
 DECAPx2_ASAP7_75t_R FILLER_15_203 ();
 FILLER_ASAP7_75t_R FILLER_15_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_211 ();
 DECAPx6_ASAP7_75t_R FILLER_15_221 ();
 FILLER_ASAP7_75t_R FILLER_15_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_243 ();
 FILLER_ASAP7_75t_R FILLER_16_26 ();
 FILLER_ASAP7_75t_R FILLER_16_37 ();
 DECAPx2_ASAP7_75t_R FILLER_16_59 ();
 DECAPx1_ASAP7_75t_R FILLER_16_78 ();
 DECAPx2_ASAP7_75t_R FILLER_16_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_119 ();
 DECAPx10_ASAP7_75t_R FILLER_16_140 ();
 DECAPx4_ASAP7_75t_R FILLER_16_162 ();
 FILLER_ASAP7_75t_R FILLER_16_172 ();
 DECAPx1_ASAP7_75t_R FILLER_16_186 ();
 FILLER_ASAP7_75t_R FILLER_16_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_198 ();
 DECAPx2_ASAP7_75t_R FILLER_16_219 ();
 FILLER_ASAP7_75t_R FILLER_16_225 ();
 DECAPx1_ASAP7_75t_R FILLER_16_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_234 ();
 FILLER_ASAP7_75t_R FILLER_16_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_14 ();
 FILLER_ASAP7_75t_R FILLER_17_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_23 ();
 FILLER_ASAP7_75t_R FILLER_17_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_46 ();
 DECAPx6_ASAP7_75t_R FILLER_17_53 ();
 FILLER_ASAP7_75t_R FILLER_17_67 ();
 DECAPx6_ASAP7_75t_R FILLER_17_75 ();
 FILLER_ASAP7_75t_R FILLER_17_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_98 ();
 DECAPx6_ASAP7_75t_R FILLER_17_117 ();
 DECAPx1_ASAP7_75t_R FILLER_17_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_135 ();
 DECAPx1_ASAP7_75t_R FILLER_17_146 ();
 DECAPx10_ASAP7_75t_R FILLER_17_182 ();
 DECAPx10_ASAP7_75t_R FILLER_17_204 ();
 DECAPx2_ASAP7_75t_R FILLER_17_226 ();
 FILLER_ASAP7_75t_R FILLER_18_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_40 ();
 DECAPx6_ASAP7_75t_R FILLER_18_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_90 ();
 DECAPx2_ASAP7_75t_R FILLER_18_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_115 ();
 DECAPx6_ASAP7_75t_R FILLER_18_139 ();
 FILLER_ASAP7_75t_R FILLER_18_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_161 ();
 DECAPx2_ASAP7_75t_R FILLER_18_168 ();
 DECAPx2_ASAP7_75t_R FILLER_18_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_237 ();
 DECAPx1_ASAP7_75t_R FILLER_19_2 ();
 FILLER_ASAP7_75t_R FILLER_19_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_55 ();
 DECAPx2_ASAP7_75t_R FILLER_19_59 ();
 FILLER_ASAP7_75t_R FILLER_19_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_67 ();
 DECAPx6_ASAP7_75t_R FILLER_19_71 ();
 FILLER_ASAP7_75t_R FILLER_19_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_87 ();
 FILLER_ASAP7_75t_R FILLER_19_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_103 ();
 FILLER_ASAP7_75t_R FILLER_19_111 ();
 DECAPx6_ASAP7_75t_R FILLER_19_138 ();
 DECAPx2_ASAP7_75t_R FILLER_19_152 ();
 DECAPx2_ASAP7_75t_R FILLER_19_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_186 ();
 DECAPx4_ASAP7_75t_R FILLER_19_207 ();
 FILLER_ASAP7_75t_R FILLER_19_217 ();
 FILLER_ASAP7_75t_R FILLER_19_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_227 ();
 DECAPx2_ASAP7_75t_R FILLER_19_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_79 ();
 DECAPx10_ASAP7_75t_R FILLER_20_83 ();
 DECAPx1_ASAP7_75t_R FILLER_20_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_114 ();
 DECAPx10_ASAP7_75t_R FILLER_20_135 ();
 DECAPx2_ASAP7_75t_R FILLER_20_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_194 ();
 DECAPx2_ASAP7_75t_R FILLER_20_218 ();
 FILLER_ASAP7_75t_R FILLER_20_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_233 ();
 DECAPx1_ASAP7_75t_R FILLER_20_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_20 ();
 FILLER_ASAP7_75t_R FILLER_21_39 ();
 DECAPx10_ASAP7_75t_R FILLER_21_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_75 ();
 DECAPx1_ASAP7_75t_R FILLER_21_106 ();
 DECAPx2_ASAP7_75t_R FILLER_21_120 ();
 FILLER_ASAP7_75t_R FILLER_21_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_134 ();
 DECAPx2_ASAP7_75t_R FILLER_21_155 ();
 FILLER_ASAP7_75t_R FILLER_21_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_169 ();
 DECAPx10_ASAP7_75t_R FILLER_21_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_198 ();
 FILLER_ASAP7_75t_R FILLER_21_219 ();
 DECAPx1_ASAP7_75t_R FILLER_21_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_228 ();
 FILLER_ASAP7_75t_R FILLER_21_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_31 ();
 FILLER_ASAP7_75t_R FILLER_22_38 ();
 FILLER_ASAP7_75t_R FILLER_22_109 ();
 DECAPx10_ASAP7_75t_R FILLER_22_131 ();
 DECAPx4_ASAP7_75t_R FILLER_22_153 ();
 DECAPx1_ASAP7_75t_R FILLER_22_169 ();
 DECAPx10_ASAP7_75t_R FILLER_22_196 ();
 FILLER_ASAP7_75t_R FILLER_22_218 ();
 DECAPx4_ASAP7_75t_R FILLER_22_232 ();
 FILLER_ASAP7_75t_R FILLER_22_242 ();
 DECAPx1_ASAP7_75t_R FILLER_23_8 ();
 DECAPx6_ASAP7_75t_R FILLER_23_44 ();
 DECAPx2_ASAP7_75t_R FILLER_23_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_64 ();
 FILLER_ASAP7_75t_R FILLER_23_79 ();
 DECAPx1_ASAP7_75t_R FILLER_23_87 ();
 DECAPx1_ASAP7_75t_R FILLER_23_97 ();
 DECAPx10_ASAP7_75t_R FILLER_23_111 ();
 DECAPx10_ASAP7_75t_R FILLER_23_133 ();
 DECAPx10_ASAP7_75t_R FILLER_23_155 ();
 DECAPx6_ASAP7_75t_R FILLER_23_177 ();
 DECAPx6_ASAP7_75t_R FILLER_23_197 ();
 DECAPx1_ASAP7_75t_R FILLER_23_240 ();
 FILLER_ASAP7_75t_R FILLER_24_26 ();
 DECAPx2_ASAP7_75t_R FILLER_24_34 ();
 FILLER_ASAP7_75t_R FILLER_24_40 ();
 FILLER_ASAP7_75t_R FILLER_24_62 ();
 FILLER_ASAP7_75t_R FILLER_24_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_74 ();
 DECAPx10_ASAP7_75t_R FILLER_24_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_103 ();
 FILLER_ASAP7_75t_R FILLER_24_124 ();
 DECAPx10_ASAP7_75t_R FILLER_24_129 ();
 FILLER_ASAP7_75t_R FILLER_24_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_179 ();
 FILLER_ASAP7_75t_R FILLER_24_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_185 ();
 DECAPx6_ASAP7_75t_R FILLER_24_192 ();
 FILLER_ASAP7_75t_R FILLER_24_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_208 ();
 DECAPx4_ASAP7_75t_R FILLER_24_215 ();
 DECAPx2_ASAP7_75t_R FILLER_24_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_2 ();
 FILLER_ASAP7_75t_R FILLER_25_9 ();
 FILLER_ASAP7_75t_R FILLER_25_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_19 ();
 FILLER_ASAP7_75t_R FILLER_25_49 ();
 DECAPx4_ASAP7_75t_R FILLER_25_61 ();
 DECAPx10_ASAP7_75t_R FILLER_25_86 ();
 FILLER_ASAP7_75t_R FILLER_25_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_110 ();
 DECAPx6_ASAP7_75t_R FILLER_25_131 ();
 DECAPx2_ASAP7_75t_R FILLER_25_145 ();
 DECAPx6_ASAP7_75t_R FILLER_25_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_191 ();
 DECAPx1_ASAP7_75t_R FILLER_25_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_231 ();
 DECAPx2_ASAP7_75t_R FILLER_25_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_25 ();
 DECAPx2_ASAP7_75t_R FILLER_26_32 ();
 DECAPx1_ASAP7_75t_R FILLER_26_44 ();
 FILLER_ASAP7_75t_R FILLER_26_58 ();
 FILLER_ASAP7_75t_R FILLER_26_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_76 ();
 DECAPx4_ASAP7_75t_R FILLER_26_97 ();
 FILLER_ASAP7_75t_R FILLER_26_107 ();
 DECAPx6_ASAP7_75t_R FILLER_26_161 ();
 FILLER_ASAP7_75t_R FILLER_26_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_189 ();
 DECAPx2_ASAP7_75t_R FILLER_26_196 ();
 FILLER_ASAP7_75t_R FILLER_26_202 ();
 DECAPx1_ASAP7_75t_R FILLER_26_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_243 ();
 DECAPx2_ASAP7_75t_R FILLER_27_2 ();
 FILLER_ASAP7_75t_R FILLER_27_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_10 ();
 FILLER_ASAP7_75t_R FILLER_27_35 ();
 DECAPx10_ASAP7_75t_R FILLER_27_43 ();
 FILLER_ASAP7_75t_R FILLER_27_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_67 ();
 FILLER_ASAP7_75t_R FILLER_27_74 ();
 DECAPx10_ASAP7_75t_R FILLER_27_91 ();
 DECAPx2_ASAP7_75t_R FILLER_27_113 ();
 DECAPx2_ASAP7_75t_R FILLER_27_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_135 ();
 DECAPx10_ASAP7_75t_R FILLER_27_142 ();
 DECAPx1_ASAP7_75t_R FILLER_27_164 ();
 FILLER_ASAP7_75t_R FILLER_27_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_173 ();
 DECAPx10_ASAP7_75t_R FILLER_27_182 ();
 DECAPx4_ASAP7_75t_R FILLER_27_210 ();
 DECAPx1_ASAP7_75t_R FILLER_28_2 ();
 FILLER_ASAP7_75t_R FILLER_28_32 ();
 DECAPx6_ASAP7_75t_R FILLER_28_43 ();
 DECAPx2_ASAP7_75t_R FILLER_28_57 ();
 DECAPx10_ASAP7_75t_R FILLER_28_104 ();
 DECAPx4_ASAP7_75t_R FILLER_28_126 ();
 FILLER_ASAP7_75t_R FILLER_28_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_158 ();
 DECAPx2_ASAP7_75t_R FILLER_28_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_171 ();
 DECAPx2_ASAP7_75t_R FILLER_28_198 ();
 FILLER_ASAP7_75t_R FILLER_28_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_206 ();
 DECAPx2_ASAP7_75t_R FILLER_28_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_219 ();
 FILLER_ASAP7_75t_R FILLER_28_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_231 ();
 DECAPx2_ASAP7_75t_R FILLER_29_2 ();
 FILLER_ASAP7_75t_R FILLER_29_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_10 ();
 FILLER_ASAP7_75t_R FILLER_29_37 ();
 FILLER_ASAP7_75t_R FILLER_29_45 ();
 DECAPx2_ASAP7_75t_R FILLER_29_53 ();
 FILLER_ASAP7_75t_R FILLER_29_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_61 ();
 DECAPx1_ASAP7_75t_R FILLER_29_67 ();
 DECAPx2_ASAP7_75t_R FILLER_29_80 ();
 FILLER_ASAP7_75t_R FILLER_29_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_88 ();
 DECAPx10_ASAP7_75t_R FILLER_29_109 ();
 FILLER_ASAP7_75t_R FILLER_29_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_133 ();
 FILLER_ASAP7_75t_R FILLER_29_186 ();
 FILLER_ASAP7_75t_R FILLER_29_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_200 ();
 FILLER_ASAP7_75t_R FILLER_29_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_223 ();
 DECAPx4_ASAP7_75t_R FILLER_29_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_2 ();
 FILLER_ASAP7_75t_R FILLER_30_15 ();
 FILLER_ASAP7_75t_R FILLER_30_35 ();
 DECAPx1_ASAP7_75t_R FILLER_30_72 ();
 DECAPx10_ASAP7_75t_R FILLER_30_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_118 ();
 DECAPx6_ASAP7_75t_R FILLER_30_139 ();
 DECAPx1_ASAP7_75t_R FILLER_30_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_157 ();
 FILLER_ASAP7_75t_R FILLER_30_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_163 ();
 DECAPx1_ASAP7_75t_R FILLER_30_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_180 ();
 FILLER_ASAP7_75t_R FILLER_30_201 ();
 FILLER_ASAP7_75t_R FILLER_30_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_225 ();
 DECAPx6_ASAP7_75t_R FILLER_30_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_243 ();
 DECAPx2_ASAP7_75t_R FILLER_31_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_64 ();
 DECAPx10_ASAP7_75t_R FILLER_31_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_90 ();
 DECAPx4_ASAP7_75t_R FILLER_31_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_111 ();
 DECAPx1_ASAP7_75t_R FILLER_31_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_122 ();
 DECAPx1_ASAP7_75t_R FILLER_31_131 ();
 DECAPx6_ASAP7_75t_R FILLER_31_186 ();
 FILLER_ASAP7_75t_R FILLER_31_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_202 ();
 DECAPx2_ASAP7_75t_R FILLER_31_232 ();
 DECAPx1_ASAP7_75t_R FILLER_32_8 ();
 DECAPx4_ASAP7_75t_R FILLER_32_21 ();
 DECAPx2_ASAP7_75t_R FILLER_32_39 ();
 DECAPx2_ASAP7_75t_R FILLER_32_65 ();
 FILLER_ASAP7_75t_R FILLER_32_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_73 ();
 DECAPx4_ASAP7_75t_R FILLER_32_84 ();
 FILLER_ASAP7_75t_R FILLER_32_94 ();
 DECAPx10_ASAP7_75t_R FILLER_32_128 ();
 DECAPx6_ASAP7_75t_R FILLER_32_150 ();
 DECAPx2_ASAP7_75t_R FILLER_32_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_194 ();
 DECAPx10_ASAP7_75t_R FILLER_32_201 ();
 DECAPx6_ASAP7_75t_R FILLER_32_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_237 ();
 FILLER_ASAP7_75t_R FILLER_33_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_31 ();
 DECAPx6_ASAP7_75t_R FILLER_33_35 ();
 FILLER_ASAP7_75t_R FILLER_33_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_51 ();
 DECAPx10_ASAP7_75t_R FILLER_33_55 ();
 DECAPx10_ASAP7_75t_R FILLER_33_77 ();
 DECAPx6_ASAP7_75t_R FILLER_33_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_119 ();
 DECAPx10_ASAP7_75t_R FILLER_33_126 ();
 DECAPx10_ASAP7_75t_R FILLER_33_148 ();
 DECAPx1_ASAP7_75t_R FILLER_33_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_190 ();
 DECAPx2_ASAP7_75t_R FILLER_33_211 ();
 DECAPx2_ASAP7_75t_R FILLER_33_226 ();
 FILLER_ASAP7_75t_R FILLER_33_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_234 ();
 FILLER_ASAP7_75t_R FILLER_34_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_23 ();
 DECAPx6_ASAP7_75t_R FILLER_34_38 ();
 DECAPx1_ASAP7_75t_R FILLER_34_52 ();
 DECAPx1_ASAP7_75t_R FILLER_34_59 ();
 DECAPx6_ASAP7_75t_R FILLER_34_81 ();
 FILLER_ASAP7_75t_R FILLER_34_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_97 ();
 DECAPx6_ASAP7_75t_R FILLER_34_104 ();
 FILLER_ASAP7_75t_R FILLER_34_118 ();
 FILLER_ASAP7_75t_R FILLER_34_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_128 ();
 DECAPx6_ASAP7_75t_R FILLER_34_161 ();
 DECAPx1_ASAP7_75t_R FILLER_34_175 ();
 DECAPx2_ASAP7_75t_R FILLER_34_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_191 ();
 FILLER_ASAP7_75t_R FILLER_34_198 ();
 DECAPx10_ASAP7_75t_R FILLER_34_220 ();
 FILLER_ASAP7_75t_R FILLER_34_242 ();
 DECAPx2_ASAP7_75t_R FILLER_35_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_35 ();
 DECAPx2_ASAP7_75t_R FILLER_35_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_96 ();
 DECAPx6_ASAP7_75t_R FILLER_35_100 ();
 FILLER_ASAP7_75t_R FILLER_35_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_116 ();
 DECAPx1_ASAP7_75t_R FILLER_35_123 ();
 DECAPx4_ASAP7_75t_R FILLER_35_133 ();
 FILLER_ASAP7_75t_R FILLER_35_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_145 ();
 DECAPx6_ASAP7_75t_R FILLER_35_154 ();
 DECAPx1_ASAP7_75t_R FILLER_35_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_172 ();
 DECAPx10_ASAP7_75t_R FILLER_35_185 ();
 DECAPx4_ASAP7_75t_R FILLER_35_207 ();
 FILLER_ASAP7_75t_R FILLER_35_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_226 ();
 DECAPx4_ASAP7_75t_R FILLER_35_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_243 ();
 DECAPx2_ASAP7_75t_R FILLER_36_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_8 ();
 DECAPx2_ASAP7_75t_R FILLER_36_15 ();
 FILLER_ASAP7_75t_R FILLER_36_56 ();
 FILLER_ASAP7_75t_R FILLER_36_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_80 ();
 FILLER_ASAP7_75t_R FILLER_36_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_103 ();
 DECAPx2_ASAP7_75t_R FILLER_36_107 ();
 FILLER_ASAP7_75t_R FILLER_36_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_115 ();
 FILLER_ASAP7_75t_R FILLER_36_122 ();
 DECAPx4_ASAP7_75t_R FILLER_36_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_142 ();
 FILLER_ASAP7_75t_R FILLER_36_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_157 ();
 DECAPx1_ASAP7_75t_R FILLER_36_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_182 ();
 DECAPx1_ASAP7_75t_R FILLER_36_189 ();
 DECAPx2_ASAP7_75t_R FILLER_36_219 ();
 FILLER_ASAP7_75t_R FILLER_36_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_227 ();
 DECAPx1_ASAP7_75t_R FILLER_36_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_46 ();
 FILLER_ASAP7_75t_R FILLER_37_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_73 ();
 DECAPx10_ASAP7_75t_R FILLER_37_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_147 ();
 FILLER_ASAP7_75t_R FILLER_37_200 ();
 DECAPx4_ASAP7_75t_R FILLER_37_225 ();
 FILLER_ASAP7_75t_R FILLER_37_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_237 ();
 DECAPx1_ASAP7_75t_R FILLER_38_14 ();
 DECAPx2_ASAP7_75t_R FILLER_38_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_54 ();
 DECAPx2_ASAP7_75t_R FILLER_38_73 ();
 DECAPx1_ASAP7_75t_R FILLER_38_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_103 ();
 DECAPx1_ASAP7_75t_R FILLER_38_130 ();
 FILLER_ASAP7_75t_R FILLER_38_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_142 ();
 DECAPx6_ASAP7_75t_R FILLER_38_155 ();
 DECAPx1_ASAP7_75t_R FILLER_38_169 ();
 DECAPx10_ASAP7_75t_R FILLER_38_197 ();
 DECAPx4_ASAP7_75t_R FILLER_38_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_21 ();
 DECAPx2_ASAP7_75t_R FILLER_39_51 ();
 FILLER_ASAP7_75t_R FILLER_39_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_59 ();
 DECAPx1_ASAP7_75t_R FILLER_39_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_70 ();
 FILLER_ASAP7_75t_R FILLER_39_103 ();
 DECAPx1_ASAP7_75t_R FILLER_39_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_136 ();
 DECAPx1_ASAP7_75t_R FILLER_39_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_153 ();
 DECAPx4_ASAP7_75t_R FILLER_39_160 ();
 FILLER_ASAP7_75t_R FILLER_39_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_190 ();
 FILLER_ASAP7_75t_R FILLER_39_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_199 ();
 DECAPx6_ASAP7_75t_R FILLER_39_223 ();
 DECAPx2_ASAP7_75t_R FILLER_39_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_243 ();
 DECAPx2_ASAP7_75t_R FILLER_40_2 ();
 FILLER_ASAP7_75t_R FILLER_40_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_10 ();
 DECAPx2_ASAP7_75t_R FILLER_40_17 ();
 DECAPx2_ASAP7_75t_R FILLER_40_29 ();
 DECAPx6_ASAP7_75t_R FILLER_40_55 ();
 DECAPx1_ASAP7_75t_R FILLER_40_69 ();
 DECAPx1_ASAP7_75t_R FILLER_40_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_101 ();
 FILLER_ASAP7_75t_R FILLER_40_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_164 ();
 DECAPx10_ASAP7_75t_R FILLER_40_168 ();
 DECAPx4_ASAP7_75t_R FILLER_40_190 ();
 FILLER_ASAP7_75t_R FILLER_40_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_202 ();
 FILLER_ASAP7_75t_R FILLER_40_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_225 ();
 DECAPx2_ASAP7_75t_R FILLER_40_229 ();
 FILLER_ASAP7_75t_R FILLER_40_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_237 ();
 DECAPx6_ASAP7_75t_R FILLER_41_2 ();
 DECAPx1_ASAP7_75t_R FILLER_41_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_20 ();
 DECAPx4_ASAP7_75t_R FILLER_41_27 ();
 FILLER_ASAP7_75t_R FILLER_41_37 ();
 DECAPx10_ASAP7_75t_R FILLER_41_85 ();
 DECAPx4_ASAP7_75t_R FILLER_41_107 ();
 FILLER_ASAP7_75t_R FILLER_41_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_123 ();
 DECAPx2_ASAP7_75t_R FILLER_41_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_156 ();
 DECAPx6_ASAP7_75t_R FILLER_41_177 ();
 DECAPx1_ASAP7_75t_R FILLER_41_191 ();
 DECAPx6_ASAP7_75t_R FILLER_41_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_229 ();
 DECAPx1_ASAP7_75t_R FILLER_41_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_243 ();
 DECAPx10_ASAP7_75t_R FILLER_42_2 ();
 DECAPx10_ASAP7_75t_R FILLER_42_24 ();
 DECAPx10_ASAP7_75t_R FILLER_42_46 ();
 DECAPx10_ASAP7_75t_R FILLER_42_68 ();
 DECAPx10_ASAP7_75t_R FILLER_42_90 ();
 DECAPx10_ASAP7_75t_R FILLER_42_112 ();
 DECAPx2_ASAP7_75t_R FILLER_42_134 ();
 FILLER_ASAP7_75t_R FILLER_42_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_142 ();
 DECAPx6_ASAP7_75t_R FILLER_42_166 ();
 FILLER_ASAP7_75t_R FILLER_42_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_182 ();
 DECAPx4_ASAP7_75t_R FILLER_42_186 ();
 FILLER_ASAP7_75t_R FILLER_42_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_198 ();
 DECAPx1_ASAP7_75t_R FILLER_42_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_223 ();
 DECAPx6_ASAP7_75t_R FILLER_42_227 ();
 FILLER_ASAP7_75t_R FILLER_42_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_243 ();
 DECAPx10_ASAP7_75t_R FILLER_43_2 ();
 DECAPx10_ASAP7_75t_R FILLER_43_24 ();
 DECAPx6_ASAP7_75t_R FILLER_43_46 ();
 DECAPx10_ASAP7_75t_R FILLER_43_63 ();
 DECAPx10_ASAP7_75t_R FILLER_43_85 ();
 DECAPx10_ASAP7_75t_R FILLER_43_107 ();
 DECAPx10_ASAP7_75t_R FILLER_43_129 ();
 DECAPx4_ASAP7_75t_R FILLER_43_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_161 ();
 DECAPx10_ASAP7_75t_R FILLER_43_165 ();
 DECAPx10_ASAP7_75t_R FILLER_43_187 ();
 DECAPx10_ASAP7_75t_R FILLER_43_209 ();
 DECAPx4_ASAP7_75t_R FILLER_43_231 ();
 FILLER_ASAP7_75t_R FILLER_43_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_243 ();
 DECAPx10_ASAP7_75t_R FILLER_44_2 ();
 DECAPx10_ASAP7_75t_R FILLER_44_24 ();
 DECAPx6_ASAP7_75t_R FILLER_44_46 ();
 FILLER_ASAP7_75t_R FILLER_44_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_62 ();
 DECAPx10_ASAP7_75t_R FILLER_44_69 ();
 DECAPx6_ASAP7_75t_R FILLER_44_91 ();
 DECAPx1_ASAP7_75t_R FILLER_44_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_109 ();
 DECAPx6_ASAP7_75t_R FILLER_44_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_130 ();
 DECAPx2_ASAP7_75t_R FILLER_44_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_143 ();
 DECAPx10_ASAP7_75t_R FILLER_44_147 ();
 DECAPx10_ASAP7_75t_R FILLER_44_169 ();
 DECAPx10_ASAP7_75t_R FILLER_44_191 ();
 DECAPx10_ASAP7_75t_R FILLER_44_213 ();
 DECAPx2_ASAP7_75t_R FILLER_44_235 ();
 FILLER_ASAP7_75t_R FILLER_44_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_243 ();
 DECAPx10_ASAP7_75t_R FILLER_45_2 ();
 DECAPx10_ASAP7_75t_R FILLER_45_24 ();
 DECAPx6_ASAP7_75t_R FILLER_45_46 ();
 DECAPx1_ASAP7_75t_R FILLER_45_60 ();
 DECAPx10_ASAP7_75t_R FILLER_45_70 ();
 DECAPx10_ASAP7_75t_R FILLER_45_92 ();
 DECAPx2_ASAP7_75t_R FILLER_45_114 ();
 FILLER_ASAP7_75t_R FILLER_45_120 ();
 DECAPx2_ASAP7_75t_R FILLER_45_134 ();
 DECAPx10_ASAP7_75t_R FILLER_45_146 ();
 DECAPx4_ASAP7_75t_R FILLER_45_168 ();
 FILLER_ASAP7_75t_R FILLER_45_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_180 ();
 DECAPx10_ASAP7_75t_R FILLER_45_187 ();
 DECAPx10_ASAP7_75t_R FILLER_45_209 ();
 DECAPx4_ASAP7_75t_R FILLER_45_231 ();
 FILLER_ASAP7_75t_R FILLER_45_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_243 ();
 DECAPx10_ASAP7_75t_R FILLER_46_2 ();
 DECAPx10_ASAP7_75t_R FILLER_46_24 ();
 DECAPx6_ASAP7_75t_R FILLER_46_46 ();
 DECAPx1_ASAP7_75t_R FILLER_46_60 ();
 DECAPx2_ASAP7_75t_R FILLER_46_88 ();
 FILLER_ASAP7_75t_R FILLER_46_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_96 ();
 DECAPx2_ASAP7_75t_R FILLER_46_103 ();
 DECAPx1_ASAP7_75t_R FILLER_46_145 ();
 DECAPx1_ASAP7_75t_R FILLER_46_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_166 ();
 DECAPx2_ASAP7_75t_R FILLER_46_179 ();
 FILLER_ASAP7_75t_R FILLER_46_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_187 ();
 DECAPx10_ASAP7_75t_R FILLER_46_194 ();
 DECAPx10_ASAP7_75t_R FILLER_46_216 ();
 DECAPx2_ASAP7_75t_R FILLER_46_238 ();
 DECAPx10_ASAP7_75t_R FILLER_47_2 ();
 DECAPx6_ASAP7_75t_R FILLER_47_24 ();
 DECAPx1_ASAP7_75t_R FILLER_47_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_42 ();
 DECAPx4_ASAP7_75t_R FILLER_47_49 ();
 FILLER_ASAP7_75t_R FILLER_47_59 ();
 FILLER_ASAP7_75t_R FILLER_47_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_81 ();
 DECAPx2_ASAP7_75t_R FILLER_47_160 ();
 FILLER_ASAP7_75t_R FILLER_47_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_168 ();
 FILLER_ASAP7_75t_R FILLER_47_175 ();
 DECAPx10_ASAP7_75t_R FILLER_47_189 ();
 DECAPx10_ASAP7_75t_R FILLER_47_211 ();
 DECAPx4_ASAP7_75t_R FILLER_47_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_243 ();
endmodule
