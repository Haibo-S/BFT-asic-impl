module t_switch (ce,
    clk,
    done,
    l_i_bp,
    l_i_v,
    l_o_bp,
    l_o_v,
    r_i_bp,
    r_i_v,
    r_o_bp,
    r_o_v,
    rst,
    u0_i_bp,
    u0_i_v,
    u0_o_bp,
    u0_o_v,
    l_i,
    l_o,
    r_i,
    r_o,
    u0_i,
    u0_o);
 input ce;
 input clk;
 output done;
 output l_i_bp;
 input l_i_v;
 input l_o_bp;
 output l_o_v;
 output r_i_bp;
 input r_i_v;
 input r_o_bp;
 output r_o_v;
 input rst;
 output u0_i_bp;
 input u0_i_v;
 input u0_o_bp;
 output u0_o_v;
 input [35:0] l_i;
 output [35:0] l_o;
 input [35:0] r_i;
 output [35:0] r_o;
 input [35:0] u0_i;
 output [35:0] u0_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 INVx1_ASAP7_75t_R _0684_ (.A(net64),
    .Y(_0342_));
 NOR2x1_ASAP7_75t_R _0685_ (.A(net66),
    .B(net65),
    .Y(_0343_));
 AND3x4_ASAP7_75t_R _0686_ (.A(net75),
    .B(_0342_),
    .C(_0343_),
    .Y(_0344_));
 BUFx6f_ASAP7_75t_R _0687_ (.A(_0005_),
    .Y(_0345_));
 BUFx6f_ASAP7_75t_R _0688_ (.A(u0_i_v),
    .Y(_0346_));
 INVx2_ASAP7_75t_R _0689_ (.A(net102),
    .Y(_0347_));
 AND2x2_ASAP7_75t_R _0690_ (.A(_0346_),
    .B(_0347_),
    .Y(_0348_));
 AO21x1_ASAP7_75t_R _0691_ (.A1(_0345_),
    .A2(_0348_),
    .B(net38),
    .Y(_0349_));
 OA21x2_ASAP7_75t_R _0692_ (.A1(net66),
    .A2(net65),
    .B(net75),
    .Y(_0350_));
 OA21x2_ASAP7_75t_R _0693_ (.A1(net28),
    .A2(net27),
    .B(net37),
    .Y(_0351_));
 AO21x1_ASAP7_75t_R _0694_ (.A1(_0345_),
    .A2(_0351_),
    .B(net113),
    .Y(_0352_));
 AND2x2_ASAP7_75t_R _0695_ (.A(_0350_),
    .B(_0352_),
    .Y(_0353_));
 AOI21x1_ASAP7_75t_R _0696_ (.A1(_0344_),
    .A2(_0349_),
    .B(_0353_),
    .Y(_0354_));
 INVx1_ASAP7_75t_R _0697_ (.A(_0354_),
    .Y(net153));
 AO21x1_ASAP7_75t_R _0698_ (.A1(_0004_),
    .A2(_0350_),
    .B(net113),
    .Y(_0355_));
 AND3x1_ASAP7_75t_R _0699_ (.A(_0346_),
    .B(net102),
    .C(_0004_),
    .Y(_0356_));
 AND2x4_ASAP7_75t_R _0700_ (.A(net37),
    .B(net26),
    .Y(_0357_));
 NOR2x1_ASAP7_75t_R _0701_ (.A(net28),
    .B(net27),
    .Y(_0358_));
 OA211x2_ASAP7_75t_R _0702_ (.A1(net76),
    .A2(_0356_),
    .B(_0357_),
    .C(_0358_),
    .Y(_0359_));
 AO21x1_ASAP7_75t_R _0703_ (.A1(_0351_),
    .A2(_0355_),
    .B(_0359_),
    .Y(_0360_));
 BUFx3_ASAP7_75t_R _0704_ (.A(_0360_),
    .Y(net115));
 AND2x2_ASAP7_75t_R _0705_ (.A(net76),
    .B(net102),
    .Y(_0361_));
 AO21x1_ASAP7_75t_R _0706_ (.A1(_0347_),
    .A2(net38),
    .B(_0361_),
    .Y(_0362_));
 BUFx6f_ASAP7_75t_R _0707_ (.A(_0006_),
    .Y(_0363_));
 AND3x1_ASAP7_75t_R _0708_ (.A(_0346_),
    .B(_0347_),
    .C(_0363_),
    .Y(_0364_));
 AND5x1_ASAP7_75t_R _0709_ (.A(_0346_),
    .B(net102),
    .C(_0363_),
    .D(_0358_),
    .E(_0357_),
    .Y(_0365_));
 AOI221x1_ASAP7_75t_R _0710_ (.A1(_0346_),
    .A2(_0362_),
    .B1(_0364_),
    .B2(_0344_),
    .C(_0365_),
    .Y(_0366_));
 INVx2_ASAP7_75t_R _0711_ (.A(_0366_),
    .Y(net191));
 BUFx6f_ASAP7_75t_R _0712_ (.A(rst),
    .Y(_0367_));
 INVx2_ASAP7_75t_R _0713_ (.A(_0367_),
    .Y(_0368_));
 BUFx6f_ASAP7_75t_R _0714_ (.A(_0368_),
    .Y(_0369_));
 OAI21x1_ASAP7_75t_R _0715_ (.A1(_0363_),
    .A2(net115),
    .B(_0004_),
    .Y(_0370_));
 NOR2x1_ASAP7_75t_R _0716_ (.A(_0367_),
    .B(net115),
    .Y(_0371_));
 NOR2x1_ASAP7_75t_R _0717_ (.A(_0345_),
    .B(net191),
    .Y(_0372_));
 AO32x1_ASAP7_75t_R _0718_ (.A1(_0369_),
    .A2(net153),
    .A3(_0370_),
    .B1(_0371_),
    .B2(_0372_),
    .Y(_0003_));
 OAI22x1_ASAP7_75t_R _0719_ (.A1(_0363_),
    .A2(net115),
    .B1(_0366_),
    .B2(_0004_),
    .Y(_0373_));
 NOR2x1_ASAP7_75t_R _0720_ (.A(_0345_),
    .B(_0367_),
    .Y(_0374_));
 AO32x1_ASAP7_75t_R _0721_ (.A1(_0369_),
    .A2(_0354_),
    .A3(_0373_),
    .B1(_0374_),
    .B2(net191),
    .Y(_0002_));
 INVx1_ASAP7_75t_R _0722_ (.A(_0004_),
    .Y(_0375_));
 AND2x2_ASAP7_75t_R _0723_ (.A(_0375_),
    .B(_0366_),
    .Y(_0376_));
 OAI21x1_ASAP7_75t_R _0724_ (.A1(_0345_),
    .A2(net191),
    .B(_0363_),
    .Y(_0377_));
 AO221x1_ASAP7_75t_R _0725_ (.A1(_0354_),
    .A2(_0376_),
    .B1(_0377_),
    .B2(net115),
    .C(_0367_),
    .Y(_0001_));
 OR3x1_ASAP7_75t_R _0726_ (.A(net37),
    .B(_0346_),
    .C(net75),
    .Y(_0378_));
 INVx1_ASAP7_75t_R _0727_ (.A(_0378_),
    .Y(_0000_));
 INVx1_ASAP7_75t_R _0728_ (.A(_0007_),
    .Y(net228));
 INVx1_ASAP7_75t_R _0729_ (.A(_0008_),
    .Y(net227));
 INVx1_ASAP7_75t_R _0730_ (.A(_0009_),
    .Y(net226));
 INVx1_ASAP7_75t_R _0731_ (.A(_0010_),
    .Y(net225));
 INVx1_ASAP7_75t_R _0732_ (.A(_0011_),
    .Y(net224));
 INVx1_ASAP7_75t_R _0733_ (.A(_0012_),
    .Y(net223));
 INVx1_ASAP7_75t_R _0734_ (.A(_0013_),
    .Y(net222));
 INVx1_ASAP7_75t_R _0735_ (.A(_0014_),
    .Y(net221));
 INVx1_ASAP7_75t_R _0736_ (.A(_0015_),
    .Y(net220));
 INVx1_ASAP7_75t_R _0737_ (.A(_0016_),
    .Y(net219));
 INVx1_ASAP7_75t_R _0738_ (.A(_0017_),
    .Y(net218));
 INVx1_ASAP7_75t_R _0739_ (.A(_0018_),
    .Y(net217));
 INVx1_ASAP7_75t_R _0740_ (.A(_0019_),
    .Y(net216));
 INVx1_ASAP7_75t_R _0741_ (.A(_0020_),
    .Y(net215));
 INVx1_ASAP7_75t_R _0742_ (.A(_0021_),
    .Y(net214));
 INVx1_ASAP7_75t_R _0743_ (.A(_0022_),
    .Y(net213));
 INVx1_ASAP7_75t_R _0744_ (.A(_0023_),
    .Y(net212));
 INVx1_ASAP7_75t_R _0745_ (.A(_0024_),
    .Y(net211));
 INVx1_ASAP7_75t_R _0746_ (.A(_0025_),
    .Y(net210));
 INVx1_ASAP7_75t_R _0747_ (.A(_0026_),
    .Y(net209));
 INVx1_ASAP7_75t_R _0748_ (.A(_0027_),
    .Y(net208));
 INVx1_ASAP7_75t_R _0749_ (.A(_0028_),
    .Y(net207));
 INVx1_ASAP7_75t_R _0750_ (.A(_0029_),
    .Y(net206));
 INVx1_ASAP7_75t_R _0751_ (.A(_0030_),
    .Y(net205));
 INVx1_ASAP7_75t_R _0752_ (.A(_0031_),
    .Y(net204));
 INVx1_ASAP7_75t_R _0753_ (.A(_0032_),
    .Y(net203));
 INVx1_ASAP7_75t_R _0754_ (.A(_0033_),
    .Y(net202));
 INVx1_ASAP7_75t_R _0755_ (.A(_0034_),
    .Y(net201));
 INVx1_ASAP7_75t_R _0756_ (.A(_0035_),
    .Y(net200));
 INVx1_ASAP7_75t_R _0757_ (.A(_0036_),
    .Y(net199));
 INVx1_ASAP7_75t_R _0758_ (.A(_0037_),
    .Y(net198));
 INVx1_ASAP7_75t_R _0759_ (.A(_0038_),
    .Y(net197));
 INVx1_ASAP7_75t_R _0760_ (.A(_0039_),
    .Y(net196));
 INVx1_ASAP7_75t_R _0761_ (.A(_0040_),
    .Y(net195));
 INVx1_ASAP7_75t_R _0762_ (.A(_0041_),
    .Y(net194));
 INVx1_ASAP7_75t_R _0763_ (.A(_0042_),
    .Y(net193));
 INVx1_ASAP7_75t_R _0764_ (.A(_0043_),
    .Y(net192));
 INVx1_ASAP7_75t_R _0765_ (.A(_0044_),
    .Y(net190));
 INVx1_ASAP7_75t_R _0766_ (.A(_0045_),
    .Y(net189));
 INVx1_ASAP7_75t_R _0767_ (.A(_0046_),
    .Y(net188));
 INVx1_ASAP7_75t_R _0768_ (.A(_0047_),
    .Y(net187));
 INVx1_ASAP7_75t_R _0769_ (.A(_0048_),
    .Y(net186));
 INVx1_ASAP7_75t_R _0770_ (.A(_0049_),
    .Y(net185));
 INVx1_ASAP7_75t_R _0771_ (.A(_0050_),
    .Y(net184));
 INVx1_ASAP7_75t_R _0772_ (.A(_0051_),
    .Y(net183));
 INVx1_ASAP7_75t_R _0773_ (.A(_0052_),
    .Y(net182));
 INVx1_ASAP7_75t_R _0774_ (.A(_0053_),
    .Y(net181));
 INVx1_ASAP7_75t_R _0775_ (.A(_0054_),
    .Y(net180));
 INVx1_ASAP7_75t_R _0776_ (.A(_0055_),
    .Y(net179));
 INVx1_ASAP7_75t_R _0777_ (.A(_0056_),
    .Y(net178));
 INVx1_ASAP7_75t_R _0778_ (.A(_0057_),
    .Y(net177));
 INVx1_ASAP7_75t_R _0779_ (.A(_0058_),
    .Y(net176));
 INVx1_ASAP7_75t_R _0780_ (.A(_0059_),
    .Y(net175));
 INVx1_ASAP7_75t_R _0781_ (.A(_0060_),
    .Y(net174));
 INVx1_ASAP7_75t_R _0782_ (.A(_0061_),
    .Y(net173));
 INVx1_ASAP7_75t_R _0783_ (.A(_0062_),
    .Y(net172));
 INVx1_ASAP7_75t_R _0784_ (.A(_0063_),
    .Y(net171));
 INVx1_ASAP7_75t_R _0785_ (.A(_0064_),
    .Y(net170));
 INVx1_ASAP7_75t_R _0786_ (.A(_0065_),
    .Y(net169));
 INVx1_ASAP7_75t_R _0787_ (.A(_0066_),
    .Y(net168));
 INVx1_ASAP7_75t_R _0788_ (.A(_0067_),
    .Y(net167));
 INVx1_ASAP7_75t_R _0789_ (.A(_0068_),
    .Y(net166));
 INVx1_ASAP7_75t_R _0790_ (.A(_0069_),
    .Y(net165));
 INVx1_ASAP7_75t_R _0791_ (.A(_0070_),
    .Y(net164));
 INVx1_ASAP7_75t_R _0792_ (.A(_0071_),
    .Y(net163));
 INVx1_ASAP7_75t_R _0793_ (.A(_0072_),
    .Y(net162));
 INVx1_ASAP7_75t_R _0794_ (.A(_0073_),
    .Y(net161));
 INVx1_ASAP7_75t_R _0795_ (.A(_0074_),
    .Y(net160));
 INVx1_ASAP7_75t_R _0796_ (.A(_0075_),
    .Y(net159));
 INVx1_ASAP7_75t_R _0797_ (.A(_0076_),
    .Y(net158));
 INVx1_ASAP7_75t_R _0798_ (.A(_0077_),
    .Y(net157));
 INVx1_ASAP7_75t_R _0799_ (.A(_0078_),
    .Y(net156));
 INVx1_ASAP7_75t_R _0800_ (.A(_0079_),
    .Y(net155));
 INVx1_ASAP7_75t_R _0801_ (.A(_0080_),
    .Y(net154));
 INVx1_ASAP7_75t_R _0802_ (.A(_0081_),
    .Y(net151));
 INVx1_ASAP7_75t_R _0803_ (.A(_0082_),
    .Y(net150));
 INVx1_ASAP7_75t_R _0804_ (.A(_0083_),
    .Y(net149));
 INVx1_ASAP7_75t_R _0805_ (.A(_0084_),
    .Y(net148));
 INVx1_ASAP7_75t_R _0806_ (.A(_0085_),
    .Y(net147));
 INVx1_ASAP7_75t_R _0807_ (.A(_0086_),
    .Y(net146));
 INVx1_ASAP7_75t_R _0808_ (.A(_0087_),
    .Y(net145));
 INVx1_ASAP7_75t_R _0809_ (.A(_0088_),
    .Y(net144));
 INVx1_ASAP7_75t_R _0810_ (.A(_0089_),
    .Y(net143));
 INVx1_ASAP7_75t_R _0811_ (.A(_0090_),
    .Y(net142));
 INVx1_ASAP7_75t_R _0812_ (.A(_0091_),
    .Y(net141));
 INVx1_ASAP7_75t_R _0813_ (.A(_0092_),
    .Y(net140));
 INVx1_ASAP7_75t_R _0814_ (.A(_0093_),
    .Y(net139));
 INVx1_ASAP7_75t_R _0815_ (.A(_0094_),
    .Y(net138));
 INVx1_ASAP7_75t_R _0816_ (.A(_0095_),
    .Y(net137));
 INVx1_ASAP7_75t_R _0817_ (.A(_0096_),
    .Y(net136));
 INVx1_ASAP7_75t_R _0818_ (.A(_0097_),
    .Y(net135));
 INVx1_ASAP7_75t_R _0819_ (.A(_0098_),
    .Y(net134));
 INVx1_ASAP7_75t_R _0820_ (.A(_0099_),
    .Y(net133));
 INVx1_ASAP7_75t_R _0821_ (.A(_0100_),
    .Y(net132));
 INVx1_ASAP7_75t_R _0822_ (.A(_0101_),
    .Y(net131));
 INVx1_ASAP7_75t_R _0823_ (.A(_0102_),
    .Y(net130));
 INVx1_ASAP7_75t_R _0824_ (.A(_0103_),
    .Y(net129));
 INVx1_ASAP7_75t_R _0825_ (.A(_0104_),
    .Y(net128));
 INVx1_ASAP7_75t_R _0826_ (.A(_0105_),
    .Y(net127));
 INVx1_ASAP7_75t_R _0827_ (.A(_0106_),
    .Y(net126));
 INVx1_ASAP7_75t_R _0828_ (.A(_0107_),
    .Y(net125));
 INVx1_ASAP7_75t_R _0829_ (.A(_0108_),
    .Y(net124));
 INVx1_ASAP7_75t_R _0830_ (.A(_0109_),
    .Y(net123));
 INVx1_ASAP7_75t_R _0831_ (.A(_0110_),
    .Y(net122));
 INVx1_ASAP7_75t_R _0832_ (.A(_0111_),
    .Y(net121));
 INVx1_ASAP7_75t_R _0833_ (.A(_0112_),
    .Y(net120));
 INVx1_ASAP7_75t_R _0834_ (.A(_0113_),
    .Y(net119));
 INVx1_ASAP7_75t_R _0835_ (.A(_0114_),
    .Y(net118));
 INVx1_ASAP7_75t_R _0836_ (.A(_0115_),
    .Y(net117));
 INVx1_ASAP7_75t_R _0837_ (.A(_0116_),
    .Y(net116));
 INVx1_ASAP7_75t_R _0838_ (.A(_0117_),
    .Y(net114));
 INVx1_ASAP7_75t_R _0839_ (.A(_0118_),
    .Y(net152));
 BUFx12f_ASAP7_75t_R _0840_ (.A(net38),
    .Y(_0379_));
 BUFx6f_ASAP7_75t_R _0841_ (.A(_0379_),
    .Y(_0380_));
 INVx1_ASAP7_75t_R _0842_ (.A(net75),
    .Y(_0381_));
 OR4x1_ASAP7_75t_R _0843_ (.A(net66),
    .B(net65),
    .C(_0381_),
    .D(net64),
    .Y(_0382_));
 BUFx6f_ASAP7_75t_R _0844_ (.A(_0382_),
    .Y(_0383_));
 INVx1_ASAP7_75t_R _0845_ (.A(_0363_),
    .Y(_0384_));
 AND2x6_ASAP7_75t_R _0846_ (.A(_0345_),
    .B(_0384_),
    .Y(_0385_));
 INVx1_ASAP7_75t_R _0847_ (.A(net38),
    .Y(_0386_));
 AND3x4_ASAP7_75t_R _0848_ (.A(_0346_),
    .B(_0347_),
    .C(_0386_),
    .Y(_0387_));
 OAI21x1_ASAP7_75t_R _0849_ (.A1(_0383_),
    .A2(_0385_),
    .B(_0387_),
    .Y(_0388_));
 BUFx6f_ASAP7_75t_R _0850_ (.A(_0388_),
    .Y(_0389_));
 BUFx6f_ASAP7_75t_R _0851_ (.A(_0383_),
    .Y(_0390_));
 BUFx6f_ASAP7_75t_R _0852_ (.A(_0385_),
    .Y(_0391_));
 BUFx3_ASAP7_75t_R _0853_ (.A(_0387_),
    .Y(_0392_));
 OA211x2_ASAP7_75t_R _0854_ (.A1(_0390_),
    .A2(_0391_),
    .B(_0392_),
    .C(net77),
    .Y(_0393_));
 AO21x1_ASAP7_75t_R _0855_ (.A1(net39),
    .A2(_0389_),
    .B(_0393_),
    .Y(_0394_));
 BUFx6f_ASAP7_75t_R _0856_ (.A(_0379_),
    .Y(_0395_));
 NAND2x1_ASAP7_75t_R _0857_ (.A(_0395_),
    .B(_0116_),
    .Y(_0396_));
 OA211x2_ASAP7_75t_R _0858_ (.A1(_0380_),
    .A2(_0394_),
    .B(_0396_),
    .C(_0369_),
    .Y(_0119_));
 OA211x2_ASAP7_75t_R _0859_ (.A1(_0390_),
    .A2(_0391_),
    .B(_0392_),
    .C(net78),
    .Y(_0397_));
 AO21x1_ASAP7_75t_R _0860_ (.A1(net40),
    .A2(_0389_),
    .B(_0397_),
    .Y(_0398_));
 NAND2x1_ASAP7_75t_R _0861_ (.A(_0395_),
    .B(_0115_),
    .Y(_0399_));
 OA211x2_ASAP7_75t_R _0862_ (.A1(_0380_),
    .A2(_0398_),
    .B(_0399_),
    .C(_0369_),
    .Y(_0120_));
 OA211x2_ASAP7_75t_R _0863_ (.A1(_0390_),
    .A2(_0391_),
    .B(_0392_),
    .C(net79),
    .Y(_0400_));
 AO21x1_ASAP7_75t_R _0864_ (.A1(net41),
    .A2(_0389_),
    .B(_0400_),
    .Y(_0401_));
 BUFx12f_ASAP7_75t_R _0865_ (.A(_0379_),
    .Y(_0402_));
 NAND2x1_ASAP7_75t_R _0866_ (.A(_0402_),
    .B(_0114_),
    .Y(_0403_));
 OA211x2_ASAP7_75t_R _0867_ (.A1(_0380_),
    .A2(_0401_),
    .B(_0403_),
    .C(_0369_),
    .Y(_0121_));
 OA211x2_ASAP7_75t_R _0868_ (.A1(_0390_),
    .A2(_0391_),
    .B(_0392_),
    .C(net80),
    .Y(_0404_));
 AO21x1_ASAP7_75t_R _0869_ (.A1(net42),
    .A2(_0389_),
    .B(_0404_),
    .Y(_0405_));
 NAND2x1_ASAP7_75t_R _0870_ (.A(_0402_),
    .B(_0113_),
    .Y(_0406_));
 OA211x2_ASAP7_75t_R _0871_ (.A1(_0380_),
    .A2(_0405_),
    .B(_0406_),
    .C(_0369_),
    .Y(_0122_));
 OA211x2_ASAP7_75t_R _0872_ (.A1(_0390_),
    .A2(_0391_),
    .B(_0392_),
    .C(net81),
    .Y(_0407_));
 AO21x1_ASAP7_75t_R _0873_ (.A1(net43),
    .A2(_0389_),
    .B(_0407_),
    .Y(_0408_));
 NAND2x1_ASAP7_75t_R _0874_ (.A(_0402_),
    .B(_0112_),
    .Y(_0409_));
 OA211x2_ASAP7_75t_R _0875_ (.A1(_0380_),
    .A2(_0408_),
    .B(_0409_),
    .C(_0369_),
    .Y(_0123_));
 OA211x2_ASAP7_75t_R _0876_ (.A1(_0390_),
    .A2(_0391_),
    .B(_0392_),
    .C(net82),
    .Y(_0410_));
 AO21x1_ASAP7_75t_R _0877_ (.A1(net44),
    .A2(_0389_),
    .B(_0410_),
    .Y(_0411_));
 NAND2x1_ASAP7_75t_R _0878_ (.A(_0402_),
    .B(_0111_),
    .Y(_0412_));
 OA211x2_ASAP7_75t_R _0879_ (.A1(_0380_),
    .A2(_0411_),
    .B(_0412_),
    .C(_0369_),
    .Y(_0124_));
 OA211x2_ASAP7_75t_R _0880_ (.A1(_0390_),
    .A2(_0391_),
    .B(_0392_),
    .C(net83),
    .Y(_0413_));
 AO21x1_ASAP7_75t_R _0881_ (.A1(net45),
    .A2(_0389_),
    .B(_0413_),
    .Y(_0414_));
 NAND2x1_ASAP7_75t_R _0882_ (.A(_0402_),
    .B(_0110_),
    .Y(_0415_));
 OA211x2_ASAP7_75t_R _0883_ (.A1(_0380_),
    .A2(_0414_),
    .B(_0415_),
    .C(_0369_),
    .Y(_0125_));
 OA211x2_ASAP7_75t_R _0884_ (.A1(_0390_),
    .A2(_0391_),
    .B(_0392_),
    .C(net84),
    .Y(_0416_));
 AO21x1_ASAP7_75t_R _0885_ (.A1(net46),
    .A2(_0389_),
    .B(_0416_),
    .Y(_0417_));
 NAND2x1_ASAP7_75t_R _0886_ (.A(_0402_),
    .B(_0109_),
    .Y(_0418_));
 BUFx6f_ASAP7_75t_R _0887_ (.A(_0368_),
    .Y(_0419_));
 BUFx3_ASAP7_75t_R _0888_ (.A(_0419_),
    .Y(_0420_));
 OA211x2_ASAP7_75t_R _0889_ (.A1(_0380_),
    .A2(_0417_),
    .B(_0418_),
    .C(_0420_),
    .Y(_0126_));
 OA211x2_ASAP7_75t_R _0890_ (.A1(_0390_),
    .A2(_0391_),
    .B(_0392_),
    .C(net85),
    .Y(_0421_));
 AO21x1_ASAP7_75t_R _0891_ (.A1(net47),
    .A2(_0389_),
    .B(_0421_),
    .Y(_0422_));
 NAND2x1_ASAP7_75t_R _0892_ (.A(_0402_),
    .B(_0108_),
    .Y(_0423_));
 OA211x2_ASAP7_75t_R _0893_ (.A1(_0380_),
    .A2(_0422_),
    .B(_0423_),
    .C(_0420_),
    .Y(_0127_));
 BUFx6f_ASAP7_75t_R _0894_ (.A(_0383_),
    .Y(_0424_));
 OA211x2_ASAP7_75t_R _0895_ (.A1(_0424_),
    .A2(_0391_),
    .B(_0392_),
    .C(net86),
    .Y(_0425_));
 AO21x1_ASAP7_75t_R _0896_ (.A1(net48),
    .A2(_0389_),
    .B(_0425_),
    .Y(_0426_));
 NAND2x1_ASAP7_75t_R _0897_ (.A(_0402_),
    .B(_0107_),
    .Y(_0427_));
 OA211x2_ASAP7_75t_R _0898_ (.A1(_0380_),
    .A2(_0426_),
    .B(_0427_),
    .C(_0420_),
    .Y(_0128_));
 BUFx6f_ASAP7_75t_R _0899_ (.A(_0379_),
    .Y(_0428_));
 BUFx6f_ASAP7_75t_R _0900_ (.A(_0388_),
    .Y(_0429_));
 BUFx6f_ASAP7_75t_R _0901_ (.A(_0385_),
    .Y(_0430_));
 BUFx3_ASAP7_75t_R _0902_ (.A(_0387_),
    .Y(_0431_));
 OA211x2_ASAP7_75t_R _0903_ (.A1(_0424_),
    .A2(_0430_),
    .B(_0431_),
    .C(net87),
    .Y(_0432_));
 AO21x1_ASAP7_75t_R _0904_ (.A1(net49),
    .A2(_0429_),
    .B(_0432_),
    .Y(_0433_));
 NAND2x1_ASAP7_75t_R _0905_ (.A(_0402_),
    .B(_0106_),
    .Y(_0434_));
 OA211x2_ASAP7_75t_R _0906_ (.A1(_0428_),
    .A2(_0433_),
    .B(_0434_),
    .C(_0420_),
    .Y(_0129_));
 OA211x2_ASAP7_75t_R _0907_ (.A1(_0424_),
    .A2(_0430_),
    .B(_0431_),
    .C(net88),
    .Y(_0435_));
 AO21x1_ASAP7_75t_R _0908_ (.A1(net50),
    .A2(_0429_),
    .B(_0435_),
    .Y(_0436_));
 NAND2x1_ASAP7_75t_R _0909_ (.A(_0402_),
    .B(_0105_),
    .Y(_0437_));
 OA211x2_ASAP7_75t_R _0910_ (.A1(_0428_),
    .A2(_0436_),
    .B(_0437_),
    .C(_0420_),
    .Y(_0130_));
 OA211x2_ASAP7_75t_R _0911_ (.A1(_0424_),
    .A2(_0430_),
    .B(_0431_),
    .C(net89),
    .Y(_0438_));
 AO21x1_ASAP7_75t_R _0912_ (.A1(net51),
    .A2(_0429_),
    .B(_0438_),
    .Y(_0439_));
 BUFx12f_ASAP7_75t_R _0913_ (.A(_0379_),
    .Y(_0440_));
 NAND2x1_ASAP7_75t_R _0914_ (.A(_0440_),
    .B(_0104_),
    .Y(_0441_));
 OA211x2_ASAP7_75t_R _0915_ (.A1(_0428_),
    .A2(_0439_),
    .B(_0441_),
    .C(_0420_),
    .Y(_0131_));
 OA211x2_ASAP7_75t_R _0916_ (.A1(_0424_),
    .A2(_0430_),
    .B(_0431_),
    .C(net90),
    .Y(_0442_));
 AO21x1_ASAP7_75t_R _0917_ (.A1(net52),
    .A2(_0429_),
    .B(_0442_),
    .Y(_0443_));
 NAND2x1_ASAP7_75t_R _0918_ (.A(_0440_),
    .B(_0103_),
    .Y(_0444_));
 OA211x2_ASAP7_75t_R _0919_ (.A1(_0428_),
    .A2(_0443_),
    .B(_0444_),
    .C(_0420_),
    .Y(_0132_));
 OA211x2_ASAP7_75t_R _0920_ (.A1(_0424_),
    .A2(_0430_),
    .B(_0431_),
    .C(net91),
    .Y(_0445_));
 AO21x1_ASAP7_75t_R _0921_ (.A1(net53),
    .A2(_0429_),
    .B(_0445_),
    .Y(_0446_));
 NAND2x1_ASAP7_75t_R _0922_ (.A(_0440_),
    .B(_0102_),
    .Y(_0447_));
 OA211x2_ASAP7_75t_R _0923_ (.A1(_0428_),
    .A2(_0446_),
    .B(_0447_),
    .C(_0420_),
    .Y(_0133_));
 OA211x2_ASAP7_75t_R _0924_ (.A1(_0424_),
    .A2(_0430_),
    .B(_0431_),
    .C(net92),
    .Y(_0448_));
 AO21x1_ASAP7_75t_R _0925_ (.A1(net54),
    .A2(_0429_),
    .B(_0448_),
    .Y(_0449_));
 NAND2x1_ASAP7_75t_R _0926_ (.A(_0440_),
    .B(_0101_),
    .Y(_0450_));
 OA211x2_ASAP7_75t_R _0927_ (.A1(_0428_),
    .A2(_0449_),
    .B(_0450_),
    .C(_0420_),
    .Y(_0134_));
 OA211x2_ASAP7_75t_R _0928_ (.A1(_0424_),
    .A2(_0430_),
    .B(_0431_),
    .C(net93),
    .Y(_0451_));
 AO21x1_ASAP7_75t_R _0929_ (.A1(net55),
    .A2(_0429_),
    .B(_0451_),
    .Y(_0452_));
 NAND2x1_ASAP7_75t_R _0930_ (.A(_0440_),
    .B(_0100_),
    .Y(_0453_));
 OA211x2_ASAP7_75t_R _0931_ (.A1(_0428_),
    .A2(_0452_),
    .B(_0453_),
    .C(_0420_),
    .Y(_0135_));
 OA211x2_ASAP7_75t_R _0932_ (.A1(_0424_),
    .A2(_0430_),
    .B(_0431_),
    .C(net94),
    .Y(_0454_));
 AO21x1_ASAP7_75t_R _0933_ (.A1(net56),
    .A2(_0429_),
    .B(_0454_),
    .Y(_0455_));
 NAND2x1_ASAP7_75t_R _0934_ (.A(_0440_),
    .B(_0099_),
    .Y(_0456_));
 BUFx6f_ASAP7_75t_R _0935_ (.A(_0419_),
    .Y(_0457_));
 OA211x2_ASAP7_75t_R _0936_ (.A1(_0428_),
    .A2(_0455_),
    .B(_0456_),
    .C(_0457_),
    .Y(_0136_));
 OA211x2_ASAP7_75t_R _0937_ (.A1(_0424_),
    .A2(_0430_),
    .B(_0431_),
    .C(net95),
    .Y(_0458_));
 AO21x1_ASAP7_75t_R _0938_ (.A1(net57),
    .A2(_0429_),
    .B(_0458_),
    .Y(_0459_));
 NAND2x1_ASAP7_75t_R _0939_ (.A(_0440_),
    .B(_0098_),
    .Y(_0460_));
 OA211x2_ASAP7_75t_R _0940_ (.A1(_0428_),
    .A2(_0459_),
    .B(_0460_),
    .C(_0457_),
    .Y(_0137_));
 BUFx6f_ASAP7_75t_R _0941_ (.A(_0383_),
    .Y(_0461_));
 OA211x2_ASAP7_75t_R _0942_ (.A1(_0461_),
    .A2(_0430_),
    .B(_0431_),
    .C(net96),
    .Y(_0462_));
 AO21x1_ASAP7_75t_R _0943_ (.A1(net58),
    .A2(_0429_),
    .B(_0462_),
    .Y(_0463_));
 NAND2x1_ASAP7_75t_R _0944_ (.A(_0440_),
    .B(_0097_),
    .Y(_0464_));
 OA211x2_ASAP7_75t_R _0945_ (.A1(_0428_),
    .A2(_0463_),
    .B(_0464_),
    .C(_0457_),
    .Y(_0138_));
 BUFx6f_ASAP7_75t_R _0946_ (.A(_0379_),
    .Y(_0465_));
 BUFx6f_ASAP7_75t_R _0947_ (.A(_0388_),
    .Y(_0466_));
 BUFx6f_ASAP7_75t_R _0948_ (.A(_0385_),
    .Y(_0467_));
 BUFx3_ASAP7_75t_R _0949_ (.A(_0387_),
    .Y(_0468_));
 OA211x2_ASAP7_75t_R _0950_ (.A1(_0461_),
    .A2(_0467_),
    .B(_0468_),
    .C(net97),
    .Y(_0469_));
 AO21x1_ASAP7_75t_R _0951_ (.A1(net59),
    .A2(_0466_),
    .B(_0469_),
    .Y(_0470_));
 NAND2x1_ASAP7_75t_R _0952_ (.A(_0440_),
    .B(_0096_),
    .Y(_0471_));
 OA211x2_ASAP7_75t_R _0953_ (.A1(_0465_),
    .A2(_0470_),
    .B(_0471_),
    .C(_0457_),
    .Y(_0139_));
 OA211x2_ASAP7_75t_R _0954_ (.A1(_0461_),
    .A2(_0467_),
    .B(_0468_),
    .C(net98),
    .Y(_0472_));
 AO21x1_ASAP7_75t_R _0955_ (.A1(net60),
    .A2(_0466_),
    .B(_0472_),
    .Y(_0473_));
 NAND2x1_ASAP7_75t_R _0956_ (.A(_0440_),
    .B(_0095_),
    .Y(_0474_));
 OA211x2_ASAP7_75t_R _0957_ (.A1(_0465_),
    .A2(_0473_),
    .B(_0474_),
    .C(_0457_),
    .Y(_0140_));
 OA211x2_ASAP7_75t_R _0958_ (.A1(_0461_),
    .A2(_0467_),
    .B(_0468_),
    .C(net99),
    .Y(_0475_));
 AO21x1_ASAP7_75t_R _0959_ (.A1(net61),
    .A2(_0466_),
    .B(_0475_),
    .Y(_0476_));
 BUFx12f_ASAP7_75t_R _0960_ (.A(_0379_),
    .Y(_0477_));
 NAND2x1_ASAP7_75t_R _0961_ (.A(_0477_),
    .B(_0094_),
    .Y(_0478_));
 OA211x2_ASAP7_75t_R _0962_ (.A1(_0465_),
    .A2(_0476_),
    .B(_0478_),
    .C(_0457_),
    .Y(_0141_));
 OA211x2_ASAP7_75t_R _0963_ (.A1(_0461_),
    .A2(_0467_),
    .B(_0468_),
    .C(net100),
    .Y(_0479_));
 AO21x1_ASAP7_75t_R _0964_ (.A1(net62),
    .A2(_0466_),
    .B(_0479_),
    .Y(_0480_));
 NAND2x1_ASAP7_75t_R _0965_ (.A(_0477_),
    .B(_0093_),
    .Y(_0481_));
 OA211x2_ASAP7_75t_R _0966_ (.A1(_0465_),
    .A2(_0480_),
    .B(_0481_),
    .C(_0457_),
    .Y(_0142_));
 OA211x2_ASAP7_75t_R _0967_ (.A1(_0461_),
    .A2(_0467_),
    .B(_0468_),
    .C(net101),
    .Y(_0482_));
 AO21x1_ASAP7_75t_R _0968_ (.A1(net63),
    .A2(_0466_),
    .B(_0482_),
    .Y(_0483_));
 NAND2x1_ASAP7_75t_R _0969_ (.A(_0477_),
    .B(_0092_),
    .Y(_0484_));
 OA211x2_ASAP7_75t_R _0970_ (.A1(_0465_),
    .A2(_0483_),
    .B(_0484_),
    .C(_0457_),
    .Y(_0143_));
 NAND2x1_ASAP7_75t_R _0971_ (.A(_0346_),
    .B(_0347_),
    .Y(_0485_));
 AND3x1_ASAP7_75t_R _0972_ (.A(net64),
    .B(_0386_),
    .C(_0485_),
    .Y(_0486_));
 AO21x1_ASAP7_75t_R _0973_ (.A1(_0395_),
    .A2(net141),
    .B(_0486_),
    .Y(_0487_));
 AND2x2_ASAP7_75t_R _0974_ (.A(_0369_),
    .B(_0487_),
    .Y(_0144_));
 OA211x2_ASAP7_75t_R _0975_ (.A1(_0461_),
    .A2(_0467_),
    .B(_0468_),
    .C(net103),
    .Y(_0488_));
 AO21x1_ASAP7_75t_R _0976_ (.A1(net65),
    .A2(_0466_),
    .B(_0488_),
    .Y(_0489_));
 NAND2x1_ASAP7_75t_R _0977_ (.A(_0477_),
    .B(_0090_),
    .Y(_0490_));
 OA211x2_ASAP7_75t_R _0978_ (.A1(_0465_),
    .A2(_0489_),
    .B(_0490_),
    .C(_0457_),
    .Y(_0145_));
 OA211x2_ASAP7_75t_R _0979_ (.A1(_0461_),
    .A2(_0467_),
    .B(_0468_),
    .C(net104),
    .Y(_0491_));
 AO21x1_ASAP7_75t_R _0980_ (.A1(net66),
    .A2(_0466_),
    .B(_0491_),
    .Y(_0492_));
 NAND2x1_ASAP7_75t_R _0981_ (.A(_0477_),
    .B(_0089_),
    .Y(_0493_));
 OA211x2_ASAP7_75t_R _0982_ (.A1(_0465_),
    .A2(_0492_),
    .B(_0493_),
    .C(_0457_),
    .Y(_0146_));
 OA211x2_ASAP7_75t_R _0983_ (.A1(_0461_),
    .A2(_0467_),
    .B(_0468_),
    .C(net105),
    .Y(_0494_));
 AO21x1_ASAP7_75t_R _0984_ (.A1(net67),
    .A2(_0466_),
    .B(_0494_),
    .Y(_0495_));
 NAND2x1_ASAP7_75t_R _0985_ (.A(_0477_),
    .B(_0088_),
    .Y(_0496_));
 BUFx6f_ASAP7_75t_R _0986_ (.A(_0419_),
    .Y(_0497_));
 OA211x2_ASAP7_75t_R _0987_ (.A1(_0465_),
    .A2(_0495_),
    .B(_0496_),
    .C(_0497_),
    .Y(_0147_));
 OA211x2_ASAP7_75t_R _0988_ (.A1(_0461_),
    .A2(_0467_),
    .B(_0468_),
    .C(net106),
    .Y(_0498_));
 AO21x1_ASAP7_75t_R _0989_ (.A1(net68),
    .A2(_0466_),
    .B(_0498_),
    .Y(_0499_));
 NAND2x1_ASAP7_75t_R _0990_ (.A(_0477_),
    .B(_0087_),
    .Y(_0500_));
 OA211x2_ASAP7_75t_R _0991_ (.A1(_0465_),
    .A2(_0499_),
    .B(_0500_),
    .C(_0497_),
    .Y(_0148_));
 OA211x2_ASAP7_75t_R _0992_ (.A1(_0383_),
    .A2(_0467_),
    .B(_0468_),
    .C(net107),
    .Y(_0501_));
 AO21x1_ASAP7_75t_R _0993_ (.A1(net69),
    .A2(_0466_),
    .B(_0501_),
    .Y(_0502_));
 NAND2x1_ASAP7_75t_R _0994_ (.A(_0477_),
    .B(_0086_),
    .Y(_0503_));
 OA211x2_ASAP7_75t_R _0995_ (.A1(_0465_),
    .A2(_0502_),
    .B(_0503_),
    .C(_0497_),
    .Y(_0149_));
 OA211x2_ASAP7_75t_R _0996_ (.A1(_0383_),
    .A2(_0385_),
    .B(_0387_),
    .C(net108),
    .Y(_0504_));
 AO21x1_ASAP7_75t_R _0997_ (.A1(net70),
    .A2(_0388_),
    .B(_0504_),
    .Y(_0505_));
 NAND2x1_ASAP7_75t_R _0998_ (.A(_0477_),
    .B(_0085_),
    .Y(_0506_));
 OA211x2_ASAP7_75t_R _0999_ (.A1(_0395_),
    .A2(_0505_),
    .B(_0506_),
    .C(_0497_),
    .Y(_0150_));
 OA211x2_ASAP7_75t_R _1000_ (.A1(_0383_),
    .A2(_0385_),
    .B(_0387_),
    .C(net109),
    .Y(_0507_));
 AO21x1_ASAP7_75t_R _1001_ (.A1(net71),
    .A2(_0388_),
    .B(_0507_),
    .Y(_0508_));
 NAND2x1_ASAP7_75t_R _1002_ (.A(_0477_),
    .B(_0084_),
    .Y(_0509_));
 OA211x2_ASAP7_75t_R _1003_ (.A1(_0395_),
    .A2(_0508_),
    .B(_0509_),
    .C(_0497_),
    .Y(_0151_));
 OA211x2_ASAP7_75t_R _1004_ (.A1(_0383_),
    .A2(_0385_),
    .B(_0387_),
    .C(net110),
    .Y(_0510_));
 AO21x1_ASAP7_75t_R _1005_ (.A1(net72),
    .A2(_0388_),
    .B(_0510_),
    .Y(_0511_));
 NAND2x1_ASAP7_75t_R _1006_ (.A(_0379_),
    .B(_0083_),
    .Y(_0512_));
 OA211x2_ASAP7_75t_R _1007_ (.A1(_0395_),
    .A2(_0511_),
    .B(_0512_),
    .C(_0497_),
    .Y(_0152_));
 OA211x2_ASAP7_75t_R _1008_ (.A1(_0383_),
    .A2(_0385_),
    .B(_0387_),
    .C(net111),
    .Y(_0513_));
 AO21x1_ASAP7_75t_R _1009_ (.A1(net73),
    .A2(_0388_),
    .B(_0513_),
    .Y(_0514_));
 NAND2x1_ASAP7_75t_R _1010_ (.A(_0379_),
    .B(_0082_),
    .Y(_0515_));
 OA211x2_ASAP7_75t_R _1011_ (.A1(_0395_),
    .A2(_0514_),
    .B(_0515_),
    .C(_0497_),
    .Y(_0153_));
 OA211x2_ASAP7_75t_R _1012_ (.A1(_0383_),
    .A2(_0385_),
    .B(_0387_),
    .C(net112),
    .Y(_0516_));
 AO21x1_ASAP7_75t_R _1013_ (.A1(net74),
    .A2(_0388_),
    .B(_0516_),
    .Y(_0517_));
 NAND2x1_ASAP7_75t_R _1014_ (.A(_0379_),
    .B(_0081_),
    .Y(_0518_));
 OA211x2_ASAP7_75t_R _1015_ (.A1(_0395_),
    .A2(_0517_),
    .B(_0518_),
    .C(_0497_),
    .Y(_0154_));
 NAND2x1_ASAP7_75t_R _1016_ (.A(_0395_),
    .B(net152),
    .Y(_0519_));
 AND3x1_ASAP7_75t_R _1017_ (.A(_0345_),
    .B(_0344_),
    .C(_0348_),
    .Y(_0520_));
 AO221x1_ASAP7_75t_R _1018_ (.A1(_0390_),
    .A2(_0485_),
    .B1(_0520_),
    .B2(_0363_),
    .C(_0395_),
    .Y(_0521_));
 AOI21x1_ASAP7_75t_R _1019_ (.A1(_0519_),
    .A2(_0521_),
    .B(_0367_),
    .Y(_0155_));
 BUFx12f_ASAP7_75t_R _1020_ (.A(net76),
    .Y(_0522_));
 BUFx6f_ASAP7_75t_R _1021_ (.A(_0522_),
    .Y(_0523_));
 OA211x2_ASAP7_75t_R _1022_ (.A1(_0375_),
    .A2(_0363_),
    .B(_0358_),
    .C(_0357_),
    .Y(_0524_));
 BUFx6f_ASAP7_75t_R _1023_ (.A(_0524_),
    .Y(_0525_));
 NAND2x1_ASAP7_75t_R _1024_ (.A(_0346_),
    .B(net102),
    .Y(_0526_));
 OR2x2_ASAP7_75t_R _1025_ (.A(net76),
    .B(_0526_),
    .Y(_0527_));
 BUFx6f_ASAP7_75t_R _1026_ (.A(_0527_),
    .Y(_0528_));
 NOR2x2_ASAP7_75t_R _1027_ (.A(_0525_),
    .B(_0528_),
    .Y(_0529_));
 BUFx6f_ASAP7_75t_R _1028_ (.A(_0529_),
    .Y(_0530_));
 BUFx6f_ASAP7_75t_R _1029_ (.A(_0525_),
    .Y(_0531_));
 BUFx6f_ASAP7_75t_R _1030_ (.A(_0528_),
    .Y(_0532_));
 OA21x2_ASAP7_75t_R _1031_ (.A1(_0531_),
    .A2(_0532_),
    .B(net1),
    .Y(_0533_));
 AO21x1_ASAP7_75t_R _1032_ (.A1(net77),
    .A2(_0530_),
    .B(_0533_),
    .Y(_0534_));
 BUFx6f_ASAP7_75t_R _1033_ (.A(net76),
    .Y(_0535_));
 NAND2x1_ASAP7_75t_R _1034_ (.A(_0535_),
    .B(_0080_),
    .Y(_0536_));
 OA211x2_ASAP7_75t_R _1035_ (.A1(_0523_),
    .A2(_0534_),
    .B(_0536_),
    .C(_0497_),
    .Y(_0156_));
 OA21x2_ASAP7_75t_R _1036_ (.A1(_0531_),
    .A2(_0532_),
    .B(net2),
    .Y(_0537_));
 AO21x1_ASAP7_75t_R _1037_ (.A1(net78),
    .A2(_0530_),
    .B(_0537_),
    .Y(_0538_));
 NAND2x1_ASAP7_75t_R _1038_ (.A(_0535_),
    .B(_0079_),
    .Y(_0539_));
 OA211x2_ASAP7_75t_R _1039_ (.A1(_0523_),
    .A2(_0538_),
    .B(_0539_),
    .C(_0497_),
    .Y(_0157_));
 OA21x2_ASAP7_75t_R _1040_ (.A1(_0531_),
    .A2(_0532_),
    .B(net3),
    .Y(_0540_));
 AO21x1_ASAP7_75t_R _1041_ (.A1(net79),
    .A2(_0530_),
    .B(_0540_),
    .Y(_0541_));
 BUFx12f_ASAP7_75t_R _1042_ (.A(_0522_),
    .Y(_0542_));
 NAND2x1_ASAP7_75t_R _1043_ (.A(_0542_),
    .B(_0078_),
    .Y(_0543_));
 BUFx3_ASAP7_75t_R _1044_ (.A(_0419_),
    .Y(_0544_));
 OA211x2_ASAP7_75t_R _1045_ (.A1(_0523_),
    .A2(_0541_),
    .B(_0543_),
    .C(_0544_),
    .Y(_0158_));
 OA21x2_ASAP7_75t_R _1046_ (.A1(_0531_),
    .A2(_0532_),
    .B(net4),
    .Y(_0545_));
 AO21x1_ASAP7_75t_R _1047_ (.A1(net80),
    .A2(_0530_),
    .B(_0545_),
    .Y(_0546_));
 NAND2x1_ASAP7_75t_R _1048_ (.A(_0542_),
    .B(_0077_),
    .Y(_0547_));
 OA211x2_ASAP7_75t_R _1049_ (.A1(_0523_),
    .A2(_0546_),
    .B(_0547_),
    .C(_0544_),
    .Y(_0159_));
 OA21x2_ASAP7_75t_R _1050_ (.A1(_0531_),
    .A2(_0532_),
    .B(net5),
    .Y(_0548_));
 AO21x1_ASAP7_75t_R _1051_ (.A1(net81),
    .A2(_0530_),
    .B(_0548_),
    .Y(_0549_));
 NAND2x1_ASAP7_75t_R _1052_ (.A(_0542_),
    .B(_0076_),
    .Y(_0550_));
 OA211x2_ASAP7_75t_R _1053_ (.A1(_0523_),
    .A2(_0549_),
    .B(_0550_),
    .C(_0544_),
    .Y(_0160_));
 OA21x2_ASAP7_75t_R _1054_ (.A1(_0531_),
    .A2(_0532_),
    .B(net6),
    .Y(_0551_));
 AO21x1_ASAP7_75t_R _1055_ (.A1(net82),
    .A2(_0530_),
    .B(_0551_),
    .Y(_0552_));
 NAND2x1_ASAP7_75t_R _1056_ (.A(_0542_),
    .B(_0075_),
    .Y(_0553_));
 OA211x2_ASAP7_75t_R _1057_ (.A1(_0523_),
    .A2(_0552_),
    .B(_0553_),
    .C(_0544_),
    .Y(_0161_));
 OA21x2_ASAP7_75t_R _1058_ (.A1(_0531_),
    .A2(_0532_),
    .B(net7),
    .Y(_0554_));
 AO21x1_ASAP7_75t_R _1059_ (.A1(net83),
    .A2(_0530_),
    .B(_0554_),
    .Y(_0555_));
 NAND2x1_ASAP7_75t_R _1060_ (.A(_0542_),
    .B(_0074_),
    .Y(_0556_));
 OA211x2_ASAP7_75t_R _1061_ (.A1(_0523_),
    .A2(_0555_),
    .B(_0556_),
    .C(_0544_),
    .Y(_0162_));
 OA21x2_ASAP7_75t_R _1062_ (.A1(_0531_),
    .A2(_0532_),
    .B(net8),
    .Y(_0557_));
 AO21x1_ASAP7_75t_R _1063_ (.A1(net84),
    .A2(_0530_),
    .B(_0557_),
    .Y(_0558_));
 NAND2x1_ASAP7_75t_R _1064_ (.A(_0542_),
    .B(_0073_),
    .Y(_0559_));
 OA211x2_ASAP7_75t_R _1065_ (.A1(_0523_),
    .A2(_0558_),
    .B(_0559_),
    .C(_0544_),
    .Y(_0163_));
 OA21x2_ASAP7_75t_R _1066_ (.A1(_0531_),
    .A2(_0532_),
    .B(net9),
    .Y(_0560_));
 AO21x1_ASAP7_75t_R _1067_ (.A1(net85),
    .A2(_0530_),
    .B(_0560_),
    .Y(_0561_));
 NAND2x1_ASAP7_75t_R _1068_ (.A(_0542_),
    .B(_0072_),
    .Y(_0562_));
 OA211x2_ASAP7_75t_R _1069_ (.A1(_0523_),
    .A2(_0561_),
    .B(_0562_),
    .C(_0544_),
    .Y(_0164_));
 OA21x2_ASAP7_75t_R _1070_ (.A1(_0531_),
    .A2(_0532_),
    .B(net10),
    .Y(_0563_));
 AO21x1_ASAP7_75t_R _1071_ (.A1(net86),
    .A2(_0530_),
    .B(_0563_),
    .Y(_0564_));
 NAND2x1_ASAP7_75t_R _1072_ (.A(_0542_),
    .B(_0071_),
    .Y(_0565_));
 OA211x2_ASAP7_75t_R _1073_ (.A1(_0523_),
    .A2(_0564_),
    .B(_0565_),
    .C(_0544_),
    .Y(_0165_));
 BUFx6f_ASAP7_75t_R _1074_ (.A(_0522_),
    .Y(_0566_));
 BUFx6f_ASAP7_75t_R _1075_ (.A(_0529_),
    .Y(_0567_));
 BUFx6f_ASAP7_75t_R _1076_ (.A(_0525_),
    .Y(_0568_));
 BUFx6f_ASAP7_75t_R _1077_ (.A(_0528_),
    .Y(_0569_));
 OA21x2_ASAP7_75t_R _1078_ (.A1(_0568_),
    .A2(_0569_),
    .B(net11),
    .Y(_0570_));
 AO21x1_ASAP7_75t_R _1079_ (.A1(net87),
    .A2(_0567_),
    .B(_0570_),
    .Y(_0571_));
 NAND2x1_ASAP7_75t_R _1080_ (.A(_0542_),
    .B(_0070_),
    .Y(_0572_));
 OA211x2_ASAP7_75t_R _1081_ (.A1(_0566_),
    .A2(_0571_),
    .B(_0572_),
    .C(_0544_),
    .Y(_0166_));
 OA21x2_ASAP7_75t_R _1082_ (.A1(_0568_),
    .A2(_0569_),
    .B(net12),
    .Y(_0573_));
 AO21x1_ASAP7_75t_R _1083_ (.A1(net88),
    .A2(_0567_),
    .B(_0573_),
    .Y(_0574_));
 NAND2x1_ASAP7_75t_R _1084_ (.A(_0542_),
    .B(_0069_),
    .Y(_0575_));
 OA211x2_ASAP7_75t_R _1085_ (.A1(_0566_),
    .A2(_0574_),
    .B(_0575_),
    .C(_0544_),
    .Y(_0167_));
 OA21x2_ASAP7_75t_R _1086_ (.A1(_0568_),
    .A2(_0569_),
    .B(net13),
    .Y(_0576_));
 AO21x1_ASAP7_75t_R _1087_ (.A1(net89),
    .A2(_0567_),
    .B(_0576_),
    .Y(_0577_));
 BUFx12f_ASAP7_75t_R _1088_ (.A(_0522_),
    .Y(_0578_));
 NAND2x1_ASAP7_75t_R _1089_ (.A(_0578_),
    .B(_0068_),
    .Y(_0579_));
 BUFx3_ASAP7_75t_R _1090_ (.A(_0419_),
    .Y(_0580_));
 OA211x2_ASAP7_75t_R _1091_ (.A1(_0566_),
    .A2(_0577_),
    .B(_0579_),
    .C(_0580_),
    .Y(_0168_));
 OA21x2_ASAP7_75t_R _1092_ (.A1(_0568_),
    .A2(_0569_),
    .B(net14),
    .Y(_0581_));
 AO21x1_ASAP7_75t_R _1093_ (.A1(net90),
    .A2(_0567_),
    .B(_0581_),
    .Y(_0582_));
 NAND2x1_ASAP7_75t_R _1094_ (.A(_0578_),
    .B(_0067_),
    .Y(_0583_));
 OA211x2_ASAP7_75t_R _1095_ (.A1(_0566_),
    .A2(_0582_),
    .B(_0583_),
    .C(_0580_),
    .Y(_0169_));
 OA21x2_ASAP7_75t_R _1096_ (.A1(_0568_),
    .A2(_0569_),
    .B(net15),
    .Y(_0584_));
 AO21x1_ASAP7_75t_R _1097_ (.A1(net91),
    .A2(_0567_),
    .B(_0584_),
    .Y(_0585_));
 NAND2x1_ASAP7_75t_R _1098_ (.A(_0578_),
    .B(_0066_),
    .Y(_0586_));
 OA211x2_ASAP7_75t_R _1099_ (.A1(_0566_),
    .A2(_0585_),
    .B(_0586_),
    .C(_0580_),
    .Y(_0170_));
 OA21x2_ASAP7_75t_R _1100_ (.A1(_0568_),
    .A2(_0569_),
    .B(net16),
    .Y(_0587_));
 AO21x1_ASAP7_75t_R _1101_ (.A1(net92),
    .A2(_0567_),
    .B(_0587_),
    .Y(_0588_));
 NAND2x1_ASAP7_75t_R _1102_ (.A(_0578_),
    .B(_0065_),
    .Y(_0589_));
 OA211x2_ASAP7_75t_R _1103_ (.A1(_0566_),
    .A2(_0588_),
    .B(_0589_),
    .C(_0580_),
    .Y(_0171_));
 OA21x2_ASAP7_75t_R _1104_ (.A1(_0568_),
    .A2(_0569_),
    .B(net17),
    .Y(_0590_));
 AO21x1_ASAP7_75t_R _1105_ (.A1(net93),
    .A2(_0567_),
    .B(_0590_),
    .Y(_0591_));
 NAND2x1_ASAP7_75t_R _1106_ (.A(_0578_),
    .B(_0064_),
    .Y(_0592_));
 OA211x2_ASAP7_75t_R _1107_ (.A1(_0566_),
    .A2(_0591_),
    .B(_0592_),
    .C(_0580_),
    .Y(_0172_));
 OA21x2_ASAP7_75t_R _1108_ (.A1(_0568_),
    .A2(_0569_),
    .B(net18),
    .Y(_0593_));
 AO21x1_ASAP7_75t_R _1109_ (.A1(net94),
    .A2(_0567_),
    .B(_0593_),
    .Y(_0594_));
 NAND2x1_ASAP7_75t_R _1110_ (.A(_0578_),
    .B(_0063_),
    .Y(_0595_));
 OA211x2_ASAP7_75t_R _1111_ (.A1(_0566_),
    .A2(_0594_),
    .B(_0595_),
    .C(_0580_),
    .Y(_0173_));
 OA21x2_ASAP7_75t_R _1112_ (.A1(_0568_),
    .A2(_0569_),
    .B(net19),
    .Y(_0596_));
 AO21x1_ASAP7_75t_R _1113_ (.A1(net95),
    .A2(_0567_),
    .B(_0596_),
    .Y(_0597_));
 NAND2x1_ASAP7_75t_R _1114_ (.A(_0578_),
    .B(_0062_),
    .Y(_0598_));
 OA211x2_ASAP7_75t_R _1115_ (.A1(_0566_),
    .A2(_0597_),
    .B(_0598_),
    .C(_0580_),
    .Y(_0174_));
 OA21x2_ASAP7_75t_R _1116_ (.A1(_0568_),
    .A2(_0569_),
    .B(net20),
    .Y(_0599_));
 AO21x1_ASAP7_75t_R _1117_ (.A1(net96),
    .A2(_0567_),
    .B(_0599_),
    .Y(_0600_));
 NAND2x1_ASAP7_75t_R _1118_ (.A(_0578_),
    .B(_0061_),
    .Y(_0601_));
 OA211x2_ASAP7_75t_R _1119_ (.A1(_0566_),
    .A2(_0600_),
    .B(_0601_),
    .C(_0580_),
    .Y(_0175_));
 BUFx6f_ASAP7_75t_R _1120_ (.A(_0522_),
    .Y(_0602_));
 BUFx6f_ASAP7_75t_R _1121_ (.A(_0529_),
    .Y(_0603_));
 BUFx6f_ASAP7_75t_R _1122_ (.A(_0525_),
    .Y(_0604_));
 BUFx6f_ASAP7_75t_R _1123_ (.A(_0528_),
    .Y(_0605_));
 OA21x2_ASAP7_75t_R _1124_ (.A1(_0604_),
    .A2(_0605_),
    .B(net21),
    .Y(_0606_));
 AO21x1_ASAP7_75t_R _1125_ (.A1(net97),
    .A2(_0603_),
    .B(_0606_),
    .Y(_0607_));
 NAND2x1_ASAP7_75t_R _1126_ (.A(_0578_),
    .B(_0060_),
    .Y(_0608_));
 OA211x2_ASAP7_75t_R _1127_ (.A1(_0602_),
    .A2(_0607_),
    .B(_0608_),
    .C(_0580_),
    .Y(_0176_));
 OA21x2_ASAP7_75t_R _1128_ (.A1(_0604_),
    .A2(_0605_),
    .B(net22),
    .Y(_0609_));
 AO21x1_ASAP7_75t_R _1129_ (.A1(net98),
    .A2(_0603_),
    .B(_0609_),
    .Y(_0610_));
 NAND2x1_ASAP7_75t_R _1130_ (.A(_0578_),
    .B(_0059_),
    .Y(_0611_));
 OA211x2_ASAP7_75t_R _1131_ (.A1(_0602_),
    .A2(_0610_),
    .B(_0611_),
    .C(_0580_),
    .Y(_0177_));
 OA21x2_ASAP7_75t_R _1132_ (.A1(_0604_),
    .A2(_0605_),
    .B(net23),
    .Y(_0612_));
 AO21x1_ASAP7_75t_R _1133_ (.A1(net99),
    .A2(_0603_),
    .B(_0612_),
    .Y(_0613_));
 BUFx12f_ASAP7_75t_R _1134_ (.A(_0522_),
    .Y(_0614_));
 NAND2x1_ASAP7_75t_R _1135_ (.A(_0614_),
    .B(_0058_),
    .Y(_0615_));
 BUFx6f_ASAP7_75t_R _1136_ (.A(_0419_),
    .Y(_0616_));
 OA211x2_ASAP7_75t_R _1137_ (.A1(_0602_),
    .A2(_0613_),
    .B(_0615_),
    .C(_0616_),
    .Y(_0178_));
 OA21x2_ASAP7_75t_R _1138_ (.A1(_0604_),
    .A2(_0605_),
    .B(net24),
    .Y(_0617_));
 AO21x1_ASAP7_75t_R _1139_ (.A1(net100),
    .A2(_0603_),
    .B(_0617_),
    .Y(_0618_));
 NAND2x1_ASAP7_75t_R _1140_ (.A(_0614_),
    .B(_0057_),
    .Y(_0619_));
 OA211x2_ASAP7_75t_R _1141_ (.A1(_0602_),
    .A2(_0618_),
    .B(_0619_),
    .C(_0616_),
    .Y(_0179_));
 OA21x2_ASAP7_75t_R _1142_ (.A1(_0604_),
    .A2(_0605_),
    .B(net25),
    .Y(_0620_));
 AO21x1_ASAP7_75t_R _1143_ (.A1(net101),
    .A2(_0603_),
    .B(_0620_),
    .Y(_0621_));
 NAND2x1_ASAP7_75t_R _1144_ (.A(_0614_),
    .B(_0056_),
    .Y(_0622_));
 OA211x2_ASAP7_75t_R _1145_ (.A1(_0602_),
    .A2(_0621_),
    .B(_0622_),
    .C(_0616_),
    .Y(_0180_));
 INVx1_ASAP7_75t_R _1146_ (.A(_0535_),
    .Y(_0623_));
 OR3x1_ASAP7_75t_R _1147_ (.A(net26),
    .B(_0522_),
    .C(_0529_),
    .Y(_0624_));
 OA211x2_ASAP7_75t_R _1148_ (.A1(_0623_),
    .A2(net179),
    .B(_0624_),
    .C(_0616_),
    .Y(_0181_));
 OA21x2_ASAP7_75t_R _1149_ (.A1(_0604_),
    .A2(_0605_),
    .B(net27),
    .Y(_0625_));
 AO21x1_ASAP7_75t_R _1150_ (.A1(net103),
    .A2(_0603_),
    .B(_0625_),
    .Y(_0626_));
 NAND2x1_ASAP7_75t_R _1151_ (.A(_0614_),
    .B(_0054_),
    .Y(_0627_));
 OA211x2_ASAP7_75t_R _1152_ (.A1(_0602_),
    .A2(_0626_),
    .B(_0627_),
    .C(_0616_),
    .Y(_0182_));
 OA21x2_ASAP7_75t_R _1153_ (.A1(_0604_),
    .A2(_0605_),
    .B(net28),
    .Y(_0628_));
 AO21x1_ASAP7_75t_R _1154_ (.A1(net104),
    .A2(_0603_),
    .B(_0628_),
    .Y(_0629_));
 NAND2x1_ASAP7_75t_R _1155_ (.A(_0614_),
    .B(_0053_),
    .Y(_0630_));
 OA211x2_ASAP7_75t_R _1156_ (.A1(_0602_),
    .A2(_0629_),
    .B(_0630_),
    .C(_0616_),
    .Y(_0183_));
 OA21x2_ASAP7_75t_R _1157_ (.A1(_0604_),
    .A2(_0605_),
    .B(net29),
    .Y(_0631_));
 AO21x1_ASAP7_75t_R _1158_ (.A1(net105),
    .A2(_0603_),
    .B(_0631_),
    .Y(_0632_));
 NAND2x1_ASAP7_75t_R _1159_ (.A(_0614_),
    .B(_0052_),
    .Y(_0633_));
 OA211x2_ASAP7_75t_R _1160_ (.A1(_0602_),
    .A2(_0632_),
    .B(_0633_),
    .C(_0616_),
    .Y(_0184_));
 OA21x2_ASAP7_75t_R _1161_ (.A1(_0604_),
    .A2(_0605_),
    .B(net30),
    .Y(_0634_));
 AO21x1_ASAP7_75t_R _1162_ (.A1(net106),
    .A2(_0603_),
    .B(_0634_),
    .Y(_0635_));
 NAND2x1_ASAP7_75t_R _1163_ (.A(_0614_),
    .B(_0051_),
    .Y(_0636_));
 OA211x2_ASAP7_75t_R _1164_ (.A1(_0602_),
    .A2(_0635_),
    .B(_0636_),
    .C(_0616_),
    .Y(_0185_));
 OA21x2_ASAP7_75t_R _1165_ (.A1(_0604_),
    .A2(_0605_),
    .B(net31),
    .Y(_0637_));
 AO21x1_ASAP7_75t_R _1166_ (.A1(net107),
    .A2(_0603_),
    .B(_0637_),
    .Y(_0638_));
 NAND2x1_ASAP7_75t_R _1167_ (.A(_0614_),
    .B(_0050_),
    .Y(_0639_));
 OA211x2_ASAP7_75t_R _1168_ (.A1(_0602_),
    .A2(_0638_),
    .B(_0639_),
    .C(_0616_),
    .Y(_0186_));
 OA21x2_ASAP7_75t_R _1169_ (.A1(_0525_),
    .A2(_0528_),
    .B(net32),
    .Y(_0640_));
 AO21x1_ASAP7_75t_R _1170_ (.A1(net108),
    .A2(_0529_),
    .B(_0640_),
    .Y(_0641_));
 NAND2x1_ASAP7_75t_R _1171_ (.A(_0614_),
    .B(_0049_),
    .Y(_0642_));
 OA211x2_ASAP7_75t_R _1172_ (.A1(_0535_),
    .A2(_0641_),
    .B(_0642_),
    .C(_0616_),
    .Y(_0187_));
 OA21x2_ASAP7_75t_R _1173_ (.A1(_0525_),
    .A2(_0528_),
    .B(net33),
    .Y(_0643_));
 AO21x1_ASAP7_75t_R _1174_ (.A1(net109),
    .A2(_0529_),
    .B(_0643_),
    .Y(_0644_));
 NAND2x1_ASAP7_75t_R _1175_ (.A(_0614_),
    .B(_0048_),
    .Y(_0645_));
 BUFx3_ASAP7_75t_R _1176_ (.A(_0419_),
    .Y(_0646_));
 OA211x2_ASAP7_75t_R _1177_ (.A1(_0535_),
    .A2(_0644_),
    .B(_0645_),
    .C(_0646_),
    .Y(_0188_));
 OA21x2_ASAP7_75t_R _1178_ (.A1(_0525_),
    .A2(_0528_),
    .B(net34),
    .Y(_0647_));
 AO21x1_ASAP7_75t_R _1179_ (.A1(net110),
    .A2(_0529_),
    .B(_0647_),
    .Y(_0648_));
 NAND2x1_ASAP7_75t_R _1180_ (.A(_0522_),
    .B(_0047_),
    .Y(_0649_));
 OA211x2_ASAP7_75t_R _1181_ (.A1(_0535_),
    .A2(_0648_),
    .B(_0649_),
    .C(_0646_),
    .Y(_0189_));
 OA21x2_ASAP7_75t_R _1182_ (.A1(_0525_),
    .A2(_0528_),
    .B(net35),
    .Y(_0650_));
 AO21x1_ASAP7_75t_R _1183_ (.A1(net111),
    .A2(_0529_),
    .B(_0650_),
    .Y(_0651_));
 NAND2x1_ASAP7_75t_R _1184_ (.A(_0522_),
    .B(_0046_),
    .Y(_0652_));
 OA211x2_ASAP7_75t_R _1185_ (.A1(_0535_),
    .A2(_0651_),
    .B(_0652_),
    .C(_0646_),
    .Y(_0190_));
 OA21x2_ASAP7_75t_R _1186_ (.A1(_0525_),
    .A2(_0528_),
    .B(net36),
    .Y(_0653_));
 AO21x1_ASAP7_75t_R _1187_ (.A1(net112),
    .A2(_0529_),
    .B(_0653_),
    .Y(_0654_));
 NAND2x1_ASAP7_75t_R _1188_ (.A(_0522_),
    .B(_0045_),
    .Y(_0655_));
 OA211x2_ASAP7_75t_R _1189_ (.A1(_0535_),
    .A2(_0654_),
    .B(_0655_),
    .C(_0646_),
    .Y(_0191_));
 NAND2x1_ASAP7_75t_R _1190_ (.A(_0535_),
    .B(net190),
    .Y(_0656_));
 NAND2x1_ASAP7_75t_R _1191_ (.A(_0358_),
    .B(_0357_),
    .Y(_0657_));
 AND3x1_ASAP7_75t_R _1192_ (.A(_0363_),
    .B(_0358_),
    .C(_0357_),
    .Y(_0658_));
 AO221x1_ASAP7_75t_R _1193_ (.A1(_0657_),
    .A2(_0526_),
    .B1(_0356_),
    .B2(_0658_),
    .C(_0535_),
    .Y(_0659_));
 AOI21x1_ASAP7_75t_R _1194_ (.A1(_0656_),
    .A2(_0659_),
    .B(_0367_),
    .Y(_0192_));
 BUFx12f_ASAP7_75t_R _1195_ (.A(net113),
    .Y(_0660_));
 BUFx6f_ASAP7_75t_R _1196_ (.A(_0660_),
    .Y(_0661_));
 OAI21x1_ASAP7_75t_R _1197_ (.A1(_0375_),
    .A2(_0345_),
    .B(_0351_),
    .Y(_0662_));
 INVx1_ASAP7_75t_R _1198_ (.A(net113),
    .Y(_0663_));
 AND2x6_ASAP7_75t_R _1199_ (.A(_0663_),
    .B(_0350_),
    .Y(_0664_));
 NAND2x2_ASAP7_75t_R _1200_ (.A(_0662_),
    .B(_0664_),
    .Y(_0665_));
 BUFx6f_ASAP7_75t_R _1201_ (.A(_0665_),
    .Y(_0666_));
 BUFx6f_ASAP7_75t_R _1202_ (.A(_0662_),
    .Y(_0667_));
 BUFx6f_ASAP7_75t_R _1203_ (.A(_0664_),
    .Y(_0668_));
 AND3x1_ASAP7_75t_R _1204_ (.A(net39),
    .B(_0667_),
    .C(_0668_),
    .Y(_0669_));
 AO21x1_ASAP7_75t_R _1205_ (.A1(net1),
    .A2(_0666_),
    .B(_0669_),
    .Y(_0670_));
 BUFx6f_ASAP7_75t_R _1206_ (.A(_0660_),
    .Y(_0671_));
 NAND2x1_ASAP7_75t_R _1207_ (.A(_0671_),
    .B(_0043_),
    .Y(_0672_));
 OA211x2_ASAP7_75t_R _1208_ (.A1(_0661_),
    .A2(_0670_),
    .B(_0672_),
    .C(_0646_),
    .Y(_0193_));
 AND3x1_ASAP7_75t_R _1209_ (.A(net40),
    .B(_0667_),
    .C(_0668_),
    .Y(_0673_));
 AO21x1_ASAP7_75t_R _1210_ (.A1(net2),
    .A2(_0666_),
    .B(_0673_),
    .Y(_0674_));
 NAND2x1_ASAP7_75t_R _1211_ (.A(_0671_),
    .B(_0042_),
    .Y(_0675_));
 OA211x2_ASAP7_75t_R _1212_ (.A1(_0661_),
    .A2(_0674_),
    .B(_0675_),
    .C(_0646_),
    .Y(_0194_));
 AND3x1_ASAP7_75t_R _1213_ (.A(net41),
    .B(_0667_),
    .C(_0668_),
    .Y(_0676_));
 AO21x1_ASAP7_75t_R _1214_ (.A1(net3),
    .A2(_0666_),
    .B(_0676_),
    .Y(_0677_));
 NAND2x1_ASAP7_75t_R _1215_ (.A(_0671_),
    .B(_0041_),
    .Y(_0678_));
 OA211x2_ASAP7_75t_R _1216_ (.A1(_0661_),
    .A2(_0677_),
    .B(_0678_),
    .C(_0646_),
    .Y(_0195_));
 AND3x1_ASAP7_75t_R _1217_ (.A(net42),
    .B(_0667_),
    .C(_0668_),
    .Y(_0679_));
 AO21x1_ASAP7_75t_R _1218_ (.A1(net4),
    .A2(_0666_),
    .B(_0679_),
    .Y(_0680_));
 NAND2x1_ASAP7_75t_R _1219_ (.A(_0671_),
    .B(_0040_),
    .Y(_0681_));
 OA211x2_ASAP7_75t_R _1220_ (.A1(_0661_),
    .A2(_0680_),
    .B(_0681_),
    .C(_0646_),
    .Y(_0196_));
 AND3x1_ASAP7_75t_R _1221_ (.A(net43),
    .B(_0667_),
    .C(_0668_),
    .Y(_0682_));
 AO21x1_ASAP7_75t_R _1222_ (.A1(net5),
    .A2(_0666_),
    .B(_0682_),
    .Y(_0683_));
 BUFx12f_ASAP7_75t_R _1223_ (.A(_0660_),
    .Y(_0230_));
 NAND2x1_ASAP7_75t_R _1224_ (.A(_0230_),
    .B(_0039_),
    .Y(_0231_));
 OA211x2_ASAP7_75t_R _1225_ (.A1(_0661_),
    .A2(_0683_),
    .B(_0231_),
    .C(_0646_),
    .Y(_0197_));
 AND3x1_ASAP7_75t_R _1226_ (.A(net44),
    .B(_0667_),
    .C(_0668_),
    .Y(_0232_));
 AO21x1_ASAP7_75t_R _1227_ (.A1(net6),
    .A2(_0666_),
    .B(_0232_),
    .Y(_0233_));
 NAND2x1_ASAP7_75t_R _1228_ (.A(_0230_),
    .B(_0038_),
    .Y(_0234_));
 OA211x2_ASAP7_75t_R _1229_ (.A1(_0661_),
    .A2(_0233_),
    .B(_0234_),
    .C(_0646_),
    .Y(_0198_));
 AND3x1_ASAP7_75t_R _1230_ (.A(net45),
    .B(_0667_),
    .C(_0668_),
    .Y(_0235_));
 AO21x1_ASAP7_75t_R _1231_ (.A1(net7),
    .A2(_0666_),
    .B(_0235_),
    .Y(_0236_));
 NAND2x1_ASAP7_75t_R _1232_ (.A(_0230_),
    .B(_0037_),
    .Y(_0237_));
 BUFx3_ASAP7_75t_R _1233_ (.A(_0419_),
    .Y(_0238_));
 OA211x2_ASAP7_75t_R _1234_ (.A1(_0661_),
    .A2(_0236_),
    .B(_0237_),
    .C(_0238_),
    .Y(_0199_));
 AND3x1_ASAP7_75t_R _1235_ (.A(net46),
    .B(_0667_),
    .C(_0668_),
    .Y(_0239_));
 AO21x1_ASAP7_75t_R _1236_ (.A1(net8),
    .A2(_0666_),
    .B(_0239_),
    .Y(_0240_));
 NAND2x1_ASAP7_75t_R _1237_ (.A(_0230_),
    .B(_0036_),
    .Y(_0241_));
 OA211x2_ASAP7_75t_R _1238_ (.A1(_0661_),
    .A2(_0240_),
    .B(_0241_),
    .C(_0238_),
    .Y(_0200_));
 AND3x1_ASAP7_75t_R _1239_ (.A(net47),
    .B(_0667_),
    .C(_0668_),
    .Y(_0242_));
 AO21x1_ASAP7_75t_R _1240_ (.A1(net9),
    .A2(_0666_),
    .B(_0242_),
    .Y(_0243_));
 NAND2x1_ASAP7_75t_R _1241_ (.A(_0230_),
    .B(_0035_),
    .Y(_0244_));
 OA211x2_ASAP7_75t_R _1242_ (.A1(_0661_),
    .A2(_0243_),
    .B(_0244_),
    .C(_0238_),
    .Y(_0201_));
 AND3x1_ASAP7_75t_R _1243_ (.A(net48),
    .B(_0667_),
    .C(_0668_),
    .Y(_0245_));
 AO21x1_ASAP7_75t_R _1244_ (.A1(net10),
    .A2(_0666_),
    .B(_0245_),
    .Y(_0246_));
 NAND2x1_ASAP7_75t_R _1245_ (.A(_0230_),
    .B(_0034_),
    .Y(_0247_));
 OA211x2_ASAP7_75t_R _1246_ (.A1(_0661_),
    .A2(_0246_),
    .B(_0247_),
    .C(_0238_),
    .Y(_0202_));
 BUFx6f_ASAP7_75t_R _1247_ (.A(_0660_),
    .Y(_0248_));
 BUFx6f_ASAP7_75t_R _1248_ (.A(_0665_),
    .Y(_0249_));
 BUFx6f_ASAP7_75t_R _1249_ (.A(_0662_),
    .Y(_0250_));
 BUFx6f_ASAP7_75t_R _1250_ (.A(_0664_),
    .Y(_0251_));
 AND3x1_ASAP7_75t_R _1251_ (.A(net49),
    .B(_0250_),
    .C(_0251_),
    .Y(_0252_));
 AO21x1_ASAP7_75t_R _1252_ (.A1(net11),
    .A2(_0249_),
    .B(_0252_),
    .Y(_0253_));
 NAND2x1_ASAP7_75t_R _1253_ (.A(_0230_),
    .B(_0033_),
    .Y(_0254_));
 OA211x2_ASAP7_75t_R _1254_ (.A1(_0248_),
    .A2(_0253_),
    .B(_0254_),
    .C(_0238_),
    .Y(_0203_));
 AND3x1_ASAP7_75t_R _1255_ (.A(net50),
    .B(_0250_),
    .C(_0251_),
    .Y(_0255_));
 AO21x1_ASAP7_75t_R _1256_ (.A1(net12),
    .A2(_0249_),
    .B(_0255_),
    .Y(_0256_));
 NAND2x1_ASAP7_75t_R _1257_ (.A(_0230_),
    .B(_0032_),
    .Y(_0257_));
 OA211x2_ASAP7_75t_R _1258_ (.A1(_0248_),
    .A2(_0256_),
    .B(_0257_),
    .C(_0238_),
    .Y(_0204_));
 AND3x1_ASAP7_75t_R _1259_ (.A(net51),
    .B(_0250_),
    .C(_0251_),
    .Y(_0258_));
 AO21x1_ASAP7_75t_R _1260_ (.A1(net13),
    .A2(_0249_),
    .B(_0258_),
    .Y(_0259_));
 NAND2x1_ASAP7_75t_R _1261_ (.A(_0230_),
    .B(_0031_),
    .Y(_0260_));
 OA211x2_ASAP7_75t_R _1262_ (.A1(_0248_),
    .A2(_0259_),
    .B(_0260_),
    .C(_0238_),
    .Y(_0205_));
 AND3x1_ASAP7_75t_R _1263_ (.A(net52),
    .B(_0250_),
    .C(_0251_),
    .Y(_0261_));
 AO21x1_ASAP7_75t_R _1264_ (.A1(net14),
    .A2(_0249_),
    .B(_0261_),
    .Y(_0262_));
 NAND2x1_ASAP7_75t_R _1265_ (.A(_0230_),
    .B(_0030_),
    .Y(_0263_));
 OA211x2_ASAP7_75t_R _1266_ (.A1(_0248_),
    .A2(_0262_),
    .B(_0263_),
    .C(_0238_),
    .Y(_0206_));
 AND3x1_ASAP7_75t_R _1267_ (.A(net53),
    .B(_0250_),
    .C(_0251_),
    .Y(_0264_));
 AO21x1_ASAP7_75t_R _1268_ (.A1(net15),
    .A2(_0249_),
    .B(_0264_),
    .Y(_0265_));
 BUFx12f_ASAP7_75t_R _1269_ (.A(_0660_),
    .Y(_0266_));
 NAND2x1_ASAP7_75t_R _1270_ (.A(_0266_),
    .B(_0029_),
    .Y(_0267_));
 OA211x2_ASAP7_75t_R _1271_ (.A1(_0248_),
    .A2(_0265_),
    .B(_0267_),
    .C(_0238_),
    .Y(_0207_));
 AND3x1_ASAP7_75t_R _1272_ (.A(net54),
    .B(_0250_),
    .C(_0251_),
    .Y(_0268_));
 AO21x1_ASAP7_75t_R _1273_ (.A1(net16),
    .A2(_0249_),
    .B(_0268_),
    .Y(_0269_));
 NAND2x1_ASAP7_75t_R _1274_ (.A(_0266_),
    .B(_0028_),
    .Y(_0270_));
 OA211x2_ASAP7_75t_R _1275_ (.A1(_0248_),
    .A2(_0269_),
    .B(_0270_),
    .C(_0238_),
    .Y(_0208_));
 AND3x1_ASAP7_75t_R _1276_ (.A(net55),
    .B(_0250_),
    .C(_0251_),
    .Y(_0271_));
 AO21x1_ASAP7_75t_R _1277_ (.A1(net17),
    .A2(_0249_),
    .B(_0271_),
    .Y(_0272_));
 NAND2x1_ASAP7_75t_R _1278_ (.A(_0266_),
    .B(_0027_),
    .Y(_0273_));
 BUFx3_ASAP7_75t_R _1279_ (.A(_0419_),
    .Y(_0274_));
 OA211x2_ASAP7_75t_R _1280_ (.A1(_0248_),
    .A2(_0272_),
    .B(_0273_),
    .C(_0274_),
    .Y(_0209_));
 AND3x1_ASAP7_75t_R _1281_ (.A(net56),
    .B(_0250_),
    .C(_0251_),
    .Y(_0275_));
 AO21x1_ASAP7_75t_R _1282_ (.A1(net18),
    .A2(_0249_),
    .B(_0275_),
    .Y(_0276_));
 NAND2x1_ASAP7_75t_R _1283_ (.A(_0266_),
    .B(_0026_),
    .Y(_0277_));
 OA211x2_ASAP7_75t_R _1284_ (.A1(_0248_),
    .A2(_0276_),
    .B(_0277_),
    .C(_0274_),
    .Y(_0210_));
 AND3x1_ASAP7_75t_R _1285_ (.A(net57),
    .B(_0250_),
    .C(_0251_),
    .Y(_0278_));
 AO21x1_ASAP7_75t_R _1286_ (.A1(net19),
    .A2(_0249_),
    .B(_0278_),
    .Y(_0279_));
 NAND2x1_ASAP7_75t_R _1287_ (.A(_0266_),
    .B(_0025_),
    .Y(_0280_));
 OA211x2_ASAP7_75t_R _1288_ (.A1(_0248_),
    .A2(_0279_),
    .B(_0280_),
    .C(_0274_),
    .Y(_0211_));
 AND3x1_ASAP7_75t_R _1289_ (.A(net58),
    .B(_0250_),
    .C(_0251_),
    .Y(_0281_));
 AO21x1_ASAP7_75t_R _1290_ (.A1(net20),
    .A2(_0249_),
    .B(_0281_),
    .Y(_0282_));
 NAND2x1_ASAP7_75t_R _1291_ (.A(_0266_),
    .B(_0024_),
    .Y(_0283_));
 OA211x2_ASAP7_75t_R _1292_ (.A1(_0248_),
    .A2(_0282_),
    .B(_0283_),
    .C(_0274_),
    .Y(_0212_));
 BUFx6f_ASAP7_75t_R _1293_ (.A(_0660_),
    .Y(_0284_));
 BUFx6f_ASAP7_75t_R _1294_ (.A(_0665_),
    .Y(_0285_));
 BUFx6f_ASAP7_75t_R _1295_ (.A(_0662_),
    .Y(_0286_));
 BUFx6f_ASAP7_75t_R _1296_ (.A(_0664_),
    .Y(_0287_));
 AND3x1_ASAP7_75t_R _1297_ (.A(net59),
    .B(_0286_),
    .C(_0287_),
    .Y(_0288_));
 AO21x1_ASAP7_75t_R _1298_ (.A1(net21),
    .A2(_0285_),
    .B(_0288_),
    .Y(_0289_));
 NAND2x1_ASAP7_75t_R _1299_ (.A(_0266_),
    .B(_0023_),
    .Y(_0290_));
 OA211x2_ASAP7_75t_R _1300_ (.A1(_0284_),
    .A2(_0289_),
    .B(_0290_),
    .C(_0274_),
    .Y(_0213_));
 AND3x1_ASAP7_75t_R _1301_ (.A(net60),
    .B(_0286_),
    .C(_0287_),
    .Y(_0291_));
 AO21x1_ASAP7_75t_R _1302_ (.A1(net22),
    .A2(_0285_),
    .B(_0291_),
    .Y(_0292_));
 NAND2x1_ASAP7_75t_R _1303_ (.A(_0266_),
    .B(_0022_),
    .Y(_0293_));
 OA211x2_ASAP7_75t_R _1304_ (.A1(_0284_),
    .A2(_0292_),
    .B(_0293_),
    .C(_0274_),
    .Y(_0214_));
 AND3x1_ASAP7_75t_R _1305_ (.A(net61),
    .B(_0286_),
    .C(_0287_),
    .Y(_0294_));
 AO21x1_ASAP7_75t_R _1306_ (.A1(net23),
    .A2(_0285_),
    .B(_0294_),
    .Y(_0295_));
 NAND2x1_ASAP7_75t_R _1307_ (.A(_0266_),
    .B(_0021_),
    .Y(_0296_));
 OA211x2_ASAP7_75t_R _1308_ (.A1(_0284_),
    .A2(_0295_),
    .B(_0296_),
    .C(_0274_),
    .Y(_0215_));
 AND3x1_ASAP7_75t_R _1309_ (.A(net62),
    .B(_0286_),
    .C(_0287_),
    .Y(_0297_));
 AO21x1_ASAP7_75t_R _1310_ (.A1(net24),
    .A2(_0285_),
    .B(_0297_),
    .Y(_0298_));
 NAND2x1_ASAP7_75t_R _1311_ (.A(_0266_),
    .B(_0020_),
    .Y(_0299_));
 OA211x2_ASAP7_75t_R _1312_ (.A1(_0284_),
    .A2(_0298_),
    .B(_0299_),
    .C(_0274_),
    .Y(_0216_));
 AND3x1_ASAP7_75t_R _1313_ (.A(net63),
    .B(_0286_),
    .C(_0287_),
    .Y(_0300_));
 AO21x1_ASAP7_75t_R _1314_ (.A1(net25),
    .A2(_0285_),
    .B(_0300_),
    .Y(_0301_));
 BUFx12f_ASAP7_75t_R _1315_ (.A(_0660_),
    .Y(_0302_));
 NAND2x1_ASAP7_75t_R _1316_ (.A(_0302_),
    .B(_0019_),
    .Y(_0303_));
 OA211x2_ASAP7_75t_R _1317_ (.A1(_0284_),
    .A2(_0301_),
    .B(_0303_),
    .C(_0274_),
    .Y(_0217_));
 AND3x1_ASAP7_75t_R _1318_ (.A(net64),
    .B(_0286_),
    .C(_0287_),
    .Y(_0304_));
 AO21x1_ASAP7_75t_R _1319_ (.A1(net26),
    .A2(_0285_),
    .B(_0304_),
    .Y(_0305_));
 NAND2x1_ASAP7_75t_R _1320_ (.A(_0302_),
    .B(_0018_),
    .Y(_0306_));
 OA211x2_ASAP7_75t_R _1321_ (.A1(_0284_),
    .A2(_0305_),
    .B(_0306_),
    .C(_0274_),
    .Y(_0218_));
 AND3x1_ASAP7_75t_R _1322_ (.A(net65),
    .B(_0286_),
    .C(_0287_),
    .Y(_0307_));
 AO21x1_ASAP7_75t_R _1323_ (.A1(net27),
    .A2(_0285_),
    .B(_0307_),
    .Y(_0308_));
 NAND2x1_ASAP7_75t_R _1324_ (.A(_0302_),
    .B(_0017_),
    .Y(_0309_));
 BUFx3_ASAP7_75t_R _1325_ (.A(_0419_),
    .Y(_0310_));
 OA211x2_ASAP7_75t_R _1326_ (.A1(_0284_),
    .A2(_0308_),
    .B(_0309_),
    .C(_0310_),
    .Y(_0219_));
 AND3x1_ASAP7_75t_R _1327_ (.A(net66),
    .B(_0286_),
    .C(_0287_),
    .Y(_0311_));
 AO21x1_ASAP7_75t_R _1328_ (.A1(net28),
    .A2(_0285_),
    .B(_0311_),
    .Y(_0312_));
 NAND2x1_ASAP7_75t_R _1329_ (.A(_0302_),
    .B(_0016_),
    .Y(_0313_));
 OA211x2_ASAP7_75t_R _1330_ (.A1(_0284_),
    .A2(_0312_),
    .B(_0313_),
    .C(_0310_),
    .Y(_0220_));
 AND3x1_ASAP7_75t_R _1331_ (.A(net67),
    .B(_0286_),
    .C(_0287_),
    .Y(_0314_));
 AO21x1_ASAP7_75t_R _1332_ (.A1(net29),
    .A2(_0285_),
    .B(_0314_),
    .Y(_0315_));
 NAND2x1_ASAP7_75t_R _1333_ (.A(_0302_),
    .B(_0015_),
    .Y(_0316_));
 OA211x2_ASAP7_75t_R _1334_ (.A1(_0284_),
    .A2(_0315_),
    .B(_0316_),
    .C(_0310_),
    .Y(_0221_));
 AND3x1_ASAP7_75t_R _1335_ (.A(net68),
    .B(_0286_),
    .C(_0287_),
    .Y(_0317_));
 AO21x1_ASAP7_75t_R _1336_ (.A1(net30),
    .A2(_0285_),
    .B(_0317_),
    .Y(_0318_));
 NAND2x1_ASAP7_75t_R _1337_ (.A(_0302_),
    .B(_0014_),
    .Y(_0319_));
 OA211x2_ASAP7_75t_R _1338_ (.A1(_0284_),
    .A2(_0318_),
    .B(_0319_),
    .C(_0310_),
    .Y(_0222_));
 AND3x1_ASAP7_75t_R _1339_ (.A(net69),
    .B(_0662_),
    .C(_0664_),
    .Y(_0320_));
 AO21x1_ASAP7_75t_R _1340_ (.A1(net31),
    .A2(_0665_),
    .B(_0320_),
    .Y(_0321_));
 NAND2x1_ASAP7_75t_R _1341_ (.A(_0302_),
    .B(_0013_),
    .Y(_0322_));
 OA211x2_ASAP7_75t_R _1342_ (.A1(_0671_),
    .A2(_0321_),
    .B(_0322_),
    .C(_0310_),
    .Y(_0223_));
 AND3x1_ASAP7_75t_R _1343_ (.A(net70),
    .B(_0662_),
    .C(_0664_),
    .Y(_0323_));
 AO21x1_ASAP7_75t_R _1344_ (.A1(net32),
    .A2(_0665_),
    .B(_0323_),
    .Y(_0324_));
 NAND2x1_ASAP7_75t_R _1345_ (.A(_0302_),
    .B(_0012_),
    .Y(_0325_));
 OA211x2_ASAP7_75t_R _1346_ (.A1(_0671_),
    .A2(_0324_),
    .B(_0325_),
    .C(_0310_),
    .Y(_0224_));
 AND3x1_ASAP7_75t_R _1347_ (.A(net71),
    .B(_0662_),
    .C(_0664_),
    .Y(_0326_));
 AO21x1_ASAP7_75t_R _1348_ (.A1(net33),
    .A2(_0665_),
    .B(_0326_),
    .Y(_0327_));
 NAND2x1_ASAP7_75t_R _1349_ (.A(_0302_),
    .B(_0011_),
    .Y(_0328_));
 OA211x2_ASAP7_75t_R _1350_ (.A1(_0671_),
    .A2(_0327_),
    .B(_0328_),
    .C(_0310_),
    .Y(_0225_));
 AND3x1_ASAP7_75t_R _1351_ (.A(net72),
    .B(_0662_),
    .C(_0664_),
    .Y(_0329_));
 AO21x1_ASAP7_75t_R _1352_ (.A1(net34),
    .A2(_0665_),
    .B(_0329_),
    .Y(_0330_));
 NAND2x1_ASAP7_75t_R _1353_ (.A(_0302_),
    .B(_0010_),
    .Y(_0331_));
 OA211x2_ASAP7_75t_R _1354_ (.A1(_0671_),
    .A2(_0330_),
    .B(_0331_),
    .C(_0310_),
    .Y(_0226_));
 AND3x1_ASAP7_75t_R _1355_ (.A(net73),
    .B(_0662_),
    .C(_0664_),
    .Y(_0332_));
 AO21x1_ASAP7_75t_R _1356_ (.A1(net35),
    .A2(_0665_),
    .B(_0332_),
    .Y(_0333_));
 NAND2x1_ASAP7_75t_R _1357_ (.A(_0660_),
    .B(_0009_),
    .Y(_0334_));
 OA211x2_ASAP7_75t_R _1358_ (.A1(_0671_),
    .A2(_0333_),
    .B(_0334_),
    .C(_0310_),
    .Y(_0227_));
 AND3x1_ASAP7_75t_R _1359_ (.A(net74),
    .B(_0662_),
    .C(_0664_),
    .Y(_0335_));
 AO21x1_ASAP7_75t_R _1360_ (.A1(net36),
    .A2(_0665_),
    .B(_0335_),
    .Y(_0336_));
 NAND2x1_ASAP7_75t_R _1361_ (.A(_0660_),
    .B(_0008_),
    .Y(_0337_));
 OA211x2_ASAP7_75t_R _1362_ (.A1(_0671_),
    .A2(_0336_),
    .B(_0337_),
    .C(_0310_),
    .Y(_0228_));
 AND4x1_ASAP7_75t_R _1363_ (.A(_0004_),
    .B(_0345_),
    .C(_0350_),
    .D(_0351_),
    .Y(_0338_));
 NOR2x1_ASAP7_75t_R _1364_ (.A(_0350_),
    .B(_0351_),
    .Y(_0339_));
 OR3x1_ASAP7_75t_R _1365_ (.A(_0660_),
    .B(_0338_),
    .C(_0339_),
    .Y(_0340_));
 OA21x2_ASAP7_75t_R _1366_ (.A1(_0663_),
    .A2(_0007_),
    .B(_0340_),
    .Y(_0341_));
 NOR2x1_ASAP7_75t_R _1367_ (.A(_0367_),
    .B(_0341_),
    .Y(_0229_));
 DFFHQNx1_ASAP7_75t_R \done_sig$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .D(_0000_),
    .QN(_0117_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[0]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0119_),
    .QN(_0116_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[10]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0120_),
    .QN(_0115_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[11]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0121_),
    .QN(_0114_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[12]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0122_),
    .QN(_0113_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[13]$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0123_),
    .QN(_0112_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[14]$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0124_),
    .QN(_0111_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[15]$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0125_),
    .QN(_0110_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[16]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0126_),
    .QN(_0109_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[17]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0127_),
    .QN(_0108_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[18]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0128_),
    .QN(_0107_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[19]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0129_),
    .QN(_0106_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[1]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0130_),
    .QN(_0105_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[20]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0131_),
    .QN(_0104_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[21]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0132_),
    .QN(_0103_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[22]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0133_),
    .QN(_0102_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[23]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0134_),
    .QN(_0101_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[24]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0135_),
    .QN(_0100_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[25]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0136_),
    .QN(_0099_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[26]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0137_),
    .QN(_0098_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[27]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0138_),
    .QN(_0097_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[28]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0139_),
    .QN(_0096_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[29]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0140_),
    .QN(_0095_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[2]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0141_),
    .QN(_0094_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[30]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0142_),
    .QN(_0093_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[31]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0143_),
    .QN(_0092_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[32]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0144_),
    .QN(_0091_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[33]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0145_),
    .QN(_0090_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[34]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0146_),
    .QN(_0089_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[35]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0147_),
    .QN(_0088_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[3]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0148_),
    .QN(_0087_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[4]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0149_),
    .QN(_0086_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[5]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0150_),
    .QN(_0085_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[6]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0151_),
    .QN(_0084_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[7]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0152_),
    .QN(_0083_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[8]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0153_),
    .QN(_0082_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[9]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0154_),
    .QN(_0081_));
 DFFHQNx1_ASAP7_75t_R \l_o_v_r$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0155_),
    .QN(_0118_));
 DFFHQNx3_ASAP7_75t_R \r.rr[0]$_DFF_P_  (.CLK(clknet_4_10_0_clk),
    .D(_0001_),
    .QN(_0004_));
 DFFHQNx1_ASAP7_75t_R \r.rr[1]$_DFF_P_  (.CLK(clknet_4_10_0_clk),
    .D(_0002_),
    .QN(_0006_));
 DFFHQNx1_ASAP7_75t_R \r.rr[2]$_DFF_P_  (.CLK(clknet_4_10_0_clk),
    .D(_0003_),
    .QN(_0005_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[0]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0156_),
    .QN(_0080_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[10]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0157_),
    .QN(_0079_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[11]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0158_),
    .QN(_0078_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[12]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0159_),
    .QN(_0077_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[13]$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0160_),
    .QN(_0076_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[14]$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0161_),
    .QN(_0075_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[15]$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0162_),
    .QN(_0074_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[16]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0163_),
    .QN(_0073_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[17]$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0164_),
    .QN(_0072_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[18]$_SDFFE_PP0N_  (.CLK(clknet_4_0_0_clk),
    .D(_0165_),
    .QN(_0071_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[19]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0166_),
    .QN(_0070_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[1]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0167_),
    .QN(_0069_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[20]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0168_),
    .QN(_0068_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[21]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0169_),
    .QN(_0067_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[22]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0170_),
    .QN(_0066_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[23]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0171_),
    .QN(_0065_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[24]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0172_),
    .QN(_0064_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[25]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0173_),
    .QN(_0063_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[26]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0174_),
    .QN(_0062_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[27]$_SDFFE_PP0N_  (.CLK(clknet_4_6_0_clk),
    .D(_0175_),
    .QN(_0061_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[28]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0176_),
    .QN(_0060_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[29]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0177_),
    .QN(_0059_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[2]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0178_),
    .QN(_0058_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[30]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0179_),
    .QN(_0057_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[31]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0180_),
    .QN(_0056_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[32]$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0181_),
    .QN(_0055_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[33]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0182_),
    .QN(_0054_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[34]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0183_),
    .QN(_0053_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[35]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0184_),
    .QN(_0052_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[3]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0185_),
    .QN(_0051_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[4]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0186_),
    .QN(_0050_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[5]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0187_),
    .QN(_0049_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[6]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0188_),
    .QN(_0048_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[7]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0189_),
    .QN(_0047_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[8]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0190_),
    .QN(_0046_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[9]$_SDFFE_PP0N_  (.CLK(clknet_4_8_0_clk),
    .D(_0191_),
    .QN(_0045_));
 DFFHQNx1_ASAP7_75t_R \r_o_v_r$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0192_),
    .QN(_0044_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[0]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0193_),
    .QN(_0043_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[10]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0194_),
    .QN(_0042_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[11]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0195_),
    .QN(_0041_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[12]$_SDFFE_PP0N_  (.CLK(clknet_4_2_0_clk),
    .D(_0196_),
    .QN(_0040_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[13]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0197_),
    .QN(_0039_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[14]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0198_),
    .QN(_0038_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[15]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0199_),
    .QN(_0037_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[16]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0200_),
    .QN(_0036_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[17]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0201_),
    .QN(_0035_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[18]$_SDFFE_PP0N_  (.CLK(clknet_4_1_0_clk),
    .D(_0202_),
    .QN(_0034_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[19]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0203_),
    .QN(_0033_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[1]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0204_),
    .QN(_0032_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[20]$_SDFFE_PP0N_  (.CLK(clknet_4_4_0_clk),
    .D(_0205_),
    .QN(_0031_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[21]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0206_),
    .QN(_0030_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[22]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0207_),
    .QN(_0029_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[23]$_SDFFE_PP0N_  (.CLK(clknet_4_5_0_clk),
    .D(_0208_),
    .QN(_0028_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[24]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0209_),
    .QN(_0027_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[25]$_SDFFE_PP0N_  (.CLK(clknet_4_13_0_clk),
    .D(_0210_),
    .QN(_0026_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[26]$_SDFFE_PP0N_  (.CLK(clknet_4_7_0_clk),
    .D(_0211_),
    .QN(_0025_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[27]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0212_),
    .QN(_0024_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[28]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0213_),
    .QN(_0023_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[29]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0214_),
    .QN(_0022_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[2]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0215_),
    .QN(_0021_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[30]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0216_),
    .QN(_0020_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[31]$_SDFFE_PP0N_  (.CLK(clknet_4_15_0_clk),
    .D(_0217_),
    .QN(_0019_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[32]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0218_),
    .QN(_0018_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[33]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0219_),
    .QN(_0017_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[34]$_SDFFE_PP0N_  (.CLK(clknet_4_11_0_clk),
    .D(_0220_),
    .QN(_0016_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[35]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0221_),
    .QN(_0015_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[3]$_SDFFE_PP0N_  (.CLK(clknet_4_14_0_clk),
    .D(_0222_),
    .QN(_0014_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[4]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0223_),
    .QN(_0013_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[5]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0224_),
    .QN(_0012_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[6]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0225_),
    .QN(_0011_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[7]$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .D(_0226_),
    .QN(_0010_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[8]$_SDFFE_PP0N_  (.CLK(clknet_4_3_0_clk),
    .D(_0227_),
    .QN(_0009_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[9]$_SDFFE_PP0N_  (.CLK(clknet_4_12_0_clk),
    .D(_0228_),
    .QN(_0008_));
 DFFHQNx1_ASAP7_75t_R \u0_o_v_r$_SDFFE_PP0N_  (.CLK(clknet_4_10_0_clk),
    .D(_0229_),
    .QN(_0007_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Left_111 ();
 BUFx3_ASAP7_75t_R input1 (.A(l_i[0]),
    .Y(net1));
 BUFx3_ASAP7_75t_R input2 (.A(l_i[10]),
    .Y(net2));
 BUFx3_ASAP7_75t_R input3 (.A(l_i[11]),
    .Y(net3));
 BUFx3_ASAP7_75t_R input4 (.A(l_i[12]),
    .Y(net4));
 BUFx3_ASAP7_75t_R input5 (.A(l_i[13]),
    .Y(net5));
 BUFx3_ASAP7_75t_R input6 (.A(l_i[14]),
    .Y(net6));
 BUFx3_ASAP7_75t_R input7 (.A(l_i[15]),
    .Y(net7));
 BUFx3_ASAP7_75t_R input8 (.A(l_i[16]),
    .Y(net8));
 BUFx3_ASAP7_75t_R input9 (.A(l_i[17]),
    .Y(net9));
 BUFx3_ASAP7_75t_R input10 (.A(l_i[18]),
    .Y(net10));
 BUFx3_ASAP7_75t_R input11 (.A(l_i[19]),
    .Y(net11));
 BUFx3_ASAP7_75t_R input12 (.A(l_i[1]),
    .Y(net12));
 BUFx3_ASAP7_75t_R input13 (.A(l_i[20]),
    .Y(net13));
 BUFx3_ASAP7_75t_R input14 (.A(l_i[21]),
    .Y(net14));
 BUFx3_ASAP7_75t_R input15 (.A(l_i[22]),
    .Y(net15));
 BUFx3_ASAP7_75t_R input16 (.A(l_i[23]),
    .Y(net16));
 BUFx3_ASAP7_75t_R input17 (.A(l_i[24]),
    .Y(net17));
 BUFx3_ASAP7_75t_R input18 (.A(l_i[25]),
    .Y(net18));
 BUFx3_ASAP7_75t_R input19 (.A(l_i[26]),
    .Y(net19));
 BUFx3_ASAP7_75t_R input20 (.A(l_i[27]),
    .Y(net20));
 BUFx3_ASAP7_75t_R input21 (.A(l_i[28]),
    .Y(net21));
 BUFx3_ASAP7_75t_R input22 (.A(l_i[29]),
    .Y(net22));
 BUFx3_ASAP7_75t_R input23 (.A(l_i[2]),
    .Y(net23));
 BUFx3_ASAP7_75t_R input24 (.A(l_i[30]),
    .Y(net24));
 BUFx3_ASAP7_75t_R input25 (.A(l_i[31]),
    .Y(net25));
 BUFx3_ASAP7_75t_R input26 (.A(l_i[32]),
    .Y(net26));
 BUFx3_ASAP7_75t_R input27 (.A(l_i[33]),
    .Y(net27));
 BUFx3_ASAP7_75t_R input28 (.A(l_i[34]),
    .Y(net28));
 BUFx3_ASAP7_75t_R input29 (.A(l_i[35]),
    .Y(net29));
 BUFx3_ASAP7_75t_R input30 (.A(l_i[3]),
    .Y(net30));
 BUFx3_ASAP7_75t_R input31 (.A(l_i[4]),
    .Y(net31));
 BUFx3_ASAP7_75t_R input32 (.A(l_i[5]),
    .Y(net32));
 BUFx3_ASAP7_75t_R input33 (.A(l_i[6]),
    .Y(net33));
 BUFx3_ASAP7_75t_R input34 (.A(l_i[7]),
    .Y(net34));
 BUFx3_ASAP7_75t_R input35 (.A(l_i[8]),
    .Y(net35));
 BUFx3_ASAP7_75t_R input36 (.A(l_i[9]),
    .Y(net36));
 BUFx3_ASAP7_75t_R input37 (.A(l_i_v),
    .Y(net37));
 BUFx3_ASAP7_75t_R input38 (.A(l_o_bp),
    .Y(net38));
 BUFx3_ASAP7_75t_R input39 (.A(r_i[0]),
    .Y(net39));
 BUFx3_ASAP7_75t_R input40 (.A(r_i[10]),
    .Y(net40));
 BUFx3_ASAP7_75t_R input41 (.A(r_i[11]),
    .Y(net41));
 BUFx3_ASAP7_75t_R input42 (.A(r_i[12]),
    .Y(net42));
 BUFx3_ASAP7_75t_R input43 (.A(r_i[13]),
    .Y(net43));
 BUFx3_ASAP7_75t_R input44 (.A(r_i[14]),
    .Y(net44));
 BUFx3_ASAP7_75t_R input45 (.A(r_i[15]),
    .Y(net45));
 BUFx3_ASAP7_75t_R input46 (.A(r_i[16]),
    .Y(net46));
 BUFx3_ASAP7_75t_R input47 (.A(r_i[17]),
    .Y(net47));
 BUFx3_ASAP7_75t_R input48 (.A(r_i[18]),
    .Y(net48));
 BUFx3_ASAP7_75t_R input49 (.A(r_i[19]),
    .Y(net49));
 BUFx3_ASAP7_75t_R input50 (.A(r_i[1]),
    .Y(net50));
 BUFx3_ASAP7_75t_R input51 (.A(r_i[20]),
    .Y(net51));
 BUFx3_ASAP7_75t_R input52 (.A(r_i[21]),
    .Y(net52));
 BUFx3_ASAP7_75t_R input53 (.A(r_i[22]),
    .Y(net53));
 BUFx3_ASAP7_75t_R input54 (.A(r_i[23]),
    .Y(net54));
 BUFx3_ASAP7_75t_R input55 (.A(r_i[24]),
    .Y(net55));
 BUFx3_ASAP7_75t_R input56 (.A(r_i[25]),
    .Y(net56));
 BUFx3_ASAP7_75t_R input57 (.A(r_i[26]),
    .Y(net57));
 BUFx3_ASAP7_75t_R input58 (.A(r_i[27]),
    .Y(net58));
 BUFx3_ASAP7_75t_R input59 (.A(r_i[28]),
    .Y(net59));
 BUFx3_ASAP7_75t_R input60 (.A(r_i[29]),
    .Y(net60));
 BUFx3_ASAP7_75t_R input61 (.A(r_i[2]),
    .Y(net61));
 BUFx3_ASAP7_75t_R input62 (.A(r_i[30]),
    .Y(net62));
 BUFx3_ASAP7_75t_R input63 (.A(r_i[31]),
    .Y(net63));
 BUFx3_ASAP7_75t_R input64 (.A(r_i[32]),
    .Y(net64));
 BUFx3_ASAP7_75t_R input65 (.A(r_i[33]),
    .Y(net65));
 BUFx3_ASAP7_75t_R input66 (.A(r_i[34]),
    .Y(net66));
 BUFx3_ASAP7_75t_R input67 (.A(r_i[35]),
    .Y(net67));
 BUFx3_ASAP7_75t_R input68 (.A(r_i[3]),
    .Y(net68));
 BUFx3_ASAP7_75t_R input69 (.A(r_i[4]),
    .Y(net69));
 BUFx3_ASAP7_75t_R input70 (.A(r_i[5]),
    .Y(net70));
 BUFx3_ASAP7_75t_R input71 (.A(r_i[6]),
    .Y(net71));
 BUFx3_ASAP7_75t_R input72 (.A(r_i[7]),
    .Y(net72));
 BUFx3_ASAP7_75t_R input73 (.A(r_i[8]),
    .Y(net73));
 BUFx3_ASAP7_75t_R input74 (.A(r_i[9]),
    .Y(net74));
 BUFx3_ASAP7_75t_R input75 (.A(r_i_v),
    .Y(net75));
 BUFx6f_ASAP7_75t_R input76 (.A(r_o_bp),
    .Y(net76));
 BUFx3_ASAP7_75t_R input77 (.A(u0_i[0]),
    .Y(net77));
 BUFx3_ASAP7_75t_R input78 (.A(u0_i[10]),
    .Y(net78));
 BUFx3_ASAP7_75t_R input79 (.A(u0_i[11]),
    .Y(net79));
 BUFx3_ASAP7_75t_R input80 (.A(u0_i[12]),
    .Y(net80));
 BUFx3_ASAP7_75t_R input81 (.A(u0_i[13]),
    .Y(net81));
 BUFx3_ASAP7_75t_R input82 (.A(u0_i[14]),
    .Y(net82));
 BUFx3_ASAP7_75t_R input83 (.A(u0_i[15]),
    .Y(net83));
 BUFx3_ASAP7_75t_R input84 (.A(u0_i[16]),
    .Y(net84));
 BUFx3_ASAP7_75t_R input85 (.A(u0_i[17]),
    .Y(net85));
 BUFx3_ASAP7_75t_R input86 (.A(u0_i[18]),
    .Y(net86));
 BUFx3_ASAP7_75t_R input87 (.A(u0_i[19]),
    .Y(net87));
 BUFx3_ASAP7_75t_R input88 (.A(u0_i[1]),
    .Y(net88));
 BUFx3_ASAP7_75t_R input89 (.A(u0_i[20]),
    .Y(net89));
 BUFx3_ASAP7_75t_R input90 (.A(u0_i[21]),
    .Y(net90));
 BUFx3_ASAP7_75t_R input91 (.A(u0_i[22]),
    .Y(net91));
 BUFx3_ASAP7_75t_R input92 (.A(u0_i[23]),
    .Y(net92));
 BUFx3_ASAP7_75t_R input93 (.A(u0_i[24]),
    .Y(net93));
 BUFx3_ASAP7_75t_R input94 (.A(u0_i[25]),
    .Y(net94));
 BUFx3_ASAP7_75t_R input95 (.A(u0_i[26]),
    .Y(net95));
 BUFx3_ASAP7_75t_R input96 (.A(u0_i[27]),
    .Y(net96));
 BUFx3_ASAP7_75t_R input97 (.A(u0_i[28]),
    .Y(net97));
 BUFx3_ASAP7_75t_R input98 (.A(u0_i[29]),
    .Y(net98));
 BUFx3_ASAP7_75t_R input99 (.A(u0_i[2]),
    .Y(net99));
 BUFx3_ASAP7_75t_R input100 (.A(u0_i[30]),
    .Y(net100));
 BUFx3_ASAP7_75t_R input101 (.A(u0_i[31]),
    .Y(net101));
 BUFx3_ASAP7_75t_R input102 (.A(u0_i[32]),
    .Y(net102));
 BUFx3_ASAP7_75t_R input103 (.A(u0_i[33]),
    .Y(net103));
 BUFx3_ASAP7_75t_R input104 (.A(u0_i[34]),
    .Y(net104));
 BUFx3_ASAP7_75t_R input105 (.A(u0_i[35]),
    .Y(net105));
 BUFx3_ASAP7_75t_R input106 (.A(u0_i[3]),
    .Y(net106));
 BUFx3_ASAP7_75t_R input107 (.A(u0_i[4]),
    .Y(net107));
 BUFx3_ASAP7_75t_R input108 (.A(u0_i[5]),
    .Y(net108));
 BUFx3_ASAP7_75t_R input109 (.A(u0_i[6]),
    .Y(net109));
 BUFx3_ASAP7_75t_R input110 (.A(u0_i[7]),
    .Y(net110));
 BUFx3_ASAP7_75t_R input111 (.A(u0_i[8]),
    .Y(net111));
 BUFx3_ASAP7_75t_R input112 (.A(u0_i[9]),
    .Y(net112));
 BUFx3_ASAP7_75t_R input113 (.A(u0_o_bp),
    .Y(net113));
 BUFx3_ASAP7_75t_R output114 (.A(net114),
    .Y(done));
 BUFx3_ASAP7_75t_R output115 (.A(net115),
    .Y(l_i_bp));
 BUFx3_ASAP7_75t_R output116 (.A(net116),
    .Y(l_o[0]));
 BUFx3_ASAP7_75t_R output117 (.A(net117),
    .Y(l_o[10]));
 BUFx3_ASAP7_75t_R output118 (.A(net118),
    .Y(l_o[11]));
 BUFx3_ASAP7_75t_R output119 (.A(net119),
    .Y(l_o[12]));
 BUFx3_ASAP7_75t_R output120 (.A(net120),
    .Y(l_o[13]));
 BUFx3_ASAP7_75t_R output121 (.A(net121),
    .Y(l_o[14]));
 BUFx3_ASAP7_75t_R output122 (.A(net122),
    .Y(l_o[15]));
 BUFx3_ASAP7_75t_R output123 (.A(net123),
    .Y(l_o[16]));
 BUFx3_ASAP7_75t_R output124 (.A(net124),
    .Y(l_o[17]));
 BUFx3_ASAP7_75t_R output125 (.A(net125),
    .Y(l_o[18]));
 BUFx3_ASAP7_75t_R output126 (.A(net126),
    .Y(l_o[19]));
 BUFx3_ASAP7_75t_R output127 (.A(net127),
    .Y(l_o[1]));
 BUFx3_ASAP7_75t_R output128 (.A(net128),
    .Y(l_o[20]));
 BUFx3_ASAP7_75t_R output129 (.A(net129),
    .Y(l_o[21]));
 BUFx3_ASAP7_75t_R output130 (.A(net130),
    .Y(l_o[22]));
 BUFx3_ASAP7_75t_R output131 (.A(net131),
    .Y(l_o[23]));
 BUFx3_ASAP7_75t_R output132 (.A(net132),
    .Y(l_o[24]));
 BUFx3_ASAP7_75t_R output133 (.A(net133),
    .Y(l_o[25]));
 BUFx3_ASAP7_75t_R output134 (.A(net134),
    .Y(l_o[26]));
 BUFx3_ASAP7_75t_R output135 (.A(net135),
    .Y(l_o[27]));
 BUFx3_ASAP7_75t_R output136 (.A(net136),
    .Y(l_o[28]));
 BUFx3_ASAP7_75t_R output137 (.A(net137),
    .Y(l_o[29]));
 BUFx3_ASAP7_75t_R output138 (.A(net138),
    .Y(l_o[2]));
 BUFx3_ASAP7_75t_R output139 (.A(net139),
    .Y(l_o[30]));
 BUFx3_ASAP7_75t_R output140 (.A(net140),
    .Y(l_o[31]));
 BUFx3_ASAP7_75t_R output141 (.A(net141),
    .Y(l_o[32]));
 BUFx3_ASAP7_75t_R output142 (.A(net142),
    .Y(l_o[33]));
 BUFx3_ASAP7_75t_R output143 (.A(net143),
    .Y(l_o[34]));
 BUFx3_ASAP7_75t_R output144 (.A(net144),
    .Y(l_o[35]));
 BUFx3_ASAP7_75t_R output145 (.A(net145),
    .Y(l_o[3]));
 BUFx3_ASAP7_75t_R output146 (.A(net146),
    .Y(l_o[4]));
 BUFx3_ASAP7_75t_R output147 (.A(net147),
    .Y(l_o[5]));
 BUFx3_ASAP7_75t_R output148 (.A(net148),
    .Y(l_o[6]));
 BUFx3_ASAP7_75t_R output149 (.A(net149),
    .Y(l_o[7]));
 BUFx3_ASAP7_75t_R output150 (.A(net150),
    .Y(l_o[8]));
 BUFx3_ASAP7_75t_R output151 (.A(net151),
    .Y(l_o[9]));
 BUFx3_ASAP7_75t_R output152 (.A(net152),
    .Y(l_o_v));
 BUFx3_ASAP7_75t_R output153 (.A(net153),
    .Y(r_i_bp));
 BUFx3_ASAP7_75t_R output154 (.A(net154),
    .Y(r_o[0]));
 BUFx3_ASAP7_75t_R output155 (.A(net155),
    .Y(r_o[10]));
 BUFx3_ASAP7_75t_R output156 (.A(net156),
    .Y(r_o[11]));
 BUFx3_ASAP7_75t_R output157 (.A(net157),
    .Y(r_o[12]));
 BUFx3_ASAP7_75t_R output158 (.A(net158),
    .Y(r_o[13]));
 BUFx3_ASAP7_75t_R output159 (.A(net159),
    .Y(r_o[14]));
 BUFx3_ASAP7_75t_R output160 (.A(net160),
    .Y(r_o[15]));
 BUFx3_ASAP7_75t_R output161 (.A(net161),
    .Y(r_o[16]));
 BUFx3_ASAP7_75t_R output162 (.A(net162),
    .Y(r_o[17]));
 BUFx3_ASAP7_75t_R output163 (.A(net163),
    .Y(r_o[18]));
 BUFx3_ASAP7_75t_R output164 (.A(net164),
    .Y(r_o[19]));
 BUFx3_ASAP7_75t_R output165 (.A(net165),
    .Y(r_o[1]));
 BUFx3_ASAP7_75t_R output166 (.A(net166),
    .Y(r_o[20]));
 BUFx3_ASAP7_75t_R output167 (.A(net167),
    .Y(r_o[21]));
 BUFx3_ASAP7_75t_R output168 (.A(net168),
    .Y(r_o[22]));
 BUFx3_ASAP7_75t_R output169 (.A(net169),
    .Y(r_o[23]));
 BUFx3_ASAP7_75t_R output170 (.A(net170),
    .Y(r_o[24]));
 BUFx3_ASAP7_75t_R output171 (.A(net171),
    .Y(r_o[25]));
 BUFx3_ASAP7_75t_R output172 (.A(net172),
    .Y(r_o[26]));
 BUFx3_ASAP7_75t_R output173 (.A(net173),
    .Y(r_o[27]));
 BUFx3_ASAP7_75t_R output174 (.A(net174),
    .Y(r_o[28]));
 BUFx3_ASAP7_75t_R output175 (.A(net175),
    .Y(r_o[29]));
 BUFx3_ASAP7_75t_R output176 (.A(net176),
    .Y(r_o[2]));
 BUFx3_ASAP7_75t_R output177 (.A(net177),
    .Y(r_o[30]));
 BUFx3_ASAP7_75t_R output178 (.A(net178),
    .Y(r_o[31]));
 BUFx3_ASAP7_75t_R output179 (.A(net179),
    .Y(r_o[32]));
 BUFx3_ASAP7_75t_R output180 (.A(net180),
    .Y(r_o[33]));
 BUFx3_ASAP7_75t_R output181 (.A(net181),
    .Y(r_o[34]));
 BUFx3_ASAP7_75t_R output182 (.A(net182),
    .Y(r_o[35]));
 BUFx3_ASAP7_75t_R output183 (.A(net183),
    .Y(r_o[3]));
 BUFx3_ASAP7_75t_R output184 (.A(net184),
    .Y(r_o[4]));
 BUFx3_ASAP7_75t_R output185 (.A(net185),
    .Y(r_o[5]));
 BUFx3_ASAP7_75t_R output186 (.A(net186),
    .Y(r_o[6]));
 BUFx3_ASAP7_75t_R output187 (.A(net187),
    .Y(r_o[7]));
 BUFx3_ASAP7_75t_R output188 (.A(net188),
    .Y(r_o[8]));
 BUFx3_ASAP7_75t_R output189 (.A(net189),
    .Y(r_o[9]));
 BUFx3_ASAP7_75t_R output190 (.A(net190),
    .Y(r_o_v));
 BUFx3_ASAP7_75t_R output191 (.A(net191),
    .Y(u0_i_bp));
 BUFx3_ASAP7_75t_R output192 (.A(net192),
    .Y(u0_o[0]));
 BUFx3_ASAP7_75t_R output193 (.A(net193),
    .Y(u0_o[10]));
 BUFx3_ASAP7_75t_R output194 (.A(net194),
    .Y(u0_o[11]));
 BUFx3_ASAP7_75t_R output195 (.A(net195),
    .Y(u0_o[12]));
 BUFx3_ASAP7_75t_R output196 (.A(net196),
    .Y(u0_o[13]));
 BUFx3_ASAP7_75t_R output197 (.A(net197),
    .Y(u0_o[14]));
 BUFx3_ASAP7_75t_R output198 (.A(net198),
    .Y(u0_o[15]));
 BUFx3_ASAP7_75t_R output199 (.A(net199),
    .Y(u0_o[16]));
 BUFx3_ASAP7_75t_R output200 (.A(net200),
    .Y(u0_o[17]));
 BUFx3_ASAP7_75t_R output201 (.A(net201),
    .Y(u0_o[18]));
 BUFx3_ASAP7_75t_R output202 (.A(net202),
    .Y(u0_o[19]));
 BUFx3_ASAP7_75t_R output203 (.A(net203),
    .Y(u0_o[1]));
 BUFx3_ASAP7_75t_R output204 (.A(net204),
    .Y(u0_o[20]));
 BUFx3_ASAP7_75t_R output205 (.A(net205),
    .Y(u0_o[21]));
 BUFx3_ASAP7_75t_R output206 (.A(net206),
    .Y(u0_o[22]));
 BUFx3_ASAP7_75t_R output207 (.A(net207),
    .Y(u0_o[23]));
 BUFx3_ASAP7_75t_R output208 (.A(net208),
    .Y(u0_o[24]));
 BUFx3_ASAP7_75t_R output209 (.A(net209),
    .Y(u0_o[25]));
 BUFx3_ASAP7_75t_R output210 (.A(net210),
    .Y(u0_o[26]));
 BUFx3_ASAP7_75t_R output211 (.A(net211),
    .Y(u0_o[27]));
 BUFx3_ASAP7_75t_R output212 (.A(net212),
    .Y(u0_o[28]));
 BUFx3_ASAP7_75t_R output213 (.A(net213),
    .Y(u0_o[29]));
 BUFx3_ASAP7_75t_R output214 (.A(net214),
    .Y(u0_o[2]));
 BUFx3_ASAP7_75t_R output215 (.A(net215),
    .Y(u0_o[30]));
 BUFx3_ASAP7_75t_R output216 (.A(net216),
    .Y(u0_o[31]));
 BUFx3_ASAP7_75t_R output217 (.A(net217),
    .Y(u0_o[32]));
 BUFx3_ASAP7_75t_R output218 (.A(net218),
    .Y(u0_o[33]));
 BUFx3_ASAP7_75t_R output219 (.A(net219),
    .Y(u0_o[34]));
 BUFx3_ASAP7_75t_R output220 (.A(net220),
    .Y(u0_o[35]));
 BUFx3_ASAP7_75t_R output221 (.A(net221),
    .Y(u0_o[3]));
 BUFx3_ASAP7_75t_R output222 (.A(net222),
    .Y(u0_o[4]));
 BUFx3_ASAP7_75t_R output223 (.A(net223),
    .Y(u0_o[5]));
 BUFx3_ASAP7_75t_R output224 (.A(net224),
    .Y(u0_o[6]));
 BUFx3_ASAP7_75t_R output225 (.A(net225),
    .Y(u0_o[7]));
 BUFx3_ASAP7_75t_R output226 (.A(net226),
    .Y(u0_o[8]));
 BUFx3_ASAP7_75t_R output227 (.A(net227),
    .Y(u0_o[9]));
 BUFx3_ASAP7_75t_R output228 (.A(net228),
    .Y(u0_o_v));
 BUFx4_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_0_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_1_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_2_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_3_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_4_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_5_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_6_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_7_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_8_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_9_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_10_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_11_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_12_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_13_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_14_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_15_0_clk));
 BUFx12_ASAP7_75t_R clkload0 (.A(clknet_4_0_0_clk));
 INVxp67_ASAP7_75t_R clkload1 (.A(clknet_4_1_0_clk));
 BUFx24_ASAP7_75t_R clkload2 (.A(clknet_4_2_0_clk));
 INVx3_ASAP7_75t_R clkload3 (.A(clknet_4_3_0_clk));
 BUFx24_ASAP7_75t_R clkload4 (.A(clknet_4_4_0_clk));
 INVx3_ASAP7_75t_R clkload5 (.A(clknet_4_5_0_clk));
 INVx6_ASAP7_75t_R clkload6 (.A(clknet_4_6_0_clk));
 BUFx24_ASAP7_75t_R clkload7 (.A(clknet_4_7_0_clk));
 BUFx12_ASAP7_75t_R clkload8 (.A(clknet_4_8_0_clk));
 BUFx24_ASAP7_75t_R clkload9 (.A(clknet_4_9_0_clk));
 INVx3_ASAP7_75t_R clkload10 (.A(clknet_4_10_0_clk));
 INVx3_ASAP7_75t_R clkload11 (.A(clknet_4_11_0_clk));
 BUFx24_ASAP7_75t_R clkload12 (.A(clknet_4_12_0_clk));
 BUFx12_ASAP7_75t_R clkload13 (.A(clknet_4_13_0_clk));
 BUFx12_ASAP7_75t_R clkload14 (.A(clknet_4_14_0_clk));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24 ();
 FILLER_ASAP7_75t_R FILLER_0_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143 ();
 FILLER_ASAP7_75t_R FILLER_0_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201 ();
 DECAPx6_ASAP7_75t_R FILLER_0_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227 ();
 DECAPx10_ASAP7_75t_R FILLER_0_234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256 ();
 FILLER_ASAP7_75t_R FILLER_0_278 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx6_ASAP7_75t_R FILLER_1_24 ();
 DECAPx2_ASAP7_75t_R FILLER_1_120 ();
 FILLER_ASAP7_75t_R FILLER_1_126 ();
 DECAPx1_ASAP7_75t_R FILLER_1_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_144 ();
 DECAPx1_ASAP7_75t_R FILLER_1_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_161 ();
 DECAPx10_ASAP7_75t_R FILLER_1_180 ();
 FILLER_ASAP7_75t_R FILLER_1_202 ();
 DECAPx10_ASAP7_75t_R FILLER_1_210 ();
 DECAPx10_ASAP7_75t_R FILLER_1_232 ();
 DECAPx10_ASAP7_75t_R FILLER_1_254 ();
 DECAPx1_ASAP7_75t_R FILLER_1_276 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx6_ASAP7_75t_R FILLER_2_24 ();
 FILLER_ASAP7_75t_R FILLER_2_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_40 ();
 FILLER_ASAP7_75t_R FILLER_2_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_72 ();
 FILLER_ASAP7_75t_R FILLER_2_79 ();
 DECAPx1_ASAP7_75t_R FILLER_2_98 ();
 FILLER_ASAP7_75t_R FILLER_2_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_107 ();
 FILLER_ASAP7_75t_R FILLER_2_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_116 ();
 DECAPx2_ASAP7_75t_R FILLER_2_123 ();
 DECAPx2_ASAP7_75t_R FILLER_2_135 ();
 FILLER_ASAP7_75t_R FILLER_2_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_143 ();
 FILLER_ASAP7_75t_R FILLER_2_156 ();
 DECAPx4_ASAP7_75t_R FILLER_2_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_180 ();
 DECAPx10_ASAP7_75t_R FILLER_2_187 ();
 DECAPx10_ASAP7_75t_R FILLER_2_209 ();
 DECAPx10_ASAP7_75t_R FILLER_2_231 ();
 DECAPx10_ASAP7_75t_R FILLER_2_253 ();
 DECAPx1_ASAP7_75t_R FILLER_2_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_279 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx2_ASAP7_75t_R FILLER_3_24 ();
 FILLER_ASAP7_75t_R FILLER_3_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_50 ();
 FILLER_ASAP7_75t_R FILLER_3_59 ();
 DECAPx6_ASAP7_75t_R FILLER_3_101 ();
 DECAPx1_ASAP7_75t_R FILLER_3_115 ();
 DECAPx10_ASAP7_75t_R FILLER_3_122 ();
 DECAPx10_ASAP7_75t_R FILLER_3_144 ();
 DECAPx10_ASAP7_75t_R FILLER_3_166 ();
 DECAPx10_ASAP7_75t_R FILLER_3_188 ();
 DECAPx10_ASAP7_75t_R FILLER_3_210 ();
 DECAPx10_ASAP7_75t_R FILLER_3_232 ();
 DECAPx10_ASAP7_75t_R FILLER_3_254 ();
 DECAPx1_ASAP7_75t_R FILLER_3_276 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx1_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_71 ();
 DECAPx1_ASAP7_75t_R FILLER_4_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_97 ();
 DECAPx4_ASAP7_75t_R FILLER_4_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_128 ();
 DECAPx6_ASAP7_75t_R FILLER_4_138 ();
 DECAPx1_ASAP7_75t_R FILLER_4_152 ();
 FILLER_ASAP7_75t_R FILLER_4_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_178 ();
 DECAPx10_ASAP7_75t_R FILLER_4_182 ();
 FILLER_ASAP7_75t_R FILLER_4_204 ();
 DECAPx10_ASAP7_75t_R FILLER_4_226 ();
 DECAPx10_ASAP7_75t_R FILLER_4_248 ();
 DECAPx4_ASAP7_75t_R FILLER_4_270 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx4_ASAP7_75t_R FILLER_5_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_34 ();
 DECAPx6_ASAP7_75t_R FILLER_5_44 ();
 DECAPx1_ASAP7_75t_R FILLER_5_58 ();
 DECAPx1_ASAP7_75t_R FILLER_5_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_98 ();
 DECAPx6_ASAP7_75t_R FILLER_5_102 ();
 DECAPx2_ASAP7_75t_R FILLER_5_136 ();
 FILLER_ASAP7_75t_R FILLER_5_142 ();
 DECAPx2_ASAP7_75t_R FILLER_5_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_192 ();
 DECAPx1_ASAP7_75t_R FILLER_5_227 ();
 DECAPx10_ASAP7_75t_R FILLER_5_237 ();
 DECAPx6_ASAP7_75t_R FILLER_5_259 ();
 DECAPx2_ASAP7_75t_R FILLER_5_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_279 ();
 DECAPx6_ASAP7_75t_R FILLER_6_2 ();
 DECAPx1_ASAP7_75t_R FILLER_6_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_20 ();
 DECAPx6_ASAP7_75t_R FILLER_6_49 ();
 DECAPx1_ASAP7_75t_R FILLER_6_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_67 ();
 FILLER_ASAP7_75t_R FILLER_6_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_76 ();
 DECAPx1_ASAP7_75t_R FILLER_6_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_105 ();
 DECAPx4_ASAP7_75t_R FILLER_6_120 ();
 DECAPx4_ASAP7_75t_R FILLER_6_133 ();
 FILLER_ASAP7_75t_R FILLER_6_143 ();
 FILLER_ASAP7_75t_R FILLER_6_159 ();
 FILLER_ASAP7_75t_R FILLER_6_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_174 ();
 FILLER_ASAP7_75t_R FILLER_6_212 ();
 DECAPx10_ASAP7_75t_R FILLER_6_240 ();
 DECAPx6_ASAP7_75t_R FILLER_6_262 ();
 DECAPx1_ASAP7_75t_R FILLER_6_276 ();
 FILLER_ASAP7_75t_R FILLER_7_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_4 ();
 DECAPx2_ASAP7_75t_R FILLER_7_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_20 ();
 DECAPx2_ASAP7_75t_R FILLER_7_29 ();
 FILLER_ASAP7_75t_R FILLER_7_35 ();
 FILLER_ASAP7_75t_R FILLER_7_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_80 ();
 FILLER_ASAP7_75t_R FILLER_7_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_91 ();
 FILLER_ASAP7_75t_R FILLER_7_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_109 ();
 DECAPx10_ASAP7_75t_R FILLER_7_119 ();
 DECAPx6_ASAP7_75t_R FILLER_7_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_155 ();
 DECAPx2_ASAP7_75t_R FILLER_7_176 ();
 DECAPx6_ASAP7_75t_R FILLER_7_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_199 ();
 DECAPx4_ASAP7_75t_R FILLER_7_203 ();
 FILLER_ASAP7_75t_R FILLER_7_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_215 ();
 DECAPx1_ASAP7_75t_R FILLER_7_224 ();
 DECAPx2_ASAP7_75t_R FILLER_7_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_237 ();
 DECAPx10_ASAP7_75t_R FILLER_7_241 ();
 DECAPx6_ASAP7_75t_R FILLER_7_263 ();
 FILLER_ASAP7_75t_R FILLER_7_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_279 ();
 DECAPx1_ASAP7_75t_R FILLER_8_2 ();
 DECAPx2_ASAP7_75t_R FILLER_8_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_40 ();
 DECAPx1_ASAP7_75t_R FILLER_8_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_52 ();
 FILLER_ASAP7_75t_R FILLER_8_61 ();
 DECAPx2_ASAP7_75t_R FILLER_8_77 ();
 DECAPx4_ASAP7_75t_R FILLER_8_123 ();
 FILLER_ASAP7_75t_R FILLER_8_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_135 ();
 DECAPx4_ASAP7_75t_R FILLER_8_139 ();
 FILLER_ASAP7_75t_R FILLER_8_149 ();
 FILLER_ASAP7_75t_R FILLER_8_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_163 ();
 DECAPx1_ASAP7_75t_R FILLER_8_172 ();
 FILLER_ASAP7_75t_R FILLER_8_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_184 ();
 DECAPx2_ASAP7_75t_R FILLER_8_205 ();
 FILLER_ASAP7_75t_R FILLER_8_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_213 ();
 FILLER_ASAP7_75t_R FILLER_8_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_224 ();
 DECAPx6_ASAP7_75t_R FILLER_8_231 ();
 DECAPx1_ASAP7_75t_R FILLER_8_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_249 ();
 DECAPx10_ASAP7_75t_R FILLER_8_256 ();
 FILLER_ASAP7_75t_R FILLER_8_278 ();
 DECAPx4_ASAP7_75t_R FILLER_9_2 ();
 FILLER_ASAP7_75t_R FILLER_9_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_20 ();
 DECAPx2_ASAP7_75t_R FILLER_9_27 ();
 FILLER_ASAP7_75t_R FILLER_9_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_35 ();
 DECAPx2_ASAP7_75t_R FILLER_9_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_54 ();
 DECAPx1_ASAP7_75t_R FILLER_9_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_66 ();
 DECAPx6_ASAP7_75t_R FILLER_9_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_110 ();
 DECAPx4_ASAP7_75t_R FILLER_9_117 ();
 FILLER_ASAP7_75t_R FILLER_9_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_158 ();
 FILLER_ASAP7_75t_R FILLER_9_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_201 ();
 DECAPx2_ASAP7_75t_R FILLER_9_205 ();
 FILLER_ASAP7_75t_R FILLER_9_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_234 ();
 DECAPx10_ASAP7_75t_R FILLER_9_255 ();
 FILLER_ASAP7_75t_R FILLER_9_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_279 ();
 DECAPx2_ASAP7_75t_R FILLER_10_2 ();
 DECAPx1_ASAP7_75t_R FILLER_10_20 ();
 FILLER_ASAP7_75t_R FILLER_10_30 ();
 FILLER_ASAP7_75t_R FILLER_10_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_48 ();
 FILLER_ASAP7_75t_R FILLER_10_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_58 ();
 FILLER_ASAP7_75t_R FILLER_10_77 ();
 FILLER_ASAP7_75t_R FILLER_10_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_101 ();
 DECAPx10_ASAP7_75t_R FILLER_10_122 ();
 FILLER_ASAP7_75t_R FILLER_10_144 ();
 DECAPx2_ASAP7_75t_R FILLER_10_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_158 ();
 FILLER_ASAP7_75t_R FILLER_10_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_181 ();
 DECAPx10_ASAP7_75t_R FILLER_10_188 ();
 DECAPx10_ASAP7_75t_R FILLER_10_210 ();
 DECAPx10_ASAP7_75t_R FILLER_10_232 ();
 DECAPx10_ASAP7_75t_R FILLER_10_254 ();
 DECAPx1_ASAP7_75t_R FILLER_10_276 ();
 FILLER_ASAP7_75t_R FILLER_11_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_27 ();
 DECAPx6_ASAP7_75t_R FILLER_11_42 ();
 FILLER_ASAP7_75t_R FILLER_11_91 ();
 DECAPx1_ASAP7_75t_R FILLER_11_101 ();
 DECAPx4_ASAP7_75t_R FILLER_11_111 ();
 FILLER_ASAP7_75t_R FILLER_11_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_129 ();
 DECAPx2_ASAP7_75t_R FILLER_11_136 ();
 FILLER_ASAP7_75t_R FILLER_11_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_182 ();
 FILLER_ASAP7_75t_R FILLER_11_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_190 ();
 DECAPx2_ASAP7_75t_R FILLER_11_203 ();
 FILLER_ASAP7_75t_R FILLER_11_209 ();
 DECAPx2_ASAP7_75t_R FILLER_11_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_230 ();
 FILLER_ASAP7_75t_R FILLER_11_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_247 ();
 DECAPx1_ASAP7_75t_R FILLER_11_254 ();
 DECAPx2_ASAP7_75t_R FILLER_11_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_267 ();
 DECAPx2_ASAP7_75t_R FILLER_11_274 ();
 FILLER_ASAP7_75t_R FILLER_12_2 ();
 DECAPx1_ASAP7_75t_R FILLER_12_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_18 ();
 FILLER_ASAP7_75t_R FILLER_12_25 ();
 DECAPx2_ASAP7_75t_R FILLER_12_41 ();
 FILLER_ASAP7_75t_R FILLER_12_47 ();
 DECAPx2_ASAP7_75t_R FILLER_12_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_62 ();
 FILLER_ASAP7_75t_R FILLER_12_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_87 ();
 DECAPx4_ASAP7_75t_R FILLER_12_114 ();
 FILLER_ASAP7_75t_R FILLER_12_127 ();
 DECAPx1_ASAP7_75t_R FILLER_12_137 ();
 DECAPx1_ASAP7_75t_R FILLER_12_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_148 ();
 DECAPx1_ASAP7_75t_R FILLER_12_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_209 ();
 DECAPx2_ASAP7_75t_R FILLER_12_236 ();
 DECAPx2_ASAP7_75t_R FILLER_12_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_254 ();
 DECAPx1_ASAP7_75t_R FILLER_12_258 ();
 DECAPx4_ASAP7_75t_R FILLER_12_268 ();
 FILLER_ASAP7_75t_R FILLER_12_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_14 ();
 FILLER_ASAP7_75t_R FILLER_13_27 ();
 DECAPx6_ASAP7_75t_R FILLER_13_35 ();
 FILLER_ASAP7_75t_R FILLER_13_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_51 ();
 FILLER_ASAP7_75t_R FILLER_13_58 ();
 DECAPx4_ASAP7_75t_R FILLER_13_80 ();
 FILLER_ASAP7_75t_R FILLER_13_90 ();
 FILLER_ASAP7_75t_R FILLER_13_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_117 ();
 DECAPx1_ASAP7_75t_R FILLER_13_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_142 ();
 DECAPx4_ASAP7_75t_R FILLER_13_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_167 ();
 DECAPx4_ASAP7_75t_R FILLER_13_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_229 ();
 DECAPx2_ASAP7_75t_R FILLER_13_250 ();
 DECAPx4_ASAP7_75t_R FILLER_13_268 ();
 FILLER_ASAP7_75t_R FILLER_13_278 ();
 DECAPx10_ASAP7_75t_R FILLER_14_30 ();
 DECAPx4_ASAP7_75t_R FILLER_14_52 ();
 FILLER_ASAP7_75t_R FILLER_14_62 ();
 DECAPx1_ASAP7_75t_R FILLER_14_67 ();
 DECAPx1_ASAP7_75t_R FILLER_14_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_89 ();
 DECAPx2_ASAP7_75t_R FILLER_14_98 ();
 FILLER_ASAP7_75t_R FILLER_14_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_106 ();
 DECAPx2_ASAP7_75t_R FILLER_14_113 ();
 FILLER_ASAP7_75t_R FILLER_14_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_121 ();
 DECAPx1_ASAP7_75t_R FILLER_14_125 ();
 DECAPx2_ASAP7_75t_R FILLER_14_135 ();
 FILLER_ASAP7_75t_R FILLER_14_141 ();
 DECAPx6_ASAP7_75t_R FILLER_14_158 ();
 DECAPx1_ASAP7_75t_R FILLER_14_172 ();
 FILLER_ASAP7_75t_R FILLER_14_190 ();
 DECAPx4_ASAP7_75t_R FILLER_14_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_223 ();
 DECAPx1_ASAP7_75t_R FILLER_14_230 ();
 DECAPx10_ASAP7_75t_R FILLER_14_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_264 ();
 FILLER_ASAP7_75t_R FILLER_14_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_279 ();
 FILLER_ASAP7_75t_R FILLER_15_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_4 ();
 FILLER_ASAP7_75t_R FILLER_15_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_35 ();
 FILLER_ASAP7_75t_R FILLER_15_42 ();
 DECAPx2_ASAP7_75t_R FILLER_15_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_90 ();
 DECAPx6_ASAP7_75t_R FILLER_15_111 ();
 DECAPx1_ASAP7_75t_R FILLER_15_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_129 ();
 DECAPx1_ASAP7_75t_R FILLER_15_138 ();
 DECAPx2_ASAP7_75t_R FILLER_15_145 ();
 FILLER_ASAP7_75t_R FILLER_15_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_153 ();
 DECAPx6_ASAP7_75t_R FILLER_15_160 ();
 FILLER_ASAP7_75t_R FILLER_15_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_196 ();
 FILLER_ASAP7_75t_R FILLER_15_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_207 ();
 FILLER_ASAP7_75t_R FILLER_15_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_238 ();
 DECAPx4_ASAP7_75t_R FILLER_15_268 ();
 FILLER_ASAP7_75t_R FILLER_15_278 ();
 FILLER_ASAP7_75t_R FILLER_16_48 ();
 DECAPx1_ASAP7_75t_R FILLER_16_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_62 ();
 DECAPx10_ASAP7_75t_R FILLER_16_70 ();
 DECAPx2_ASAP7_75t_R FILLER_16_92 ();
 FILLER_ASAP7_75t_R FILLER_16_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_100 ();
 DECAPx10_ASAP7_75t_R FILLER_16_104 ();
 FILLER_ASAP7_75t_R FILLER_16_126 ();
 DECAPx4_ASAP7_75t_R FILLER_16_180 ();
 FILLER_ASAP7_75t_R FILLER_16_190 ();
 DECAPx2_ASAP7_75t_R FILLER_16_268 ();
 DECAPx2_ASAP7_75t_R FILLER_17_14 ();
 DECAPx1_ASAP7_75t_R FILLER_17_34 ();
 FILLER_ASAP7_75t_R FILLER_17_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_47 ();
 FILLER_ASAP7_75t_R FILLER_17_60 ();
 FILLER_ASAP7_75t_R FILLER_17_82 ();
 FILLER_ASAP7_75t_R FILLER_17_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_92 ();
 DECAPx2_ASAP7_75t_R FILLER_17_107 ();
 DECAPx10_ASAP7_75t_R FILLER_17_137 ();
 DECAPx2_ASAP7_75t_R FILLER_17_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_190 ();
 DECAPx4_ASAP7_75t_R FILLER_17_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_231 ();
 DECAPx1_ASAP7_75t_R FILLER_17_244 ();
 DECAPx6_ASAP7_75t_R FILLER_17_251 ();
 FILLER_ASAP7_75t_R FILLER_17_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_11 ();
 FILLER_ASAP7_75t_R FILLER_18_38 ();
 DECAPx6_ASAP7_75t_R FILLER_18_52 ();
 FILLER_ASAP7_75t_R FILLER_18_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_103 ();
 DECAPx10_ASAP7_75t_R FILLER_18_114 ();
 DECAPx10_ASAP7_75t_R FILLER_18_136 ();
 DECAPx2_ASAP7_75t_R FILLER_18_158 ();
 FILLER_ASAP7_75t_R FILLER_18_164 ();
 FILLER_ASAP7_75t_R FILLER_18_174 ();
 DECAPx2_ASAP7_75t_R FILLER_18_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_228 ();
 DECAPx6_ASAP7_75t_R FILLER_18_260 ();
 DECAPx2_ASAP7_75t_R FILLER_19_8 ();
 FILLER_ASAP7_75t_R FILLER_19_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_34 ();
 DECAPx6_ASAP7_75t_R FILLER_19_43 ();
 DECAPx1_ASAP7_75t_R FILLER_19_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_71 ();
 DECAPx6_ASAP7_75t_R FILLER_19_115 ();
 FILLER_ASAP7_75t_R FILLER_19_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_131 ();
 DECAPx2_ASAP7_75t_R FILLER_19_152 ();
 FILLER_ASAP7_75t_R FILLER_19_158 ();
 DECAPx6_ASAP7_75t_R FILLER_19_170 ();
 DECAPx1_ASAP7_75t_R FILLER_19_184 ();
 DECAPx1_ASAP7_75t_R FILLER_19_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_218 ();
 DECAPx10_ASAP7_75t_R FILLER_19_226 ();
 DECAPx6_ASAP7_75t_R FILLER_19_248 ();
 DECAPx1_ASAP7_75t_R FILLER_19_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_279 ();
 DECAPx1_ASAP7_75t_R FILLER_20_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_12 ();
 DECAPx1_ASAP7_75t_R FILLER_20_31 ();
 DECAPx6_ASAP7_75t_R FILLER_20_48 ();
 FILLER_ASAP7_75t_R FILLER_20_62 ();
 DECAPx1_ASAP7_75t_R FILLER_20_82 ();
 DECAPx10_ASAP7_75t_R FILLER_20_103 ();
 DECAPx6_ASAP7_75t_R FILLER_20_125 ();
 FILLER_ASAP7_75t_R FILLER_20_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_141 ();
 DECAPx10_ASAP7_75t_R FILLER_20_152 ();
 DECAPx6_ASAP7_75t_R FILLER_20_174 ();
 FILLER_ASAP7_75t_R FILLER_20_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_190 ();
 DECAPx4_ASAP7_75t_R FILLER_20_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_224 ();
 FILLER_ASAP7_75t_R FILLER_20_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_233 ();
 DECAPx2_ASAP7_75t_R FILLER_20_248 ();
 DECAPx2_ASAP7_75t_R FILLER_20_266 ();
 FILLER_ASAP7_75t_R FILLER_20_278 ();
 DECAPx1_ASAP7_75t_R FILLER_21_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_12 ();
 FILLER_ASAP7_75t_R FILLER_21_29 ();
 FILLER_ASAP7_75t_R FILLER_21_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_95 ();
 FILLER_ASAP7_75t_R FILLER_21_104 ();
 DECAPx1_ASAP7_75t_R FILLER_21_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_116 ();
 DECAPx10_ASAP7_75t_R FILLER_21_127 ();
 DECAPx10_ASAP7_75t_R FILLER_21_149 ();
 DECAPx6_ASAP7_75t_R FILLER_21_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_185 ();
 DECAPx6_ASAP7_75t_R FILLER_21_199 ();
 DECAPx1_ASAP7_75t_R FILLER_21_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_217 ();
 DECAPx1_ASAP7_75t_R FILLER_21_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_235 ();
 DECAPx2_ASAP7_75t_R FILLER_21_259 ();
 FILLER_ASAP7_75t_R FILLER_21_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_279 ();
 FILLER_ASAP7_75t_R FILLER_22_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_22 ();
 FILLER_ASAP7_75t_R FILLER_22_31 ();
 DECAPx6_ASAP7_75t_R FILLER_22_51 ();
 FILLER_ASAP7_75t_R FILLER_22_65 ();
 DECAPx10_ASAP7_75t_R FILLER_22_117 ();
 DECAPx2_ASAP7_75t_R FILLER_22_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_145 ();
 DECAPx10_ASAP7_75t_R FILLER_22_156 ();
 DECAPx10_ASAP7_75t_R FILLER_22_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_200 ();
 FILLER_ASAP7_75t_R FILLER_22_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_233 ();
 DECAPx1_ASAP7_75t_R FILLER_22_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_252 ();
 DECAPx2_ASAP7_75t_R FILLER_22_259 ();
 FILLER_ASAP7_75t_R FILLER_22_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_267 ();
 FILLER_ASAP7_75t_R FILLER_23_31 ();
 DECAPx2_ASAP7_75t_R FILLER_23_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_47 ();
 FILLER_ASAP7_75t_R FILLER_23_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_56 ();
 DECAPx10_ASAP7_75t_R FILLER_23_77 ();
 DECAPx10_ASAP7_75t_R FILLER_23_99 ();
 DECAPx6_ASAP7_75t_R FILLER_23_121 ();
 FILLER_ASAP7_75t_R FILLER_23_135 ();
 DECAPx1_ASAP7_75t_R FILLER_23_147 ();
 DECAPx6_ASAP7_75t_R FILLER_23_161 ();
 DECAPx2_ASAP7_75t_R FILLER_23_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_181 ();
 DECAPx2_ASAP7_75t_R FILLER_23_202 ();
 FILLER_ASAP7_75t_R FILLER_23_214 ();
 DECAPx2_ASAP7_75t_R FILLER_23_228 ();
 FILLER_ASAP7_75t_R FILLER_23_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_236 ();
 FILLER_ASAP7_75t_R FILLER_23_266 ();
 DECAPx10_ASAP7_75t_R FILLER_24_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_30 ();
 DECAPx6_ASAP7_75t_R FILLER_24_37 ();
 DECAPx2_ASAP7_75t_R FILLER_24_51 ();
 FILLER_ASAP7_75t_R FILLER_24_77 ();
 DECAPx2_ASAP7_75t_R FILLER_24_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_91 ();
 DECAPx4_ASAP7_75t_R FILLER_24_100 ();
 DECAPx4_ASAP7_75t_R FILLER_24_120 ();
 DECAPx10_ASAP7_75t_R FILLER_24_156 ();
 DECAPx2_ASAP7_75t_R FILLER_24_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_184 ();
 DECAPx6_ASAP7_75t_R FILLER_24_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_211 ();
 DECAPx1_ASAP7_75t_R FILLER_24_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_222 ();
 FILLER_ASAP7_75t_R FILLER_24_229 ();
 DECAPx2_ASAP7_75t_R FILLER_24_251 ();
 FILLER_ASAP7_75t_R FILLER_24_263 ();
 FILLER_ASAP7_75t_R FILLER_24_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_17 ();
 DECAPx1_ASAP7_75t_R FILLER_25_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_28 ();
 DECAPx6_ASAP7_75t_R FILLER_25_43 ();
 DECAPx2_ASAP7_75t_R FILLER_25_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_63 ();
 DECAPx2_ASAP7_75t_R FILLER_25_78 ();
 DECAPx6_ASAP7_75t_R FILLER_25_97 ();
 DECAPx2_ASAP7_75t_R FILLER_25_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_138 ();
 DECAPx1_ASAP7_75t_R FILLER_25_142 ();
 DECAPx10_ASAP7_75t_R FILLER_25_156 ();
 DECAPx4_ASAP7_75t_R FILLER_25_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_206 ();
 DECAPx2_ASAP7_75t_R FILLER_25_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_243 ();
 FILLER_ASAP7_75t_R FILLER_25_250 ();
 DECAPx10_ASAP7_75t_R FILLER_25_255 ();
 FILLER_ASAP7_75t_R FILLER_25_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_279 ();
 DECAPx6_ASAP7_75t_R FILLER_26_8 ();
 DECAPx1_ASAP7_75t_R FILLER_26_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_26 ();
 DECAPx1_ASAP7_75t_R FILLER_26_30 ();
 DECAPx4_ASAP7_75t_R FILLER_26_54 ();
 FILLER_ASAP7_75t_R FILLER_26_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_66 ();
 DECAPx6_ASAP7_75t_R FILLER_26_102 ();
 DECAPx2_ASAP7_75t_R FILLER_26_124 ();
 DECAPx1_ASAP7_75t_R FILLER_26_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_140 ();
 DECAPx4_ASAP7_75t_R FILLER_26_151 ();
 FILLER_ASAP7_75t_R FILLER_26_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_163 ();
 DECAPx10_ASAP7_75t_R FILLER_26_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_192 ();
 DECAPx6_ASAP7_75t_R FILLER_26_199 ();
 DECAPx1_ASAP7_75t_R FILLER_26_236 ();
 DECAPx4_ASAP7_75t_R FILLER_26_249 ();
 FILLER_ASAP7_75t_R FILLER_26_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_261 ();
 DECAPx2_ASAP7_75t_R FILLER_26_268 ();
 DECAPx2_ASAP7_75t_R FILLER_27_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_14 ();
 DECAPx1_ASAP7_75t_R FILLER_27_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_25 ();
 FILLER_ASAP7_75t_R FILLER_27_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_46 ();
 DECAPx2_ASAP7_75t_R FILLER_27_55 ();
 FILLER_ASAP7_75t_R FILLER_27_61 ();
 DECAPx10_ASAP7_75t_R FILLER_27_79 ();
 DECAPx6_ASAP7_75t_R FILLER_27_101 ();
 DECAPx1_ASAP7_75t_R FILLER_27_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_119 ();
 DECAPx2_ASAP7_75t_R FILLER_27_131 ();
 FILLER_ASAP7_75t_R FILLER_27_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_139 ();
 DECAPx10_ASAP7_75t_R FILLER_27_150 ();
 DECAPx6_ASAP7_75t_R FILLER_27_172 ();
 DECAPx1_ASAP7_75t_R FILLER_27_186 ();
 DECAPx2_ASAP7_75t_R FILLER_27_210 ();
 DECAPx1_ASAP7_75t_R FILLER_27_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_226 ();
 FILLER_ASAP7_75t_R FILLER_27_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_266 ();
 DECAPx2_ASAP7_75t_R FILLER_27_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_279 ();
 DECAPx1_ASAP7_75t_R FILLER_28_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_38 ();
 FILLER_ASAP7_75t_R FILLER_28_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_68 ();
 FILLER_ASAP7_75t_R FILLER_28_75 ();
 FILLER_ASAP7_75t_R FILLER_28_88 ();
 DECAPx1_ASAP7_75t_R FILLER_28_96 ();
 DECAPx10_ASAP7_75t_R FILLER_28_135 ();
 DECAPx6_ASAP7_75t_R FILLER_28_157 ();
 FILLER_ASAP7_75t_R FILLER_28_171 ();
 DECAPx4_ASAP7_75t_R FILLER_28_183 ();
 FILLER_ASAP7_75t_R FILLER_28_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_195 ();
 DECAPx10_ASAP7_75t_R FILLER_28_224 ();
 DECAPx6_ASAP7_75t_R FILLER_28_246 ();
 DECAPx1_ASAP7_75t_R FILLER_28_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_264 ();
 DECAPx10_ASAP7_75t_R FILLER_29_2 ();
 DECAPx1_ASAP7_75t_R FILLER_29_30 ();
 DECAPx1_ASAP7_75t_R FILLER_29_40 ();
 FILLER_ASAP7_75t_R FILLER_29_50 ();
 FILLER_ASAP7_75t_R FILLER_29_72 ();
 DECAPx1_ASAP7_75t_R FILLER_29_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_107 ();
 FILLER_ASAP7_75t_R FILLER_29_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_122 ();
 DECAPx10_ASAP7_75t_R FILLER_29_143 ();
 DECAPx6_ASAP7_75t_R FILLER_29_165 ();
 DECAPx2_ASAP7_75t_R FILLER_29_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_185 ();
 DECAPx4_ASAP7_75t_R FILLER_29_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_222 ();
 FILLER_ASAP7_75t_R FILLER_29_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_228 ();
 DECAPx1_ASAP7_75t_R FILLER_29_237 ();
 DECAPx6_ASAP7_75t_R FILLER_29_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_261 ();
 DECAPx2_ASAP7_75t_R FILLER_29_274 ();
 DECAPx2_ASAP7_75t_R FILLER_30_2 ();
 FILLER_ASAP7_75t_R FILLER_30_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_22 ();
 DECAPx2_ASAP7_75t_R FILLER_30_32 ();
 DECAPx10_ASAP7_75t_R FILLER_30_46 ();
 DECAPx10_ASAP7_75t_R FILLER_30_68 ();
 DECAPx10_ASAP7_75t_R FILLER_30_90 ();
 DECAPx1_ASAP7_75t_R FILLER_30_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_116 ();
 DECAPx6_ASAP7_75t_R FILLER_30_120 ();
 DECAPx2_ASAP7_75t_R FILLER_30_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_140 ();
 DECAPx4_ASAP7_75t_R FILLER_30_161 ();
 DECAPx2_ASAP7_75t_R FILLER_30_174 ();
 DECAPx10_ASAP7_75t_R FILLER_30_186 ();
 DECAPx10_ASAP7_75t_R FILLER_30_208 ();
 FILLER_ASAP7_75t_R FILLER_30_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_252 ();
 DECAPx4_ASAP7_75t_R FILLER_30_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_273 ();
 DECAPx2_ASAP7_75t_R FILLER_31_8 ();
 FILLER_ASAP7_75t_R FILLER_31_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_16 ();
 DECAPx2_ASAP7_75t_R FILLER_31_23 ();
 FILLER_ASAP7_75t_R FILLER_31_29 ();
 DECAPx4_ASAP7_75t_R FILLER_31_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_67 ();
 DECAPx2_ASAP7_75t_R FILLER_31_74 ();
 DECAPx10_ASAP7_75t_R FILLER_31_107 ();
 DECAPx4_ASAP7_75t_R FILLER_31_129 ();
 FILLER_ASAP7_75t_R FILLER_31_139 ();
 DECAPx2_ASAP7_75t_R FILLER_31_149 ();
 DECAPx2_ASAP7_75t_R FILLER_31_161 ();
 FILLER_ASAP7_75t_R FILLER_31_167 ();
 DECAPx10_ASAP7_75t_R FILLER_31_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_207 ();
 DECAPx10_ASAP7_75t_R FILLER_31_214 ();
 DECAPx4_ASAP7_75t_R FILLER_31_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_246 ();
 DECAPx10_ASAP7_75t_R FILLER_31_256 ();
 FILLER_ASAP7_75t_R FILLER_31_278 ();
 DECAPx2_ASAP7_75t_R FILLER_32_2 ();
 FILLER_ASAP7_75t_R FILLER_32_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_10 ();
 DECAPx10_ASAP7_75t_R FILLER_32_17 ();
 DECAPx2_ASAP7_75t_R FILLER_32_39 ();
 FILLER_ASAP7_75t_R FILLER_32_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_77 ();
 FILLER_ASAP7_75t_R FILLER_32_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_92 ();
 FILLER_ASAP7_75t_R FILLER_32_99 ();
 DECAPx1_ASAP7_75t_R FILLER_32_109 ();
 DECAPx1_ASAP7_75t_R FILLER_32_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_123 ();
 DECAPx2_ASAP7_75t_R FILLER_32_132 ();
 DECAPx6_ASAP7_75t_R FILLER_32_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_158 ();
 DECAPx6_ASAP7_75t_R FILLER_32_162 ();
 DECAPx2_ASAP7_75t_R FILLER_32_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_182 ();
 DECAPx2_ASAP7_75t_R FILLER_32_201 ();
 DECAPx6_ASAP7_75t_R FILLER_32_233 ();
 DECAPx6_ASAP7_75t_R FILLER_32_250 ();
 DECAPx1_ASAP7_75t_R FILLER_32_264 ();
 DECAPx2_ASAP7_75t_R FILLER_32_274 ();
 DECAPx1_ASAP7_75t_R FILLER_33_2 ();
 FILLER_ASAP7_75t_R FILLER_33_12 ();
 DECAPx1_ASAP7_75t_R FILLER_33_20 ();
 FILLER_ASAP7_75t_R FILLER_33_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_32 ();
 FILLER_ASAP7_75t_R FILLER_33_56 ();
 FILLER_ASAP7_75t_R FILLER_33_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_71 ();
 DECAPx1_ASAP7_75t_R FILLER_33_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_82 ();
 DECAPx4_ASAP7_75t_R FILLER_33_89 ();
 FILLER_ASAP7_75t_R FILLER_33_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_101 ();
 DECAPx2_ASAP7_75t_R FILLER_33_181 ();
 DECAPx6_ASAP7_75t_R FILLER_33_190 ();
 DECAPx1_ASAP7_75t_R FILLER_33_204 ();
 DECAPx1_ASAP7_75t_R FILLER_33_224 ();
 DECAPx4_ASAP7_75t_R FILLER_33_248 ();
 DECAPx6_ASAP7_75t_R FILLER_33_264 ();
 FILLER_ASAP7_75t_R FILLER_33_278 ();
 DECAPx10_ASAP7_75t_R FILLER_34_2 ();
 DECAPx2_ASAP7_75t_R FILLER_34_24 ();
 FILLER_ASAP7_75t_R FILLER_34_30 ();
 DECAPx1_ASAP7_75t_R FILLER_34_62 ();
 DECAPx1_ASAP7_75t_R FILLER_34_79 ();
 FILLER_ASAP7_75t_R FILLER_34_91 ();
 DECAPx1_ASAP7_75t_R FILLER_34_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_100 ();
 FILLER_ASAP7_75t_R FILLER_34_107 ();
 FILLER_ASAP7_75t_R FILLER_34_115 ();
 DECAPx2_ASAP7_75t_R FILLER_34_125 ();
 DECAPx4_ASAP7_75t_R FILLER_34_137 ();
 FILLER_ASAP7_75t_R FILLER_34_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_149 ();
 DECAPx10_ASAP7_75t_R FILLER_34_170 ();
 DECAPx10_ASAP7_75t_R FILLER_34_192 ();
 DECAPx10_ASAP7_75t_R FILLER_34_214 ();
 DECAPx10_ASAP7_75t_R FILLER_34_236 ();
 DECAPx10_ASAP7_75t_R FILLER_34_258 ();
 DECAPx1_ASAP7_75t_R FILLER_35_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_6 ();
 DECAPx10_ASAP7_75t_R FILLER_35_36 ();
 DECAPx1_ASAP7_75t_R FILLER_35_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_100 ();
 DECAPx1_ASAP7_75t_R FILLER_35_115 ();
 DECAPx2_ASAP7_75t_R FILLER_35_139 ();
 FILLER_ASAP7_75t_R FILLER_35_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_147 ();
 DECAPx2_ASAP7_75t_R FILLER_35_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_162 ();
 DECAPx2_ASAP7_75t_R FILLER_35_187 ();
 DECAPx4_ASAP7_75t_R FILLER_35_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_219 ();
 DECAPx10_ASAP7_75t_R FILLER_35_226 ();
 DECAPx1_ASAP7_75t_R FILLER_35_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_255 ();
 DECAPx6_ASAP7_75t_R FILLER_35_262 ();
 DECAPx1_ASAP7_75t_R FILLER_35_276 ();
 DECAPx10_ASAP7_75t_R FILLER_36_2 ();
 FILLER_ASAP7_75t_R FILLER_36_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_26 ();
 DECAPx10_ASAP7_75t_R FILLER_36_39 ();
 DECAPx6_ASAP7_75t_R FILLER_36_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_75 ();
 FILLER_ASAP7_75t_R FILLER_36_92 ();
 DECAPx4_ASAP7_75t_R FILLER_36_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_141 ();
 DECAPx1_ASAP7_75t_R FILLER_36_155 ();
 FILLER_ASAP7_75t_R FILLER_36_199 ();
 DECAPx1_ASAP7_75t_R FILLER_36_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_213 ();
 DECAPx10_ASAP7_75t_R FILLER_36_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_260 ();
 DECAPx2_ASAP7_75t_R FILLER_36_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_279 ();
 DECAPx10_ASAP7_75t_R FILLER_37_2 ();
 DECAPx2_ASAP7_75t_R FILLER_37_24 ();
 FILLER_ASAP7_75t_R FILLER_37_30 ();
 DECAPx2_ASAP7_75t_R FILLER_37_52 ();
 FILLER_ASAP7_75t_R FILLER_37_58 ();
 DECAPx2_ASAP7_75t_R FILLER_37_70 ();
 FILLER_ASAP7_75t_R FILLER_37_90 ();
 DECAPx2_ASAP7_75t_R FILLER_37_112 ();
 FILLER_ASAP7_75t_R FILLER_37_134 ();
 DECAPx2_ASAP7_75t_R FILLER_37_152 ();
 FILLER_ASAP7_75t_R FILLER_37_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_168 ();
 FILLER_ASAP7_75t_R FILLER_37_207 ();
 DECAPx1_ASAP7_75t_R FILLER_37_223 ();
 FILLER_ASAP7_75t_R FILLER_37_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_255 ();
 DECAPx2_ASAP7_75t_R FILLER_37_268 ();
 DECAPx2_ASAP7_75t_R FILLER_38_8 ();
 DECAPx2_ASAP7_75t_R FILLER_38_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_26 ();
 DECAPx2_ASAP7_75t_R FILLER_38_37 ();
 FILLER_ASAP7_75t_R FILLER_38_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_45 ();
 FILLER_ASAP7_75t_R FILLER_38_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_97 ();
 FILLER_ASAP7_75t_R FILLER_38_126 ();
 FILLER_ASAP7_75t_R FILLER_38_141 ();
 DECAPx1_ASAP7_75t_R FILLER_38_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_153 ();
 FILLER_ASAP7_75t_R FILLER_38_160 ();
 FILLER_ASAP7_75t_R FILLER_38_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_184 ();
 FILLER_ASAP7_75t_R FILLER_38_198 ();
 DECAPx1_ASAP7_75t_R FILLER_38_220 ();
 DECAPx10_ASAP7_75t_R FILLER_38_232 ();
 DECAPx4_ASAP7_75t_R FILLER_38_254 ();
 FILLER_ASAP7_75t_R FILLER_38_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_266 ();
 DECAPx2_ASAP7_75t_R FILLER_38_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_279 ();
 DECAPx10_ASAP7_75t_R FILLER_39_2 ();
 FILLER_ASAP7_75t_R FILLER_39_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_26 ();
 DECAPx6_ASAP7_75t_R FILLER_39_35 ();
 DECAPx1_ASAP7_75t_R FILLER_39_49 ();
 DECAPx2_ASAP7_75t_R FILLER_39_69 ();
 FILLER_ASAP7_75t_R FILLER_39_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_85 ();
 DECAPx10_ASAP7_75t_R FILLER_39_95 ();
 DECAPx2_ASAP7_75t_R FILLER_39_117 ();
 FILLER_ASAP7_75t_R FILLER_39_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_125 ();
 DECAPx2_ASAP7_75t_R FILLER_39_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_138 ();
 DECAPx1_ASAP7_75t_R FILLER_39_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_151 ();
 DECAPx4_ASAP7_75t_R FILLER_39_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_169 ();
 DECAPx10_ASAP7_75t_R FILLER_39_176 ();
 DECAPx1_ASAP7_75t_R FILLER_39_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_202 ();
 DECAPx2_ASAP7_75t_R FILLER_39_216 ();
 DECAPx10_ASAP7_75t_R FILLER_39_242 ();
 DECAPx4_ASAP7_75t_R FILLER_39_264 ();
 DECAPx4_ASAP7_75t_R FILLER_40_2 ();
 FILLER_ASAP7_75t_R FILLER_40_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_14 ();
 FILLER_ASAP7_75t_R FILLER_40_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_40 ();
 DECAPx2_ASAP7_75t_R FILLER_40_66 ();
 FILLER_ASAP7_75t_R FILLER_40_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_74 ();
 DECAPx10_ASAP7_75t_R FILLER_40_85 ();
 DECAPx6_ASAP7_75t_R FILLER_40_107 ();
 FILLER_ASAP7_75t_R FILLER_40_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_123 ();
 FILLER_ASAP7_75t_R FILLER_40_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_134 ();
 DECAPx6_ASAP7_75t_R FILLER_40_151 ();
 DECAPx1_ASAP7_75t_R FILLER_40_165 ();
 DECAPx2_ASAP7_75t_R FILLER_40_199 ();
 DECAPx1_ASAP7_75t_R FILLER_40_212 ();
 DECAPx2_ASAP7_75t_R FILLER_40_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_228 ();
 DECAPx1_ASAP7_75t_R FILLER_40_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_259 ();
 DECAPx1_ASAP7_75t_R FILLER_40_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_273 ();
 FILLER_ASAP7_75t_R FILLER_41_2 ();
 DECAPx10_ASAP7_75t_R FILLER_41_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_42 ();
 DECAPx2_ASAP7_75t_R FILLER_41_49 ();
 FILLER_ASAP7_75t_R FILLER_41_55 ();
 DECAPx1_ASAP7_75t_R FILLER_41_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_79 ();
 DECAPx4_ASAP7_75t_R FILLER_41_94 ();
 DECAPx4_ASAP7_75t_R FILLER_41_133 ();
 DECAPx2_ASAP7_75t_R FILLER_41_153 ();
 FILLER_ASAP7_75t_R FILLER_41_179 ();
 DECAPx2_ASAP7_75t_R FILLER_41_204 ();
 FILLER_ASAP7_75t_R FILLER_41_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_212 ();
 DECAPx2_ASAP7_75t_R FILLER_41_233 ();
 FILLER_ASAP7_75t_R FILLER_41_239 ();
 DECAPx2_ASAP7_75t_R FILLER_41_247 ();
 DECAPx10_ASAP7_75t_R FILLER_41_256 ();
 FILLER_ASAP7_75t_R FILLER_41_278 ();
 DECAPx10_ASAP7_75t_R FILLER_42_2 ();
 DECAPx4_ASAP7_75t_R FILLER_42_24 ();
 FILLER_ASAP7_75t_R FILLER_42_34 ();
 DECAPx10_ASAP7_75t_R FILLER_42_53 ();
 DECAPx1_ASAP7_75t_R FILLER_42_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_79 ();
 DECAPx1_ASAP7_75t_R FILLER_42_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_117 ();
 FILLER_ASAP7_75t_R FILLER_42_130 ();
 DECAPx1_ASAP7_75t_R FILLER_42_135 ();
 DECAPx4_ASAP7_75t_R FILLER_42_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_155 ();
 DECAPx1_ASAP7_75t_R FILLER_42_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_191 ();
 DECAPx6_ASAP7_75t_R FILLER_42_206 ();
 DECAPx1_ASAP7_75t_R FILLER_42_220 ();
 DECAPx4_ASAP7_75t_R FILLER_42_268 ();
 FILLER_ASAP7_75t_R FILLER_42_278 ();
 DECAPx1_ASAP7_75t_R FILLER_43_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_6 ();
 DECAPx4_ASAP7_75t_R FILLER_43_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_32 ();
 FILLER_ASAP7_75t_R FILLER_43_39 ();
 DECAPx4_ASAP7_75t_R FILLER_43_47 ();
 FILLER_ASAP7_75t_R FILLER_43_57 ();
 FILLER_ASAP7_75t_R FILLER_43_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_67 ();
 DECAPx6_ASAP7_75t_R FILLER_43_78 ();
 FILLER_ASAP7_75t_R FILLER_43_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_94 ();
 DECAPx2_ASAP7_75t_R FILLER_43_114 ();
 DECAPx2_ASAP7_75t_R FILLER_43_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_161 ();
 FILLER_ASAP7_75t_R FILLER_43_192 ();
 DECAPx2_ASAP7_75t_R FILLER_43_214 ();
 DECAPx1_ASAP7_75t_R FILLER_43_240 ();
 DECAPx4_ASAP7_75t_R FILLER_43_250 ();
 FILLER_ASAP7_75t_R FILLER_43_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_262 ();
 FILLER_ASAP7_75t_R FILLER_43_266 ();
 DECAPx2_ASAP7_75t_R FILLER_43_274 ();
 DECAPx4_ASAP7_75t_R FILLER_44_2 ();
 FILLER_ASAP7_75t_R FILLER_44_12 ();
 DECAPx1_ASAP7_75t_R FILLER_44_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_41 ();
 DECAPx2_ASAP7_75t_R FILLER_44_52 ();
 FILLER_ASAP7_75t_R FILLER_44_78 ();
 FILLER_ASAP7_75t_R FILLER_44_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_88 ();
 FILLER_ASAP7_75t_R FILLER_44_99 ();
 DECAPx4_ASAP7_75t_R FILLER_44_114 ();
 FILLER_ASAP7_75t_R FILLER_44_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_134 ();
 DECAPx2_ASAP7_75t_R FILLER_44_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_190 ();
 DECAPx6_ASAP7_75t_R FILLER_44_202 ();
 FILLER_ASAP7_75t_R FILLER_44_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_218 ();
 FILLER_ASAP7_75t_R FILLER_44_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_229 ();
 DECAPx10_ASAP7_75t_R FILLER_44_258 ();
 DECAPx4_ASAP7_75t_R FILLER_45_2 ();
 FILLER_ASAP7_75t_R FILLER_45_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_14 ();
 DECAPx6_ASAP7_75t_R FILLER_45_21 ();
 DECAPx2_ASAP7_75t_R FILLER_45_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_47 ();
 FILLER_ASAP7_75t_R FILLER_45_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_78 ();
 FILLER_ASAP7_75t_R FILLER_45_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_93 ();
 DECAPx4_ASAP7_75t_R FILLER_45_110 ();
 FILLER_ASAP7_75t_R FILLER_45_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_122 ();
 DECAPx1_ASAP7_75t_R FILLER_45_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_133 ();
 DECAPx6_ASAP7_75t_R FILLER_45_140 ();
 DECAPx2_ASAP7_75t_R FILLER_45_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_169 ();
 DECAPx6_ASAP7_75t_R FILLER_45_176 ();
 FILLER_ASAP7_75t_R FILLER_45_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_192 ();
 DECAPx2_ASAP7_75t_R FILLER_45_199 ();
 FILLER_ASAP7_75t_R FILLER_45_212 ();
 DECAPx10_ASAP7_75t_R FILLER_45_226 ();
 DECAPx10_ASAP7_75t_R FILLER_45_248 ();
 DECAPx4_ASAP7_75t_R FILLER_45_270 ();
 DECAPx6_ASAP7_75t_R FILLER_46_2 ();
 FILLER_ASAP7_75t_R FILLER_46_16 ();
 DECAPx2_ASAP7_75t_R FILLER_46_24 ();
 FILLER_ASAP7_75t_R FILLER_46_40 ();
 FILLER_ASAP7_75t_R FILLER_46_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_50 ();
 DECAPx1_ASAP7_75t_R FILLER_46_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_69 ();
 DECAPx1_ASAP7_75t_R FILLER_46_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_82 ();
 DECAPx1_ASAP7_75t_R FILLER_46_90 ();
 FILLER_ASAP7_75t_R FILLER_46_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_113 ();
 FILLER_ASAP7_75t_R FILLER_46_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_132 ();
 DECAPx2_ASAP7_75t_R FILLER_46_139 ();
 FILLER_ASAP7_75t_R FILLER_46_145 ();
 DECAPx10_ASAP7_75t_R FILLER_46_160 ();
 DECAPx6_ASAP7_75t_R FILLER_46_182 ();
 FILLER_ASAP7_75t_R FILLER_46_196 ();
 FILLER_ASAP7_75t_R FILLER_46_211 ();
 DECAPx2_ASAP7_75t_R FILLER_46_219 ();
 FILLER_ASAP7_75t_R FILLER_46_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_227 ();
 DECAPx10_ASAP7_75t_R FILLER_46_236 ();
 DECAPx4_ASAP7_75t_R FILLER_46_258 ();
 DECAPx2_ASAP7_75t_R FILLER_46_274 ();
 DECAPx10_ASAP7_75t_R FILLER_47_2 ();
 DECAPx6_ASAP7_75t_R FILLER_47_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_52 ();
 DECAPx2_ASAP7_75t_R FILLER_47_62 ();
 FILLER_ASAP7_75t_R FILLER_47_68 ();
 DECAPx4_ASAP7_75t_R FILLER_47_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_86 ();
 DECAPx4_ASAP7_75t_R FILLER_47_106 ();
 FILLER_ASAP7_75t_R FILLER_47_116 ();
 DECAPx4_ASAP7_75t_R FILLER_47_128 ();
 FILLER_ASAP7_75t_R FILLER_47_146 ();
 DECAPx2_ASAP7_75t_R FILLER_47_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_168 ();
 DECAPx1_ASAP7_75t_R FILLER_47_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_193 ();
 FILLER_ASAP7_75t_R FILLER_47_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_224 ();
 DECAPx10_ASAP7_75t_R FILLER_47_251 ();
 DECAPx2_ASAP7_75t_R FILLER_47_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_279 ();
 DECAPx6_ASAP7_75t_R FILLER_48_2 ();
 DECAPx2_ASAP7_75t_R FILLER_48_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_22 ();
 DECAPx6_ASAP7_75t_R FILLER_48_33 ();
 FILLER_ASAP7_75t_R FILLER_48_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_49 ();
 DECAPx4_ASAP7_75t_R FILLER_48_54 ();
 FILLER_ASAP7_75t_R FILLER_48_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_66 ();
 DECAPx4_ASAP7_75t_R FILLER_48_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_83 ();
 DECAPx10_ASAP7_75t_R FILLER_48_90 ();
 DECAPx4_ASAP7_75t_R FILLER_48_112 ();
 FILLER_ASAP7_75t_R FILLER_48_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_152 ();
 DECAPx2_ASAP7_75t_R FILLER_48_161 ();
 FILLER_ASAP7_75t_R FILLER_48_167 ();
 DECAPx6_ASAP7_75t_R FILLER_48_183 ();
 DECAPx1_ASAP7_75t_R FILLER_48_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_215 ();
 DECAPx2_ASAP7_75t_R FILLER_48_222 ();
 DECAPx2_ASAP7_75t_R FILLER_48_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_242 ();
 DECAPx10_ASAP7_75t_R FILLER_48_246 ();
 DECAPx4_ASAP7_75t_R FILLER_48_268 ();
 FILLER_ASAP7_75t_R FILLER_48_278 ();
 DECAPx2_ASAP7_75t_R FILLER_49_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_8 ();
 FILLER_ASAP7_75t_R FILLER_49_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_83 ();
 DECAPx1_ASAP7_75t_R FILLER_49_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_112 ();
 DECAPx1_ASAP7_75t_R FILLER_49_142 ();
 FILLER_ASAP7_75t_R FILLER_49_152 ();
 FILLER_ASAP7_75t_R FILLER_49_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_168 ();
 DECAPx4_ASAP7_75t_R FILLER_49_175 ();
 FILLER_ASAP7_75t_R FILLER_49_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_187 ();
 DECAPx4_ASAP7_75t_R FILLER_49_194 ();
 DECAPx2_ASAP7_75t_R FILLER_49_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_216 ();
 FILLER_ASAP7_75t_R FILLER_49_223 ();
 DECAPx4_ASAP7_75t_R FILLER_49_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_261 ();
 DECAPx2_ASAP7_75t_R FILLER_49_271 ();
 FILLER_ASAP7_75t_R FILLER_49_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_279 ();
 DECAPx6_ASAP7_75t_R FILLER_50_2 ();
 DECAPx1_ASAP7_75t_R FILLER_50_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_20 ();
 FILLER_ASAP7_75t_R FILLER_50_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_45 ();
 FILLER_ASAP7_75t_R FILLER_50_54 ();
 DECAPx6_ASAP7_75t_R FILLER_50_72 ();
 FILLER_ASAP7_75t_R FILLER_50_86 ();
 DECAPx4_ASAP7_75t_R FILLER_50_91 ();
 FILLER_ASAP7_75t_R FILLER_50_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_103 ();
 DECAPx1_ASAP7_75t_R FILLER_50_127 ();
 DECAPx4_ASAP7_75t_R FILLER_50_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_153 ();
 DECAPx1_ASAP7_75t_R FILLER_50_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_180 ();
 DECAPx1_ASAP7_75t_R FILLER_50_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_188 ();
 DECAPx4_ASAP7_75t_R FILLER_50_197 ();
 FILLER_ASAP7_75t_R FILLER_50_207 ();
 DECAPx10_ASAP7_75t_R FILLER_50_229 ();
 DECAPx4_ASAP7_75t_R FILLER_50_251 ();
 DECAPx6_ASAP7_75t_R FILLER_50_264 ();
 FILLER_ASAP7_75t_R FILLER_50_278 ();
 DECAPx2_ASAP7_75t_R FILLER_51_2 ();
 FILLER_ASAP7_75t_R FILLER_51_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_10 ();
 DECAPx10_ASAP7_75t_R FILLER_51_21 ();
 DECAPx1_ASAP7_75t_R FILLER_51_43 ();
 DECAPx6_ASAP7_75t_R FILLER_51_57 ();
 DECAPx1_ASAP7_75t_R FILLER_51_71 ();
 DECAPx2_ASAP7_75t_R FILLER_51_81 ();
 FILLER_ASAP7_75t_R FILLER_51_87 ();
 DECAPx1_ASAP7_75t_R FILLER_51_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_185 ();
 FILLER_ASAP7_75t_R FILLER_51_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_222 ();
 FILLER_ASAP7_75t_R FILLER_51_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_236 ();
 DECAPx10_ASAP7_75t_R FILLER_51_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_279 ();
 DECAPx10_ASAP7_75t_R FILLER_52_2 ();
 DECAPx2_ASAP7_75t_R FILLER_52_24 ();
 DECAPx10_ASAP7_75t_R FILLER_52_50 ();
 FILLER_ASAP7_75t_R FILLER_52_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_127 ();
 DECAPx1_ASAP7_75t_R FILLER_52_163 ();
 DECAPx4_ASAP7_75t_R FILLER_52_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_204 ();
 DECAPx1_ASAP7_75t_R FILLER_52_220 ();
 DECAPx10_ASAP7_75t_R FILLER_52_236 ();
 DECAPx10_ASAP7_75t_R FILLER_52_258 ();
 DECAPx10_ASAP7_75t_R FILLER_53_2 ();
 DECAPx10_ASAP7_75t_R FILLER_53_24 ();
 DECAPx2_ASAP7_75t_R FILLER_53_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_52 ();
 FILLER_ASAP7_75t_R FILLER_53_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_77 ();
 FILLER_ASAP7_75t_R FILLER_53_84 ();
 DECAPx2_ASAP7_75t_R FILLER_53_119 ();
 DECAPx1_ASAP7_75t_R FILLER_53_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_179 ();
 DECAPx2_ASAP7_75t_R FILLER_53_188 ();
 FILLER_ASAP7_75t_R FILLER_53_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_196 ();
 FILLER_ASAP7_75t_R FILLER_53_203 ();
 FILLER_ASAP7_75t_R FILLER_53_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_227 ();
 DECAPx10_ASAP7_75t_R FILLER_53_231 ();
 DECAPx10_ASAP7_75t_R FILLER_53_253 ();
 DECAPx1_ASAP7_75t_R FILLER_53_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_279 ();
 DECAPx10_ASAP7_75t_R FILLER_54_2 ();
 DECAPx10_ASAP7_75t_R FILLER_54_24 ();
 DECAPx10_ASAP7_75t_R FILLER_54_46 ();
 DECAPx4_ASAP7_75t_R FILLER_54_68 ();
 FILLER_ASAP7_75t_R FILLER_54_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_156 ();
 FILLER_ASAP7_75t_R FILLER_54_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_199 ();
 DECAPx10_ASAP7_75t_R FILLER_54_241 ();
 DECAPx6_ASAP7_75t_R FILLER_54_263 ();
 FILLER_ASAP7_75t_R FILLER_54_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_279 ();
 DECAPx10_ASAP7_75t_R FILLER_55_2 ();
 DECAPx10_ASAP7_75t_R FILLER_55_24 ();
 DECAPx10_ASAP7_75t_R FILLER_55_46 ();
 DECAPx6_ASAP7_75t_R FILLER_55_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_82 ();
 DECAPx1_ASAP7_75t_R FILLER_55_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_243 ();
 DECAPx10_ASAP7_75t_R FILLER_55_250 ();
 DECAPx2_ASAP7_75t_R FILLER_55_272 ();
 FILLER_ASAP7_75t_R FILLER_55_278 ();
endmodule
