module pi_switch (ce,
    clk,
    done,
    rst,
    l_i,
    l_o,
    r_i,
    r_o,
    u0_i,
    u0_o,
    u1_i,
    u1_o);
 input ce;
 input clk;
 output done;
 input rst;
 input [36:0] l_i;
 output [36:0] l_o;
 input [36:0] r_i;
 output [36:0] r_o;
 input [36:0] u0_i;
 output [36:0] u0_o;
 input [36:0] u1_i;
 output [36:0] u1_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire clknet_0_clk;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 BUFx6f_ASAP7_75t_R _0580_ (.A(r_i[36]),
    .Y(_0358_));
 BUFx6f_ASAP7_75t_R _0581_ (.A(u1_i[36]),
    .Y(_0359_));
 BUFx12f_ASAP7_75t_R _0582_ (.A(u0_i[36]),
    .Y(_0360_));
 BUFx6f_ASAP7_75t_R _0583_ (.A(_0360_),
    .Y(_0361_));
 BUFx6f_ASAP7_75t_R _0584_ (.A(_0361_),
    .Y(_0362_));
 OR4x1_ASAP7_75t_R _0585_ (.A(_0358_),
    .B(net29),
    .C(_0359_),
    .D(_0362_),
    .Y(_0363_));
 INVx1_ASAP7_75t_R _0586_ (.A(_0363_),
    .Y(_0000_));
 INVx1_ASAP7_75t_R _0587_ (.A(_0001_),
    .Y(net286));
 INVx1_ASAP7_75t_R _0588_ (.A(_0002_),
    .Y(net285));
 INVx1_ASAP7_75t_R _0589_ (.A(_0003_),
    .Y(net284));
 INVx1_ASAP7_75t_R _0590_ (.A(_0004_),
    .Y(net283));
 INVx1_ASAP7_75t_R _0591_ (.A(_0005_),
    .Y(net282));
 INVx1_ASAP7_75t_R _0592_ (.A(_0006_),
    .Y(net281));
 INVx1_ASAP7_75t_R _0593_ (.A(_0007_),
    .Y(net280));
 INVx1_ASAP7_75t_R _0594_ (.A(_0008_),
    .Y(net279));
 INVx1_ASAP7_75t_R _0595_ (.A(_0009_),
    .Y(net278));
 INVx1_ASAP7_75t_R _0596_ (.A(_0010_),
    .Y(net277));
 INVx1_ASAP7_75t_R _0597_ (.A(_0011_),
    .Y(net276));
 INVx1_ASAP7_75t_R _0598_ (.A(_0012_),
    .Y(net275));
 INVx1_ASAP7_75t_R _0599_ (.A(_0013_),
    .Y(net274));
 INVx1_ASAP7_75t_R _0600_ (.A(_0014_),
    .Y(net273));
 INVx1_ASAP7_75t_R _0601_ (.A(_0015_),
    .Y(net272));
 INVx1_ASAP7_75t_R _0602_ (.A(_0016_),
    .Y(net271));
 INVx1_ASAP7_75t_R _0603_ (.A(_0017_),
    .Y(net270));
 INVx1_ASAP7_75t_R _0604_ (.A(_0018_),
    .Y(net269));
 INVx1_ASAP7_75t_R _0605_ (.A(_0019_),
    .Y(net268));
 INVx1_ASAP7_75t_R _0606_ (.A(_0020_),
    .Y(net267));
 INVx1_ASAP7_75t_R _0607_ (.A(_0021_),
    .Y(net266));
 INVx1_ASAP7_75t_R _0608_ (.A(_0022_),
    .Y(net265));
 INVx1_ASAP7_75t_R _0609_ (.A(_0023_),
    .Y(net264));
 INVx1_ASAP7_75t_R _0610_ (.A(_0024_),
    .Y(net263));
 INVx1_ASAP7_75t_R _0611_ (.A(_0025_),
    .Y(net262));
 INVx1_ASAP7_75t_R _0612_ (.A(_0026_),
    .Y(net261));
 INVx1_ASAP7_75t_R _0613_ (.A(_0027_),
    .Y(net260));
 INVx1_ASAP7_75t_R _0614_ (.A(_0028_),
    .Y(net259));
 INVx1_ASAP7_75t_R _0615_ (.A(_0029_),
    .Y(net258));
 INVx1_ASAP7_75t_R _0616_ (.A(_0030_),
    .Y(net257));
 INVx1_ASAP7_75t_R _0617_ (.A(_0031_),
    .Y(net256));
 INVx1_ASAP7_75t_R _0618_ (.A(_0032_),
    .Y(net255));
 INVx1_ASAP7_75t_R _0619_ (.A(_0033_),
    .Y(net254));
 INVx1_ASAP7_75t_R _0620_ (.A(_0034_),
    .Y(net253));
 INVx1_ASAP7_75t_R _0621_ (.A(_0035_),
    .Y(net252));
 INVx1_ASAP7_75t_R _0622_ (.A(_0036_),
    .Y(net251));
 INVx1_ASAP7_75t_R _0623_ (.A(_0037_),
    .Y(net250));
 INVx1_ASAP7_75t_R _0624_ (.A(_0038_),
    .Y(net249));
 INVx1_ASAP7_75t_R _0625_ (.A(_0039_),
    .Y(net248));
 INVx1_ASAP7_75t_R _0626_ (.A(_0040_),
    .Y(net247));
 INVx1_ASAP7_75t_R _0627_ (.A(_0041_),
    .Y(net246));
 INVx1_ASAP7_75t_R _0628_ (.A(_0042_),
    .Y(net245));
 INVx1_ASAP7_75t_R _0629_ (.A(_0043_),
    .Y(net244));
 INVx1_ASAP7_75t_R _0630_ (.A(_0044_),
    .Y(net243));
 INVx1_ASAP7_75t_R _0631_ (.A(_0045_),
    .Y(net242));
 INVx1_ASAP7_75t_R _0632_ (.A(_0046_),
    .Y(net241));
 INVx1_ASAP7_75t_R _0633_ (.A(_0047_),
    .Y(net240));
 INVx1_ASAP7_75t_R _0634_ (.A(_0048_),
    .Y(net239));
 INVx1_ASAP7_75t_R _0635_ (.A(_0049_),
    .Y(net238));
 INVx1_ASAP7_75t_R _0636_ (.A(_0050_),
    .Y(net237));
 INVx1_ASAP7_75t_R _0637_ (.A(_0051_),
    .Y(net236));
 INVx1_ASAP7_75t_R _0638_ (.A(_0052_),
    .Y(net235));
 INVx1_ASAP7_75t_R _0639_ (.A(_0053_),
    .Y(net234));
 INVx1_ASAP7_75t_R _0640_ (.A(_0054_),
    .Y(net233));
 INVx1_ASAP7_75t_R _0641_ (.A(_0055_),
    .Y(net232));
 INVx1_ASAP7_75t_R _0642_ (.A(_0056_),
    .Y(net231));
 INVx1_ASAP7_75t_R _0643_ (.A(_0057_),
    .Y(net230));
 INVx1_ASAP7_75t_R _0644_ (.A(_0058_),
    .Y(net229));
 INVx1_ASAP7_75t_R _0645_ (.A(_0059_),
    .Y(net228));
 INVx1_ASAP7_75t_R _0646_ (.A(_0060_),
    .Y(net227));
 INVx1_ASAP7_75t_R _0647_ (.A(_0061_),
    .Y(net226));
 INVx1_ASAP7_75t_R _0648_ (.A(_0062_),
    .Y(net225));
 INVx1_ASAP7_75t_R _0649_ (.A(_0063_),
    .Y(net224));
 INVx1_ASAP7_75t_R _0650_ (.A(_0064_),
    .Y(net223));
 INVx1_ASAP7_75t_R _0651_ (.A(_0065_),
    .Y(net222));
 INVx1_ASAP7_75t_R _0652_ (.A(_0066_),
    .Y(net221));
 INVx1_ASAP7_75t_R _0653_ (.A(_0067_),
    .Y(net220));
 INVx1_ASAP7_75t_R _0654_ (.A(_0068_),
    .Y(net219));
 INVx1_ASAP7_75t_R _0655_ (.A(_0069_),
    .Y(net218));
 INVx1_ASAP7_75t_R _0656_ (.A(_0070_),
    .Y(net217));
 INVx1_ASAP7_75t_R _0657_ (.A(_0071_),
    .Y(net216));
 INVx1_ASAP7_75t_R _0658_ (.A(_0072_),
    .Y(net215));
 INVx1_ASAP7_75t_R _0659_ (.A(_0073_),
    .Y(net214));
 INVx1_ASAP7_75t_R _0660_ (.A(_0074_),
    .Y(net213));
 INVx1_ASAP7_75t_R _0661_ (.A(_0075_),
    .Y(net212));
 INVx1_ASAP7_75t_R _0662_ (.A(_0076_),
    .Y(net211));
 INVx1_ASAP7_75t_R _0663_ (.A(_0077_),
    .Y(net210));
 INVx1_ASAP7_75t_R _0664_ (.A(_0078_),
    .Y(net209));
 INVx1_ASAP7_75t_R _0665_ (.A(_0079_),
    .Y(net208));
 INVx1_ASAP7_75t_R _0666_ (.A(_0080_),
    .Y(net207));
 INVx1_ASAP7_75t_R _0667_ (.A(_0081_),
    .Y(net206));
 INVx1_ASAP7_75t_R _0668_ (.A(_0082_),
    .Y(net205));
 INVx1_ASAP7_75t_R _0669_ (.A(_0083_),
    .Y(net204));
 INVx1_ASAP7_75t_R _0670_ (.A(_0084_),
    .Y(net203));
 INVx1_ASAP7_75t_R _0671_ (.A(_0085_),
    .Y(net202));
 INVx1_ASAP7_75t_R _0672_ (.A(_0086_),
    .Y(net201));
 INVx1_ASAP7_75t_R _0673_ (.A(_0087_),
    .Y(net200));
 INVx1_ASAP7_75t_R _0674_ (.A(_0088_),
    .Y(net199));
 INVx1_ASAP7_75t_R _0675_ (.A(_0089_),
    .Y(net198));
 INVx1_ASAP7_75t_R _0676_ (.A(_0090_),
    .Y(net197));
 INVx1_ASAP7_75t_R _0677_ (.A(_0091_),
    .Y(net196));
 INVx1_ASAP7_75t_R _0678_ (.A(_0092_),
    .Y(net195));
 INVx1_ASAP7_75t_R _0679_ (.A(_0093_),
    .Y(net194));
 INVx1_ASAP7_75t_R _0680_ (.A(_0094_),
    .Y(net193));
 INVx1_ASAP7_75t_R _0681_ (.A(_0095_),
    .Y(net192));
 INVx1_ASAP7_75t_R _0682_ (.A(_0096_),
    .Y(net191));
 INVx1_ASAP7_75t_R _0683_ (.A(_0097_),
    .Y(net190));
 INVx1_ASAP7_75t_R _0684_ (.A(_0098_),
    .Y(net189));
 INVx1_ASAP7_75t_R _0685_ (.A(_0099_),
    .Y(net188));
 INVx1_ASAP7_75t_R _0686_ (.A(_0100_),
    .Y(net187));
 INVx1_ASAP7_75t_R _0687_ (.A(_0101_),
    .Y(net186));
 INVx1_ASAP7_75t_R _0688_ (.A(_0102_),
    .Y(net185));
 INVx1_ASAP7_75t_R _0689_ (.A(_0103_),
    .Y(net184));
 INVx1_ASAP7_75t_R _0690_ (.A(_0104_),
    .Y(net183));
 INVx1_ASAP7_75t_R _0691_ (.A(_0105_),
    .Y(net182));
 INVx1_ASAP7_75t_R _0692_ (.A(_0106_),
    .Y(net181));
 INVx1_ASAP7_75t_R _0693_ (.A(_0107_),
    .Y(net180));
 INVx1_ASAP7_75t_R _0694_ (.A(_0108_),
    .Y(net179));
 INVx1_ASAP7_75t_R _0695_ (.A(_0109_),
    .Y(net178));
 INVx1_ASAP7_75t_R _0696_ (.A(_0110_),
    .Y(net177));
 INVx1_ASAP7_75t_R _0697_ (.A(_0111_),
    .Y(net176));
 INVx1_ASAP7_75t_R _0698_ (.A(_0112_),
    .Y(net175));
 INVx1_ASAP7_75t_R _0699_ (.A(_0113_),
    .Y(net174));
 INVx1_ASAP7_75t_R _0700_ (.A(_0114_),
    .Y(net173));
 INVx1_ASAP7_75t_R _0701_ (.A(_0115_),
    .Y(net172));
 INVx1_ASAP7_75t_R _0702_ (.A(_0116_),
    .Y(net171));
 INVx1_ASAP7_75t_R _0703_ (.A(_0117_),
    .Y(net170));
 INVx1_ASAP7_75t_R _0704_ (.A(_0118_),
    .Y(net169));
 INVx1_ASAP7_75t_R _0705_ (.A(_0119_),
    .Y(net168));
 INVx1_ASAP7_75t_R _0706_ (.A(_0120_),
    .Y(net167));
 INVx1_ASAP7_75t_R _0707_ (.A(_0121_),
    .Y(net166));
 INVx1_ASAP7_75t_R _0708_ (.A(_0122_),
    .Y(net165));
 INVx1_ASAP7_75t_R _0709_ (.A(_0123_),
    .Y(net164));
 INVx1_ASAP7_75t_R _0710_ (.A(_0124_),
    .Y(net163));
 INVx1_ASAP7_75t_R _0711_ (.A(_0125_),
    .Y(net162));
 INVx1_ASAP7_75t_R _0712_ (.A(_0126_),
    .Y(net161));
 INVx1_ASAP7_75t_R _0713_ (.A(_0127_),
    .Y(net160));
 INVx1_ASAP7_75t_R _0714_ (.A(_0128_),
    .Y(net159));
 INVx1_ASAP7_75t_R _0715_ (.A(_0129_),
    .Y(net158));
 INVx1_ASAP7_75t_R _0716_ (.A(_0130_),
    .Y(net157));
 INVx1_ASAP7_75t_R _0717_ (.A(_0131_),
    .Y(net156));
 INVx1_ASAP7_75t_R _0718_ (.A(_0132_),
    .Y(net155));
 INVx1_ASAP7_75t_R _0719_ (.A(_0133_),
    .Y(net154));
 INVx1_ASAP7_75t_R _0720_ (.A(_0134_),
    .Y(net153));
 INVx1_ASAP7_75t_R _0721_ (.A(_0135_),
    .Y(net152));
 INVx1_ASAP7_75t_R _0722_ (.A(_0136_),
    .Y(net151));
 INVx1_ASAP7_75t_R _0723_ (.A(_0137_),
    .Y(net150));
 INVx1_ASAP7_75t_R _0724_ (.A(_0138_),
    .Y(net149));
 INVx1_ASAP7_75t_R _0725_ (.A(_0139_),
    .Y(net148));
 INVx1_ASAP7_75t_R _0726_ (.A(_0140_),
    .Y(net147));
 INVx1_ASAP7_75t_R _0727_ (.A(_0141_),
    .Y(net146));
 INVx1_ASAP7_75t_R _0728_ (.A(_0142_),
    .Y(net145));
 INVx1_ASAP7_75t_R _0729_ (.A(_0143_),
    .Y(net144));
 INVx1_ASAP7_75t_R _0730_ (.A(_0144_),
    .Y(net143));
 INVx1_ASAP7_75t_R _0731_ (.A(_0145_),
    .Y(net142));
 AND2x4_ASAP7_75t_R _0732_ (.A(_0359_),
    .B(_0360_),
    .Y(_0364_));
 BUFx3_ASAP7_75t_R _0733_ (.A(u1_i[32]),
    .Y(_0365_));
 INVx1_ASAP7_75t_R _0734_ (.A(_0365_),
    .Y(_0366_));
 NOR3x1_ASAP7_75t_R _0735_ (.A(net64),
    .B(net63),
    .C(net62),
    .Y(_0367_));
 AO21x1_ASAP7_75t_R _0736_ (.A1(_0358_),
    .A2(_0367_),
    .B(net98),
    .Y(_0368_));
 OR2x6_ASAP7_75t_R _0737_ (.A(net28),
    .B(net27),
    .Y(_0369_));
 NAND2x1_ASAP7_75t_R _0738_ (.A(net29),
    .B(net26),
    .Y(_0370_));
 OA21x2_ASAP7_75t_R _0739_ (.A1(_0369_),
    .A2(_0370_),
    .B(net98),
    .Y(_0371_));
 AO21x1_ASAP7_75t_R _0740_ (.A1(_0366_),
    .A2(_0368_),
    .B(_0371_),
    .Y(_0372_));
 NOR2x2_ASAP7_75t_R _0741_ (.A(net28),
    .B(net27),
    .Y(_0373_));
 AND2x4_ASAP7_75t_R _0742_ (.A(net29),
    .B(net26),
    .Y(_0374_));
 AND2x4_ASAP7_75t_R _0743_ (.A(_0373_),
    .B(_0374_),
    .Y(_0375_));
 AND2x2_ASAP7_75t_R _0744_ (.A(_0359_),
    .B(_0366_),
    .Y(_0376_));
 NAND2x1_ASAP7_75t_R _0745_ (.A(_0358_),
    .B(_0367_),
    .Y(_0377_));
 AO21x1_ASAP7_75t_R _0746_ (.A1(_0375_),
    .A2(_0376_),
    .B(_0377_),
    .Y(_0378_));
 INVx2_ASAP7_75t_R _0747_ (.A(_0360_),
    .Y(_0379_));
 AND2x2_ASAP7_75t_R _0748_ (.A(_0371_),
    .B(_0377_),
    .Y(_0380_));
 AO221x1_ASAP7_75t_R _0749_ (.A1(_0364_),
    .A2(_0372_),
    .B1(_0378_),
    .B2(_0379_),
    .C(_0380_),
    .Y(_0381_));
 BUFx6f_ASAP7_75t_R _0750_ (.A(_0381_),
    .Y(_0382_));
 BUFx6f_ASAP7_75t_R _0751_ (.A(_0382_),
    .Y(_0383_));
 INVx2_ASAP7_75t_R _0752_ (.A(_0359_),
    .Y(_0384_));
 AND3x1_ASAP7_75t_R _0753_ (.A(_0384_),
    .B(_0373_),
    .C(_0374_),
    .Y(_0385_));
 INVx1_ASAP7_75t_R _0754_ (.A(_0358_),
    .Y(_0386_));
 OR3x1_ASAP7_75t_R _0755_ (.A(net64),
    .B(net63),
    .C(net62),
    .Y(_0387_));
 AND2x2_ASAP7_75t_R _0756_ (.A(_0359_),
    .B(_0365_),
    .Y(_0388_));
 OR3x1_ASAP7_75t_R _0757_ (.A(_0386_),
    .B(_0387_),
    .C(_0388_),
    .Y(_0389_));
 INVx2_ASAP7_75t_R _0758_ (.A(net98),
    .Y(_0390_));
 OA21x2_ASAP7_75t_R _0759_ (.A1(_0390_),
    .A2(_0388_),
    .B(_0360_),
    .Y(_0391_));
 AO21x1_ASAP7_75t_R _0760_ (.A1(_0373_),
    .A2(_0374_),
    .B(_0390_),
    .Y(_0392_));
 OA211x2_ASAP7_75t_R _0761_ (.A1(_0385_),
    .A2(_0389_),
    .B(_0391_),
    .C(_0392_),
    .Y(_0393_));
 OA211x2_ASAP7_75t_R _0762_ (.A1(_0369_),
    .A2(_0370_),
    .B(_0365_),
    .C(_0379_),
    .Y(_0394_));
 OA21x2_ASAP7_75t_R _0763_ (.A1(_0384_),
    .A2(_0394_),
    .B(_0377_),
    .Y(_0395_));
 NOR2x2_ASAP7_75t_R _0764_ (.A(_0393_),
    .B(_0395_),
    .Y(_0396_));
 AND2x2_ASAP7_75t_R _0765_ (.A(net37),
    .B(_0396_),
    .Y(_0397_));
 OR2x2_ASAP7_75t_R _0766_ (.A(_0393_),
    .B(_0395_),
    .Y(_0398_));
 BUFx6f_ASAP7_75t_R _0767_ (.A(_0398_),
    .Y(_0399_));
 AND2x2_ASAP7_75t_R _0768_ (.A(net73),
    .B(_0399_),
    .Y(_0400_));
 AOI221x1_ASAP7_75t_R _0769_ (.A1(_0364_),
    .A2(_0372_),
    .B1(_0378_),
    .B2(_0379_),
    .C(_0380_),
    .Y(_0401_));
 INVx5_ASAP7_75t_R _0770_ (.A(net72),
    .Y(_0402_));
 BUFx12f_ASAP7_75t_R _0771_ (.A(_0402_),
    .Y(_0403_));
 OA21x2_ASAP7_75t_R _0772_ (.A1(net108),
    .A2(_0401_),
    .B(_0403_),
    .Y(_0404_));
 OA31x2_ASAP7_75t_R _0773_ (.A1(_0383_),
    .A2(_0397_),
    .A3(_0400_),
    .B1(_0404_),
    .Y(_0146_));
 BUFx6f_ASAP7_75t_R _0774_ (.A(_0399_),
    .Y(_0405_));
 AND2x2_ASAP7_75t_R _0775_ (.A(net74),
    .B(_0405_),
    .Y(_0406_));
 BUFx6f_ASAP7_75t_R _0776_ (.A(_0396_),
    .Y(_0407_));
 AO21x1_ASAP7_75t_R _0777_ (.A1(net38),
    .A2(_0407_),
    .B(_0383_),
    .Y(_0408_));
 BUFx6f_ASAP7_75t_R _0778_ (.A(_0401_),
    .Y(_0409_));
 BUFx6f_ASAP7_75t_R _0779_ (.A(_0402_),
    .Y(_0410_));
 OA21x2_ASAP7_75t_R _0780_ (.A1(net109),
    .A2(_0409_),
    .B(_0410_),
    .Y(_0411_));
 OA21x2_ASAP7_75t_R _0781_ (.A1(_0406_),
    .A2(_0408_),
    .B(_0411_),
    .Y(_0147_));
 AND2x2_ASAP7_75t_R _0782_ (.A(net75),
    .B(_0405_),
    .Y(_0412_));
 AO21x1_ASAP7_75t_R _0783_ (.A1(net39),
    .A2(_0407_),
    .B(_0383_),
    .Y(_0413_));
 OA21x2_ASAP7_75t_R _0784_ (.A1(net110),
    .A2(_0409_),
    .B(_0410_),
    .Y(_0414_));
 OA21x2_ASAP7_75t_R _0785_ (.A1(_0412_),
    .A2(_0413_),
    .B(_0414_),
    .Y(_0148_));
 AND2x2_ASAP7_75t_R _0786_ (.A(net76),
    .B(_0405_),
    .Y(_0415_));
 AO21x1_ASAP7_75t_R _0787_ (.A1(net40),
    .A2(_0407_),
    .B(_0383_),
    .Y(_0416_));
 OA21x2_ASAP7_75t_R _0788_ (.A1(net111),
    .A2(_0409_),
    .B(_0410_),
    .Y(_0417_));
 OA21x2_ASAP7_75t_R _0789_ (.A1(_0415_),
    .A2(_0416_),
    .B(_0417_),
    .Y(_0149_));
 AND2x2_ASAP7_75t_R _0790_ (.A(net77),
    .B(_0405_),
    .Y(_0418_));
 AO21x1_ASAP7_75t_R _0791_ (.A1(net41),
    .A2(_0407_),
    .B(_0383_),
    .Y(_0419_));
 OA21x2_ASAP7_75t_R _0792_ (.A1(net112),
    .A2(_0409_),
    .B(_0410_),
    .Y(_0420_));
 OA21x2_ASAP7_75t_R _0793_ (.A1(_0418_),
    .A2(_0419_),
    .B(_0420_),
    .Y(_0150_));
 AND2x2_ASAP7_75t_R _0794_ (.A(net78),
    .B(_0405_),
    .Y(_0421_));
 AO21x1_ASAP7_75t_R _0795_ (.A1(net42),
    .A2(_0407_),
    .B(_0383_),
    .Y(_0422_));
 OA21x2_ASAP7_75t_R _0796_ (.A1(net113),
    .A2(_0409_),
    .B(_0410_),
    .Y(_0423_));
 OA21x2_ASAP7_75t_R _0797_ (.A1(_0421_),
    .A2(_0422_),
    .B(_0423_),
    .Y(_0151_));
 AND2x2_ASAP7_75t_R _0798_ (.A(net79),
    .B(_0405_),
    .Y(_0424_));
 AO21x1_ASAP7_75t_R _0799_ (.A1(net43),
    .A2(_0407_),
    .B(_0383_),
    .Y(_0425_));
 OA21x2_ASAP7_75t_R _0800_ (.A1(net114),
    .A2(_0409_),
    .B(_0410_),
    .Y(_0426_));
 OA21x2_ASAP7_75t_R _0801_ (.A1(_0424_),
    .A2(_0425_),
    .B(_0426_),
    .Y(_0152_));
 AND2x2_ASAP7_75t_R _0802_ (.A(net80),
    .B(_0405_),
    .Y(_0427_));
 AO21x1_ASAP7_75t_R _0803_ (.A1(net44),
    .A2(_0407_),
    .B(_0383_),
    .Y(_0428_));
 OA21x2_ASAP7_75t_R _0804_ (.A1(net115),
    .A2(_0409_),
    .B(_0410_),
    .Y(_0429_));
 OA21x2_ASAP7_75t_R _0805_ (.A1(_0427_),
    .A2(_0428_),
    .B(_0429_),
    .Y(_0153_));
 AND2x2_ASAP7_75t_R _0806_ (.A(net81),
    .B(_0405_),
    .Y(_0430_));
 AO21x1_ASAP7_75t_R _0807_ (.A1(net45),
    .A2(_0407_),
    .B(_0383_),
    .Y(_0431_));
 OA21x2_ASAP7_75t_R _0808_ (.A1(net116),
    .A2(_0409_),
    .B(_0410_),
    .Y(_0432_));
 OA21x2_ASAP7_75t_R _0809_ (.A1(_0430_),
    .A2(_0431_),
    .B(_0432_),
    .Y(_0154_));
 AND2x2_ASAP7_75t_R _0810_ (.A(net82),
    .B(_0405_),
    .Y(_0433_));
 AO21x1_ASAP7_75t_R _0811_ (.A1(net46),
    .A2(_0407_),
    .B(_0383_),
    .Y(_0434_));
 OA21x2_ASAP7_75t_R _0812_ (.A1(net117),
    .A2(_0409_),
    .B(_0410_),
    .Y(_0435_));
 OA21x2_ASAP7_75t_R _0813_ (.A1(_0433_),
    .A2(_0434_),
    .B(_0435_),
    .Y(_0155_));
 AND2x2_ASAP7_75t_R _0814_ (.A(net83),
    .B(_0405_),
    .Y(_0436_));
 BUFx6f_ASAP7_75t_R _0815_ (.A(_0382_),
    .Y(_0437_));
 AO21x1_ASAP7_75t_R _0816_ (.A1(net47),
    .A2(_0407_),
    .B(_0437_),
    .Y(_0438_));
 BUFx6f_ASAP7_75t_R _0817_ (.A(_0402_),
    .Y(_0439_));
 OA21x2_ASAP7_75t_R _0818_ (.A1(net118),
    .A2(_0409_),
    .B(_0439_),
    .Y(_0440_));
 OA21x2_ASAP7_75t_R _0819_ (.A1(_0436_),
    .A2(_0438_),
    .B(_0440_),
    .Y(_0156_));
 BUFx6f_ASAP7_75t_R _0820_ (.A(_0399_),
    .Y(_0441_));
 AND2x2_ASAP7_75t_R _0821_ (.A(net84),
    .B(_0441_),
    .Y(_0442_));
 BUFx6f_ASAP7_75t_R _0822_ (.A(_0396_),
    .Y(_0443_));
 AO21x1_ASAP7_75t_R _0823_ (.A1(net48),
    .A2(_0443_),
    .B(_0437_),
    .Y(_0444_));
 BUFx6f_ASAP7_75t_R _0824_ (.A(_0401_),
    .Y(_0445_));
 OA21x2_ASAP7_75t_R _0825_ (.A1(net119),
    .A2(_0445_),
    .B(_0439_),
    .Y(_0446_));
 OA21x2_ASAP7_75t_R _0826_ (.A1(_0442_),
    .A2(_0444_),
    .B(_0446_),
    .Y(_0157_));
 AND2x2_ASAP7_75t_R _0827_ (.A(net85),
    .B(_0441_),
    .Y(_0447_));
 AO21x1_ASAP7_75t_R _0828_ (.A1(net49),
    .A2(_0443_),
    .B(_0437_),
    .Y(_0448_));
 OA21x2_ASAP7_75t_R _0829_ (.A1(net120),
    .A2(_0445_),
    .B(_0439_),
    .Y(_0449_));
 OA21x2_ASAP7_75t_R _0830_ (.A1(_0447_),
    .A2(_0448_),
    .B(_0449_),
    .Y(_0158_));
 AND2x2_ASAP7_75t_R _0831_ (.A(net86),
    .B(_0441_),
    .Y(_0450_));
 AO21x1_ASAP7_75t_R _0832_ (.A1(net50),
    .A2(_0443_),
    .B(_0437_),
    .Y(_0451_));
 OA21x2_ASAP7_75t_R _0833_ (.A1(net121),
    .A2(_0445_),
    .B(_0439_),
    .Y(_0452_));
 OA21x2_ASAP7_75t_R _0834_ (.A1(_0450_),
    .A2(_0451_),
    .B(_0452_),
    .Y(_0159_));
 AND2x2_ASAP7_75t_R _0835_ (.A(net87),
    .B(_0441_),
    .Y(_0453_));
 AO21x1_ASAP7_75t_R _0836_ (.A1(net51),
    .A2(_0443_),
    .B(_0437_),
    .Y(_0454_));
 OA21x2_ASAP7_75t_R _0837_ (.A1(net122),
    .A2(_0445_),
    .B(_0439_),
    .Y(_0455_));
 OA21x2_ASAP7_75t_R _0838_ (.A1(_0453_),
    .A2(_0454_),
    .B(_0455_),
    .Y(_0160_));
 AND2x2_ASAP7_75t_R _0839_ (.A(net88),
    .B(_0441_),
    .Y(_0456_));
 AO21x1_ASAP7_75t_R _0840_ (.A1(net52),
    .A2(_0443_),
    .B(_0437_),
    .Y(_0457_));
 OA21x2_ASAP7_75t_R _0841_ (.A1(net123),
    .A2(_0445_),
    .B(_0439_),
    .Y(_0458_));
 OA21x2_ASAP7_75t_R _0842_ (.A1(_0456_),
    .A2(_0457_),
    .B(_0458_),
    .Y(_0161_));
 AND2x2_ASAP7_75t_R _0843_ (.A(net89),
    .B(_0441_),
    .Y(_0459_));
 AO21x1_ASAP7_75t_R _0844_ (.A1(net53),
    .A2(_0443_),
    .B(_0437_),
    .Y(_0460_));
 OA21x2_ASAP7_75t_R _0845_ (.A1(net124),
    .A2(_0445_),
    .B(_0439_),
    .Y(_0461_));
 OA21x2_ASAP7_75t_R _0846_ (.A1(_0459_),
    .A2(_0460_),
    .B(_0461_),
    .Y(_0162_));
 AND2x2_ASAP7_75t_R _0847_ (.A(net90),
    .B(_0441_),
    .Y(_0462_));
 AO21x1_ASAP7_75t_R _0848_ (.A1(net54),
    .A2(_0443_),
    .B(_0437_),
    .Y(_0463_));
 OA21x2_ASAP7_75t_R _0849_ (.A1(net125),
    .A2(_0445_),
    .B(_0439_),
    .Y(_0464_));
 OA21x2_ASAP7_75t_R _0850_ (.A1(_0462_),
    .A2(_0463_),
    .B(_0464_),
    .Y(_0163_));
 AND2x2_ASAP7_75t_R _0851_ (.A(net91),
    .B(_0441_),
    .Y(_0465_));
 AO21x1_ASAP7_75t_R _0852_ (.A1(net55),
    .A2(_0443_),
    .B(_0437_),
    .Y(_0466_));
 OA21x2_ASAP7_75t_R _0853_ (.A1(net126),
    .A2(_0445_),
    .B(_0439_),
    .Y(_0467_));
 OA21x2_ASAP7_75t_R _0854_ (.A1(_0465_),
    .A2(_0466_),
    .B(_0467_),
    .Y(_0164_));
 AND2x2_ASAP7_75t_R _0855_ (.A(net92),
    .B(_0441_),
    .Y(_0468_));
 AO21x1_ASAP7_75t_R _0856_ (.A1(net56),
    .A2(_0443_),
    .B(_0437_),
    .Y(_0469_));
 OA21x2_ASAP7_75t_R _0857_ (.A1(net127),
    .A2(_0445_),
    .B(_0439_),
    .Y(_0470_));
 OA21x2_ASAP7_75t_R _0858_ (.A1(_0468_),
    .A2(_0469_),
    .B(_0470_),
    .Y(_0165_));
 AND2x2_ASAP7_75t_R _0859_ (.A(net93),
    .B(_0441_),
    .Y(_0471_));
 BUFx6f_ASAP7_75t_R _0860_ (.A(_0382_),
    .Y(_0472_));
 AO21x1_ASAP7_75t_R _0861_ (.A1(net57),
    .A2(_0443_),
    .B(_0472_),
    .Y(_0473_));
 BUFx6f_ASAP7_75t_R _0862_ (.A(_0402_),
    .Y(_0474_));
 OA21x2_ASAP7_75t_R _0863_ (.A1(net128),
    .A2(_0445_),
    .B(_0474_),
    .Y(_0475_));
 OA21x2_ASAP7_75t_R _0864_ (.A1(_0471_),
    .A2(_0473_),
    .B(_0475_),
    .Y(_0166_));
 BUFx6f_ASAP7_75t_R _0865_ (.A(_0399_),
    .Y(_0476_));
 AND2x2_ASAP7_75t_R _0866_ (.A(net94),
    .B(_0476_),
    .Y(_0477_));
 BUFx6f_ASAP7_75t_R _0867_ (.A(_0396_),
    .Y(_0478_));
 AO21x1_ASAP7_75t_R _0868_ (.A1(net58),
    .A2(_0478_),
    .B(_0472_),
    .Y(_0479_));
 BUFx6f_ASAP7_75t_R _0869_ (.A(_0401_),
    .Y(_0480_));
 OA21x2_ASAP7_75t_R _0870_ (.A1(net129),
    .A2(_0480_),
    .B(_0474_),
    .Y(_0481_));
 OA21x2_ASAP7_75t_R _0871_ (.A1(_0477_),
    .A2(_0479_),
    .B(_0481_),
    .Y(_0167_));
 AND2x2_ASAP7_75t_R _0872_ (.A(net95),
    .B(_0476_),
    .Y(_0482_));
 AO21x1_ASAP7_75t_R _0873_ (.A1(net59),
    .A2(_0478_),
    .B(_0472_),
    .Y(_0483_));
 OA21x2_ASAP7_75t_R _0874_ (.A1(net130),
    .A2(_0480_),
    .B(_0474_),
    .Y(_0484_));
 OA21x2_ASAP7_75t_R _0875_ (.A1(_0482_),
    .A2(_0483_),
    .B(_0484_),
    .Y(_0168_));
 AND2x2_ASAP7_75t_R _0876_ (.A(net96),
    .B(_0476_),
    .Y(_0485_));
 AO21x1_ASAP7_75t_R _0877_ (.A1(net60),
    .A2(_0478_),
    .B(_0472_),
    .Y(_0486_));
 OA21x2_ASAP7_75t_R _0878_ (.A1(net131),
    .A2(_0480_),
    .B(_0474_),
    .Y(_0487_));
 OA21x2_ASAP7_75t_R _0879_ (.A1(_0485_),
    .A2(_0486_),
    .B(_0487_),
    .Y(_0169_));
 AND2x2_ASAP7_75t_R _0880_ (.A(net97),
    .B(_0476_),
    .Y(_0488_));
 AO21x1_ASAP7_75t_R _0881_ (.A1(net61),
    .A2(_0478_),
    .B(_0472_),
    .Y(_0489_));
 OA21x2_ASAP7_75t_R _0882_ (.A1(net132),
    .A2(_0480_),
    .B(_0474_),
    .Y(_0490_));
 OA21x2_ASAP7_75t_R _0883_ (.A1(_0488_),
    .A2(_0489_),
    .B(_0490_),
    .Y(_0170_));
 AND2x2_ASAP7_75t_R _0884_ (.A(_0365_),
    .B(_0382_),
    .Y(_0491_));
 AND3x1_ASAP7_75t_R _0885_ (.A(net98),
    .B(_0401_),
    .C(_0399_),
    .Y(_0492_));
 BUFx6f_ASAP7_75t_R _0886_ (.A(_0403_),
    .Y(_0493_));
 OA21x2_ASAP7_75t_R _0887_ (.A1(_0491_),
    .A2(_0492_),
    .B(_0493_),
    .Y(_0171_));
 AND2x2_ASAP7_75t_R _0888_ (.A(net133),
    .B(_0382_),
    .Y(_0494_));
 AND3x1_ASAP7_75t_R _0889_ (.A(net99),
    .B(_0401_),
    .C(_0399_),
    .Y(_0495_));
 OA21x2_ASAP7_75t_R _0890_ (.A1(_0494_),
    .A2(_0495_),
    .B(_0493_),
    .Y(_0172_));
 AND2x2_ASAP7_75t_R _0891_ (.A(net134),
    .B(_0382_),
    .Y(_0496_));
 AND3x1_ASAP7_75t_R _0892_ (.A(net100),
    .B(_0401_),
    .C(_0399_),
    .Y(_0497_));
 OA21x2_ASAP7_75t_R _0893_ (.A1(_0496_),
    .A2(_0497_),
    .B(_0493_),
    .Y(_0173_));
 OA21x2_ASAP7_75t_R _0894_ (.A1(_0379_),
    .A2(_0371_),
    .B(_0384_),
    .Y(_0498_));
 OA21x2_ASAP7_75t_R _0895_ (.A1(_0394_),
    .A2(_0498_),
    .B(_0377_),
    .Y(_0499_));
 NOR2x1_ASAP7_75t_R _0896_ (.A(net72),
    .B(_0499_),
    .Y(_0174_));
 AND2x2_ASAP7_75t_R _0897_ (.A(net101),
    .B(_0476_),
    .Y(_0500_));
 AO21x1_ASAP7_75t_R _0898_ (.A1(net65),
    .A2(_0478_),
    .B(_0472_),
    .Y(_0501_));
 OA21x2_ASAP7_75t_R _0899_ (.A1(net135),
    .A2(_0480_),
    .B(_0474_),
    .Y(_0502_));
 OA21x2_ASAP7_75t_R _0900_ (.A1(_0500_),
    .A2(_0501_),
    .B(_0502_),
    .Y(_0175_));
 AND2x2_ASAP7_75t_R _0901_ (.A(net102),
    .B(_0476_),
    .Y(_0503_));
 AO21x1_ASAP7_75t_R _0902_ (.A1(net66),
    .A2(_0478_),
    .B(_0472_),
    .Y(_0504_));
 OA21x2_ASAP7_75t_R _0903_ (.A1(net136),
    .A2(_0480_),
    .B(_0474_),
    .Y(_0505_));
 OA21x2_ASAP7_75t_R _0904_ (.A1(_0503_),
    .A2(_0504_),
    .B(_0505_),
    .Y(_0176_));
 AND2x2_ASAP7_75t_R _0905_ (.A(net103),
    .B(_0476_),
    .Y(_0506_));
 AO21x1_ASAP7_75t_R _0906_ (.A1(net67),
    .A2(_0478_),
    .B(_0472_),
    .Y(_0507_));
 OA21x2_ASAP7_75t_R _0907_ (.A1(net137),
    .A2(_0480_),
    .B(_0474_),
    .Y(_0508_));
 OA21x2_ASAP7_75t_R _0908_ (.A1(_0506_),
    .A2(_0507_),
    .B(_0508_),
    .Y(_0177_));
 AND2x2_ASAP7_75t_R _0909_ (.A(net104),
    .B(_0476_),
    .Y(_0509_));
 AO21x1_ASAP7_75t_R _0910_ (.A1(net68),
    .A2(_0478_),
    .B(_0472_),
    .Y(_0510_));
 OA21x2_ASAP7_75t_R _0911_ (.A1(net138),
    .A2(_0480_),
    .B(_0474_),
    .Y(_0511_));
 OA21x2_ASAP7_75t_R _0912_ (.A1(_0509_),
    .A2(_0510_),
    .B(_0511_),
    .Y(_0178_));
 AND2x2_ASAP7_75t_R _0913_ (.A(net105),
    .B(_0476_),
    .Y(_0512_));
 AO21x1_ASAP7_75t_R _0914_ (.A1(net69),
    .A2(_0478_),
    .B(_0472_),
    .Y(_0513_));
 OA21x2_ASAP7_75t_R _0915_ (.A1(net139),
    .A2(_0480_),
    .B(_0474_),
    .Y(_0514_));
 OA21x2_ASAP7_75t_R _0916_ (.A1(_0512_),
    .A2(_0513_),
    .B(_0514_),
    .Y(_0179_));
 AND2x2_ASAP7_75t_R _0917_ (.A(net106),
    .B(_0476_),
    .Y(_0515_));
 AO21x1_ASAP7_75t_R _0918_ (.A1(net70),
    .A2(_0478_),
    .B(_0382_),
    .Y(_0516_));
 OA21x2_ASAP7_75t_R _0919_ (.A1(net140),
    .A2(_0480_),
    .B(_0403_),
    .Y(_0517_));
 OA21x2_ASAP7_75t_R _0920_ (.A1(_0515_),
    .A2(_0516_),
    .B(_0517_),
    .Y(_0180_));
 AND2x2_ASAP7_75t_R _0921_ (.A(net107),
    .B(_0399_),
    .Y(_0518_));
 AO21x1_ASAP7_75t_R _0922_ (.A1(net71),
    .A2(_0396_),
    .B(_0382_),
    .Y(_0519_));
 OA21x2_ASAP7_75t_R _0923_ (.A1(net141),
    .A2(_0401_),
    .B(_0403_),
    .Y(_0520_));
 OA21x2_ASAP7_75t_R _0924_ (.A1(_0518_),
    .A2(_0519_),
    .B(_0520_),
    .Y(_0181_));
 OR3x1_ASAP7_75t_R _0925_ (.A(_0365_),
    .B(_0369_),
    .C(_0370_),
    .Y(_0521_));
 AND3x1_ASAP7_75t_R _0926_ (.A(_0358_),
    .B(_0379_),
    .C(_0367_),
    .Y(_0522_));
 AO21x1_ASAP7_75t_R _0927_ (.A1(_0521_),
    .A2(_0522_),
    .B(_0394_),
    .Y(_0523_));
 OA211x2_ASAP7_75t_R _0928_ (.A1(_0386_),
    .A2(_0387_),
    .B(_0390_),
    .C(_0360_),
    .Y(_0524_));
 AND4x1_ASAP7_75t_R _0929_ (.A(_0365_),
    .B(_0360_),
    .C(_0373_),
    .D(_0374_),
    .Y(_0525_));
 AND4x1_ASAP7_75t_R _0930_ (.A(_0358_),
    .B(_0365_),
    .C(_0390_),
    .D(_0367_),
    .Y(_0526_));
 OR3x1_ASAP7_75t_R _0931_ (.A(_0524_),
    .B(_0525_),
    .C(_0526_),
    .Y(_0527_));
 OAI21x1_ASAP7_75t_R _0932_ (.A1(_0523_),
    .A2(_0527_),
    .B(_0359_),
    .Y(_0528_));
 BUFx6f_ASAP7_75t_R _0933_ (.A(_0528_),
    .Y(_0529_));
 OR3x1_ASAP7_75t_R _0934_ (.A(net98),
    .B(_0369_),
    .C(_0370_),
    .Y(_0530_));
 AND3x1_ASAP7_75t_R _0935_ (.A(_0358_),
    .B(_0384_),
    .C(_0367_),
    .Y(_0531_));
 AO221x1_ASAP7_75t_R _0936_ (.A1(_0368_),
    .A2(_0376_),
    .B1(_0530_),
    .B2(_0531_),
    .C(_0371_),
    .Y(_0532_));
 BUFx6f_ASAP7_75t_R _0937_ (.A(_0532_),
    .Y(_0533_));
 NAND2x2_ASAP7_75t_R _0938_ (.A(_0360_),
    .B(_0533_),
    .Y(_0534_));
 BUFx3_ASAP7_75t_R _0939_ (.A(_0534_),
    .Y(_0535_));
 AND2x2_ASAP7_75t_R _0940_ (.A(_0362_),
    .B(net73),
    .Y(_0536_));
 BUFx6f_ASAP7_75t_R _0941_ (.A(_0533_),
    .Y(_0537_));
 OA21x2_ASAP7_75t_R _0942_ (.A1(_0523_),
    .A2(_0527_),
    .B(_0359_),
    .Y(_0538_));
 BUFx6f_ASAP7_75t_R _0943_ (.A(_0538_),
    .Y(_0539_));
 AO221x1_ASAP7_75t_R _0944_ (.A1(net1),
    .A2(_0535_),
    .B1(_0536_),
    .B2(_0537_),
    .C(_0539_),
    .Y(_0540_));
 BUFx6f_ASAP7_75t_R _0945_ (.A(_0403_),
    .Y(_0541_));
 OA211x2_ASAP7_75t_R _0946_ (.A1(net108),
    .A2(_0529_),
    .B(_0540_),
    .C(_0541_),
    .Y(_0182_));
 AND2x2_ASAP7_75t_R _0947_ (.A(_0362_),
    .B(net74),
    .Y(_0542_));
 AO221x1_ASAP7_75t_R _0948_ (.A1(net2),
    .A2(_0535_),
    .B1(_0542_),
    .B2(_0537_),
    .C(_0539_),
    .Y(_0543_));
 OA211x2_ASAP7_75t_R _0949_ (.A1(net109),
    .A2(_0529_),
    .B(_0543_),
    .C(_0541_),
    .Y(_0183_));
 AND2x2_ASAP7_75t_R _0950_ (.A(_0362_),
    .B(net75),
    .Y(_0544_));
 AO221x1_ASAP7_75t_R _0951_ (.A1(net3),
    .A2(_0535_),
    .B1(_0544_),
    .B2(_0537_),
    .C(_0539_),
    .Y(_0545_));
 OA211x2_ASAP7_75t_R _0952_ (.A1(net110),
    .A2(_0529_),
    .B(_0545_),
    .C(_0541_),
    .Y(_0184_));
 AND2x2_ASAP7_75t_R _0953_ (.A(_0362_),
    .B(net76),
    .Y(_0546_));
 AO221x1_ASAP7_75t_R _0954_ (.A1(net4),
    .A2(_0535_),
    .B1(_0546_),
    .B2(_0537_),
    .C(_0539_),
    .Y(_0547_));
 OA211x2_ASAP7_75t_R _0955_ (.A1(net111),
    .A2(_0529_),
    .B(_0547_),
    .C(_0541_),
    .Y(_0185_));
 AND2x2_ASAP7_75t_R _0956_ (.A(_0362_),
    .B(net77),
    .Y(_0548_));
 AO221x1_ASAP7_75t_R _0957_ (.A1(net5),
    .A2(_0535_),
    .B1(_0548_),
    .B2(_0537_),
    .C(_0539_),
    .Y(_0549_));
 BUFx3_ASAP7_75t_R _0958_ (.A(_0402_),
    .Y(_0550_));
 OA211x2_ASAP7_75t_R _0959_ (.A1(net112),
    .A2(_0529_),
    .B(_0549_),
    .C(_0550_),
    .Y(_0186_));
 AND2x2_ASAP7_75t_R _0960_ (.A(_0362_),
    .B(net78),
    .Y(_0551_));
 AO221x1_ASAP7_75t_R _0961_ (.A1(net6),
    .A2(_0535_),
    .B1(_0551_),
    .B2(_0537_),
    .C(_0539_),
    .Y(_0552_));
 OA211x2_ASAP7_75t_R _0962_ (.A1(net113),
    .A2(_0529_),
    .B(_0552_),
    .C(_0550_),
    .Y(_0187_));
 BUFx6f_ASAP7_75t_R _0963_ (.A(_0360_),
    .Y(_0553_));
 AND2x2_ASAP7_75t_R _0964_ (.A(_0553_),
    .B(net79),
    .Y(_0554_));
 AO221x1_ASAP7_75t_R _0965_ (.A1(net7),
    .A2(_0535_),
    .B1(_0554_),
    .B2(_0537_),
    .C(_0539_),
    .Y(_0555_));
 OA211x2_ASAP7_75t_R _0966_ (.A1(net114),
    .A2(_0529_),
    .B(_0555_),
    .C(_0550_),
    .Y(_0188_));
 AND2x2_ASAP7_75t_R _0967_ (.A(_0553_),
    .B(net80),
    .Y(_0556_));
 AO221x1_ASAP7_75t_R _0968_ (.A1(net8),
    .A2(_0535_),
    .B1(_0556_),
    .B2(_0537_),
    .C(_0539_),
    .Y(_0557_));
 OA211x2_ASAP7_75t_R _0969_ (.A1(net115),
    .A2(_0529_),
    .B(_0557_),
    .C(_0550_),
    .Y(_0189_));
 AND2x2_ASAP7_75t_R _0970_ (.A(_0553_),
    .B(net81),
    .Y(_0558_));
 AO221x1_ASAP7_75t_R _0971_ (.A1(net9),
    .A2(_0535_),
    .B1(_0558_),
    .B2(_0537_),
    .C(_0539_),
    .Y(_0559_));
 OA211x2_ASAP7_75t_R _0972_ (.A1(net116),
    .A2(_0529_),
    .B(_0559_),
    .C(_0550_),
    .Y(_0190_));
 AND2x2_ASAP7_75t_R _0973_ (.A(_0553_),
    .B(net82),
    .Y(_0560_));
 AO221x1_ASAP7_75t_R _0974_ (.A1(net10),
    .A2(_0535_),
    .B1(_0560_),
    .B2(_0537_),
    .C(_0539_),
    .Y(_0561_));
 OA211x2_ASAP7_75t_R _0975_ (.A1(net117),
    .A2(_0529_),
    .B(_0561_),
    .C(_0550_),
    .Y(_0191_));
 BUFx6f_ASAP7_75t_R _0976_ (.A(_0528_),
    .Y(_0562_));
 BUFx6f_ASAP7_75t_R _0977_ (.A(_0534_),
    .Y(_0563_));
 AND2x2_ASAP7_75t_R _0978_ (.A(_0553_),
    .B(net83),
    .Y(_0564_));
 BUFx6f_ASAP7_75t_R _0979_ (.A(_0533_),
    .Y(_0565_));
 BUFx6f_ASAP7_75t_R _0980_ (.A(_0538_),
    .Y(_0566_));
 AO221x1_ASAP7_75t_R _0981_ (.A1(net11),
    .A2(_0563_),
    .B1(_0564_),
    .B2(_0565_),
    .C(_0566_),
    .Y(_0567_));
 OA211x2_ASAP7_75t_R _0982_ (.A1(net118),
    .A2(_0562_),
    .B(_0567_),
    .C(_0550_),
    .Y(_0192_));
 AND2x2_ASAP7_75t_R _0983_ (.A(_0553_),
    .B(net84),
    .Y(_0568_));
 AO221x1_ASAP7_75t_R _0984_ (.A1(net12),
    .A2(_0563_),
    .B1(_0568_),
    .B2(_0565_),
    .C(_0566_),
    .Y(_0569_));
 OA211x2_ASAP7_75t_R _0985_ (.A1(net119),
    .A2(_0562_),
    .B(_0569_),
    .C(_0550_),
    .Y(_0193_));
 AND2x2_ASAP7_75t_R _0986_ (.A(_0553_),
    .B(net85),
    .Y(_0570_));
 AO221x1_ASAP7_75t_R _0987_ (.A1(net13),
    .A2(_0563_),
    .B1(_0570_),
    .B2(_0565_),
    .C(_0566_),
    .Y(_0571_));
 OA211x2_ASAP7_75t_R _0988_ (.A1(net120),
    .A2(_0562_),
    .B(_0571_),
    .C(_0550_),
    .Y(_0194_));
 AND2x2_ASAP7_75t_R _0989_ (.A(_0553_),
    .B(net86),
    .Y(_0572_));
 AO221x1_ASAP7_75t_R _0990_ (.A1(net14),
    .A2(_0563_),
    .B1(_0572_),
    .B2(_0565_),
    .C(_0566_),
    .Y(_0573_));
 OA211x2_ASAP7_75t_R _0991_ (.A1(net121),
    .A2(_0562_),
    .B(_0573_),
    .C(_0550_),
    .Y(_0195_));
 AND2x2_ASAP7_75t_R _0992_ (.A(_0553_),
    .B(net87),
    .Y(_0574_));
 AO221x1_ASAP7_75t_R _0993_ (.A1(net15),
    .A2(_0563_),
    .B1(_0574_),
    .B2(_0565_),
    .C(_0566_),
    .Y(_0575_));
 BUFx3_ASAP7_75t_R _0994_ (.A(_0402_),
    .Y(_0576_));
 OA211x2_ASAP7_75t_R _0995_ (.A1(net122),
    .A2(_0562_),
    .B(_0575_),
    .C(_0576_),
    .Y(_0196_));
 AND2x2_ASAP7_75t_R _0996_ (.A(_0553_),
    .B(net88),
    .Y(_0577_));
 AO221x1_ASAP7_75t_R _0997_ (.A1(net16),
    .A2(_0563_),
    .B1(_0577_),
    .B2(_0565_),
    .C(_0566_),
    .Y(_0578_));
 OA211x2_ASAP7_75t_R _0998_ (.A1(net123),
    .A2(_0562_),
    .B(_0578_),
    .C(_0576_),
    .Y(_0197_));
 BUFx6f_ASAP7_75t_R _0999_ (.A(_0360_),
    .Y(_0290_));
 AND2x2_ASAP7_75t_R _1000_ (.A(_0290_),
    .B(net89),
    .Y(_0291_));
 AO221x1_ASAP7_75t_R _1001_ (.A1(net17),
    .A2(_0563_),
    .B1(_0291_),
    .B2(_0565_),
    .C(_0566_),
    .Y(_0292_));
 OA211x2_ASAP7_75t_R _1002_ (.A1(net124),
    .A2(_0562_),
    .B(_0292_),
    .C(_0576_),
    .Y(_0198_));
 AND2x2_ASAP7_75t_R _1003_ (.A(_0290_),
    .B(net90),
    .Y(_0293_));
 AO221x1_ASAP7_75t_R _1004_ (.A1(net18),
    .A2(_0563_),
    .B1(_0293_),
    .B2(_0565_),
    .C(_0566_),
    .Y(_0294_));
 OA211x2_ASAP7_75t_R _1005_ (.A1(net125),
    .A2(_0562_),
    .B(_0294_),
    .C(_0576_),
    .Y(_0199_));
 AND2x2_ASAP7_75t_R _1006_ (.A(_0290_),
    .B(net91),
    .Y(_0295_));
 AO221x1_ASAP7_75t_R _1007_ (.A1(net19),
    .A2(_0563_),
    .B1(_0295_),
    .B2(_0565_),
    .C(_0566_),
    .Y(_0296_));
 OA211x2_ASAP7_75t_R _1008_ (.A1(net126),
    .A2(_0562_),
    .B(_0296_),
    .C(_0576_),
    .Y(_0200_));
 AND2x2_ASAP7_75t_R _1009_ (.A(_0290_),
    .B(net92),
    .Y(_0297_));
 AO221x1_ASAP7_75t_R _1010_ (.A1(net20),
    .A2(_0563_),
    .B1(_0297_),
    .B2(_0565_),
    .C(_0566_),
    .Y(_0298_));
 OA211x2_ASAP7_75t_R _1011_ (.A1(net127),
    .A2(_0562_),
    .B(_0298_),
    .C(_0576_),
    .Y(_0201_));
 BUFx6f_ASAP7_75t_R _1012_ (.A(_0528_),
    .Y(_0299_));
 BUFx6f_ASAP7_75t_R _1013_ (.A(_0534_),
    .Y(_0300_));
 AND2x2_ASAP7_75t_R _1014_ (.A(_0290_),
    .B(net93),
    .Y(_0301_));
 BUFx6f_ASAP7_75t_R _1015_ (.A(_0533_),
    .Y(_0302_));
 BUFx6f_ASAP7_75t_R _1016_ (.A(_0538_),
    .Y(_0303_));
 AO221x1_ASAP7_75t_R _1017_ (.A1(net21),
    .A2(_0300_),
    .B1(_0301_),
    .B2(_0302_),
    .C(_0303_),
    .Y(_0304_));
 OA211x2_ASAP7_75t_R _1018_ (.A1(net128),
    .A2(_0299_),
    .B(_0304_),
    .C(_0576_),
    .Y(_0202_));
 AND2x2_ASAP7_75t_R _1019_ (.A(_0290_),
    .B(net94),
    .Y(_0305_));
 AO221x1_ASAP7_75t_R _1020_ (.A1(net22),
    .A2(_0300_),
    .B1(_0305_),
    .B2(_0302_),
    .C(_0303_),
    .Y(_0306_));
 OA211x2_ASAP7_75t_R _1021_ (.A1(net129),
    .A2(_0299_),
    .B(_0306_),
    .C(_0576_),
    .Y(_0203_));
 AND2x2_ASAP7_75t_R _1022_ (.A(_0290_),
    .B(net95),
    .Y(_0307_));
 AO221x1_ASAP7_75t_R _1023_ (.A1(net23),
    .A2(_0300_),
    .B1(_0307_),
    .B2(_0302_),
    .C(_0303_),
    .Y(_0308_));
 OA211x2_ASAP7_75t_R _1024_ (.A1(net130),
    .A2(_0299_),
    .B(_0308_),
    .C(_0576_),
    .Y(_0204_));
 AND2x2_ASAP7_75t_R _1025_ (.A(_0290_),
    .B(net96),
    .Y(_0309_));
 AO221x1_ASAP7_75t_R _1026_ (.A1(net24),
    .A2(_0300_),
    .B1(_0309_),
    .B2(_0302_),
    .C(_0303_),
    .Y(_0310_));
 OA211x2_ASAP7_75t_R _1027_ (.A1(net131),
    .A2(_0299_),
    .B(_0310_),
    .C(_0576_),
    .Y(_0205_));
 AND2x2_ASAP7_75t_R _1028_ (.A(_0290_),
    .B(net97),
    .Y(_0311_));
 AO221x1_ASAP7_75t_R _1029_ (.A1(net25),
    .A2(_0300_),
    .B1(_0311_),
    .B2(_0302_),
    .C(_0303_),
    .Y(_0312_));
 BUFx3_ASAP7_75t_R _1030_ (.A(_0402_),
    .Y(_0313_));
 OA211x2_ASAP7_75t_R _1031_ (.A1(net132),
    .A2(_0299_),
    .B(_0312_),
    .C(_0313_),
    .Y(_0206_));
 NAND2x1_ASAP7_75t_R _1032_ (.A(_0373_),
    .B(_0374_),
    .Y(_0314_));
 AND2x4_ASAP7_75t_R _1033_ (.A(_0358_),
    .B(_0367_),
    .Y(_0315_));
 AND3x1_ASAP7_75t_R _1034_ (.A(_0379_),
    .B(_0314_),
    .C(_0315_),
    .Y(_0316_));
 AO21x1_ASAP7_75t_R _1035_ (.A1(_0362_),
    .A2(_0377_),
    .B(_0316_),
    .Y(_0317_));
 AO21x1_ASAP7_75t_R _1036_ (.A1(_0361_),
    .A2(net98),
    .B(_0388_),
    .Y(_0318_));
 OA21x2_ASAP7_75t_R _1037_ (.A1(_0314_),
    .A2(_0315_),
    .B(_0318_),
    .Y(_0319_));
 AO221x1_ASAP7_75t_R _1038_ (.A1(net26),
    .A2(_0300_),
    .B1(_0317_),
    .B2(_0359_),
    .C(_0319_),
    .Y(_0320_));
 OA211x2_ASAP7_75t_R _1039_ (.A1(_0365_),
    .A2(_0299_),
    .B(_0320_),
    .C(_0313_),
    .Y(_0207_));
 AND2x2_ASAP7_75t_R _1040_ (.A(_0290_),
    .B(net99),
    .Y(_0321_));
 AO221x1_ASAP7_75t_R _1041_ (.A1(net27),
    .A2(_0300_),
    .B1(_0321_),
    .B2(_0302_),
    .C(_0303_),
    .Y(_0322_));
 OA211x2_ASAP7_75t_R _1042_ (.A1(net133),
    .A2(_0299_),
    .B(_0322_),
    .C(_0313_),
    .Y(_0208_));
 AND2x2_ASAP7_75t_R _1043_ (.A(_0361_),
    .B(net100),
    .Y(_0323_));
 AO221x1_ASAP7_75t_R _1044_ (.A1(net28),
    .A2(_0300_),
    .B1(_0323_),
    .B2(_0302_),
    .C(_0303_),
    .Y(_0324_));
 OA211x2_ASAP7_75t_R _1045_ (.A1(net134),
    .A2(_0299_),
    .B(_0324_),
    .C(_0313_),
    .Y(_0209_));
 OR3x1_ASAP7_75t_R _1046_ (.A(_0365_),
    .B(_0362_),
    .C(_0315_),
    .Y(_0325_));
 AO21x1_ASAP7_75t_R _1047_ (.A1(_0362_),
    .A2(_0368_),
    .B(_0359_),
    .Y(_0326_));
 AO21x1_ASAP7_75t_R _1048_ (.A1(_0325_),
    .A2(_0326_),
    .B(_0375_),
    .Y(_0327_));
 AND2x2_ASAP7_75t_R _1049_ (.A(_0493_),
    .B(_0327_),
    .Y(_0210_));
 AND2x2_ASAP7_75t_R _1050_ (.A(_0361_),
    .B(net101),
    .Y(_0328_));
 AO221x1_ASAP7_75t_R _1051_ (.A1(net30),
    .A2(_0300_),
    .B1(_0328_),
    .B2(_0302_),
    .C(_0303_),
    .Y(_0329_));
 OA211x2_ASAP7_75t_R _1052_ (.A1(net135),
    .A2(_0299_),
    .B(_0329_),
    .C(_0313_),
    .Y(_0211_));
 AND2x2_ASAP7_75t_R _1053_ (.A(_0361_),
    .B(net102),
    .Y(_0330_));
 AO221x1_ASAP7_75t_R _1054_ (.A1(net31),
    .A2(_0300_),
    .B1(_0330_),
    .B2(_0302_),
    .C(_0303_),
    .Y(_0331_));
 OA211x2_ASAP7_75t_R _1055_ (.A1(net136),
    .A2(_0299_),
    .B(_0331_),
    .C(_0313_),
    .Y(_0212_));
 AND2x2_ASAP7_75t_R _1056_ (.A(_0361_),
    .B(net103),
    .Y(_0332_));
 AO221x1_ASAP7_75t_R _1057_ (.A1(net32),
    .A2(_0534_),
    .B1(_0332_),
    .B2(_0302_),
    .C(_0303_),
    .Y(_0333_));
 OA211x2_ASAP7_75t_R _1058_ (.A1(net137),
    .A2(_0528_),
    .B(_0333_),
    .C(_0313_),
    .Y(_0213_));
 AND2x2_ASAP7_75t_R _1059_ (.A(_0361_),
    .B(net104),
    .Y(_0334_));
 AO221x1_ASAP7_75t_R _1060_ (.A1(net33),
    .A2(_0534_),
    .B1(_0334_),
    .B2(_0533_),
    .C(_0538_),
    .Y(_0335_));
 OA211x2_ASAP7_75t_R _1061_ (.A1(net138),
    .A2(_0528_),
    .B(_0335_),
    .C(_0313_),
    .Y(_0214_));
 AND2x2_ASAP7_75t_R _1062_ (.A(_0361_),
    .B(net105),
    .Y(_0336_));
 AO221x1_ASAP7_75t_R _1063_ (.A1(net34),
    .A2(_0534_),
    .B1(_0336_),
    .B2(_0533_),
    .C(_0538_),
    .Y(_0337_));
 OA211x2_ASAP7_75t_R _1064_ (.A1(net139),
    .A2(_0528_),
    .B(_0337_),
    .C(_0313_),
    .Y(_0215_));
 AND2x2_ASAP7_75t_R _1065_ (.A(_0361_),
    .B(net106),
    .Y(_0338_));
 AO221x1_ASAP7_75t_R _1066_ (.A1(net35),
    .A2(_0534_),
    .B1(_0338_),
    .B2(_0533_),
    .C(_0538_),
    .Y(_0339_));
 OA211x2_ASAP7_75t_R _1067_ (.A1(net140),
    .A2(_0528_),
    .B(_0339_),
    .C(_0313_),
    .Y(_0216_));
 AND2x2_ASAP7_75t_R _1068_ (.A(_0361_),
    .B(net107),
    .Y(_0340_));
 AO221x1_ASAP7_75t_R _1069_ (.A1(net36),
    .A2(_0534_),
    .B1(_0340_),
    .B2(_0533_),
    .C(_0538_),
    .Y(_0341_));
 OA211x2_ASAP7_75t_R _1070_ (.A1(net141),
    .A2(_0528_),
    .B(_0341_),
    .C(_0410_),
    .Y(_0217_));
 AND2x2_ASAP7_75t_R _1071_ (.A(_0493_),
    .B(net1),
    .Y(_0218_));
 AND2x2_ASAP7_75t_R _1072_ (.A(_0493_),
    .B(net2),
    .Y(_0219_));
 AND2x2_ASAP7_75t_R _1073_ (.A(_0493_),
    .B(net3),
    .Y(_0220_));
 BUFx6f_ASAP7_75t_R _1074_ (.A(_0403_),
    .Y(_0342_));
 AND2x2_ASAP7_75t_R _1075_ (.A(_0342_),
    .B(net4),
    .Y(_0221_));
 AND2x2_ASAP7_75t_R _1076_ (.A(_0342_),
    .B(net5),
    .Y(_0222_));
 AND2x2_ASAP7_75t_R _1077_ (.A(_0342_),
    .B(net6),
    .Y(_0223_));
 AND2x2_ASAP7_75t_R _1078_ (.A(_0342_),
    .B(net7),
    .Y(_0224_));
 AND2x2_ASAP7_75t_R _1079_ (.A(_0342_),
    .B(net8),
    .Y(_0225_));
 AND2x2_ASAP7_75t_R _1080_ (.A(_0342_),
    .B(net9),
    .Y(_0226_));
 AND2x2_ASAP7_75t_R _1081_ (.A(_0342_),
    .B(net10),
    .Y(_0227_));
 AND2x2_ASAP7_75t_R _1082_ (.A(_0342_),
    .B(net11),
    .Y(_0228_));
 AND2x2_ASAP7_75t_R _1083_ (.A(_0342_),
    .B(net12),
    .Y(_0229_));
 AND2x2_ASAP7_75t_R _1084_ (.A(_0342_),
    .B(net13),
    .Y(_0230_));
 BUFx6f_ASAP7_75t_R _1085_ (.A(_0403_),
    .Y(_0343_));
 AND2x2_ASAP7_75t_R _1086_ (.A(_0343_),
    .B(net14),
    .Y(_0231_));
 AND2x2_ASAP7_75t_R _1087_ (.A(_0343_),
    .B(net15),
    .Y(_0232_));
 AND2x2_ASAP7_75t_R _1088_ (.A(_0343_),
    .B(net16),
    .Y(_0233_));
 AND2x2_ASAP7_75t_R _1089_ (.A(_0343_),
    .B(net17),
    .Y(_0234_));
 AND2x2_ASAP7_75t_R _1090_ (.A(_0343_),
    .B(net18),
    .Y(_0235_));
 AND2x2_ASAP7_75t_R _1091_ (.A(_0343_),
    .B(net19),
    .Y(_0236_));
 AND2x2_ASAP7_75t_R _1092_ (.A(_0343_),
    .B(net20),
    .Y(_0237_));
 AND2x2_ASAP7_75t_R _1093_ (.A(_0343_),
    .B(net21),
    .Y(_0238_));
 AND2x2_ASAP7_75t_R _1094_ (.A(_0343_),
    .B(net22),
    .Y(_0239_));
 AND2x2_ASAP7_75t_R _1095_ (.A(_0343_),
    .B(net23),
    .Y(_0240_));
 BUFx6f_ASAP7_75t_R _1096_ (.A(_0403_),
    .Y(_0344_));
 AND2x2_ASAP7_75t_R _1097_ (.A(_0344_),
    .B(net24),
    .Y(_0241_));
 AND2x2_ASAP7_75t_R _1098_ (.A(_0344_),
    .B(net25),
    .Y(_0242_));
 AND2x2_ASAP7_75t_R _1099_ (.A(net26),
    .B(_0493_),
    .Y(_0243_));
 AND2x2_ASAP7_75t_R _1100_ (.A(net27),
    .B(_0493_),
    .Y(_0244_));
 AND2x2_ASAP7_75t_R _1101_ (.A(net28),
    .B(_0493_),
    .Y(_0245_));
 INVx1_ASAP7_75t_R _1102_ (.A(net26),
    .Y(_0345_));
 OR3x1_ASAP7_75t_R _1103_ (.A(_0345_),
    .B(_0364_),
    .C(_0369_),
    .Y(_0346_));
 AO32x1_ASAP7_75t_R _1104_ (.A1(_0375_),
    .A2(_0315_),
    .A3(_0318_),
    .B1(_0346_),
    .B2(net29),
    .Y(_0347_));
 AND2x2_ASAP7_75t_R _1105_ (.A(_0344_),
    .B(_0347_),
    .Y(_0246_));
 AND2x2_ASAP7_75t_R _1106_ (.A(_0344_),
    .B(net30),
    .Y(_0247_));
 AND2x2_ASAP7_75t_R _1107_ (.A(_0344_),
    .B(net31),
    .Y(_0248_));
 AND2x2_ASAP7_75t_R _1108_ (.A(_0344_),
    .B(net32),
    .Y(_0249_));
 AND2x2_ASAP7_75t_R _1109_ (.A(_0344_),
    .B(net33),
    .Y(_0250_));
 AND2x2_ASAP7_75t_R _1110_ (.A(_0344_),
    .B(net34),
    .Y(_0251_));
 AND2x2_ASAP7_75t_R _1111_ (.A(_0344_),
    .B(net35),
    .Y(_0252_));
 AND2x2_ASAP7_75t_R _1112_ (.A(_0344_),
    .B(net36),
    .Y(_0253_));
 BUFx6f_ASAP7_75t_R _1113_ (.A(_0403_),
    .Y(_0348_));
 AO21x1_ASAP7_75t_R _1114_ (.A1(_0360_),
    .A2(_0390_),
    .B(_0376_),
    .Y(_0349_));
 OR2x2_ASAP7_75t_R _1115_ (.A(_0364_),
    .B(_0387_),
    .Y(_0350_));
 AO32x1_ASAP7_75t_R _1116_ (.A1(_0375_),
    .A2(_0315_),
    .A3(_0349_),
    .B1(_0350_),
    .B2(_0358_),
    .Y(_0351_));
 BUFx6f_ASAP7_75t_R _1117_ (.A(_0351_),
    .Y(_0352_));
 BUFx6f_ASAP7_75t_R _1118_ (.A(_0352_),
    .Y(_0353_));
 AND3x1_ASAP7_75t_R _1119_ (.A(_0348_),
    .B(net37),
    .C(_0353_),
    .Y(_0254_));
 AND3x1_ASAP7_75t_R _1120_ (.A(_0348_),
    .B(net38),
    .C(_0353_),
    .Y(_0255_));
 AND3x1_ASAP7_75t_R _1121_ (.A(_0348_),
    .B(net39),
    .C(_0353_),
    .Y(_0256_));
 AND3x1_ASAP7_75t_R _1122_ (.A(_0348_),
    .B(net40),
    .C(_0353_),
    .Y(_0257_));
 AND3x1_ASAP7_75t_R _1123_ (.A(_0348_),
    .B(net41),
    .C(_0353_),
    .Y(_0258_));
 AND3x1_ASAP7_75t_R _1124_ (.A(_0348_),
    .B(net42),
    .C(_0353_),
    .Y(_0259_));
 AND3x1_ASAP7_75t_R _1125_ (.A(_0348_),
    .B(net43),
    .C(_0353_),
    .Y(_0260_));
 AND3x1_ASAP7_75t_R _1126_ (.A(_0348_),
    .B(net44),
    .C(_0353_),
    .Y(_0261_));
 AND3x1_ASAP7_75t_R _1127_ (.A(_0348_),
    .B(net45),
    .C(_0353_),
    .Y(_0262_));
 BUFx6f_ASAP7_75t_R _1128_ (.A(_0403_),
    .Y(_0354_));
 BUFx6f_ASAP7_75t_R _1129_ (.A(_0352_),
    .Y(_0355_));
 AND3x1_ASAP7_75t_R _1130_ (.A(_0354_),
    .B(net46),
    .C(_0355_),
    .Y(_0263_));
 AND3x1_ASAP7_75t_R _1131_ (.A(_0354_),
    .B(net47),
    .C(_0355_),
    .Y(_0264_));
 AND3x1_ASAP7_75t_R _1132_ (.A(_0354_),
    .B(net48),
    .C(_0355_),
    .Y(_0265_));
 AND3x1_ASAP7_75t_R _1133_ (.A(_0354_),
    .B(net49),
    .C(_0355_),
    .Y(_0266_));
 AND3x1_ASAP7_75t_R _1134_ (.A(_0354_),
    .B(net50),
    .C(_0355_),
    .Y(_0267_));
 AND3x1_ASAP7_75t_R _1135_ (.A(_0354_),
    .B(net51),
    .C(_0355_),
    .Y(_0268_));
 AND3x1_ASAP7_75t_R _1136_ (.A(_0354_),
    .B(net52),
    .C(_0355_),
    .Y(_0269_));
 AND3x1_ASAP7_75t_R _1137_ (.A(_0354_),
    .B(net53),
    .C(_0355_),
    .Y(_0270_));
 AND3x1_ASAP7_75t_R _1138_ (.A(_0354_),
    .B(net54),
    .C(_0355_),
    .Y(_0271_));
 AND3x1_ASAP7_75t_R _1139_ (.A(_0354_),
    .B(net55),
    .C(_0355_),
    .Y(_0272_));
 BUFx6f_ASAP7_75t_R _1140_ (.A(_0402_),
    .Y(_0356_));
 BUFx6f_ASAP7_75t_R _1141_ (.A(_0352_),
    .Y(_0357_));
 AND3x1_ASAP7_75t_R _1142_ (.A(_0356_),
    .B(net56),
    .C(_0357_),
    .Y(_0273_));
 AND3x1_ASAP7_75t_R _1143_ (.A(_0356_),
    .B(net57),
    .C(_0357_),
    .Y(_0274_));
 AND3x1_ASAP7_75t_R _1144_ (.A(_0356_),
    .B(net58),
    .C(_0357_),
    .Y(_0275_));
 AND3x1_ASAP7_75t_R _1145_ (.A(_0356_),
    .B(net59),
    .C(_0357_),
    .Y(_0276_));
 AND3x1_ASAP7_75t_R _1146_ (.A(_0356_),
    .B(net60),
    .C(_0357_),
    .Y(_0277_));
 AND3x1_ASAP7_75t_R _1147_ (.A(_0356_),
    .B(net61),
    .C(_0357_),
    .Y(_0278_));
 AND3x1_ASAP7_75t_R _1148_ (.A(net62),
    .B(_0541_),
    .C(_0357_),
    .Y(_0279_));
 AND3x1_ASAP7_75t_R _1149_ (.A(net63),
    .B(_0541_),
    .C(_0357_),
    .Y(_0280_));
 AND3x1_ASAP7_75t_R _1150_ (.A(net64),
    .B(_0541_),
    .C(_0357_),
    .Y(_0281_));
 AND2x2_ASAP7_75t_R _1151_ (.A(_0348_),
    .B(_0353_),
    .Y(_0282_));
 AND3x1_ASAP7_75t_R _1152_ (.A(_0356_),
    .B(net65),
    .C(_0357_),
    .Y(_0283_));
 AND3x1_ASAP7_75t_R _1153_ (.A(_0356_),
    .B(net66),
    .C(_0352_),
    .Y(_0284_));
 AND3x1_ASAP7_75t_R _1154_ (.A(_0356_),
    .B(net67),
    .C(_0352_),
    .Y(_0285_));
 AND3x1_ASAP7_75t_R _1155_ (.A(_0356_),
    .B(net68),
    .C(_0352_),
    .Y(_0286_));
 AND3x1_ASAP7_75t_R _1156_ (.A(_0541_),
    .B(net69),
    .C(_0352_),
    .Y(_0287_));
 AND3x1_ASAP7_75t_R _1157_ (.A(_0541_),
    .B(net70),
    .C(_0352_),
    .Y(_0288_));
 AND3x1_ASAP7_75t_R _1158_ (.A(_0541_),
    .B(net71),
    .C(_0352_),
    .Y(_0289_));
 BUFx4_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx2_ASAP7_75t_R _1160_ (.A(net287),
    .Y(l_o[35]));
 BUFx2_ASAP7_75t_R _1161_ (.A(net288),
    .Y(r_o[35]));
 BUFx2_ASAP7_75t_R _1162_ (.A(net289),
    .Y(u0_o[35]));
 BUFx2_ASAP7_75t_R _1163_ (.A(net290),
    .Y(u1_o[35]));
 DFFHQNx1_ASAP7_75t_R \done_sig$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .D(_0000_),
    .QN(_0145_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .D(_0146_),
    .QN(_0144_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[10]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .D(_0147_),
    .QN(_0143_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[11]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .D(_0148_),
    .QN(_0142_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[12]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .D(_0149_),
    .QN(_0141_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[13]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0150_),
    .QN(_0140_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[14]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0151_),
    .QN(_0139_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[15]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0152_),
    .QN(_0138_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[16]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .D(_0153_),
    .QN(_0137_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[17]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0154_),
    .QN(_0136_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[18]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .D(_0155_),
    .QN(_0135_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[19]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .D(_0156_),
    .QN(_0134_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .D(_0157_),
    .QN(_0133_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[20]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .D(_0158_),
    .QN(_0132_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[21]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .D(_0159_),
    .QN(_0131_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[22]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .D(_0160_),
    .QN(_0130_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[23]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .D(_0161_),
    .QN(_0129_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[24]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0162_),
    .QN(_0128_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[25]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0163_),
    .QN(_0127_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[26]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0164_),
    .QN(_0126_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[27]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .D(_0165_),
    .QN(_0125_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[28]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .D(_0166_),
    .QN(_0124_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[29]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .D(_0167_),
    .QN(_0123_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .D(_0168_),
    .QN(_0122_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[30]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .D(_0169_),
    .QN(_0121_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .D(_0170_),
    .QN(_0120_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_4_0_0_clk),
    .D(_0171_),
    .QN(_0119_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_4_3_0_clk),
    .D(_0172_),
    .QN(_0118_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_4_3_0_clk),
    .D(_0173_),
    .QN(_0117_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_4_0_0_clk),
    .D(_0174_),
    .QN(_0116_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .D(_0175_),
    .QN(_0115_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .D(_0176_),
    .QN(_0114_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[5]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .D(_0177_),
    .QN(_0113_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[6]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .D(_0178_),
    .QN(_0112_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[7]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .D(_0179_),
    .QN(_0111_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[8]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .D(_0180_),
    .QN(_0110_));
 DFFHQNx1_ASAP7_75t_R \l_o_r[9]$_SDFF_PP0_  (.CLK(clknet_4_3_0_clk),
    .D(_0181_),
    .QN(_0109_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .D(_0182_),
    .QN(_0108_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[10]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .D(_0183_),
    .QN(_0107_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[11]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .D(_0184_),
    .QN(_0106_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[12]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0185_),
    .QN(_0105_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[13]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0186_),
    .QN(_0104_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[14]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0187_),
    .QN(_0103_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[15]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0188_),
    .QN(_0102_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[16]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .D(_0189_),
    .QN(_0101_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[17]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .D(_0190_),
    .QN(_0100_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[18]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .D(_0191_),
    .QN(_0099_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[19]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .D(_0192_),
    .QN(_0098_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .D(_0193_),
    .QN(_0097_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[20]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .D(_0194_),
    .QN(_0096_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[21]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .D(_0195_),
    .QN(_0095_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[22]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0196_),
    .QN(_0094_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[23]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .D(_0197_),
    .QN(_0093_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[24]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0198_),
    .QN(_0092_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[25]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0199_),
    .QN(_0091_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[26]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0200_),
    .QN(_0090_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[27]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .D(_0201_),
    .QN(_0089_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[28]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .D(_0202_),
    .QN(_0088_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[29]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .D(_0203_),
    .QN(_0087_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .D(_0204_),
    .QN(_0086_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[30]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .D(_0205_),
    .QN(_0085_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .D(_0206_),
    .QN(_0084_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .D(_0207_),
    .QN(_0083_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_4_3_0_clk),
    .D(_0208_),
    .QN(_0082_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_4_3_0_clk),
    .D(_0209_),
    .QN(_0081_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_4_0_0_clk),
    .D(_0210_),
    .QN(_0080_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .D(_0211_),
    .QN(_0079_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .D(_0212_),
    .QN(_0078_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[5]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .D(_0213_),
    .QN(_0077_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[6]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .D(_0214_),
    .QN(_0076_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[7]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .D(_0215_),
    .QN(_0075_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[8]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .D(_0216_),
    .QN(_0074_));
 DFFHQNx1_ASAP7_75t_R \r_o_r[9]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .D(_0217_),
    .QN(_0073_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .D(_0218_),
    .QN(_0072_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[10]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .D(_0219_),
    .QN(_0071_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[11]$_SDFF_PP0_  (.CLK(clknet_4_0_0_clk),
    .D(_0220_),
    .QN(_0070_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[12]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .D(_0221_),
    .QN(_0069_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[13]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0222_),
    .QN(_0068_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[14]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0223_),
    .QN(_0067_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[15]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0224_),
    .QN(_0066_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[16]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .D(_0225_),
    .QN(_0065_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[17]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .D(_0226_),
    .QN(_0064_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[18]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .D(_0227_),
    .QN(_0063_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[19]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .D(_0228_),
    .QN(_0062_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .D(_0229_),
    .QN(_0061_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[20]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .D(_0230_),
    .QN(_0060_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[21]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .D(_0231_),
    .QN(_0059_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[22]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .D(_0232_),
    .QN(_0058_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[23]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .D(_0233_),
    .QN(_0057_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[24]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0234_),
    .QN(_0056_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[25]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .D(_0235_),
    .QN(_0055_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[26]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0236_),
    .QN(_0054_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[27]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .D(_0237_),
    .QN(_0053_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[28]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .D(_0238_),
    .QN(_0052_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[29]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .D(_0239_),
    .QN(_0051_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .D(_0240_),
    .QN(_0050_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[30]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .D(_0241_),
    .QN(_0049_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .D(_0242_),
    .QN(_0048_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_4_0_0_clk),
    .D(_0243_),
    .QN(_0047_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .D(_0244_),
    .QN(_0046_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .D(_0245_),
    .QN(_0045_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_4_0_0_clk),
    .D(_0246_),
    .QN(_0044_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .D(_0247_),
    .QN(_0043_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .D(_0248_),
    .QN(_0042_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[5]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .D(_0249_),
    .QN(_0041_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[6]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .D(_0250_),
    .QN(_0040_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[7]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .D(_0251_),
    .QN(_0039_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[8]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .D(_0252_),
    .QN(_0038_));
 DFFHQNx1_ASAP7_75t_R \u0_o_r[9]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .D(_0253_),
    .QN(_0037_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[0]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .D(_0254_),
    .QN(_0036_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[10]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .D(_0255_),
    .QN(_0035_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[11]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .D(_0256_),
    .QN(_0034_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[12]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .D(_0257_),
    .QN(_0033_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[13]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0258_),
    .QN(_0032_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[14]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0259_),
    .QN(_0031_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[15]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0260_),
    .QN(_0030_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[16]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .D(_0261_),
    .QN(_0029_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[17]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .D(_0262_),
    .QN(_0028_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[18]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .D(_0263_),
    .QN(_0027_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[19]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .D(_0264_),
    .QN(_0026_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[1]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .D(_0265_),
    .QN(_0025_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[20]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .D(_0266_),
    .QN(_0024_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[21]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .D(_0267_),
    .QN(_0023_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[22]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .D(_0268_),
    .QN(_0022_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[23]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .D(_0269_),
    .QN(_0021_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[24]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0270_),
    .QN(_0020_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[25]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0271_),
    .QN(_0019_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[26]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .D(_0272_),
    .QN(_0018_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[27]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .D(_0273_),
    .QN(_0017_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[28]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .D(_0274_),
    .QN(_0016_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[29]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .D(_0275_),
    .QN(_0015_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[2]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .D(_0276_),
    .QN(_0014_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[30]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .D(_0277_),
    .QN(_0013_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[31]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .D(_0278_),
    .QN(_0012_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[32]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .D(_0279_),
    .QN(_0011_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[33]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .D(_0280_),
    .QN(_0010_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[34]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .D(_0281_),
    .QN(_0009_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[36]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .D(_0282_),
    .QN(_0008_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[3]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .D(_0283_),
    .QN(_0007_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[4]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .D(_0284_),
    .QN(_0006_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[5]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .D(_0285_),
    .QN(_0005_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[6]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .D(_0286_),
    .QN(_0004_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[7]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .D(_0287_),
    .QN(_0003_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[8]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .D(_0288_),
    .QN(_0002_));
 DFFHQNx1_ASAP7_75t_R \u1_o_r[9]$_SDFF_PP0_  (.CLK(clknet_4_3_0_clk),
    .D(_0289_),
    .QN(_0001_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_109 ();
 BUFx3_ASAP7_75t_R input1 (.A(l_i[0]),
    .Y(net1));
 BUFx3_ASAP7_75t_R input2 (.A(l_i[10]),
    .Y(net2));
 BUFx3_ASAP7_75t_R input3 (.A(l_i[11]),
    .Y(net3));
 BUFx3_ASAP7_75t_R input4 (.A(l_i[12]),
    .Y(net4));
 BUFx3_ASAP7_75t_R input5 (.A(l_i[13]),
    .Y(net5));
 BUFx3_ASAP7_75t_R input6 (.A(l_i[14]),
    .Y(net6));
 BUFx3_ASAP7_75t_R input7 (.A(l_i[15]),
    .Y(net7));
 BUFx3_ASAP7_75t_R input8 (.A(l_i[16]),
    .Y(net8));
 BUFx3_ASAP7_75t_R input9 (.A(l_i[17]),
    .Y(net9));
 BUFx3_ASAP7_75t_R input10 (.A(l_i[18]),
    .Y(net10));
 BUFx3_ASAP7_75t_R input11 (.A(l_i[19]),
    .Y(net11));
 BUFx3_ASAP7_75t_R input12 (.A(l_i[1]),
    .Y(net12));
 BUFx3_ASAP7_75t_R input13 (.A(l_i[20]),
    .Y(net13));
 BUFx3_ASAP7_75t_R input14 (.A(l_i[21]),
    .Y(net14));
 BUFx3_ASAP7_75t_R input15 (.A(l_i[22]),
    .Y(net15));
 BUFx3_ASAP7_75t_R input16 (.A(l_i[23]),
    .Y(net16));
 BUFx3_ASAP7_75t_R input17 (.A(l_i[24]),
    .Y(net17));
 BUFx3_ASAP7_75t_R input18 (.A(l_i[25]),
    .Y(net18));
 BUFx3_ASAP7_75t_R input19 (.A(l_i[26]),
    .Y(net19));
 BUFx3_ASAP7_75t_R input20 (.A(l_i[27]),
    .Y(net20));
 BUFx3_ASAP7_75t_R input21 (.A(l_i[28]),
    .Y(net21));
 BUFx3_ASAP7_75t_R input22 (.A(l_i[29]),
    .Y(net22));
 BUFx3_ASAP7_75t_R input23 (.A(l_i[2]),
    .Y(net23));
 BUFx3_ASAP7_75t_R input24 (.A(l_i[30]),
    .Y(net24));
 BUFx3_ASAP7_75t_R input25 (.A(l_i[31]),
    .Y(net25));
 BUFx3_ASAP7_75t_R input26 (.A(l_i[32]),
    .Y(net26));
 BUFx3_ASAP7_75t_R input27 (.A(l_i[33]),
    .Y(net27));
 BUFx3_ASAP7_75t_R input28 (.A(l_i[34]),
    .Y(net28));
 BUFx3_ASAP7_75t_R input29 (.A(l_i[36]),
    .Y(net29));
 BUFx3_ASAP7_75t_R input30 (.A(l_i[3]),
    .Y(net30));
 BUFx3_ASAP7_75t_R input31 (.A(l_i[4]),
    .Y(net31));
 BUFx3_ASAP7_75t_R input32 (.A(l_i[5]),
    .Y(net32));
 BUFx3_ASAP7_75t_R input33 (.A(l_i[6]),
    .Y(net33));
 BUFx3_ASAP7_75t_R input34 (.A(l_i[7]),
    .Y(net34));
 BUFx3_ASAP7_75t_R input35 (.A(l_i[8]),
    .Y(net35));
 BUFx3_ASAP7_75t_R input36 (.A(l_i[9]),
    .Y(net36));
 BUFx3_ASAP7_75t_R input37 (.A(r_i[0]),
    .Y(net37));
 BUFx3_ASAP7_75t_R input38 (.A(r_i[10]),
    .Y(net38));
 BUFx3_ASAP7_75t_R input39 (.A(r_i[11]),
    .Y(net39));
 BUFx3_ASAP7_75t_R input40 (.A(r_i[12]),
    .Y(net40));
 BUFx3_ASAP7_75t_R input41 (.A(r_i[13]),
    .Y(net41));
 BUFx3_ASAP7_75t_R input42 (.A(r_i[14]),
    .Y(net42));
 BUFx3_ASAP7_75t_R input43 (.A(r_i[15]),
    .Y(net43));
 BUFx3_ASAP7_75t_R input44 (.A(r_i[16]),
    .Y(net44));
 BUFx3_ASAP7_75t_R input45 (.A(r_i[17]),
    .Y(net45));
 BUFx3_ASAP7_75t_R input46 (.A(r_i[18]),
    .Y(net46));
 BUFx3_ASAP7_75t_R input47 (.A(r_i[19]),
    .Y(net47));
 BUFx3_ASAP7_75t_R input48 (.A(r_i[1]),
    .Y(net48));
 BUFx3_ASAP7_75t_R input49 (.A(r_i[20]),
    .Y(net49));
 BUFx3_ASAP7_75t_R input50 (.A(r_i[21]),
    .Y(net50));
 BUFx3_ASAP7_75t_R input51 (.A(r_i[22]),
    .Y(net51));
 BUFx3_ASAP7_75t_R input52 (.A(r_i[23]),
    .Y(net52));
 BUFx3_ASAP7_75t_R input53 (.A(r_i[24]),
    .Y(net53));
 BUFx3_ASAP7_75t_R input54 (.A(r_i[25]),
    .Y(net54));
 BUFx3_ASAP7_75t_R input55 (.A(r_i[26]),
    .Y(net55));
 BUFx3_ASAP7_75t_R input56 (.A(r_i[27]),
    .Y(net56));
 BUFx3_ASAP7_75t_R input57 (.A(r_i[28]),
    .Y(net57));
 BUFx3_ASAP7_75t_R input58 (.A(r_i[29]),
    .Y(net58));
 BUFx3_ASAP7_75t_R input59 (.A(r_i[2]),
    .Y(net59));
 BUFx3_ASAP7_75t_R input60 (.A(r_i[30]),
    .Y(net60));
 BUFx3_ASAP7_75t_R input61 (.A(r_i[31]),
    .Y(net61));
 BUFx3_ASAP7_75t_R input62 (.A(r_i[32]),
    .Y(net62));
 BUFx3_ASAP7_75t_R input63 (.A(r_i[33]),
    .Y(net63));
 BUFx3_ASAP7_75t_R input64 (.A(r_i[34]),
    .Y(net64));
 BUFx3_ASAP7_75t_R input65 (.A(r_i[3]),
    .Y(net65));
 BUFx3_ASAP7_75t_R input66 (.A(r_i[4]),
    .Y(net66));
 BUFx3_ASAP7_75t_R input67 (.A(r_i[5]),
    .Y(net67));
 BUFx3_ASAP7_75t_R input68 (.A(r_i[6]),
    .Y(net68));
 BUFx3_ASAP7_75t_R input69 (.A(r_i[7]),
    .Y(net69));
 BUFx3_ASAP7_75t_R input70 (.A(r_i[8]),
    .Y(net70));
 BUFx3_ASAP7_75t_R input71 (.A(r_i[9]),
    .Y(net71));
 BUFx3_ASAP7_75t_R input72 (.A(rst),
    .Y(net72));
 BUFx3_ASAP7_75t_R input73 (.A(u0_i[0]),
    .Y(net73));
 BUFx3_ASAP7_75t_R input74 (.A(u0_i[10]),
    .Y(net74));
 BUFx3_ASAP7_75t_R input75 (.A(u0_i[11]),
    .Y(net75));
 BUFx3_ASAP7_75t_R input76 (.A(u0_i[12]),
    .Y(net76));
 BUFx3_ASAP7_75t_R input77 (.A(u0_i[13]),
    .Y(net77));
 BUFx3_ASAP7_75t_R input78 (.A(u0_i[14]),
    .Y(net78));
 BUFx3_ASAP7_75t_R input79 (.A(u0_i[15]),
    .Y(net79));
 BUFx3_ASAP7_75t_R input80 (.A(u0_i[16]),
    .Y(net80));
 BUFx3_ASAP7_75t_R input81 (.A(u0_i[17]),
    .Y(net81));
 BUFx3_ASAP7_75t_R input82 (.A(u0_i[18]),
    .Y(net82));
 BUFx3_ASAP7_75t_R input83 (.A(u0_i[19]),
    .Y(net83));
 BUFx3_ASAP7_75t_R input84 (.A(u0_i[1]),
    .Y(net84));
 BUFx3_ASAP7_75t_R input85 (.A(u0_i[20]),
    .Y(net85));
 BUFx3_ASAP7_75t_R input86 (.A(u0_i[21]),
    .Y(net86));
 BUFx3_ASAP7_75t_R input87 (.A(u0_i[22]),
    .Y(net87));
 BUFx3_ASAP7_75t_R input88 (.A(u0_i[23]),
    .Y(net88));
 BUFx3_ASAP7_75t_R input89 (.A(u0_i[24]),
    .Y(net89));
 BUFx3_ASAP7_75t_R input90 (.A(u0_i[25]),
    .Y(net90));
 BUFx3_ASAP7_75t_R input91 (.A(u0_i[26]),
    .Y(net91));
 BUFx3_ASAP7_75t_R input92 (.A(u0_i[27]),
    .Y(net92));
 BUFx3_ASAP7_75t_R input93 (.A(u0_i[28]),
    .Y(net93));
 BUFx3_ASAP7_75t_R input94 (.A(u0_i[29]),
    .Y(net94));
 BUFx3_ASAP7_75t_R input95 (.A(u0_i[2]),
    .Y(net95));
 BUFx3_ASAP7_75t_R input96 (.A(u0_i[30]),
    .Y(net96));
 BUFx3_ASAP7_75t_R input97 (.A(u0_i[31]),
    .Y(net97));
 BUFx3_ASAP7_75t_R input98 (.A(u0_i[32]),
    .Y(net98));
 BUFx3_ASAP7_75t_R input99 (.A(u0_i[33]),
    .Y(net99));
 BUFx3_ASAP7_75t_R input100 (.A(u0_i[34]),
    .Y(net100));
 BUFx3_ASAP7_75t_R input101 (.A(u0_i[3]),
    .Y(net101));
 BUFx3_ASAP7_75t_R input102 (.A(u0_i[4]),
    .Y(net102));
 BUFx3_ASAP7_75t_R input103 (.A(u0_i[5]),
    .Y(net103));
 BUFx3_ASAP7_75t_R input104 (.A(u0_i[6]),
    .Y(net104));
 BUFx3_ASAP7_75t_R input105 (.A(u0_i[7]),
    .Y(net105));
 BUFx3_ASAP7_75t_R input106 (.A(u0_i[8]),
    .Y(net106));
 BUFx3_ASAP7_75t_R input107 (.A(u0_i[9]),
    .Y(net107));
 BUFx3_ASAP7_75t_R input108 (.A(u1_i[0]),
    .Y(net108));
 BUFx3_ASAP7_75t_R input109 (.A(u1_i[10]),
    .Y(net109));
 BUFx3_ASAP7_75t_R input110 (.A(u1_i[11]),
    .Y(net110));
 BUFx3_ASAP7_75t_R input111 (.A(u1_i[12]),
    .Y(net111));
 BUFx3_ASAP7_75t_R input112 (.A(u1_i[13]),
    .Y(net112));
 BUFx3_ASAP7_75t_R input113 (.A(u1_i[14]),
    .Y(net113));
 BUFx3_ASAP7_75t_R input114 (.A(u1_i[15]),
    .Y(net114));
 BUFx3_ASAP7_75t_R input115 (.A(u1_i[16]),
    .Y(net115));
 BUFx3_ASAP7_75t_R input116 (.A(u1_i[17]),
    .Y(net116));
 BUFx3_ASAP7_75t_R input117 (.A(u1_i[18]),
    .Y(net117));
 BUFx3_ASAP7_75t_R input118 (.A(u1_i[19]),
    .Y(net118));
 BUFx3_ASAP7_75t_R input119 (.A(u1_i[1]),
    .Y(net119));
 BUFx3_ASAP7_75t_R input120 (.A(u1_i[20]),
    .Y(net120));
 BUFx3_ASAP7_75t_R input121 (.A(u1_i[21]),
    .Y(net121));
 BUFx3_ASAP7_75t_R input122 (.A(u1_i[22]),
    .Y(net122));
 BUFx3_ASAP7_75t_R input123 (.A(u1_i[23]),
    .Y(net123));
 BUFx3_ASAP7_75t_R input124 (.A(u1_i[24]),
    .Y(net124));
 BUFx3_ASAP7_75t_R input125 (.A(u1_i[25]),
    .Y(net125));
 BUFx3_ASAP7_75t_R input126 (.A(u1_i[26]),
    .Y(net126));
 BUFx3_ASAP7_75t_R input127 (.A(u1_i[27]),
    .Y(net127));
 BUFx3_ASAP7_75t_R input128 (.A(u1_i[28]),
    .Y(net128));
 BUFx3_ASAP7_75t_R input129 (.A(u1_i[29]),
    .Y(net129));
 BUFx3_ASAP7_75t_R input130 (.A(u1_i[2]),
    .Y(net130));
 BUFx3_ASAP7_75t_R input131 (.A(u1_i[30]),
    .Y(net131));
 BUFx3_ASAP7_75t_R input132 (.A(u1_i[31]),
    .Y(net132));
 BUFx3_ASAP7_75t_R input133 (.A(u1_i[33]),
    .Y(net133));
 BUFx3_ASAP7_75t_R input134 (.A(u1_i[34]),
    .Y(net134));
 BUFx3_ASAP7_75t_R input135 (.A(u1_i[3]),
    .Y(net135));
 BUFx3_ASAP7_75t_R input136 (.A(u1_i[4]),
    .Y(net136));
 BUFx3_ASAP7_75t_R input137 (.A(u1_i[5]),
    .Y(net137));
 BUFx3_ASAP7_75t_R input138 (.A(u1_i[6]),
    .Y(net138));
 BUFx3_ASAP7_75t_R input139 (.A(u1_i[7]),
    .Y(net139));
 BUFx3_ASAP7_75t_R input140 (.A(u1_i[8]),
    .Y(net140));
 BUFx3_ASAP7_75t_R input141 (.A(u1_i[9]),
    .Y(net141));
 BUFx3_ASAP7_75t_R output142 (.A(net142),
    .Y(done));
 BUFx3_ASAP7_75t_R output143 (.A(net143),
    .Y(l_o[0]));
 BUFx3_ASAP7_75t_R output144 (.A(net144),
    .Y(l_o[10]));
 BUFx3_ASAP7_75t_R output145 (.A(net145),
    .Y(l_o[11]));
 BUFx3_ASAP7_75t_R output146 (.A(net146),
    .Y(l_o[12]));
 BUFx3_ASAP7_75t_R output147 (.A(net147),
    .Y(l_o[13]));
 BUFx3_ASAP7_75t_R output148 (.A(net148),
    .Y(l_o[14]));
 BUFx3_ASAP7_75t_R output149 (.A(net149),
    .Y(l_o[15]));
 BUFx3_ASAP7_75t_R output150 (.A(net150),
    .Y(l_o[16]));
 BUFx3_ASAP7_75t_R output151 (.A(net151),
    .Y(l_o[17]));
 BUFx3_ASAP7_75t_R output152 (.A(net152),
    .Y(l_o[18]));
 BUFx3_ASAP7_75t_R output153 (.A(net153),
    .Y(l_o[19]));
 BUFx3_ASAP7_75t_R output154 (.A(net154),
    .Y(l_o[1]));
 BUFx3_ASAP7_75t_R output155 (.A(net155),
    .Y(l_o[20]));
 BUFx3_ASAP7_75t_R output156 (.A(net156),
    .Y(l_o[21]));
 BUFx3_ASAP7_75t_R output157 (.A(net157),
    .Y(l_o[22]));
 BUFx3_ASAP7_75t_R output158 (.A(net158),
    .Y(l_o[23]));
 BUFx3_ASAP7_75t_R output159 (.A(net159),
    .Y(l_o[24]));
 BUFx3_ASAP7_75t_R output160 (.A(net160),
    .Y(l_o[25]));
 BUFx3_ASAP7_75t_R output161 (.A(net161),
    .Y(l_o[26]));
 BUFx3_ASAP7_75t_R output162 (.A(net162),
    .Y(l_o[27]));
 BUFx3_ASAP7_75t_R output163 (.A(net163),
    .Y(l_o[28]));
 BUFx3_ASAP7_75t_R output164 (.A(net164),
    .Y(l_o[29]));
 BUFx3_ASAP7_75t_R output165 (.A(net165),
    .Y(l_o[2]));
 BUFx3_ASAP7_75t_R output166 (.A(net166),
    .Y(l_o[30]));
 BUFx3_ASAP7_75t_R output167 (.A(net167),
    .Y(l_o[31]));
 BUFx3_ASAP7_75t_R output168 (.A(net168),
    .Y(l_o[32]));
 BUFx3_ASAP7_75t_R output169 (.A(net169),
    .Y(l_o[33]));
 BUFx3_ASAP7_75t_R output170 (.A(net170),
    .Y(l_o[34]));
 BUFx3_ASAP7_75t_R output171 (.A(net171),
    .Y(l_o[36]));
 BUFx3_ASAP7_75t_R output172 (.A(net172),
    .Y(l_o[3]));
 BUFx3_ASAP7_75t_R output173 (.A(net173),
    .Y(l_o[4]));
 BUFx3_ASAP7_75t_R output174 (.A(net174),
    .Y(l_o[5]));
 BUFx3_ASAP7_75t_R output175 (.A(net175),
    .Y(l_o[6]));
 BUFx3_ASAP7_75t_R output176 (.A(net176),
    .Y(l_o[7]));
 BUFx3_ASAP7_75t_R output177 (.A(net177),
    .Y(l_o[8]));
 BUFx3_ASAP7_75t_R output178 (.A(net178),
    .Y(l_o[9]));
 BUFx3_ASAP7_75t_R output179 (.A(net179),
    .Y(r_o[0]));
 BUFx3_ASAP7_75t_R output180 (.A(net180),
    .Y(r_o[10]));
 BUFx3_ASAP7_75t_R output181 (.A(net181),
    .Y(r_o[11]));
 BUFx3_ASAP7_75t_R output182 (.A(net182),
    .Y(r_o[12]));
 BUFx3_ASAP7_75t_R output183 (.A(net183),
    .Y(r_o[13]));
 BUFx3_ASAP7_75t_R output184 (.A(net184),
    .Y(r_o[14]));
 BUFx3_ASAP7_75t_R output185 (.A(net185),
    .Y(r_o[15]));
 BUFx3_ASAP7_75t_R output186 (.A(net186),
    .Y(r_o[16]));
 BUFx3_ASAP7_75t_R output187 (.A(net187),
    .Y(r_o[17]));
 BUFx3_ASAP7_75t_R output188 (.A(net188),
    .Y(r_o[18]));
 BUFx3_ASAP7_75t_R output189 (.A(net189),
    .Y(r_o[19]));
 BUFx3_ASAP7_75t_R output190 (.A(net190),
    .Y(r_o[1]));
 BUFx3_ASAP7_75t_R output191 (.A(net191),
    .Y(r_o[20]));
 BUFx3_ASAP7_75t_R output192 (.A(net192),
    .Y(r_o[21]));
 BUFx3_ASAP7_75t_R output193 (.A(net193),
    .Y(r_o[22]));
 BUFx3_ASAP7_75t_R output194 (.A(net194),
    .Y(r_o[23]));
 BUFx3_ASAP7_75t_R output195 (.A(net195),
    .Y(r_o[24]));
 BUFx3_ASAP7_75t_R output196 (.A(net196),
    .Y(r_o[25]));
 BUFx3_ASAP7_75t_R output197 (.A(net197),
    .Y(r_o[26]));
 BUFx3_ASAP7_75t_R output198 (.A(net198),
    .Y(r_o[27]));
 BUFx3_ASAP7_75t_R output199 (.A(net199),
    .Y(r_o[28]));
 BUFx3_ASAP7_75t_R output200 (.A(net200),
    .Y(r_o[29]));
 BUFx3_ASAP7_75t_R output201 (.A(net201),
    .Y(r_o[2]));
 BUFx3_ASAP7_75t_R output202 (.A(net202),
    .Y(r_o[30]));
 BUFx3_ASAP7_75t_R output203 (.A(net203),
    .Y(r_o[31]));
 BUFx3_ASAP7_75t_R output204 (.A(net204),
    .Y(r_o[32]));
 BUFx3_ASAP7_75t_R output205 (.A(net205),
    .Y(r_o[33]));
 BUFx3_ASAP7_75t_R output206 (.A(net206),
    .Y(r_o[34]));
 BUFx3_ASAP7_75t_R output207 (.A(net207),
    .Y(r_o[36]));
 BUFx3_ASAP7_75t_R output208 (.A(net208),
    .Y(r_o[3]));
 BUFx3_ASAP7_75t_R output209 (.A(net209),
    .Y(r_o[4]));
 BUFx3_ASAP7_75t_R output210 (.A(net210),
    .Y(r_o[5]));
 BUFx3_ASAP7_75t_R output211 (.A(net211),
    .Y(r_o[6]));
 BUFx3_ASAP7_75t_R output212 (.A(net212),
    .Y(r_o[7]));
 BUFx3_ASAP7_75t_R output213 (.A(net213),
    .Y(r_o[8]));
 BUFx3_ASAP7_75t_R output214 (.A(net214),
    .Y(r_o[9]));
 BUFx3_ASAP7_75t_R output215 (.A(net215),
    .Y(u0_o[0]));
 BUFx3_ASAP7_75t_R output216 (.A(net216),
    .Y(u0_o[10]));
 BUFx3_ASAP7_75t_R output217 (.A(net217),
    .Y(u0_o[11]));
 BUFx3_ASAP7_75t_R output218 (.A(net218),
    .Y(u0_o[12]));
 BUFx3_ASAP7_75t_R output219 (.A(net219),
    .Y(u0_o[13]));
 BUFx3_ASAP7_75t_R output220 (.A(net220),
    .Y(u0_o[14]));
 BUFx3_ASAP7_75t_R output221 (.A(net221),
    .Y(u0_o[15]));
 BUFx3_ASAP7_75t_R output222 (.A(net222),
    .Y(u0_o[16]));
 BUFx3_ASAP7_75t_R output223 (.A(net223),
    .Y(u0_o[17]));
 BUFx3_ASAP7_75t_R output224 (.A(net224),
    .Y(u0_o[18]));
 BUFx3_ASAP7_75t_R output225 (.A(net225),
    .Y(u0_o[19]));
 BUFx3_ASAP7_75t_R output226 (.A(net226),
    .Y(u0_o[1]));
 BUFx3_ASAP7_75t_R output227 (.A(net227),
    .Y(u0_o[20]));
 BUFx3_ASAP7_75t_R output228 (.A(net228),
    .Y(u0_o[21]));
 BUFx3_ASAP7_75t_R output229 (.A(net229),
    .Y(u0_o[22]));
 BUFx3_ASAP7_75t_R output230 (.A(net230),
    .Y(u0_o[23]));
 BUFx3_ASAP7_75t_R output231 (.A(net231),
    .Y(u0_o[24]));
 BUFx3_ASAP7_75t_R output232 (.A(net232),
    .Y(u0_o[25]));
 BUFx3_ASAP7_75t_R output233 (.A(net233),
    .Y(u0_o[26]));
 BUFx3_ASAP7_75t_R output234 (.A(net234),
    .Y(u0_o[27]));
 BUFx3_ASAP7_75t_R output235 (.A(net235),
    .Y(u0_o[28]));
 BUFx3_ASAP7_75t_R output236 (.A(net236),
    .Y(u0_o[29]));
 BUFx3_ASAP7_75t_R output237 (.A(net237),
    .Y(u0_o[2]));
 BUFx3_ASAP7_75t_R output238 (.A(net238),
    .Y(u0_o[30]));
 BUFx3_ASAP7_75t_R output239 (.A(net239),
    .Y(u0_o[31]));
 BUFx3_ASAP7_75t_R output240 (.A(net240),
    .Y(u0_o[32]));
 BUFx3_ASAP7_75t_R output241 (.A(net241),
    .Y(u0_o[33]));
 BUFx3_ASAP7_75t_R output242 (.A(net242),
    .Y(u0_o[34]));
 BUFx3_ASAP7_75t_R output243 (.A(net243),
    .Y(u0_o[36]));
 BUFx3_ASAP7_75t_R output244 (.A(net244),
    .Y(u0_o[3]));
 BUFx3_ASAP7_75t_R output245 (.A(net245),
    .Y(u0_o[4]));
 BUFx3_ASAP7_75t_R output246 (.A(net246),
    .Y(u0_o[5]));
 BUFx3_ASAP7_75t_R output247 (.A(net247),
    .Y(u0_o[6]));
 BUFx3_ASAP7_75t_R output248 (.A(net248),
    .Y(u0_o[7]));
 BUFx3_ASAP7_75t_R output249 (.A(net249),
    .Y(u0_o[8]));
 BUFx3_ASAP7_75t_R output250 (.A(net250),
    .Y(u0_o[9]));
 BUFx3_ASAP7_75t_R output251 (.A(net251),
    .Y(u1_o[0]));
 BUFx3_ASAP7_75t_R output252 (.A(net252),
    .Y(u1_o[10]));
 BUFx3_ASAP7_75t_R output253 (.A(net253),
    .Y(u1_o[11]));
 BUFx3_ASAP7_75t_R output254 (.A(net254),
    .Y(u1_o[12]));
 BUFx3_ASAP7_75t_R output255 (.A(net255),
    .Y(u1_o[13]));
 BUFx3_ASAP7_75t_R output256 (.A(net256),
    .Y(u1_o[14]));
 BUFx3_ASAP7_75t_R output257 (.A(net257),
    .Y(u1_o[15]));
 BUFx3_ASAP7_75t_R output258 (.A(net258),
    .Y(u1_o[16]));
 BUFx3_ASAP7_75t_R output259 (.A(net259),
    .Y(u1_o[17]));
 BUFx3_ASAP7_75t_R output260 (.A(net260),
    .Y(u1_o[18]));
 BUFx3_ASAP7_75t_R output261 (.A(net261),
    .Y(u1_o[19]));
 BUFx3_ASAP7_75t_R output262 (.A(net262),
    .Y(u1_o[1]));
 BUFx3_ASAP7_75t_R output263 (.A(net263),
    .Y(u1_o[20]));
 BUFx3_ASAP7_75t_R output264 (.A(net264),
    .Y(u1_o[21]));
 BUFx3_ASAP7_75t_R output265 (.A(net265),
    .Y(u1_o[22]));
 BUFx3_ASAP7_75t_R output266 (.A(net266),
    .Y(u1_o[23]));
 BUFx3_ASAP7_75t_R output267 (.A(net267),
    .Y(u1_o[24]));
 BUFx3_ASAP7_75t_R output268 (.A(net268),
    .Y(u1_o[25]));
 BUFx3_ASAP7_75t_R output269 (.A(net269),
    .Y(u1_o[26]));
 BUFx3_ASAP7_75t_R output270 (.A(net270),
    .Y(u1_o[27]));
 BUFx3_ASAP7_75t_R output271 (.A(net271),
    .Y(u1_o[28]));
 BUFx3_ASAP7_75t_R output272 (.A(net272),
    .Y(u1_o[29]));
 BUFx3_ASAP7_75t_R output273 (.A(net273),
    .Y(u1_o[2]));
 BUFx3_ASAP7_75t_R output274 (.A(net274),
    .Y(u1_o[30]));
 BUFx3_ASAP7_75t_R output275 (.A(net275),
    .Y(u1_o[31]));
 BUFx3_ASAP7_75t_R output276 (.A(net276),
    .Y(u1_o[32]));
 BUFx3_ASAP7_75t_R output277 (.A(net277),
    .Y(u1_o[33]));
 BUFx3_ASAP7_75t_R output278 (.A(net278),
    .Y(u1_o[34]));
 BUFx3_ASAP7_75t_R output279 (.A(net279),
    .Y(u1_o[36]));
 BUFx3_ASAP7_75t_R output280 (.A(net280),
    .Y(u1_o[3]));
 BUFx3_ASAP7_75t_R output281 (.A(net281),
    .Y(u1_o[4]));
 BUFx3_ASAP7_75t_R output282 (.A(net282),
    .Y(u1_o[5]));
 BUFx3_ASAP7_75t_R output283 (.A(net283),
    .Y(u1_o[6]));
 BUFx3_ASAP7_75t_R output284 (.A(net284),
    .Y(u1_o[7]));
 BUFx3_ASAP7_75t_R output285 (.A(net285),
    .Y(u1_o[8]));
 BUFx3_ASAP7_75t_R output286 (.A(net286),
    .Y(u1_o[9]));
 TIELOx1_ASAP7_75t_R _1160__287 (.L(net287));
 TIELOx1_ASAP7_75t_R _1161__288 (.L(net288));
 TIELOx1_ASAP7_75t_R _1162__289 (.L(net289));
 TIELOx1_ASAP7_75t_R _1163__290 (.L(net290));
 BUFx10_ASAP7_75t_R clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_0_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_1_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_2_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_3_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_4_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_5_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_6_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_7_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_8_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_9_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_10_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_11_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_12_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_13_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_14_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Y(clknet_4_15_0_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload0 (.A(clknet_4_0_0_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload1 (.A(clknet_4_1_0_clk));
 INVx3_ASAP7_75t_R clkload2 (.A(clknet_4_2_0_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload3 (.A(clknet_4_3_0_clk));
 BUFx24_ASAP7_75t_R clkload4 (.A(clknet_4_4_0_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload5 (.A(clknet_4_6_0_clk));
 BUFx24_ASAP7_75t_R clkload6 (.A(clknet_4_7_0_clk));
 INVx3_ASAP7_75t_R clkload7 (.A(clknet_4_8_0_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload8 (.A(clknet_4_9_0_clk));
 BUFx24_ASAP7_75t_R clkload9 (.A(clknet_4_10_0_clk));
 INVx6_ASAP7_75t_R clkload10 (.A(clknet_4_11_0_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload11 (.A(clknet_4_12_0_clk));
 BUFx24_ASAP7_75t_R clkload12 (.A(clknet_4_13_0_clk));
 INVx5_ASAP7_75t_R clkload13 (.A(clknet_4_14_0_clk));
 BUFx12_ASAP7_75t_R clkload14 (.A(clknet_4_15_0_clk));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 FILLER_ASAP7_75t_R FILLER_0_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_54 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72 ();
 FILLER_ASAP7_75t_R FILLER_0_85 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243 ();
 DECAPx4_ASAP7_75t_R FILLER_0_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx6_ASAP7_75t_R FILLER_1_68 ();
 FILLER_ASAP7_75t_R FILLER_1_82 ();
 DECAPx4_ASAP7_75t_R FILLER_1_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_245 ();
 DECAPx6_ASAP7_75t_R FILLER_1_258 ();
 DECAPx1_ASAP7_75t_R FILLER_1_272 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_2_46 ();
 DECAPx6_ASAP7_75t_R FILLER_2_68 ();
 FILLER_ASAP7_75t_R FILLER_2_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_91 ();
 FILLER_ASAP7_75t_R FILLER_2_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_183 ();
 DECAPx2_ASAP7_75t_R FILLER_2_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_242 ();
 DECAPx10_ASAP7_75t_R FILLER_2_249 ();
 DECAPx1_ASAP7_75t_R FILLER_2_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_275 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_68 ();
 FILLER_ASAP7_75t_R FILLER_3_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_92 ();
 FILLER_ASAP7_75t_R FILLER_3_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_107 ();
 FILLER_ASAP7_75t_R FILLER_3_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_151 ();
 FILLER_ASAP7_75t_R FILLER_3_158 ();
 DECAPx1_ASAP7_75t_R FILLER_3_250 ();
 DECAPx2_ASAP7_75t_R FILLER_3_260 ();
 FILLER_ASAP7_75t_R FILLER_3_266 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_68 ();
 DECAPx2_ASAP7_75t_R FILLER_4_90 ();
 FILLER_ASAP7_75t_R FILLER_4_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_98 ();
 FILLER_ASAP7_75t_R FILLER_4_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_107 ();
 FILLER_ASAP7_75t_R FILLER_4_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_137 ();
 DECAPx1_ASAP7_75t_R FILLER_4_151 ();
 FILLER_ASAP7_75t_R FILLER_4_161 ();
 FILLER_ASAP7_75t_R FILLER_4_169 ();
 DECAPx2_ASAP7_75t_R FILLER_4_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_196 ();
 FILLER_ASAP7_75t_R FILLER_4_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_211 ();
 DECAPx6_ASAP7_75t_R FILLER_4_247 ();
 DECAPx2_ASAP7_75t_R FILLER_4_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_267 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 FILLER_ASAP7_75t_R FILLER_5_24 ();
 FILLER_ASAP7_75t_R FILLER_5_46 ();
 DECAPx6_ASAP7_75t_R FILLER_5_51 ();
 DECAPx1_ASAP7_75t_R FILLER_5_65 ();
 DECAPx2_ASAP7_75t_R FILLER_5_95 ();
 FILLER_ASAP7_75t_R FILLER_5_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_103 ();
 DECAPx6_ASAP7_75t_R FILLER_5_107 ();
 FILLER_ASAP7_75t_R FILLER_5_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_162 ();
 DECAPx6_ASAP7_75t_R FILLER_5_169 ();
 FILLER_ASAP7_75t_R FILLER_5_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_185 ();
 DECAPx1_ASAP7_75t_R FILLER_5_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_216 ();
 FILLER_ASAP7_75t_R FILLER_5_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_226 ();
 DECAPx6_ASAP7_75t_R FILLER_5_250 ();
 FILLER_ASAP7_75t_R FILLER_5_267 ();
 FILLER_ASAP7_75t_R FILLER_5_274 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx6_ASAP7_75t_R FILLER_6_24 ();
 FILLER_ASAP7_75t_R FILLER_6_38 ();
 DECAPx10_ASAP7_75t_R FILLER_6_43 ();
 DECAPx1_ASAP7_75t_R FILLER_6_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_101 ();
 FILLER_ASAP7_75t_R FILLER_6_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_128 ();
 DECAPx1_ASAP7_75t_R FILLER_6_135 ();
 DECAPx2_ASAP7_75t_R FILLER_6_192 ();
 DECAPx10_ASAP7_75t_R FILLER_6_231 ();
 DECAPx6_ASAP7_75t_R FILLER_6_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_275 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx1_ASAP7_75t_R FILLER_7_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_28 ();
 DECAPx6_ASAP7_75t_R FILLER_7_52 ();
 DECAPx1_ASAP7_75t_R FILLER_7_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_70 ();
 DECAPx4_ASAP7_75t_R FILLER_7_77 ();
 DECAPx6_ASAP7_75t_R FILLER_7_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_168 ();
 DECAPx2_ASAP7_75t_R FILLER_7_176 ();
 FILLER_ASAP7_75t_R FILLER_7_182 ();
 DECAPx2_ASAP7_75t_R FILLER_7_204 ();
 DECAPx10_ASAP7_75t_R FILLER_7_224 ();
 DECAPx10_ASAP7_75t_R FILLER_7_246 ();
 FILLER_ASAP7_75t_R FILLER_7_268 ();
 DECAPx6_ASAP7_75t_R FILLER_8_2 ();
 DECAPx6_ASAP7_75t_R FILLER_8_26 ();
 FILLER_ASAP7_75t_R FILLER_8_40 ();
 DECAPx1_ASAP7_75t_R FILLER_8_48 ();
 DECAPx1_ASAP7_75t_R FILLER_8_70 ();
 DECAPx10_ASAP7_75t_R FILLER_8_97 ();
 DECAPx4_ASAP7_75t_R FILLER_8_119 ();
 FILLER_ASAP7_75t_R FILLER_8_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_131 ();
 DECAPx6_ASAP7_75t_R FILLER_8_150 ();
 DECAPx2_ASAP7_75t_R FILLER_8_175 ();
 FILLER_ASAP7_75t_R FILLER_8_181 ();
 DECAPx4_ASAP7_75t_R FILLER_8_189 ();
 FILLER_ASAP7_75t_R FILLER_8_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_201 ();
 DECAPx1_ASAP7_75t_R FILLER_8_205 ();
 FILLER_ASAP7_75t_R FILLER_8_215 ();
 FILLER_ASAP7_75t_R FILLER_8_235 ();
 DECAPx1_ASAP7_75t_R FILLER_8_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_261 ();
 DECAPx1_ASAP7_75t_R FILLER_8_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_269 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx1_ASAP7_75t_R FILLER_9_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_46 ();
 DECAPx1_ASAP7_75t_R FILLER_9_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_64 ();
 DECAPx1_ASAP7_75t_R FILLER_9_71 ();
 DECAPx6_ASAP7_75t_R FILLER_9_88 ();
 DECAPx2_ASAP7_75t_R FILLER_9_102 ();
 DECAPx6_ASAP7_75t_R FILLER_9_111 ();
 DECAPx2_ASAP7_75t_R FILLER_9_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_131 ();
 DECAPx6_ASAP7_75t_R FILLER_9_150 ();
 DECAPx1_ASAP7_75t_R FILLER_9_164 ();
 DECAPx6_ASAP7_75t_R FILLER_9_188 ();
 FILLER_ASAP7_75t_R FILLER_9_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_216 ();
 FILLER_ASAP7_75t_R FILLER_9_235 ();
 FILLER_ASAP7_75t_R FILLER_9_257 ();
 DECAPx1_ASAP7_75t_R FILLER_9_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_266 ();
 DECAPx6_ASAP7_75t_R FILLER_10_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_27 ();
 FILLER_ASAP7_75t_R FILLER_10_44 ();
 FILLER_ASAP7_75t_R FILLER_10_80 ();
 DECAPx4_ASAP7_75t_R FILLER_10_92 ();
 FILLER_ASAP7_75t_R FILLER_10_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_104 ();
 DECAPx2_ASAP7_75t_R FILLER_10_115 ();
 DECAPx10_ASAP7_75t_R FILLER_10_124 ();
 DECAPx6_ASAP7_75t_R FILLER_10_146 ();
 FILLER_ASAP7_75t_R FILLER_10_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_162 ();
 DECAPx10_ASAP7_75t_R FILLER_10_185 ();
 DECAPx6_ASAP7_75t_R FILLER_10_207 ();
 DECAPx1_ASAP7_75t_R FILLER_10_221 ();
 DECAPx2_ASAP7_75t_R FILLER_10_231 ();
 FILLER_ASAP7_75t_R FILLER_10_237 ();
 FILLER_ASAP7_75t_R FILLER_10_262 ();
 DECAPx4_ASAP7_75t_R FILLER_11_2 ();
 DECAPx2_ASAP7_75t_R FILLER_11_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_24 ();
 FILLER_ASAP7_75t_R FILLER_11_68 ();
 DECAPx4_ASAP7_75t_R FILLER_11_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_94 ();
 DECAPx2_ASAP7_75t_R FILLER_11_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_141 ();
 DECAPx6_ASAP7_75t_R FILLER_11_145 ();
 DECAPx4_ASAP7_75t_R FILLER_11_195 ();
 DECAPx1_ASAP7_75t_R FILLER_11_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_226 ();
 DECAPx4_ASAP7_75t_R FILLER_11_235 ();
 DECAPx4_ASAP7_75t_R FILLER_11_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_275 ();
 DECAPx4_ASAP7_75t_R FILLER_12_2 ();
 FILLER_ASAP7_75t_R FILLER_12_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_14 ();
 DECAPx1_ASAP7_75t_R FILLER_12_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_25 ();
 FILLER_ASAP7_75t_R FILLER_12_36 ();
 FILLER_ASAP7_75t_R FILLER_12_56 ();
 FILLER_ASAP7_75t_R FILLER_12_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_108 ();
 FILLER_ASAP7_75t_R FILLER_12_123 ();
 FILLER_ASAP7_75t_R FILLER_12_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_143 ();
 FILLER_ASAP7_75t_R FILLER_12_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_166 ();
 DECAPx6_ASAP7_75t_R FILLER_12_213 ();
 DECAPx1_ASAP7_75t_R FILLER_12_227 ();
 FILLER_ASAP7_75t_R FILLER_12_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_269 ();
 DECAPx10_ASAP7_75t_R FILLER_13_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_24 ();
 FILLER_ASAP7_75t_R FILLER_13_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_72 ();
 FILLER_ASAP7_75t_R FILLER_13_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_140 ();
 FILLER_ASAP7_75t_R FILLER_13_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_151 ();
 FILLER_ASAP7_75t_R FILLER_13_175 ();
 DECAPx2_ASAP7_75t_R FILLER_13_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_197 ();
 DECAPx4_ASAP7_75t_R FILLER_13_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_263 ();
 DECAPx1_ASAP7_75t_R FILLER_14_2 ();
 DECAPx4_ASAP7_75t_R FILLER_14_12 ();
 FILLER_ASAP7_75t_R FILLER_14_22 ();
 FILLER_ASAP7_75t_R FILLER_14_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_55 ();
 FILLER_ASAP7_75t_R FILLER_14_99 ();
 FILLER_ASAP7_75t_R FILLER_14_111 ();
 DECAPx1_ASAP7_75t_R FILLER_14_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_154 ();
 DECAPx6_ASAP7_75t_R FILLER_14_161 ();
 DECAPx2_ASAP7_75t_R FILLER_14_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_181 ();
 DECAPx1_ASAP7_75t_R FILLER_14_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_192 ();
 FILLER_ASAP7_75t_R FILLER_14_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_201 ();
 FILLER_ASAP7_75t_R FILLER_14_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_224 ();
 DECAPx1_ASAP7_75t_R FILLER_14_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_275 ();
 DECAPx4_ASAP7_75t_R FILLER_15_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_12 ();
 DECAPx2_ASAP7_75t_R FILLER_15_24 ();
 FILLER_ASAP7_75t_R FILLER_15_30 ();
 DECAPx2_ASAP7_75t_R FILLER_15_61 ();
 FILLER_ASAP7_75t_R FILLER_15_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_69 ();
 FILLER_ASAP7_75t_R FILLER_15_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_99 ();
 DECAPx10_ASAP7_75t_R FILLER_15_120 ();
 DECAPx2_ASAP7_75t_R FILLER_15_142 ();
 FILLER_ASAP7_75t_R FILLER_15_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_150 ();
 DECAPx2_ASAP7_75t_R FILLER_15_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_207 ();
 DECAPx2_ASAP7_75t_R FILLER_15_259 ();
 FILLER_ASAP7_75t_R FILLER_15_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_17 ();
 FILLER_ASAP7_75t_R FILLER_16_51 ();
 DECAPx6_ASAP7_75t_R FILLER_16_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_71 ();
 DECAPx10_ASAP7_75t_R FILLER_16_76 ();
 DECAPx1_ASAP7_75t_R FILLER_16_98 ();
 DECAPx6_ASAP7_75t_R FILLER_16_108 ();
 DECAPx2_ASAP7_75t_R FILLER_16_122 ();
 DECAPx2_ASAP7_75t_R FILLER_16_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_144 ();
 DECAPx10_ASAP7_75t_R FILLER_16_148 ();
 DECAPx10_ASAP7_75t_R FILLER_16_170 ();
 DECAPx2_ASAP7_75t_R FILLER_16_192 ();
 FILLER_ASAP7_75t_R FILLER_16_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_216 ();
 DECAPx1_ASAP7_75t_R FILLER_16_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_231 ();
 FILLER_ASAP7_75t_R FILLER_16_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_260 ();
 DECAPx2_ASAP7_75t_R FILLER_16_264 ();
 FILLER_ASAP7_75t_R FILLER_17_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_4 ();
 DECAPx4_ASAP7_75t_R FILLER_17_25 ();
 DECAPx1_ASAP7_75t_R FILLER_17_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_60 ();
 DECAPx1_ASAP7_75t_R FILLER_17_84 ();
 DECAPx4_ASAP7_75t_R FILLER_17_95 ();
 FILLER_ASAP7_75t_R FILLER_17_105 ();
 DECAPx2_ASAP7_75t_R FILLER_17_113 ();
 FILLER_ASAP7_75t_R FILLER_17_119 ();
 DECAPx2_ASAP7_75t_R FILLER_17_151 ();
 DECAPx10_ASAP7_75t_R FILLER_17_167 ();
 DECAPx6_ASAP7_75t_R FILLER_17_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_203 ();
 FILLER_ASAP7_75t_R FILLER_17_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_238 ();
 FILLER_ASAP7_75t_R FILLER_17_262 ();
 DECAPx2_ASAP7_75t_R FILLER_17_270 ();
 FILLER_ASAP7_75t_R FILLER_18_2 ();
 DECAPx2_ASAP7_75t_R FILLER_18_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_26 ();
 DECAPx2_ASAP7_75t_R FILLER_18_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_39 ();
 DECAPx2_ASAP7_75t_R FILLER_18_57 ();
 FILLER_ASAP7_75t_R FILLER_18_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_65 ();
 DECAPx4_ASAP7_75t_R FILLER_18_87 ();
 FILLER_ASAP7_75t_R FILLER_18_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_132 ();
 DECAPx6_ASAP7_75t_R FILLER_18_143 ();
 FILLER_ASAP7_75t_R FILLER_18_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_159 ();
 DECAPx10_ASAP7_75t_R FILLER_18_166 ();
 DECAPx4_ASAP7_75t_R FILLER_18_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_234 ();
 DECAPx6_ASAP7_75t_R FILLER_18_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_269 ();
 FILLER_ASAP7_75t_R FILLER_19_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_4 ();
 DECAPx1_ASAP7_75t_R FILLER_19_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_52 ();
 DECAPx2_ASAP7_75t_R FILLER_19_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_71 ();
 DECAPx4_ASAP7_75t_R FILLER_19_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_96 ();
 DECAPx1_ASAP7_75t_R FILLER_19_121 ();
 FILLER_ASAP7_75t_R FILLER_19_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_140 ();
 DECAPx10_ASAP7_75t_R FILLER_19_144 ();
 DECAPx10_ASAP7_75t_R FILLER_19_166 ();
 DECAPx4_ASAP7_75t_R FILLER_19_188 ();
 DECAPx2_ASAP7_75t_R FILLER_19_246 ();
 FILLER_ASAP7_75t_R FILLER_19_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_275 ();
 DECAPx2_ASAP7_75t_R FILLER_20_26 ();
 FILLER_ASAP7_75t_R FILLER_20_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_34 ();
 DECAPx2_ASAP7_75t_R FILLER_20_41 ();
 DECAPx10_ASAP7_75t_R FILLER_20_73 ();
 FILLER_ASAP7_75t_R FILLER_20_95 ();
 DECAPx2_ASAP7_75t_R FILLER_20_107 ();
 DECAPx1_ASAP7_75t_R FILLER_20_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_156 ();
 DECAPx10_ASAP7_75t_R FILLER_20_167 ();
 DECAPx2_ASAP7_75t_R FILLER_20_189 ();
 FILLER_ASAP7_75t_R FILLER_20_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_197 ();
 FILLER_ASAP7_75t_R FILLER_20_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_214 ();
 DECAPx6_ASAP7_75t_R FILLER_20_235 ();
 DECAPx2_ASAP7_75t_R FILLER_20_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_264 ();
 DECAPx1_ASAP7_75t_R FILLER_20_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_8 ();
 DECAPx2_ASAP7_75t_R FILLER_21_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_27 ();
 FILLER_ASAP7_75t_R FILLER_21_62 ();
 DECAPx6_ASAP7_75t_R FILLER_21_67 ();
 DECAPx1_ASAP7_75t_R FILLER_21_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_130 ();
 DECAPx10_ASAP7_75t_R FILLER_21_141 ();
 DECAPx6_ASAP7_75t_R FILLER_21_163 ();
 DECAPx2_ASAP7_75t_R FILLER_21_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_183 ();
 DECAPx1_ASAP7_75t_R FILLER_21_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_198 ();
 DECAPx1_ASAP7_75t_R FILLER_21_219 ();
 DECAPx4_ASAP7_75t_R FILLER_21_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_253 ();
 DECAPx2_ASAP7_75t_R FILLER_21_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_14 ();
 DECAPx1_ASAP7_75t_R FILLER_22_50 ();
 DECAPx2_ASAP7_75t_R FILLER_22_64 ();
 FILLER_ASAP7_75t_R FILLER_22_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_72 ();
 DECAPx4_ASAP7_75t_R FILLER_22_97 ();
 FILLER_ASAP7_75t_R FILLER_22_107 ();
 DECAPx2_ASAP7_75t_R FILLER_22_115 ();
 FILLER_ASAP7_75t_R FILLER_22_121 ();
 DECAPx10_ASAP7_75t_R FILLER_22_157 ();
 DECAPx10_ASAP7_75t_R FILLER_22_179 ();
 DECAPx1_ASAP7_75t_R FILLER_22_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_205 ();
 DECAPx10_ASAP7_75t_R FILLER_22_212 ();
 DECAPx4_ASAP7_75t_R FILLER_22_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_244 ();
 DECAPx6_ASAP7_75t_R FILLER_22_248 ();
 FILLER_ASAP7_75t_R FILLER_22_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_40 ();
 DECAPx6_ASAP7_75t_R FILLER_23_47 ();
 DECAPx2_ASAP7_75t_R FILLER_23_61 ();
 DECAPx1_ASAP7_75t_R FILLER_23_120 ();
 DECAPx10_ASAP7_75t_R FILLER_23_157 ();
 DECAPx6_ASAP7_75t_R FILLER_23_179 ();
 FILLER_ASAP7_75t_R FILLER_23_193 ();
 DECAPx10_ASAP7_75t_R FILLER_23_201 ();
 DECAPx4_ASAP7_75t_R FILLER_23_223 ();
 FILLER_ASAP7_75t_R FILLER_23_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_235 ();
 DECAPx1_ASAP7_75t_R FILLER_23_248 ();
 FILLER_ASAP7_75t_R FILLER_23_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_260 ();
 DECAPx2_ASAP7_75t_R FILLER_23_267 ();
 FILLER_ASAP7_75t_R FILLER_23_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_275 ();
 DECAPx6_ASAP7_75t_R FILLER_24_8 ();
 DECAPx2_ASAP7_75t_R FILLER_24_48 ();
 FILLER_ASAP7_75t_R FILLER_24_54 ();
 DECAPx6_ASAP7_75t_R FILLER_24_114 ();
 DECAPx2_ASAP7_75t_R FILLER_24_128 ();
 DECAPx10_ASAP7_75t_R FILLER_24_144 ();
 DECAPx10_ASAP7_75t_R FILLER_24_166 ();
 DECAPx4_ASAP7_75t_R FILLER_24_188 ();
 FILLER_ASAP7_75t_R FILLER_24_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_213 ();
 DECAPx6_ASAP7_75t_R FILLER_24_234 ();
 DECAPx2_ASAP7_75t_R FILLER_24_248 ();
 DECAPx1_ASAP7_75t_R FILLER_24_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_2 ();
 DECAPx2_ASAP7_75t_R FILLER_25_26 ();
 FILLER_ASAP7_75t_R FILLER_25_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_77 ();
 DECAPx10_ASAP7_75t_R FILLER_25_86 ();
 DECAPx10_ASAP7_75t_R FILLER_25_108 ();
 DECAPx6_ASAP7_75t_R FILLER_25_140 ();
 FILLER_ASAP7_75t_R FILLER_25_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_156 ();
 DECAPx4_ASAP7_75t_R FILLER_25_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_177 ();
 DECAPx2_ASAP7_75t_R FILLER_25_188 ();
 DECAPx1_ASAP7_75t_R FILLER_25_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_14 ();
 DECAPx2_ASAP7_75t_R FILLER_26_49 ();
 FILLER_ASAP7_75t_R FILLER_26_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_57 ();
 DECAPx10_ASAP7_75t_R FILLER_26_64 ();
 DECAPx10_ASAP7_75t_R FILLER_26_86 ();
 DECAPx6_ASAP7_75t_R FILLER_26_108 ();
 DECAPx1_ASAP7_75t_R FILLER_26_122 ();
 DECAPx10_ASAP7_75t_R FILLER_26_133 ();
 DECAPx10_ASAP7_75t_R FILLER_26_155 ();
 FILLER_ASAP7_75t_R FILLER_26_177 ();
 DECAPx6_ASAP7_75t_R FILLER_26_195 ();
 FILLER_ASAP7_75t_R FILLER_26_209 ();
 DECAPx2_ASAP7_75t_R FILLER_26_220 ();
 FILLER_ASAP7_75t_R FILLER_26_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_228 ();
 DECAPx2_ASAP7_75t_R FILLER_26_232 ();
 FILLER_ASAP7_75t_R FILLER_26_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_240 ();
 DECAPx4_ASAP7_75t_R FILLER_26_247 ();
 FILLER_ASAP7_75t_R FILLER_26_257 ();
 DECAPx1_ASAP7_75t_R FILLER_26_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_269 ();
 FILLER_ASAP7_75t_R FILLER_27_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_43 ();
 DECAPx2_ASAP7_75t_R FILLER_27_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_58 ();
 DECAPx6_ASAP7_75t_R FILLER_27_65 ();
 FILLER_ASAP7_75t_R FILLER_27_79 ();
 DECAPx2_ASAP7_75t_R FILLER_27_110 ();
 FILLER_ASAP7_75t_R FILLER_27_116 ();
 DECAPx4_ASAP7_75t_R FILLER_27_138 ();
 FILLER_ASAP7_75t_R FILLER_27_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_150 ();
 DECAPx6_ASAP7_75t_R FILLER_27_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_204 ();
 DECAPx1_ASAP7_75t_R FILLER_27_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_269 ();
 FILLER_ASAP7_75t_R FILLER_28_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_16 ();
 DECAPx4_ASAP7_75t_R FILLER_28_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_96 ();
 DECAPx1_ASAP7_75t_R FILLER_28_107 ();
 DECAPx6_ASAP7_75t_R FILLER_28_117 ();
 DECAPx2_ASAP7_75t_R FILLER_28_151 ();
 FILLER_ASAP7_75t_R FILLER_28_157 ();
 DECAPx4_ASAP7_75t_R FILLER_28_169 ();
 FILLER_ASAP7_75t_R FILLER_28_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_181 ();
 DECAPx2_ASAP7_75t_R FILLER_28_192 ();
 FILLER_ASAP7_75t_R FILLER_28_198 ();
 DECAPx10_ASAP7_75t_R FILLER_28_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_269 ();
 DECAPx2_ASAP7_75t_R FILLER_29_2 ();
 FILLER_ASAP7_75t_R FILLER_29_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_28 ();
 DECAPx1_ASAP7_75t_R FILLER_29_36 ();
 FILLER_ASAP7_75t_R FILLER_29_50 ();
 FILLER_ASAP7_75t_R FILLER_29_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_62 ();
 FILLER_ASAP7_75t_R FILLER_29_103 ();
 FILLER_ASAP7_75t_R FILLER_29_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_137 ();
 DECAPx10_ASAP7_75t_R FILLER_29_148 ();
 DECAPx4_ASAP7_75t_R FILLER_29_170 ();
 FILLER_ASAP7_75t_R FILLER_29_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_182 ();
 DECAPx4_ASAP7_75t_R FILLER_29_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_205 ();
 DECAPx6_ASAP7_75t_R FILLER_29_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_243 ();
 DECAPx2_ASAP7_75t_R FILLER_29_250 ();
 FILLER_ASAP7_75t_R FILLER_29_256 ();
 FILLER_ASAP7_75t_R FILLER_29_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_14 ();
 DECAPx2_ASAP7_75t_R FILLER_30_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_27 ();
 DECAPx2_ASAP7_75t_R FILLER_30_40 ();
 DECAPx6_ASAP7_75t_R FILLER_30_54 ();
 DECAPx2_ASAP7_75t_R FILLER_30_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_74 ();
 FILLER_ASAP7_75t_R FILLER_30_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_94 ();
 FILLER_ASAP7_75t_R FILLER_30_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_123 ();
 DECAPx10_ASAP7_75t_R FILLER_30_134 ();
 DECAPx2_ASAP7_75t_R FILLER_30_156 ();
 DECAPx2_ASAP7_75t_R FILLER_30_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_191 ();
 DECAPx6_ASAP7_75t_R FILLER_30_210 ();
 FILLER_ASAP7_75t_R FILLER_30_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_226 ();
 DECAPx2_ASAP7_75t_R FILLER_30_247 ();
 FILLER_ASAP7_75t_R FILLER_30_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_267 ();
 FILLER_ASAP7_75t_R FILLER_30_274 ();
 FILLER_ASAP7_75t_R FILLER_31_2 ();
 FILLER_ASAP7_75t_R FILLER_31_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_38 ();
 FILLER_ASAP7_75t_R FILLER_31_46 ();
 DECAPx1_ASAP7_75t_R FILLER_31_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_95 ();
 DECAPx6_ASAP7_75t_R FILLER_31_106 ();
 FILLER_ASAP7_75t_R FILLER_31_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_122 ();
 DECAPx10_ASAP7_75t_R FILLER_31_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_155 ();
 DECAPx1_ASAP7_75t_R FILLER_31_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_166 ();
 DECAPx4_ASAP7_75t_R FILLER_31_174 ();
 FILLER_ASAP7_75t_R FILLER_31_184 ();
 DECAPx10_ASAP7_75t_R FILLER_31_202 ();
 DECAPx10_ASAP7_75t_R FILLER_31_224 ();
 DECAPx2_ASAP7_75t_R FILLER_31_246 ();
 FILLER_ASAP7_75t_R FILLER_31_252 ();
 FILLER_ASAP7_75t_R FILLER_31_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_275 ();
 DECAPx2_ASAP7_75t_R FILLER_32_54 ();
 FILLER_ASAP7_75t_R FILLER_32_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_62 ();
 DECAPx6_ASAP7_75t_R FILLER_32_66 ();
 DECAPx2_ASAP7_75t_R FILLER_32_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_86 ();
 DECAPx4_ASAP7_75t_R FILLER_32_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_117 ();
 DECAPx2_ASAP7_75t_R FILLER_32_128 ();
 FILLER_ASAP7_75t_R FILLER_32_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_136 ();
 FILLER_ASAP7_75t_R FILLER_32_157 ();
 FILLER_ASAP7_75t_R FILLER_32_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_181 ();
 FILLER_ASAP7_75t_R FILLER_32_185 ();
 FILLER_ASAP7_75t_R FILLER_32_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_217 ();
 DECAPx4_ASAP7_75t_R FILLER_32_238 ();
 DECAPx4_ASAP7_75t_R FILLER_32_251 ();
 FILLER_ASAP7_75t_R FILLER_32_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_263 ();
 FILLER_ASAP7_75t_R FILLER_33_2 ();
 FILLER_ASAP7_75t_R FILLER_33_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_38 ();
 FILLER_ASAP7_75t_R FILLER_33_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_50 ();
 DECAPx6_ASAP7_75t_R FILLER_33_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_91 ();
 DECAPx6_ASAP7_75t_R FILLER_33_98 ();
 DECAPx2_ASAP7_75t_R FILLER_33_112 ();
 DECAPx10_ASAP7_75t_R FILLER_33_128 ();
 FILLER_ASAP7_75t_R FILLER_33_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_159 ();
 FILLER_ASAP7_75t_R FILLER_33_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_199 ();
 DECAPx4_ASAP7_75t_R FILLER_33_214 ();
 FILLER_ASAP7_75t_R FILLER_33_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_246 ();
 DECAPx1_ASAP7_75t_R FILLER_33_253 ();
 DECAPx1_ASAP7_75t_R FILLER_33_266 ();
 DECAPx1_ASAP7_75t_R FILLER_34_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_6 ();
 DECAPx2_ASAP7_75t_R FILLER_34_25 ();
 FILLER_ASAP7_75t_R FILLER_34_44 ();
 DECAPx4_ASAP7_75t_R FILLER_34_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_83 ();
 DECAPx1_ASAP7_75t_R FILLER_34_98 ();
 DECAPx10_ASAP7_75t_R FILLER_34_118 ();
 DECAPx6_ASAP7_75t_R FILLER_34_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_154 ();
 DECAPx4_ASAP7_75t_R FILLER_34_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_184 ();
 DECAPx10_ASAP7_75t_R FILLER_34_191 ();
 DECAPx10_ASAP7_75t_R FILLER_34_213 ();
 DECAPx10_ASAP7_75t_R FILLER_34_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_257 ();
 DECAPx2_ASAP7_75t_R FILLER_34_270 ();
 DECAPx2_ASAP7_75t_R FILLER_35_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_49 ();
 DECAPx2_ASAP7_75t_R FILLER_35_78 ();
 DECAPx1_ASAP7_75t_R FILLER_35_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_112 ();
 DECAPx1_ASAP7_75t_R FILLER_35_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_130 ();
 DECAPx10_ASAP7_75t_R FILLER_35_151 ();
 FILLER_ASAP7_75t_R FILLER_35_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_175 ();
 DECAPx2_ASAP7_75t_R FILLER_35_212 ();
 FILLER_ASAP7_75t_R FILLER_35_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_220 ();
 DECAPx1_ASAP7_75t_R FILLER_35_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_255 ();
 DECAPx1_ASAP7_75t_R FILLER_35_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_275 ();
 FILLER_ASAP7_75t_R FILLER_36_2 ();
 DECAPx1_ASAP7_75t_R FILLER_36_24 ();
 DECAPx6_ASAP7_75t_R FILLER_36_41 ();
 DECAPx1_ASAP7_75t_R FILLER_36_55 ();
 DECAPx4_ASAP7_75t_R FILLER_36_64 ();
 DECAPx10_ASAP7_75t_R FILLER_36_77 ();
 DECAPx1_ASAP7_75t_R FILLER_36_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_124 ();
 DECAPx2_ASAP7_75t_R FILLER_36_131 ();
 FILLER_ASAP7_75t_R FILLER_36_140 ();
 DECAPx6_ASAP7_75t_R FILLER_36_145 ();
 DECAPx2_ASAP7_75t_R FILLER_36_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_165 ();
 FILLER_ASAP7_75t_R FILLER_36_215 ();
 FILLER_ASAP7_75t_R FILLER_36_220 ();
 DECAPx2_ASAP7_75t_R FILLER_36_228 ();
 DECAPx1_ASAP7_75t_R FILLER_36_254 ();
 DECAPx1_ASAP7_75t_R FILLER_36_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_14 ();
 FILLER_ASAP7_75t_R FILLER_37_21 ();
 DECAPx10_ASAP7_75t_R FILLER_37_46 ();
 DECAPx2_ASAP7_75t_R FILLER_37_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_74 ();
 DECAPx6_ASAP7_75t_R FILLER_37_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_95 ();
 DECAPx6_ASAP7_75t_R FILLER_37_133 ();
 FILLER_ASAP7_75t_R FILLER_37_147 ();
 DECAPx1_ASAP7_75t_R FILLER_37_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_159 ();
 FILLER_ASAP7_75t_R FILLER_37_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_190 ();
 DECAPx2_ASAP7_75t_R FILLER_37_262 ();
 FILLER_ASAP7_75t_R FILLER_37_268 ();
 DECAPx2_ASAP7_75t_R FILLER_38_14 ();
 FILLER_ASAP7_75t_R FILLER_38_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_22 ();
 DECAPx4_ASAP7_75t_R FILLER_38_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_39 ();
 DECAPx2_ASAP7_75t_R FILLER_38_43 ();
 DECAPx6_ASAP7_75t_R FILLER_38_55 ();
 DECAPx1_ASAP7_75t_R FILLER_38_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_73 ();
 FILLER_ASAP7_75t_R FILLER_38_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_96 ();
 DECAPx4_ASAP7_75t_R FILLER_38_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_121 ();
 DECAPx6_ASAP7_75t_R FILLER_38_145 ();
 FILLER_ASAP7_75t_R FILLER_38_159 ();
 FILLER_ASAP7_75t_R FILLER_38_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_180 ();
 DECAPx1_ASAP7_75t_R FILLER_38_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_217 ();
 DECAPx2_ASAP7_75t_R FILLER_38_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_244 ();
 FILLER_ASAP7_75t_R FILLER_38_251 ();
 DECAPx6_ASAP7_75t_R FILLER_38_256 ();
 DECAPx2_ASAP7_75t_R FILLER_38_270 ();
 DECAPx6_ASAP7_75t_R FILLER_39_8 ();
 FILLER_ASAP7_75t_R FILLER_39_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_24 ();
 FILLER_ASAP7_75t_R FILLER_39_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_33 ();
 DECAPx6_ASAP7_75t_R FILLER_39_70 ();
 FILLER_ASAP7_75t_R FILLER_39_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_86 ();
 DECAPx10_ASAP7_75t_R FILLER_39_98 ();
 FILLER_ASAP7_75t_R FILLER_39_120 ();
 DECAPx1_ASAP7_75t_R FILLER_39_128 ();
 DECAPx2_ASAP7_75t_R FILLER_39_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_141 ();
 FILLER_ASAP7_75t_R FILLER_39_168 ();
 DECAPx1_ASAP7_75t_R FILLER_39_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_205 ();
 FILLER_ASAP7_75t_R FILLER_39_238 ();
 DECAPx2_ASAP7_75t_R FILLER_39_249 ();
 FILLER_ASAP7_75t_R FILLER_39_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_257 ();
 DECAPx1_ASAP7_75t_R FILLER_40_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_42 ();
 FILLER_ASAP7_75t_R FILLER_40_53 ();
 FILLER_ASAP7_75t_R FILLER_40_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_99 ();
 DECAPx10_ASAP7_75t_R FILLER_40_103 ();
 DECAPx10_ASAP7_75t_R FILLER_40_125 ();
 DECAPx10_ASAP7_75t_R FILLER_40_147 ();
 FILLER_ASAP7_75t_R FILLER_40_169 ();
 DECAPx1_ASAP7_75t_R FILLER_40_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_191 ();
 DECAPx10_ASAP7_75t_R FILLER_40_223 ();
 DECAPx10_ASAP7_75t_R FILLER_40_245 ();
 FILLER_ASAP7_75t_R FILLER_40_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_8 ();
 FILLER_ASAP7_75t_R FILLER_41_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_17 ();
 DECAPx1_ASAP7_75t_R FILLER_41_41 ();
 DECAPx6_ASAP7_75t_R FILLER_41_105 ();
 DECAPx1_ASAP7_75t_R FILLER_41_119 ();
 FILLER_ASAP7_75t_R FILLER_41_129 ();
 DECAPx6_ASAP7_75t_R FILLER_41_151 ();
 FILLER_ASAP7_75t_R FILLER_41_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_190 ();
 DECAPx2_ASAP7_75t_R FILLER_41_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_237 ();
 DECAPx2_ASAP7_75t_R FILLER_41_244 ();
 DECAPx6_ASAP7_75t_R FILLER_41_256 ();
 DECAPx2_ASAP7_75t_R FILLER_41_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_21 ();
 DECAPx2_ASAP7_75t_R FILLER_42_28 ();
 FILLER_ASAP7_75t_R FILLER_42_34 ();
 DECAPx1_ASAP7_75t_R FILLER_42_39 ();
 FILLER_ASAP7_75t_R FILLER_42_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_59 ();
 FILLER_ASAP7_75t_R FILLER_42_66 ();
 DECAPx1_ASAP7_75t_R FILLER_42_112 ();
 DECAPx2_ASAP7_75t_R FILLER_42_136 ();
 FILLER_ASAP7_75t_R FILLER_42_142 ();
 DECAPx2_ASAP7_75t_R FILLER_42_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_153 ();
 FILLER_ASAP7_75t_R FILLER_42_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_159 ();
 DECAPx4_ASAP7_75t_R FILLER_42_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_184 ();
 FILLER_ASAP7_75t_R FILLER_42_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_215 ();
 DECAPx4_ASAP7_75t_R FILLER_42_236 ();
 FILLER_ASAP7_75t_R FILLER_42_246 ();
 DECAPx4_ASAP7_75t_R FILLER_42_251 ();
 FILLER_ASAP7_75t_R FILLER_42_261 ();
 DECAPx2_ASAP7_75t_R FILLER_42_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_275 ();
 DECAPx6_ASAP7_75t_R FILLER_43_2 ();
 DECAPx1_ASAP7_75t_R FILLER_43_16 ();
 DECAPx6_ASAP7_75t_R FILLER_43_26 ();
 DECAPx1_ASAP7_75t_R FILLER_43_40 ();
 DECAPx2_ASAP7_75t_R FILLER_43_51 ();
 FILLER_ASAP7_75t_R FILLER_43_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_59 ();
 DECAPx1_ASAP7_75t_R FILLER_43_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_92 ();
 DECAPx1_ASAP7_75t_R FILLER_43_111 ();
 DECAPx2_ASAP7_75t_R FILLER_43_141 ();
 FILLER_ASAP7_75t_R FILLER_43_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_149 ();
 DECAPx2_ASAP7_75t_R FILLER_43_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_159 ();
 DECAPx6_ASAP7_75t_R FILLER_43_167 ();
 DECAPx1_ASAP7_75t_R FILLER_43_181 ();
 FILLER_ASAP7_75t_R FILLER_43_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_201 ();
 FILLER_ASAP7_75t_R FILLER_43_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_216 ();
 DECAPx6_ASAP7_75t_R FILLER_43_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_251 ();
 DECAPx2_ASAP7_75t_R FILLER_43_264 ();
 FILLER_ASAP7_75t_R FILLER_44_2 ();
 DECAPx2_ASAP7_75t_R FILLER_44_10 ();
 DECAPx4_ASAP7_75t_R FILLER_44_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_32 ();
 FILLER_ASAP7_75t_R FILLER_44_46 ();
 FILLER_ASAP7_75t_R FILLER_44_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_70 ();
 DECAPx2_ASAP7_75t_R FILLER_44_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_80 ();
 FILLER_ASAP7_75t_R FILLER_44_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_102 ();
 DECAPx10_ASAP7_75t_R FILLER_44_110 ();
 DECAPx1_ASAP7_75t_R FILLER_44_132 ();
 DECAPx1_ASAP7_75t_R FILLER_44_169 ();
 FILLER_ASAP7_75t_R FILLER_44_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_200 ();
 DECAPx2_ASAP7_75t_R FILLER_44_220 ();
 DECAPx4_ASAP7_75t_R FILLER_44_246 ();
 FILLER_ASAP7_75t_R FILLER_44_256 ();
 DECAPx2_ASAP7_75t_R FILLER_44_264 ();
 FILLER_ASAP7_75t_R FILLER_45_2 ();
 DECAPx6_ASAP7_75t_R FILLER_45_10 ();
 DECAPx1_ASAP7_75t_R FILLER_45_24 ();
 DECAPx2_ASAP7_75t_R FILLER_45_34 ();
 DECAPx2_ASAP7_75t_R FILLER_45_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_87 ();
 FILLER_ASAP7_75t_R FILLER_45_94 ();
 FILLER_ASAP7_75t_R FILLER_45_103 ();
 FILLER_ASAP7_75t_R FILLER_45_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_136 ();
 DECAPx4_ASAP7_75t_R FILLER_45_154 ();
 DECAPx1_ASAP7_75t_R FILLER_45_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_196 ();
 FILLER_ASAP7_75t_R FILLER_45_211 ();
 DECAPx6_ASAP7_75t_R FILLER_45_233 ();
 FILLER_ASAP7_75t_R FILLER_45_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_249 ();
 DECAPx4_ASAP7_75t_R FILLER_45_256 ();
 FILLER_ASAP7_75t_R FILLER_45_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_275 ();
 DECAPx4_ASAP7_75t_R FILLER_46_2 ();
 FILLER_ASAP7_75t_R FILLER_46_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_14 ();
 DECAPx6_ASAP7_75t_R FILLER_46_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_35 ();
 DECAPx6_ASAP7_75t_R FILLER_46_48 ();
 FILLER_ASAP7_75t_R FILLER_46_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_64 ();
 DECAPx6_ASAP7_75t_R FILLER_46_74 ();
 FILLER_ASAP7_75t_R FILLER_46_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_90 ();
 DECAPx1_ASAP7_75t_R FILLER_46_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_148 ();
 DECAPx6_ASAP7_75t_R FILLER_46_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_171 ();
 FILLER_ASAP7_75t_R FILLER_46_210 ();
 DECAPx4_ASAP7_75t_R FILLER_46_232 ();
 FILLER_ASAP7_75t_R FILLER_46_242 ();
 DECAPx1_ASAP7_75t_R FILLER_46_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_251 ();
 DECAPx6_ASAP7_75t_R FILLER_46_258 ();
 DECAPx1_ASAP7_75t_R FILLER_46_272 ();
 DECAPx10_ASAP7_75t_R FILLER_47_2 ();
 DECAPx4_ASAP7_75t_R FILLER_47_24 ();
 FILLER_ASAP7_75t_R FILLER_47_34 ();
 FILLER_ASAP7_75t_R FILLER_47_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_87 ();
 DECAPx1_ASAP7_75t_R FILLER_47_91 ();
 DECAPx6_ASAP7_75t_R FILLER_47_107 ();
 DECAPx1_ASAP7_75t_R FILLER_47_121 ();
 DECAPx2_ASAP7_75t_R FILLER_47_131 ();
 FILLER_ASAP7_75t_R FILLER_47_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_139 ();
 FILLER_ASAP7_75t_R FILLER_47_149 ();
 FILLER_ASAP7_75t_R FILLER_47_171 ();
 FILLER_ASAP7_75t_R FILLER_47_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_188 ();
 DECAPx10_ASAP7_75t_R FILLER_47_197 ();
 DECAPx10_ASAP7_75t_R FILLER_47_219 ();
 DECAPx10_ASAP7_75t_R FILLER_47_241 ();
 DECAPx4_ASAP7_75t_R FILLER_47_263 ();
 FILLER_ASAP7_75t_R FILLER_47_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_275 ();
 DECAPx10_ASAP7_75t_R FILLER_48_2 ();
 DECAPx10_ASAP7_75t_R FILLER_48_24 ();
 DECAPx10_ASAP7_75t_R FILLER_48_46 ();
 DECAPx10_ASAP7_75t_R FILLER_48_68 ();
 DECAPx1_ASAP7_75t_R FILLER_48_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_100 ();
 DECAPx1_ASAP7_75t_R FILLER_48_124 ();
 DECAPx10_ASAP7_75t_R FILLER_48_131 ();
 DECAPx10_ASAP7_75t_R FILLER_48_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_175 ();
 DECAPx10_ASAP7_75t_R FILLER_48_188 ();
 DECAPx10_ASAP7_75t_R FILLER_48_210 ();
 DECAPx10_ASAP7_75t_R FILLER_48_232 ();
 DECAPx10_ASAP7_75t_R FILLER_48_254 ();
 DECAPx10_ASAP7_75t_R FILLER_49_2 ();
 DECAPx10_ASAP7_75t_R FILLER_49_24 ();
 DECAPx10_ASAP7_75t_R FILLER_49_46 ();
 DECAPx10_ASAP7_75t_R FILLER_49_68 ();
 FILLER_ASAP7_75t_R FILLER_49_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_92 ();
 DECAPx2_ASAP7_75t_R FILLER_49_113 ();
 FILLER_ASAP7_75t_R FILLER_49_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_121 ();
 DECAPx2_ASAP7_75t_R FILLER_49_125 ();
 FILLER_ASAP7_75t_R FILLER_49_154 ();
 DECAPx4_ASAP7_75t_R FILLER_49_162 ();
 FILLER_ASAP7_75t_R FILLER_49_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_174 ();
 DECAPx6_ASAP7_75t_R FILLER_49_221 ();
 DECAPx10_ASAP7_75t_R FILLER_49_238 ();
 DECAPx6_ASAP7_75t_R FILLER_49_260 ();
 FILLER_ASAP7_75t_R FILLER_49_274 ();
 DECAPx10_ASAP7_75t_R FILLER_50_2 ();
 DECAPx10_ASAP7_75t_R FILLER_50_24 ();
 DECAPx10_ASAP7_75t_R FILLER_50_46 ();
 DECAPx10_ASAP7_75t_R FILLER_50_68 ();
 DECAPx4_ASAP7_75t_R FILLER_50_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_100 ();
 DECAPx6_ASAP7_75t_R FILLER_50_107 ();
 FILLER_ASAP7_75t_R FILLER_50_121 ();
 DECAPx10_ASAP7_75t_R FILLER_50_126 ();
 DECAPx10_ASAP7_75t_R FILLER_50_148 ();
 FILLER_ASAP7_75t_R FILLER_50_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_172 ();
 FILLER_ASAP7_75t_R FILLER_50_193 ();
 DECAPx4_ASAP7_75t_R FILLER_50_198 ();
 FILLER_ASAP7_75t_R FILLER_50_231 ();
 DECAPx10_ASAP7_75t_R FILLER_50_236 ();
 DECAPx6_ASAP7_75t_R FILLER_50_258 ();
 DECAPx1_ASAP7_75t_R FILLER_50_272 ();
 DECAPx10_ASAP7_75t_R FILLER_51_2 ();
 DECAPx10_ASAP7_75t_R FILLER_51_24 ();
 DECAPx10_ASAP7_75t_R FILLER_51_46 ();
 DECAPx4_ASAP7_75t_R FILLER_51_68 ();
 DECAPx4_ASAP7_75t_R FILLER_51_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_94 ();
 DECAPx2_ASAP7_75t_R FILLER_51_113 ();
 DECAPx6_ASAP7_75t_R FILLER_51_137 ();
 DECAPx1_ASAP7_75t_R FILLER_51_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_155 ();
 DECAPx6_ASAP7_75t_R FILLER_51_196 ();
 DECAPx2_ASAP7_75t_R FILLER_51_210 ();
 DECAPx2_ASAP7_75t_R FILLER_51_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_242 ();
 DECAPx10_ASAP7_75t_R FILLER_51_246 ();
 DECAPx2_ASAP7_75t_R FILLER_51_268 ();
 FILLER_ASAP7_75t_R FILLER_51_274 ();
 DECAPx10_ASAP7_75t_R FILLER_52_2 ();
 DECAPx10_ASAP7_75t_R FILLER_52_24 ();
 FILLER_ASAP7_75t_R FILLER_52_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_48 ();
 DECAPx4_ASAP7_75t_R FILLER_52_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_72 ();
 DECAPx2_ASAP7_75t_R FILLER_52_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_98 ();
 DECAPx1_ASAP7_75t_R FILLER_52_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_109 ();
 DECAPx4_ASAP7_75t_R FILLER_52_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_168 ();
 DECAPx6_ASAP7_75t_R FILLER_52_178 ();
 DECAPx2_ASAP7_75t_R FILLER_52_192 ();
 DECAPx10_ASAP7_75t_R FILLER_52_204 ();
 DECAPx10_ASAP7_75t_R FILLER_52_226 ();
 DECAPx10_ASAP7_75t_R FILLER_52_248 ();
 DECAPx2_ASAP7_75t_R FILLER_52_270 ();
 DECAPx10_ASAP7_75t_R FILLER_53_2 ();
 DECAPx10_ASAP7_75t_R FILLER_53_24 ();
 DECAPx4_ASAP7_75t_R FILLER_53_46 ();
 FILLER_ASAP7_75t_R FILLER_53_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_88 ();
 DECAPx1_ASAP7_75t_R FILLER_53_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_111 ();
 DECAPx2_ASAP7_75t_R FILLER_53_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_124 ();
 FILLER_ASAP7_75t_R FILLER_53_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_181 ();
 DECAPx2_ASAP7_75t_R FILLER_53_200 ();
 FILLER_ASAP7_75t_R FILLER_53_206 ();
 DECAPx10_ASAP7_75t_R FILLER_53_214 ();
 DECAPx10_ASAP7_75t_R FILLER_53_236 ();
 DECAPx6_ASAP7_75t_R FILLER_53_258 ();
 DECAPx1_ASAP7_75t_R FILLER_53_272 ();
 DECAPx10_ASAP7_75t_R FILLER_54_2 ();
 DECAPx6_ASAP7_75t_R FILLER_54_24 ();
 FILLER_ASAP7_75t_R FILLER_54_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_40 ();
 FILLER_ASAP7_75t_R FILLER_54_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_68 ();
 DECAPx2_ASAP7_75t_R FILLER_54_87 ();
 FILLER_ASAP7_75t_R FILLER_54_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_206 ();
 DECAPx10_ASAP7_75t_R FILLER_54_219 ();
 DECAPx10_ASAP7_75t_R FILLER_54_241 ();
 DECAPx4_ASAP7_75t_R FILLER_54_263 ();
 FILLER_ASAP7_75t_R FILLER_54_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_275 ();
endmodule
