module bft (ce,
    clk,
    done_all,
    rst,
    cmd,
    in,
    out);
 input ce;
 input clk;
 output done_all;
 input rst;
 input [5:0] cmd;
 input [39:0] in;
 output [1279:0] out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire clknet_leaf_0_clk;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire \peo[0][0] ;
 wire \peo[0][32] ;
 wire \peo[0][33] ;
 wire \peo[0][34] ;
 wire \peo[0][35] ;
 wire \peo[0][36] ;
 wire \peo[0][39] ;
 wire \peo[10][0] ;
 wire \peo[10][11] ;
 wire \peo[10][32] ;
 wire \peo[10][33] ;
 wire \peo[10][34] ;
 wire \peo[10][35] ;
 wire \peo[10][36] ;
 wire \peo[10][39] ;
 wire \peo[11][0] ;
 wire \peo[11][10] ;
 wire \peo[12][0] ;
 wire \peo[12][12] ;
 wire \peo[12][32] ;
 wire \peo[12][33] ;
 wire \peo[12][34] ;
 wire \peo[12][35] ;
 wire \peo[12][36] ;
 wire \peo[12][39] ;
 wire \peo[13][0] ;
 wire \peo[13][10] ;
 wire \peo[14][0] ;
 wire \peo[14][11] ;
 wire \peo[14][32] ;
 wire \peo[14][33] ;
 wire \peo[14][34] ;
 wire \peo[14][35] ;
 wire \peo[14][36] ;
 wire \peo[14][39] ;
 wire \peo[15][0] ;
 wire \peo[15][10] ;
 wire \peo[16][0] ;
 wire \peo[16][14] ;
 wire \peo[16][32] ;
 wire \peo[16][33] ;
 wire \peo[16][34] ;
 wire \peo[16][35] ;
 wire \peo[16][36] ;
 wire \peo[16][39] ;
 wire \peo[17][0] ;
 wire \peo[17][10] ;
 wire \peo[18][0] ;
 wire \peo[18][11] ;
 wire \peo[18][32] ;
 wire \peo[18][33] ;
 wire \peo[18][34] ;
 wire \peo[18][35] ;
 wire \peo[18][36] ;
 wire \peo[18][39] ;
 wire \peo[19][0] ;
 wire \peo[19][10] ;
 wire \peo[19][32] ;
 wire \peo[19][33] ;
 wire \peo[19][34] ;
 wire \peo[19][35] ;
 wire \peo[19][36] ;
 wire \peo[19][39] ;
 wire \peo[1][0] ;
 wire \peo[1][10] ;
 wire \peo[1][32] ;
 wire \peo[20][0] ;
 wire \peo[20][12] ;
 wire \peo[20][32] ;
 wire \peo[20][33] ;
 wire \peo[20][34] ;
 wire \peo[20][35] ;
 wire \peo[20][36] ;
 wire \peo[20][39] ;
 wire \peo[21][0] ;
 wire \peo[21][10] ;
 wire \peo[21][32] ;
 wire \peo[22][0] ;
 wire \peo[22][11] ;
 wire \peo[22][32] ;
 wire \peo[22][33] ;
 wire \peo[22][34] ;
 wire \peo[22][35] ;
 wire \peo[22][36] ;
 wire \peo[22][39] ;
 wire \peo[23][0] ;
 wire \peo[23][10] ;
 wire \peo[23][32] ;
 wire \peo[24][0] ;
 wire \peo[24][13] ;
 wire \peo[24][32] ;
 wire \peo[24][33] ;
 wire \peo[24][34] ;
 wire \peo[24][35] ;
 wire \peo[24][36] ;
 wire \peo[24][39] ;
 wire \peo[25][0] ;
 wire \peo[25][10] ;
 wire \peo[25][32] ;
 wire \peo[26][0] ;
 wire \peo[26][11] ;
 wire \peo[26][32] ;
 wire \peo[26][33] ;
 wire \peo[26][34] ;
 wire \peo[26][35] ;
 wire \peo[26][36] ;
 wire \peo[26][39] ;
 wire \peo[27][0] ;
 wire \peo[27][10] ;
 wire \peo[27][32] ;
 wire \peo[28][0] ;
 wire \peo[28][12] ;
 wire \peo[28][32] ;
 wire \peo[28][33] ;
 wire \peo[28][34] ;
 wire \peo[28][35] ;
 wire \peo[28][36] ;
 wire \peo[28][39] ;
 wire \peo[29][0] ;
 wire \peo[29][10] ;
 wire \peo[29][32] ;
 wire \peo[2][0] ;
 wire \peo[2][11] ;
 wire \peo[2][32] ;
 wire \peo[2][33] ;
 wire \peo[2][34] ;
 wire \peo[2][35] ;
 wire \peo[2][36] ;
 wire \peo[2][39] ;
 wire \peo[30][0] ;
 wire \peo[30][11] ;
 wire \peo[30][32] ;
 wire \peo[30][33] ;
 wire \peo[30][34] ;
 wire \peo[30][35] ;
 wire \peo[30][36] ;
 wire \peo[30][39] ;
 wire \peo[31][0] ;
 wire \peo[31][10] ;
 wire \peo[31][32] ;
 wire \peo[3][0] ;
 wire \peo[4][0] ;
 wire \peo[4][12] ;
 wire \peo[4][32] ;
 wire \peo[4][33] ;
 wire \peo[4][34] ;
 wire \peo[4][35] ;
 wire \peo[4][36] ;
 wire \peo[4][39] ;
 wire \peo[5][0] ;
 wire \peo[5][10] ;
 wire \peo[6][0] ;
 wire \peo[6][11] ;
 wire \peo[6][32] ;
 wire \peo[6][33] ;
 wire \peo[6][34] ;
 wire \peo[6][35] ;
 wire \peo[6][36] ;
 wire \peo[6][39] ;
 wire \peo[7][0] ;
 wire \peo[7][10] ;
 wire \peo[8][0] ;
 wire \peo[8][13] ;
 wire \peo[8][32] ;
 wire \peo[8][33] ;
 wire \peo[8][34] ;
 wire \peo[8][35] ;
 wire \peo[8][36] ;
 wire \peo[8][39] ;
 wire \peo[9][0] ;
 wire \peo[9][10] ;
 wire \xs[0].cli0.r[0] ;
 wire \xs[0].cli0.r[1] ;
 wire \xs[0].cli1.i[33] ;
 wire \xs[0].cli1.i[34] ;
 wire \xs[0].cli1.i[35] ;
 wire \xs[0].cli1.i[36] ;
 wire \xs[0].cli1.i[39] ;
 wire \xs[0].cli1.r[0] ;
 wire \xs[0].cli1.r[1] ;
 wire \xs[10].cli0.r[0] ;
 wire \xs[10].cli0.r[1] ;
 wire \xs[10].cli1.i[33] ;
 wire \xs[10].cli1.i[34] ;
 wire \xs[10].cli1.i[35] ;
 wire \xs[10].cli1.i[36] ;
 wire \xs[10].cli1.i[39] ;
 wire \xs[10].cli1.r[0] ;
 wire \xs[10].cli1.r[1] ;
 wire \xs[11].cli0.r[0] ;
 wire \xs[11].cli0.r[1] ;
 wire \xs[11].cli1.i[33] ;
 wire \xs[11].cli1.i[34] ;
 wire \xs[11].cli1.i[35] ;
 wire \xs[11].cli1.i[36] ;
 wire \xs[11].cli1.i[39] ;
 wire \xs[11].cli1.r[0] ;
 wire \xs[11].cli1.r[1] ;
 wire \xs[12].cli0.r[0] ;
 wire \xs[12].cli0.r[1] ;
 wire \xs[12].cli1.i[33] ;
 wire \xs[12].cli1.i[34] ;
 wire \xs[12].cli1.i[35] ;
 wire \xs[12].cli1.i[36] ;
 wire \xs[12].cli1.i[39] ;
 wire \xs[12].cli1.r[0] ;
 wire \xs[12].cli1.r[1] ;
 wire \xs[13].cli0.r[0] ;
 wire \xs[13].cli0.r[1] ;
 wire \xs[13].cli1.i[33] ;
 wire \xs[13].cli1.i[34] ;
 wire \xs[13].cli1.i[35] ;
 wire \xs[13].cli1.i[36] ;
 wire \xs[13].cli1.i[39] ;
 wire \xs[13].cli1.r[0] ;
 wire \xs[13].cli1.r[1] ;
 wire \xs[14].cli0.r[0] ;
 wire \xs[14].cli0.r[1] ;
 wire \xs[14].cli1.i[33] ;
 wire \xs[14].cli1.i[34] ;
 wire \xs[14].cli1.i[35] ;
 wire \xs[14].cli1.i[36] ;
 wire \xs[14].cli1.i[39] ;
 wire \xs[14].cli1.r[0] ;
 wire \xs[14].cli1.r[1] ;
 wire \xs[15].cli0.r[0] ;
 wire \xs[15].cli0.r[1] ;
 wire \xs[15].cli1.i[33] ;
 wire \xs[15].cli1.i[34] ;
 wire \xs[15].cli1.i[35] ;
 wire \xs[15].cli1.i[36] ;
 wire \xs[15].cli1.i[39] ;
 wire \xs[15].cli1.r[0] ;
 wire \xs[15].cli1.r[1] ;
 wire \xs[1].cli0.r[0] ;
 wire \xs[1].cli0.r[1] ;
 wire \xs[1].cli1.i[10] ;
 wire \xs[1].cli1.i[32] ;
 wire \xs[1].cli1.i[33] ;
 wire \xs[1].cli1.i[34] ;
 wire \xs[1].cli1.i[35] ;
 wire \xs[1].cli1.i[36] ;
 wire \xs[1].cli1.i[39] ;
 wire \xs[1].cli1.r[0] ;
 wire \xs[1].cli1.r[1] ;
 wire \xs[2].cli0.r[0] ;
 wire \xs[2].cli0.r[1] ;
 wire \xs[2].cli1.i[32] ;
 wire \xs[2].cli1.i[33] ;
 wire \xs[2].cli1.i[34] ;
 wire \xs[2].cli1.i[35] ;
 wire \xs[2].cli1.i[36] ;
 wire \xs[2].cli1.i[39] ;
 wire \xs[2].cli1.r[0] ;
 wire \xs[2].cli1.r[1] ;
 wire \xs[3].cli0.r[0] ;
 wire \xs[3].cli0.r[1] ;
 wire \xs[3].cli1.i[32] ;
 wire \xs[3].cli1.i[33] ;
 wire \xs[3].cli1.i[34] ;
 wire \xs[3].cli1.i[35] ;
 wire \xs[3].cli1.i[36] ;
 wire \xs[3].cli1.i[39] ;
 wire \xs[3].cli1.r[0] ;
 wire \xs[3].cli1.r[1] ;
 wire \xs[4].cli0.r[0] ;
 wire \xs[4].cli0.r[1] ;
 wire \xs[4].cli1.i[32] ;
 wire \xs[4].cli1.i[33] ;
 wire \xs[4].cli1.i[34] ;
 wire \xs[4].cli1.i[35] ;
 wire \xs[4].cli1.i[36] ;
 wire \xs[4].cli1.i[39] ;
 wire \xs[4].cli1.r[0] ;
 wire \xs[4].cli1.r[1] ;
 wire \xs[5].cli0.r[0] ;
 wire \xs[5].cli0.r[1] ;
 wire \xs[5].cli1.i[32] ;
 wire \xs[5].cli1.i[33] ;
 wire \xs[5].cli1.i[34] ;
 wire \xs[5].cli1.i[35] ;
 wire \xs[5].cli1.i[36] ;
 wire \xs[5].cli1.i[39] ;
 wire \xs[5].cli1.r[0] ;
 wire \xs[5].cli1.r[1] ;
 wire \xs[6].cli0.r[0] ;
 wire \xs[6].cli0.r[1] ;
 wire \xs[6].cli1.i[32] ;
 wire \xs[6].cli1.i[33] ;
 wire \xs[6].cli1.i[34] ;
 wire \xs[6].cli1.i[35] ;
 wire \xs[6].cli1.i[36] ;
 wire \xs[6].cli1.i[39] ;
 wire \xs[6].cli1.r[0] ;
 wire \xs[6].cli1.r[1] ;
 wire \xs[7].cli0.r[0] ;
 wire \xs[7].cli0.r[1] ;
 wire \xs[7].cli1.i[32] ;
 wire \xs[7].cli1.i[33] ;
 wire \xs[7].cli1.i[34] ;
 wire \xs[7].cli1.i[35] ;
 wire \xs[7].cli1.i[36] ;
 wire \xs[7].cli1.i[39] ;
 wire \xs[7].cli1.r[0] ;
 wire \xs[7].cli1.r[1] ;
 wire \xs[8].cli0.r[0] ;
 wire \xs[8].cli0.r[1] ;
 wire \xs[8].cli1.i[32] ;
 wire \xs[8].cli1.i[33] ;
 wire \xs[8].cli1.i[34] ;
 wire \xs[8].cli1.i[35] ;
 wire \xs[8].cli1.i[36] ;
 wire \xs[8].cli1.i[39] ;
 wire \xs[8].cli1.r[0] ;
 wire \xs[8].cli1.r[1] ;
 wire \xs[9].cli0.r[0] ;
 wire \xs[9].cli0.r[1] ;
 wire \xs[9].cli1.r[0] ;
 wire \xs[9].cli1.r[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;

 BUFx6f_ASAP7_75t_R _11642_ (.A(_00536_),
    .Y(_08525_));
 INVx2_ASAP7_75t_R _11643_ (.A(_08525_),
    .Y(\xs[5].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11644_ (.A(_00541_),
    .Y(\xs[5].cli1.i[32] ));
 INVx1_ASAP7_75t_R _11645_ (.A(_00540_),
    .Y(\xs[5].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11646_ (.A(_00539_),
    .Y(\xs[5].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11647_ (.A(_00537_),
    .Y(\xs[5].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11648_ (.A(_00538_),
    .Y(\xs[5].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11649_ (.A(_00575_),
    .Y(\peo[10][39] ));
 INVx1_ASAP7_75t_R _11650_ (.A(_00580_),
    .Y(\peo[10][32] ));
 INVx1_ASAP7_75t_R _11651_ (.A(_00579_),
    .Y(\peo[10][33] ));
 INVx1_ASAP7_75t_R _11652_ (.A(_00578_),
    .Y(\peo[10][34] ));
 INVx1_ASAP7_75t_R _11653_ (.A(_00576_),
    .Y(\peo[10][36] ));
 INVx1_ASAP7_75t_R _11654_ (.A(_00577_),
    .Y(\peo[10][35] ));
 INVx1_ASAP7_75t_R _11655_ (.A(_01687_),
    .Y(\peo[1][0] ));
 INVx1_ASAP7_75t_R _11656_ (.A(_01725_),
    .Y(\peo[0][0] ));
 INVx1_ASAP7_75t_R _11657_ (.A(_01685_),
    .Y(\peo[1][32] ));
 INVx1_ASAP7_75t_R _11658_ (.A(_01724_),
    .Y(\peo[0][32] ));
 INVx1_ASAP7_75t_R _11659_ (.A(_01684_),
    .Y(\xs[0].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11660_ (.A(_01723_),
    .Y(\peo[0][33] ));
 INVx1_ASAP7_75t_R _11661_ (.A(_01683_),
    .Y(\xs[0].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11662_ (.A(_01722_),
    .Y(\peo[0][34] ));
 INVx1_ASAP7_75t_R _11663_ (.A(_01682_),
    .Y(\xs[0].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11664_ (.A(_01721_),
    .Y(\peo[0][35] ));
 INVx1_ASAP7_75t_R _11665_ (.A(_01681_),
    .Y(\xs[0].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11666_ (.A(_01720_),
    .Y(\peo[0][36] ));
 INVx1_ASAP7_75t_R _11667_ (.A(_01583_),
    .Y(\peo[21][0] ));
 INVx1_ASAP7_75t_R _11668_ (.A(_01622_),
    .Y(\peo[20][0] ));
 INVx1_ASAP7_75t_R _11669_ (.A(_01581_),
    .Y(\peo[21][32] ));
 INVx1_ASAP7_75t_R _11670_ (.A(_01620_),
    .Y(\peo[20][32] ));
 INVx1_ASAP7_75t_R _11671_ (.A(_01580_),
    .Y(\xs[10].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11672_ (.A(_01619_),
    .Y(\peo[20][33] ));
 INVx1_ASAP7_75t_R _11673_ (.A(_01579_),
    .Y(\xs[10].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11674_ (.A(_01618_),
    .Y(\peo[20][34] ));
 INVx1_ASAP7_75t_R _11675_ (.A(_01578_),
    .Y(\xs[10].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11676_ (.A(_01617_),
    .Y(\peo[20][35] ));
 INVx1_ASAP7_75t_R _11677_ (.A(_01577_),
    .Y(\xs[10].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11678_ (.A(_01616_),
    .Y(\peo[20][36] ));
 INVx2_ASAP7_75t_R _11679_ (.A(_01479_),
    .Y(\peo[23][0] ));
 INVx1_ASAP7_75t_R _11680_ (.A(_01518_),
    .Y(\peo[22][0] ));
 INVx1_ASAP7_75t_R _11681_ (.A(_01477_),
    .Y(\peo[23][32] ));
 INVx1_ASAP7_75t_R _11682_ (.A(_01516_),
    .Y(\peo[22][32] ));
 INVx1_ASAP7_75t_R _11683_ (.A(_01476_),
    .Y(\xs[11].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11684_ (.A(_01515_),
    .Y(\peo[22][33] ));
 INVx1_ASAP7_75t_R _11685_ (.A(_01475_),
    .Y(\xs[11].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11686_ (.A(_01514_),
    .Y(\peo[22][34] ));
 INVx2_ASAP7_75t_R _11687_ (.A(_01474_),
    .Y(\xs[11].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11688_ (.A(_01513_),
    .Y(\peo[22][35] ));
 INVx1_ASAP7_75t_R _11689_ (.A(_01473_),
    .Y(\xs[11].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11690_ (.A(_01512_),
    .Y(\peo[22][36] ));
 INVx1_ASAP7_75t_R _11691_ (.A(_01375_),
    .Y(\peo[25][0] ));
 INVx1_ASAP7_75t_R _11692_ (.A(_01414_),
    .Y(\peo[24][0] ));
 INVx1_ASAP7_75t_R _11693_ (.A(_01373_),
    .Y(\peo[25][32] ));
 INVx1_ASAP7_75t_R _11694_ (.A(_01412_),
    .Y(\peo[24][32] ));
 INVx1_ASAP7_75t_R _11695_ (.A(_01372_),
    .Y(\xs[12].cli1.i[33] ));
 INVx2_ASAP7_75t_R _11696_ (.A(_01411_),
    .Y(\peo[24][33] ));
 INVx1_ASAP7_75t_R _11697_ (.A(_01371_),
    .Y(\xs[12].cli1.i[34] ));
 INVx2_ASAP7_75t_R _11698_ (.A(_01410_),
    .Y(\peo[24][34] ));
 INVx1_ASAP7_75t_R _11699_ (.A(_01370_),
    .Y(\xs[12].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11700_ (.A(_01409_),
    .Y(\peo[24][35] ));
 INVx1_ASAP7_75t_R _11701_ (.A(_01369_),
    .Y(\xs[12].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11702_ (.A(_01408_),
    .Y(\peo[24][36] ));
 INVx1_ASAP7_75t_R _11703_ (.A(_01310_),
    .Y(\peo[26][0] ));
 INVx1_ASAP7_75t_R _11704_ (.A(_01271_),
    .Y(\peo[27][0] ));
 INVx1_ASAP7_75t_R _11705_ (.A(_01308_),
    .Y(\peo[26][32] ));
 INVx1_ASAP7_75t_R _11706_ (.A(_01269_),
    .Y(\peo[27][32] ));
 INVx2_ASAP7_75t_R _11707_ (.A(_01307_),
    .Y(\peo[26][33] ));
 INVx2_ASAP7_75t_R _11708_ (.A(_01268_),
    .Y(\xs[13].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11709_ (.A(_01306_),
    .Y(\peo[26][34] ));
 INVx2_ASAP7_75t_R _11710_ (.A(_01267_),
    .Y(\xs[13].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11711_ (.A(_01305_),
    .Y(\peo[26][35] ));
 INVx1_ASAP7_75t_R _11712_ (.A(_01266_),
    .Y(\xs[13].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11713_ (.A(_01304_),
    .Y(\peo[26][36] ));
 INVx1_ASAP7_75t_R _11714_ (.A(_01265_),
    .Y(\xs[13].cli1.i[36] ));
 INVx2_ASAP7_75t_R _11715_ (.A(_01167_),
    .Y(\peo[29][0] ));
 INVx1_ASAP7_75t_R _11716_ (.A(_01206_),
    .Y(\peo[28][0] ));
 INVx1_ASAP7_75t_R _11717_ (.A(_01165_),
    .Y(\peo[29][32] ));
 INVx1_ASAP7_75t_R _11718_ (.A(_01204_),
    .Y(\peo[28][32] ));
 INVx2_ASAP7_75t_R _11719_ (.A(_01164_),
    .Y(\xs[14].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11720_ (.A(_01203_),
    .Y(\peo[28][33] ));
 INVx1_ASAP7_75t_R _11721_ (.A(_01163_),
    .Y(\xs[14].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11722_ (.A(_01202_),
    .Y(\peo[28][34] ));
 INVx1_ASAP7_75t_R _11723_ (.A(_01162_),
    .Y(\xs[14].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11724_ (.A(_01201_),
    .Y(\peo[28][35] ));
 INVx1_ASAP7_75t_R _11725_ (.A(_01161_),
    .Y(\xs[14].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11726_ (.A(_01200_),
    .Y(\peo[28][36] ));
 INVx1_ASAP7_75t_R _11727_ (.A(_01102_),
    .Y(\peo[30][0] ));
 INVx1_ASAP7_75t_R _11728_ (.A(_01063_),
    .Y(\peo[31][0] ));
 INVx1_ASAP7_75t_R _11729_ (.A(_01100_),
    .Y(\peo[30][32] ));
 INVx2_ASAP7_75t_R _11730_ (.A(_01061_),
    .Y(\peo[31][32] ));
 INVx1_ASAP7_75t_R _11731_ (.A(_01099_),
    .Y(\peo[30][33] ));
 INVx1_ASAP7_75t_R _11732_ (.A(_01060_),
    .Y(\xs[15].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11733_ (.A(_01098_),
    .Y(\peo[30][34] ));
 INVx1_ASAP7_75t_R _11734_ (.A(_01059_),
    .Y(\xs[15].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11735_ (.A(_01097_),
    .Y(\peo[30][35] ));
 INVx1_ASAP7_75t_R _11736_ (.A(_01058_),
    .Y(\xs[15].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11737_ (.A(_01096_),
    .Y(\peo[30][36] ));
 INVx1_ASAP7_75t_R _11738_ (.A(_01057_),
    .Y(\xs[15].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11739_ (.A(_00959_),
    .Y(\peo[3][0] ));
 INVx1_ASAP7_75t_R _11740_ (.A(_00998_),
    .Y(\peo[2][0] ));
 INVx2_ASAP7_75t_R _11741_ (.A(_00957_),
    .Y(\xs[1].cli1.i[32] ));
 INVx1_ASAP7_75t_R _11742_ (.A(_00996_),
    .Y(\peo[2][32] ));
 INVx2_ASAP7_75t_R _11743_ (.A(_00956_),
    .Y(\xs[1].cli1.i[33] ));
 INVx2_ASAP7_75t_R _11744_ (.A(_00995_),
    .Y(\peo[2][33] ));
 INVx1_ASAP7_75t_R _11745_ (.A(_00955_),
    .Y(\xs[1].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11746_ (.A(_00994_),
    .Y(\peo[2][34] ));
 INVx1_ASAP7_75t_R _11747_ (.A(_00954_),
    .Y(\xs[1].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11748_ (.A(_00993_),
    .Y(\peo[2][35] ));
 INVx1_ASAP7_75t_R _11749_ (.A(_00953_),
    .Y(\xs[1].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11750_ (.A(_00992_),
    .Y(\peo[2][36] ));
 INVx1_ASAP7_75t_R _11751_ (.A(_00855_),
    .Y(\peo[5][0] ));
 INVx1_ASAP7_75t_R _11752_ (.A(_00894_),
    .Y(\peo[4][0] ));
 INVx1_ASAP7_75t_R _11753_ (.A(_00853_),
    .Y(\xs[2].cli1.i[32] ));
 INVx1_ASAP7_75t_R _11754_ (.A(_00892_),
    .Y(\peo[4][32] ));
 INVx1_ASAP7_75t_R _11755_ (.A(_00852_),
    .Y(\xs[2].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11756_ (.A(_00891_),
    .Y(\peo[4][33] ));
 INVx1_ASAP7_75t_R _11757_ (.A(_00851_),
    .Y(\xs[2].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11758_ (.A(_00890_),
    .Y(\peo[4][34] ));
 INVx1_ASAP7_75t_R _11759_ (.A(_00850_),
    .Y(\xs[2].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11760_ (.A(_00889_),
    .Y(\peo[4][35] ));
 INVx1_ASAP7_75t_R _11761_ (.A(_00849_),
    .Y(\xs[2].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11762_ (.A(_00888_),
    .Y(\peo[4][36] ));
 INVx1_ASAP7_75t_R _11763_ (.A(_00751_),
    .Y(\peo[7][0] ));
 INVx1_ASAP7_75t_R _11764_ (.A(_00790_),
    .Y(\peo[6][0] ));
 INVx1_ASAP7_75t_R _11765_ (.A(_00749_),
    .Y(\xs[3].cli1.i[32] ));
 INVx1_ASAP7_75t_R _11766_ (.A(_00788_),
    .Y(\peo[6][32] ));
 INVx1_ASAP7_75t_R _11767_ (.A(_00748_),
    .Y(\xs[3].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11768_ (.A(_00787_),
    .Y(\peo[6][33] ));
 INVx1_ASAP7_75t_R _11769_ (.A(_00747_),
    .Y(\xs[3].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11770_ (.A(_00786_),
    .Y(\peo[6][34] ));
 INVx1_ASAP7_75t_R _11771_ (.A(_00746_),
    .Y(\xs[3].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11772_ (.A(_00785_),
    .Y(\peo[6][35] ));
 INVx1_ASAP7_75t_R _11773_ (.A(_00745_),
    .Y(\xs[3].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11774_ (.A(_00784_),
    .Y(\peo[6][36] ));
 INVx1_ASAP7_75t_R _11775_ (.A(_00647_),
    .Y(\peo[9][0] ));
 INVx1_ASAP7_75t_R _11776_ (.A(_00686_),
    .Y(\peo[8][0] ));
 INVx1_ASAP7_75t_R _11777_ (.A(_00645_),
    .Y(\xs[4].cli1.i[32] ));
 INVx1_ASAP7_75t_R _11778_ (.A(_00684_),
    .Y(\peo[8][32] ));
 INVx1_ASAP7_75t_R _11779_ (.A(_00644_),
    .Y(\xs[4].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11780_ (.A(_00683_),
    .Y(\peo[8][33] ));
 INVx1_ASAP7_75t_R _11781_ (.A(_00643_),
    .Y(\xs[4].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11782_ (.A(_00682_),
    .Y(\peo[8][34] ));
 INVx1_ASAP7_75t_R _11783_ (.A(_00642_),
    .Y(\xs[4].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11784_ (.A(_00681_),
    .Y(\peo[8][35] ));
 INVx1_ASAP7_75t_R _11785_ (.A(_00641_),
    .Y(\xs[4].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11786_ (.A(_00680_),
    .Y(\peo[8][36] ));
 INVx1_ASAP7_75t_R _11787_ (.A(_00543_),
    .Y(\peo[11][0] ));
 INVx1_ASAP7_75t_R _11788_ (.A(_00582_),
    .Y(\peo[10][0] ));
 INVx1_ASAP7_75t_R _11789_ (.A(_00439_),
    .Y(\peo[13][0] ));
 INVx1_ASAP7_75t_R _11790_ (.A(_00478_),
    .Y(\peo[12][0] ));
 INVx1_ASAP7_75t_R _11791_ (.A(_00437_),
    .Y(\xs[6].cli1.i[32] ));
 INVx1_ASAP7_75t_R _11792_ (.A(_00476_),
    .Y(\peo[12][32] ));
 INVx1_ASAP7_75t_R _11793_ (.A(_00436_),
    .Y(\xs[6].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11794_ (.A(_00475_),
    .Y(\peo[12][33] ));
 INVx1_ASAP7_75t_R _11795_ (.A(_00435_),
    .Y(\xs[6].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11796_ (.A(_00474_),
    .Y(\peo[12][34] ));
 INVx1_ASAP7_75t_R _11797_ (.A(_00434_),
    .Y(\xs[6].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11798_ (.A(_00473_),
    .Y(\peo[12][35] ));
 INVx1_ASAP7_75t_R _11799_ (.A(_00433_),
    .Y(\xs[6].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11800_ (.A(_00472_),
    .Y(\peo[12][36] ));
 INVx1_ASAP7_75t_R _11801_ (.A(_00374_),
    .Y(\peo[14][0] ));
 INVx2_ASAP7_75t_R _11802_ (.A(_00335_),
    .Y(\peo[15][0] ));
 INVx1_ASAP7_75t_R _11803_ (.A(_00372_),
    .Y(\peo[14][32] ));
 INVx1_ASAP7_75t_R _11804_ (.A(_00333_),
    .Y(\xs[7].cli1.i[32] ));
 INVx1_ASAP7_75t_R _11805_ (.A(_00371_),
    .Y(\peo[14][33] ));
 INVx1_ASAP7_75t_R _11806_ (.A(_00332_),
    .Y(\xs[7].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11807_ (.A(_00370_),
    .Y(\peo[14][34] ));
 INVx1_ASAP7_75t_R _11808_ (.A(_00331_),
    .Y(\xs[7].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11809_ (.A(_00369_),
    .Y(\peo[14][35] ));
 INVx1_ASAP7_75t_R _11810_ (.A(_00330_),
    .Y(\xs[7].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11811_ (.A(_00368_),
    .Y(\peo[14][36] ));
 INVx2_ASAP7_75t_R _11812_ (.A(_00329_),
    .Y(\xs[7].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11813_ (.A(_00231_),
    .Y(\peo[17][0] ));
 INVx1_ASAP7_75t_R _11814_ (.A(_00270_),
    .Y(\peo[16][0] ));
 INVx1_ASAP7_75t_R _11815_ (.A(_00229_),
    .Y(\xs[8].cli1.i[32] ));
 INVx1_ASAP7_75t_R _11816_ (.A(_00268_),
    .Y(\peo[16][32] ));
 INVx1_ASAP7_75t_R _11817_ (.A(_00228_),
    .Y(\xs[8].cli1.i[33] ));
 INVx1_ASAP7_75t_R _11818_ (.A(_00267_),
    .Y(\peo[16][33] ));
 INVx1_ASAP7_75t_R _11819_ (.A(_00227_),
    .Y(\xs[8].cli1.i[34] ));
 INVx1_ASAP7_75t_R _11820_ (.A(_00266_),
    .Y(\peo[16][34] ));
 INVx1_ASAP7_75t_R _11821_ (.A(_00226_),
    .Y(\xs[8].cli1.i[35] ));
 INVx1_ASAP7_75t_R _11822_ (.A(_00265_),
    .Y(\peo[16][35] ));
 INVx2_ASAP7_75t_R _11823_ (.A(_00225_),
    .Y(\xs[8].cli1.i[36] ));
 INVx1_ASAP7_75t_R _11824_ (.A(_00264_),
    .Y(\peo[16][36] ));
 INVx1_ASAP7_75t_R _11825_ (.A(_00127_),
    .Y(\peo[19][0] ));
 INVx1_ASAP7_75t_R _11826_ (.A(_00166_),
    .Y(\peo[18][0] ));
 INVx1_ASAP7_75t_R _11827_ (.A(_00125_),
    .Y(\peo[19][32] ));
 INVx1_ASAP7_75t_R _11828_ (.A(_00164_),
    .Y(\peo[18][32] ));
 INVx1_ASAP7_75t_R _11829_ (.A(_00124_),
    .Y(\peo[19][33] ));
 INVx1_ASAP7_75t_R _11830_ (.A(_00163_),
    .Y(\peo[18][33] ));
 INVx1_ASAP7_75t_R _11831_ (.A(_00123_),
    .Y(\peo[19][34] ));
 INVx1_ASAP7_75t_R _11832_ (.A(_00162_),
    .Y(\peo[18][34] ));
 INVx1_ASAP7_75t_R _11833_ (.A(_00122_),
    .Y(\peo[19][35] ));
 INVx1_ASAP7_75t_R _11834_ (.A(_00161_),
    .Y(\peo[18][35] ));
 INVx1_ASAP7_75t_R _11835_ (.A(_00121_),
    .Y(\peo[19][36] ));
 INVx1_ASAP7_75t_R _11836_ (.A(_00160_),
    .Y(\peo[18][36] ));
 INVx1_ASAP7_75t_R _11837_ (.A(_00213_),
    .Y(\xs[8].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11838_ (.A(_00060_),
    .Y(\xs[8].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11839_ (.A(_01253_),
    .Y(\xs[13].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11840_ (.A(_00040_),
    .Y(\xs[13].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11841_ (.A(_00980_),
    .Y(\xs[1].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11842_ (.A(_00045_),
    .Y(\xs[1].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11843_ (.A(_01045_),
    .Y(\xs[15].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11844_ (.A(_00044_),
    .Y(\xs[15].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11845_ (.A(_00525_),
    .Y(\xs[5].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11846_ (.A(_00054_),
    .Y(\xs[5].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11847_ (.A(_00460_),
    .Y(\xs[6].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11848_ (.A(_00055_),
    .Y(\xs[6].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11849_ (.A(_01669_),
    .Y(\xs[0].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11850_ (.A(_00032_),
    .Y(\xs[0].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11851_ (.A(_01357_),
    .Y(\xs[12].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11852_ (.A(_00038_),
    .Y(\xs[12].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11853_ (.A(_01604_),
    .Y(\xs[10].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11854_ (.A(_00033_),
    .Y(\xs[10].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11855_ (.A(_01084_),
    .Y(\xs[15].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11856_ (.A(_00043_),
    .Y(\xs[15].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11857_ (.A(_01708_),
    .Y(\xs[0].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11858_ (.A(_00031_),
    .Y(\xs[0].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11859_ (.A(_01149_),
    .Y(\xs[14].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11860_ (.A(_00042_),
    .Y(\xs[14].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11861_ (.A(_01565_),
    .Y(\xs[10].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11862_ (.A(_00034_),
    .Y(\xs[10].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11863_ (.A(_01500_),
    .Y(\xs[11].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11864_ (.A(_00035_),
    .Y(\xs[11].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11865_ (.A(_00421_),
    .Y(\xs[6].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11866_ (.A(_00056_),
    .Y(\xs[6].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11867_ (.A(_00629_),
    .Y(\xs[4].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11868_ (.A(_00052_),
    .Y(\xs[4].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11869_ (.A(_01461_),
    .Y(\xs[11].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11870_ (.A(_00036_),
    .Y(\xs[11].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11871_ (.A(_01292_),
    .Y(\xs[13].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11872_ (.A(_00039_),
    .Y(\xs[13].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11873_ (.A(_00148_),
    .Y(\xs[9].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11874_ (.A(_00061_),
    .Y(\xs[9].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11875_ (.A(_00564_),
    .Y(\xs[5].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11876_ (.A(_00053_),
    .Y(\xs[5].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11877_ (.A(_00356_),
    .Y(\xs[7].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11878_ (.A(_00057_),
    .Y(\xs[7].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11879_ (.A(_00109_),
    .Y(\xs[9].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11880_ (.A(_00062_),
    .Y(\xs[9].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11881_ (.A(_01396_),
    .Y(\xs[12].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11882_ (.A(_00037_),
    .Y(\xs[12].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11883_ (.A(_00772_),
    .Y(\xs[3].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11884_ (.A(_00049_),
    .Y(\xs[3].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11885_ (.A(_00941_),
    .Y(\xs[1].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11886_ (.A(_00046_),
    .Y(\xs[1].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11887_ (.A(_00668_),
    .Y(\xs[4].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11888_ (.A(_00051_),
    .Y(\xs[4].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11889_ (.A(_01188_),
    .Y(\xs[14].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11890_ (.A(_00041_),
    .Y(\xs[14].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11891_ (.A(_00317_),
    .Y(\xs[7].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11892_ (.A(_00058_),
    .Y(\xs[7].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11893_ (.A(_00733_),
    .Y(\xs[3].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11894_ (.A(_00050_),
    .Y(\xs[3].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11895_ (.A(_00876_),
    .Y(\xs[2].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11896_ (.A(_00047_),
    .Y(\xs[2].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11897_ (.A(_00252_),
    .Y(\xs[8].cli0.r[1] ));
 INVx1_ASAP7_75t_R _11898_ (.A(_00059_),
    .Y(\xs[8].cli0.r[0] ));
 INVx1_ASAP7_75t_R _11899_ (.A(_00837_),
    .Y(\xs[2].cli1.r[1] ));
 INVx1_ASAP7_75t_R _11900_ (.A(_00048_),
    .Y(\xs[2].cli1.r[0] ));
 INVx1_ASAP7_75t_R _11901_ (.A(_00952_),
    .Y(\xs[1].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11902_ (.A(_00991_),
    .Y(\peo[2][39] ));
 INVx1_ASAP7_75t_R _11903_ (.A(_00848_),
    .Y(\xs[2].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11904_ (.A(_00887_),
    .Y(\peo[4][39] ));
 INVx2_ASAP7_75t_R _11905_ (.A(_01056_),
    .Y(\xs[15].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11906_ (.A(_01095_),
    .Y(\peo[30][39] ));
 INVx1_ASAP7_75t_R _11907_ (.A(_01680_),
    .Y(\xs[0].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11908_ (.A(_01719_),
    .Y(\peo[0][39] ));
 INVx2_ASAP7_75t_R _11909_ (.A(_01160_),
    .Y(\xs[14].cli1.i[39] ));
 INVx2_ASAP7_75t_R _11910_ (.A(_01199_),
    .Y(\peo[28][39] ));
 INVx1_ASAP7_75t_R _11911_ (.A(_01264_),
    .Y(\xs[13].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11912_ (.A(_01303_),
    .Y(\peo[26][39] ));
 INVx2_ASAP7_75t_R _11913_ (.A(_01368_),
    .Y(\xs[12].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11914_ (.A(_01407_),
    .Y(\peo[24][39] ));
 INVx1_ASAP7_75t_R _11915_ (.A(_01472_),
    .Y(\xs[11].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11916_ (.A(_01511_),
    .Y(\peo[22][39] ));
 INVx3_ASAP7_75t_R _11917_ (.A(_01576_),
    .Y(\xs[10].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11918_ (.A(_01615_),
    .Y(\peo[20][39] ));
 INVx1_ASAP7_75t_R _11919_ (.A(_00744_),
    .Y(\xs[3].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11920_ (.A(_00783_),
    .Y(\peo[6][39] ));
 INVx1_ASAP7_75t_R _11921_ (.A(_00328_),
    .Y(\xs[7].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11922_ (.A(_00367_),
    .Y(\peo[14][39] ));
 INVx1_ASAP7_75t_R _11923_ (.A(_00224_),
    .Y(\xs[8].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11924_ (.A(_00263_),
    .Y(\peo[16][39] ));
 INVx1_ASAP7_75t_R _11925_ (.A(_00432_),
    .Y(\xs[6].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11926_ (.A(_00471_),
    .Y(\peo[12][39] ));
 INVx2_ASAP7_75t_R _11927_ (.A(_00120_),
    .Y(\peo[19][39] ));
 INVx2_ASAP7_75t_R _11928_ (.A(_00159_),
    .Y(\peo[18][39] ));
 INVx1_ASAP7_75t_R _11929_ (.A(_00640_),
    .Y(\xs[4].cli1.i[39] ));
 INVx1_ASAP7_75t_R _11930_ (.A(_00679_),
    .Y(\peo[8][39] ));
 INVx1_ASAP7_75t_R _11931_ (.A(_00126_),
    .Y(\peo[19][10] ));
 INVx1_ASAP7_75t_R _11932_ (.A(_00165_),
    .Y(\peo[18][11] ));
 INVx1_ASAP7_75t_R _11933_ (.A(_00230_),
    .Y(\peo[17][10] ));
 INVx1_ASAP7_75t_R _11934_ (.A(_00269_),
    .Y(\peo[16][14] ));
 INVx1_ASAP7_75t_R _11935_ (.A(_00334_),
    .Y(\peo[15][10] ));
 INVx1_ASAP7_75t_R _11936_ (.A(_00373_),
    .Y(\peo[14][11] ));
 INVx1_ASAP7_75t_R _11937_ (.A(_00438_),
    .Y(\peo[13][10] ));
 INVx1_ASAP7_75t_R _11938_ (.A(_00477_),
    .Y(\peo[12][12] ));
 INVx1_ASAP7_75t_R _11939_ (.A(_00542_),
    .Y(\peo[11][10] ));
 INVx1_ASAP7_75t_R _11940_ (.A(_00581_),
    .Y(\peo[10][11] ));
 INVx1_ASAP7_75t_R _11941_ (.A(_00646_),
    .Y(\peo[9][10] ));
 INVx1_ASAP7_75t_R _11942_ (.A(_00685_),
    .Y(\peo[8][13] ));
 INVx1_ASAP7_75t_R _11943_ (.A(_00750_),
    .Y(\peo[7][10] ));
 INVx1_ASAP7_75t_R _11944_ (.A(_00789_),
    .Y(\peo[6][11] ));
 INVx1_ASAP7_75t_R _11945_ (.A(_00854_),
    .Y(\peo[5][10] ));
 INVx1_ASAP7_75t_R _11946_ (.A(_00893_),
    .Y(\peo[4][12] ));
 INVx1_ASAP7_75t_R _11947_ (.A(_00958_),
    .Y(\xs[1].cli1.i[10] ));
 INVx1_ASAP7_75t_R _11948_ (.A(_00997_),
    .Y(\peo[2][11] ));
 INVx1_ASAP7_75t_R _11949_ (.A(_01062_),
    .Y(\peo[31][10] ));
 INVx1_ASAP7_75t_R _11950_ (.A(_01101_),
    .Y(\peo[30][11] ));
 INVx1_ASAP7_75t_R _11951_ (.A(_01166_),
    .Y(\peo[29][10] ));
 INVx1_ASAP7_75t_R _11952_ (.A(_01205_),
    .Y(\peo[28][12] ));
 INVx1_ASAP7_75t_R _11953_ (.A(_01270_),
    .Y(\peo[27][10] ));
 INVx1_ASAP7_75t_R _11954_ (.A(_01309_),
    .Y(\peo[26][11] ));
 INVx1_ASAP7_75t_R _11955_ (.A(_01374_),
    .Y(\peo[25][10] ));
 INVx1_ASAP7_75t_R _11956_ (.A(_01413_),
    .Y(\peo[24][13] ));
 INVx1_ASAP7_75t_R _11957_ (.A(_01478_),
    .Y(\peo[23][10] ));
 INVx1_ASAP7_75t_R _11958_ (.A(_01517_),
    .Y(\peo[22][11] ));
 INVx1_ASAP7_75t_R _11959_ (.A(_01582_),
    .Y(\peo[21][10] ));
 INVx1_ASAP7_75t_R _11960_ (.A(_01621_),
    .Y(\peo[20][12] ));
 INVx1_ASAP7_75t_R _11961_ (.A(_01686_),
    .Y(\peo[1][10] ));
 INVx1_ASAP7_75t_R _11962_ (.A(_01726_),
    .Y(net325));
 INVx2_ASAP7_75t_R _11963_ (.A(_02357_),
    .Y(net22));
 INVx2_ASAP7_75t_R _11964_ (.A(_02358_),
    .Y(net23));
 INVx3_ASAP7_75t_R _11965_ (.A(_02359_),
    .Y(net26));
 INVx2_ASAP7_75t_R _11966_ (.A(_02360_),
    .Y(net27));
 INVx1_ASAP7_75t_R _11967_ (.A(_02361_),
    .Y(net28));
 INVx1_ASAP7_75t_R _11968_ (.A(_02362_),
    .Y(net29));
 INVx2_ASAP7_75t_R _11969_ (.A(_02363_),
    .Y(net30));
 INVx2_ASAP7_75t_R _11970_ (.A(_02364_),
    .Y(net31));
 INVx2_ASAP7_75t_R _11971_ (.A(_02365_),
    .Y(net32));
 INVx1_ASAP7_75t_R _11972_ (.A(_02366_),
    .Y(net33));
 INVx2_ASAP7_75t_R _11973_ (.A(_02367_),
    .Y(net36));
 INVx1_ASAP7_75t_R _11974_ (.A(_02368_),
    .Y(net37));
 INVx1_ASAP7_75t_R _11975_ (.A(_02369_),
    .Y(net38));
 INVx1_ASAP7_75t_R _11976_ (.A(_02370_),
    .Y(net39));
 INVx1_ASAP7_75t_R _11977_ (.A(_02371_),
    .Y(net40));
 INVx1_ASAP7_75t_R _11978_ (.A(_02372_),
    .Y(net41));
 INVx1_ASAP7_75t_R _11979_ (.A(_02373_),
    .Y(net42));
 INVx1_ASAP7_75t_R _11980_ (.A(_02374_),
    .Y(net43));
 INVx2_ASAP7_75t_R _11981_ (.A(_02375_),
    .Y(net47));
 INVx1_ASAP7_75t_R _11982_ (.A(_02376_),
    .Y(net48));
 INVx1_ASAP7_75t_R _11983_ (.A(_02377_),
    .Y(net49));
 INVx1_ASAP7_75t_R _11984_ (.A(_02378_),
    .Y(net50));
 INVx1_ASAP7_75t_R _11985_ (.A(_02379_),
    .Y(net51));
 INVx1_ASAP7_75t_R _11986_ (.A(_02380_),
    .Y(net52));
 INVx1_ASAP7_75t_R _11987_ (.A(_02381_),
    .Y(net53));
 INVx1_ASAP7_75t_R _11988_ (.A(_02382_),
    .Y(net54));
 INVx2_ASAP7_75t_R _11989_ (.A(_02383_),
    .Y(net55));
 INVx3_ASAP7_75t_R _11990_ (.A(_02384_),
    .Y(net58));
 INVx2_ASAP7_75t_R _11991_ (.A(_02385_),
    .Y(net59));
 INVx2_ASAP7_75t_R _11992_ (.A(_02386_),
    .Y(net60));
 INVx1_ASAP7_75t_R _11993_ (.A(_02387_),
    .Y(net61));
 INVx1_ASAP7_75t_R _11994_ (.A(_02388_),
    .Y(net62));
 INVx1_ASAP7_75t_R _11995_ (.A(_02389_),
    .Y(net63));
 INVx1_ASAP7_75t_R _11996_ (.A(_02390_),
    .Y(net64));
 INVx1_ASAP7_75t_R _11997_ (.A(_02391_),
    .Y(net65));
 INVx1_ASAP7_75t_R _11998_ (.A(_02392_),
    .Y(net66));
 INVx1_ASAP7_75t_R _11999_ (.A(_02393_),
    .Y(net67));
 INVx1_ASAP7_75t_R _12000_ (.A(_02394_),
    .Y(net68));
 INVx2_ASAP7_75t_R _12001_ (.A(_02395_),
    .Y(net69));
 INVx3_ASAP7_75t_R _12002_ (.A(_02396_),
    .Y(net73));
 INVx1_ASAP7_75t_R _12003_ (.A(_02397_),
    .Y(net74));
 INVx1_ASAP7_75t_R _12004_ (.A(_02398_),
    .Y(net75));
 INVx1_ASAP7_75t_R _12005_ (.A(_02399_),
    .Y(net76));
 INVx1_ASAP7_75t_R _12006_ (.A(_02400_),
    .Y(net77));
 INVx1_ASAP7_75t_R _12007_ (.A(_02401_),
    .Y(net78));
 INVx1_ASAP7_75t_R _12008_ (.A(_02402_),
    .Y(net79));
 INVx2_ASAP7_75t_R _12009_ (.A(_02403_),
    .Y(net80));
 INVx1_ASAP7_75t_R _12010_ (.A(_02404_),
    .Y(net81));
 INVx2_ASAP7_75t_R _12011_ (.A(_02405_),
    .Y(net82));
 INVx3_ASAP7_75t_R _12012_ (.A(_02406_),
    .Y(net86));
 INVx1_ASAP7_75t_R _12013_ (.A(_02407_),
    .Y(net87));
 INVx2_ASAP7_75t_R _12014_ (.A(_02408_),
    .Y(net88));
 INVx2_ASAP7_75t_R _12015_ (.A(_02409_),
    .Y(net89));
 INVx2_ASAP7_75t_R _12016_ (.A(_02410_),
    .Y(net90));
 INVx2_ASAP7_75t_R _12017_ (.A(_02411_),
    .Y(net91));
 INVx1_ASAP7_75t_R _12018_ (.A(_02412_),
    .Y(net92));
 INVx1_ASAP7_75t_R _12019_ (.A(_02413_),
    .Y(net93));
 INVx2_ASAP7_75t_R _12020_ (.A(_02414_),
    .Y(net98));
 INVx1_ASAP7_75t_R _12021_ (.A(_02415_),
    .Y(net99));
 INVx2_ASAP7_75t_R _12022_ (.A(_02416_),
    .Y(net100));
 INVx2_ASAP7_75t_R _12023_ (.A(_02417_),
    .Y(net101));
 INVx2_ASAP7_75t_R _12024_ (.A(_02418_),
    .Y(net102));
 INVx2_ASAP7_75t_R _12025_ (.A(_02419_),
    .Y(net103));
 INVx1_ASAP7_75t_R _12026_ (.A(_02420_),
    .Y(net104));
 INVx2_ASAP7_75t_R _12027_ (.A(_02421_),
    .Y(net106));
 INVx2_ASAP7_75t_R _12028_ (.A(_02422_),
    .Y(net107));
 INVx2_ASAP7_75t_R _12029_ (.A(_02423_),
    .Y(net108));
 INVx2_ASAP7_75t_R _12030_ (.A(_02424_),
    .Y(net109));
 INVx2_ASAP7_75t_R _12031_ (.A(_02425_),
    .Y(net110));
 INVx2_ASAP7_75t_R _12032_ (.A(_02426_),
    .Y(net111));
 INVx2_ASAP7_75t_R _12033_ (.A(_02427_),
    .Y(net112));
 INVx2_ASAP7_75t_R _12034_ (.A(_02428_),
    .Y(net113));
 INVx1_ASAP7_75t_R _12035_ (.A(_02429_),
    .Y(net114));
 INVx2_ASAP7_75t_R _12036_ (.A(_02430_),
    .Y(net115));
 INVx2_ASAP7_75t_R _12037_ (.A(_02431_),
    .Y(net116));
 INVx2_ASAP7_75t_R _12038_ (.A(_02432_),
    .Y(net117));
 INVx2_ASAP7_75t_R _12039_ (.A(_02433_),
    .Y(net118));
 INVx2_ASAP7_75t_R _12040_ (.A(_02434_),
    .Y(net119));
 INVx2_ASAP7_75t_R _12041_ (.A(_02435_),
    .Y(net120));
 INVx2_ASAP7_75t_R _12042_ (.A(_02436_),
    .Y(net121));
 INVx2_ASAP7_75t_R _12043_ (.A(_02437_),
    .Y(net123));
 INVx2_ASAP7_75t_R _12044_ (.A(_02438_),
    .Y(net124));
 INVx2_ASAP7_75t_R _12045_ (.A(_02439_),
    .Y(net125));
 INVx2_ASAP7_75t_R _12046_ (.A(_02440_),
    .Y(net126));
 INVx2_ASAP7_75t_R _12047_ (.A(_02441_),
    .Y(net127));
 INVx2_ASAP7_75t_R _12048_ (.A(_02442_),
    .Y(net128));
 INVx2_ASAP7_75t_R _12049_ (.A(_02443_),
    .Y(net129));
 INVx2_ASAP7_75t_R _12050_ (.A(_02444_),
    .Y(net130));
 INVx2_ASAP7_75t_R _12051_ (.A(_02445_),
    .Y(net132));
 INVx2_ASAP7_75t_R _12052_ (.A(_02446_),
    .Y(net133));
 INVx2_ASAP7_75t_R _12053_ (.A(_02447_),
    .Y(net134));
 INVx2_ASAP7_75t_R _12054_ (.A(_02448_),
    .Y(net135));
 INVx2_ASAP7_75t_R _12055_ (.A(_02449_),
    .Y(net136));
 INVx2_ASAP7_75t_R _12056_ (.A(_02450_),
    .Y(net137));
 INVx2_ASAP7_75t_R _12057_ (.A(_02451_),
    .Y(net138));
 INVx2_ASAP7_75t_R _12058_ (.A(_02452_),
    .Y(net139));
 INVx2_ASAP7_75t_R _12059_ (.A(_02453_),
    .Y(net142));
 INVx2_ASAP7_75t_R _12060_ (.A(_02454_),
    .Y(net143));
 INVx2_ASAP7_75t_R _12061_ (.A(_02455_),
    .Y(net144));
 INVx2_ASAP7_75t_R _12062_ (.A(_02456_),
    .Y(net145));
 INVx2_ASAP7_75t_R _12063_ (.A(_02457_),
    .Y(net146));
 INVx2_ASAP7_75t_R _12064_ (.A(_02458_),
    .Y(net147));
 INVx2_ASAP7_75t_R _12065_ (.A(_02459_),
    .Y(net148));
 INVx1_ASAP7_75t_R _12066_ (.A(_02460_),
    .Y(net149));
 INVx2_ASAP7_75t_R _12067_ (.A(_02461_),
    .Y(net150));
 INVx1_ASAP7_75t_R _12068_ (.A(_02462_),
    .Y(net151));
 INVx2_ASAP7_75t_R _12069_ (.A(_02463_),
    .Y(net152));
 INVx2_ASAP7_75t_R _12070_ (.A(_02464_),
    .Y(net153));
 INVx1_ASAP7_75t_R _12071_ (.A(_02465_),
    .Y(net154));
 INVx2_ASAP7_75t_R _12072_ (.A(_02466_),
    .Y(net155));
 INVx2_ASAP7_75t_R _12073_ (.A(_02467_),
    .Y(net156));
 INVx1_ASAP7_75t_R _12074_ (.A(_02468_),
    .Y(net157));
 INVx1_ASAP7_75t_R _12075_ (.A(_02469_),
    .Y(net158));
 INVx1_ASAP7_75t_R _12076_ (.A(_02470_),
    .Y(net159));
 INVx2_ASAP7_75t_R _12077_ (.A(_02471_),
    .Y(net160));
 INVx1_ASAP7_75t_R _12078_ (.A(_02472_),
    .Y(net161));
 INVx2_ASAP7_75t_R _12079_ (.A(_02473_),
    .Y(net162));
 INVx2_ASAP7_75t_R _12080_ (.A(_02474_),
    .Y(net164));
 INVx1_ASAP7_75t_R _12081_ (.A(_02475_),
    .Y(net165));
 INVx1_ASAP7_75t_R _12082_ (.A(_02476_),
    .Y(net166));
 INVx1_ASAP7_75t_R _12083_ (.A(_02477_),
    .Y(net167));
 INVx1_ASAP7_75t_R _12084_ (.A(_02478_),
    .Y(net168));
 INVx1_ASAP7_75t_R _12085_ (.A(_02479_),
    .Y(net169));
 INVx1_ASAP7_75t_R _12086_ (.A(_02480_),
    .Y(net170));
 INVx2_ASAP7_75t_R _12087_ (.A(_02481_),
    .Y(net171));
 INVx1_ASAP7_75t_R _12088_ (.A(_02482_),
    .Y(net172));
 INVx2_ASAP7_75t_R _12089_ (.A(_02483_),
    .Y(net173));
 INVx1_ASAP7_75t_R _12090_ (.A(_02484_),
    .Y(net175));
 INVx1_ASAP7_75t_R _12091_ (.A(_02485_),
    .Y(net176));
 INVx1_ASAP7_75t_R _12092_ (.A(_02486_),
    .Y(net177));
 INVx1_ASAP7_75t_R _12093_ (.A(_02487_),
    .Y(net178));
 INVx1_ASAP7_75t_R _12094_ (.A(_02488_),
    .Y(net179));
 INVx1_ASAP7_75t_R _12095_ (.A(_02489_),
    .Y(net180));
 INVx1_ASAP7_75t_R _12096_ (.A(_02490_),
    .Y(net181));
 INVx1_ASAP7_75t_R _12097_ (.A(_02491_),
    .Y(net182));
 INVx2_ASAP7_75t_R _12098_ (.A(_02492_),
    .Y(net185));
 INVx1_ASAP7_75t_R _12099_ (.A(_02493_),
    .Y(net186));
 INVx1_ASAP7_75t_R _12100_ (.A(_02494_),
    .Y(net187));
 INVx1_ASAP7_75t_R _12101_ (.A(_02495_),
    .Y(net188));
 INVx1_ASAP7_75t_R _12102_ (.A(_02496_),
    .Y(net189));
 INVx1_ASAP7_75t_R _12103_ (.A(_02497_),
    .Y(net190));
 INVx1_ASAP7_75t_R _12104_ (.A(_02498_),
    .Y(net191));
 INVx1_ASAP7_75t_R _12105_ (.A(_02499_),
    .Y(net192));
 INVx1_ASAP7_75t_R _12106_ (.A(_02500_),
    .Y(net194));
 INVx2_ASAP7_75t_R _12107_ (.A(_02501_),
    .Y(net195));
 INVx1_ASAP7_75t_R _12108_ (.A(_02502_),
    .Y(net196));
 INVx1_ASAP7_75t_R _12109_ (.A(_02503_),
    .Y(net197));
 INVx1_ASAP7_75t_R _12110_ (.A(_02504_),
    .Y(net198));
 INVx1_ASAP7_75t_R _12111_ (.A(_02505_),
    .Y(net199));
 INVx1_ASAP7_75t_R _12112_ (.A(_02506_),
    .Y(net200));
 INVx1_ASAP7_75t_R _12113_ (.A(_02507_),
    .Y(net201));
 INVx2_ASAP7_75t_R _12114_ (.A(_02508_),
    .Y(net202));
 INVx2_ASAP7_75t_R _12115_ (.A(_02509_),
    .Y(net205));
 INVx1_ASAP7_75t_R _12116_ (.A(_02510_),
    .Y(net206));
 INVx1_ASAP7_75t_R _12117_ (.A(_02511_),
    .Y(net207));
 INVx1_ASAP7_75t_R _12118_ (.A(_02512_),
    .Y(net208));
 INVx1_ASAP7_75t_R _12119_ (.A(_02513_),
    .Y(net209));
 INVx2_ASAP7_75t_R _12120_ (.A(_02514_),
    .Y(net210));
 INVx2_ASAP7_75t_R _12121_ (.A(_02515_),
    .Y(net211));
 INVx2_ASAP7_75t_R _12122_ (.A(_02516_),
    .Y(net212));
 INVx1_ASAP7_75t_R _12123_ (.A(_02517_),
    .Y(net215));
 INVx1_ASAP7_75t_R _12124_ (.A(_02518_),
    .Y(net216));
 INVx1_ASAP7_75t_R _12125_ (.A(_02519_),
    .Y(net217));
 INVx1_ASAP7_75t_R _12126_ (.A(_02520_),
    .Y(net218));
 INVx1_ASAP7_75t_R _12127_ (.A(_02521_),
    .Y(net219));
 INVx1_ASAP7_75t_R _12128_ (.A(_02522_),
    .Y(net220));
 INVx1_ASAP7_75t_R _12129_ (.A(_02523_),
    .Y(net221));
 INVx1_ASAP7_75t_R _12130_ (.A(_02524_),
    .Y(net222));
 INVx2_ASAP7_75t_R _12131_ (.A(_02525_),
    .Y(net226));
 INVx1_ASAP7_75t_R _12132_ (.A(_02526_),
    .Y(net227));
 INVx1_ASAP7_75t_R _12133_ (.A(_02527_),
    .Y(net228));
 INVx1_ASAP7_75t_R _12134_ (.A(_02528_),
    .Y(net229));
 INVx1_ASAP7_75t_R _12135_ (.A(_02529_),
    .Y(net230));
 INVx1_ASAP7_75t_R _12136_ (.A(_02530_),
    .Y(net231));
 INVx1_ASAP7_75t_R _12137_ (.A(_02531_),
    .Y(net232));
 INVx1_ASAP7_75t_R _12138_ (.A(_02532_),
    .Y(net233));
 INVx1_ASAP7_75t_R _12139_ (.A(_02533_),
    .Y(net234));
 INVx1_ASAP7_75t_R _12140_ (.A(_02534_),
    .Y(net235));
 INVx1_ASAP7_75t_R _12141_ (.A(_02535_),
    .Y(net236));
 INVx1_ASAP7_75t_R _12142_ (.A(_02536_),
    .Y(net237));
 INVx1_ASAP7_75t_R _12143_ (.A(_02537_),
    .Y(net238));
 INVx1_ASAP7_75t_R _12144_ (.A(_02538_),
    .Y(net239));
 INVx1_ASAP7_75t_R _12145_ (.A(_02539_),
    .Y(net240));
 INVx1_ASAP7_75t_R _12146_ (.A(_02540_),
    .Y(net241));
 INVx1_ASAP7_75t_R _12147_ (.A(_02541_),
    .Y(net243));
 INVx1_ASAP7_75t_R _12148_ (.A(_02542_),
    .Y(net244));
 INVx1_ASAP7_75t_R _12149_ (.A(_02543_),
    .Y(net245));
 INVx1_ASAP7_75t_R _12150_ (.A(_02544_),
    .Y(net246));
 INVx1_ASAP7_75t_R _12151_ (.A(_02545_),
    .Y(net247));
 INVx1_ASAP7_75t_R _12152_ (.A(_02546_),
    .Y(net248));
 INVx1_ASAP7_75t_R _12153_ (.A(_02547_),
    .Y(net249));
 INVx1_ASAP7_75t_R _12154_ (.A(_02548_),
    .Y(net250));
 INVx2_ASAP7_75t_R _12155_ (.A(_02549_),
    .Y(net251));
 INVx2_ASAP7_75t_R _12156_ (.A(_02550_),
    .Y(net253));
 INVx2_ASAP7_75t_R _12157_ (.A(_02551_),
    .Y(net254));
 INVx2_ASAP7_75t_R _12158_ (.A(_02552_),
    .Y(net255));
 INVx1_ASAP7_75t_R _12159_ (.A(_02553_),
    .Y(net256));
 INVx1_ASAP7_75t_R _12160_ (.A(_02554_),
    .Y(net257));
 INVx1_ASAP7_75t_R _12161_ (.A(_02555_),
    .Y(net258));
 INVx1_ASAP7_75t_R _12162_ (.A(_02556_),
    .Y(net259));
 INVx1_ASAP7_75t_R _12163_ (.A(_02557_),
    .Y(net260));
 INVx1_ASAP7_75t_R _12164_ (.A(_02558_),
    .Y(net261));
 INVx2_ASAP7_75t_R _12165_ (.A(_02559_),
    .Y(net262));
 INVx1_ASAP7_75t_R _12166_ (.A(_02560_),
    .Y(net263));
 INVx2_ASAP7_75t_R _12167_ (.A(_02561_),
    .Y(net264));
 INVx1_ASAP7_75t_R _12168_ (.A(_02562_),
    .Y(net267));
 INVx1_ASAP7_75t_R _12169_ (.A(_02563_),
    .Y(net268));
 INVx1_ASAP7_75t_R _12170_ (.A(_02564_),
    .Y(net269));
 INVx1_ASAP7_75t_R _12171_ (.A(_02565_),
    .Y(net270));
 INVx1_ASAP7_75t_R _12172_ (.A(_02566_),
    .Y(net271));
 INVx1_ASAP7_75t_R _12173_ (.A(_02567_),
    .Y(net272));
 INVx1_ASAP7_75t_R _12174_ (.A(_02568_),
    .Y(net273));
 INVx2_ASAP7_75t_R _12175_ (.A(_02569_),
    .Y(net274));
 INVx2_ASAP7_75t_R _12176_ (.A(_02570_),
    .Y(net275));
 INVx2_ASAP7_75t_R _12177_ (.A(_02571_),
    .Y(net276));
 INVx1_ASAP7_75t_R _12178_ (.A(_02572_),
    .Y(net278));
 INVx2_ASAP7_75t_R _12179_ (.A(_02573_),
    .Y(net279));
 INVx1_ASAP7_75t_R _12180_ (.A(_02574_),
    .Y(net280));
 INVx2_ASAP7_75t_R _12181_ (.A(_02575_),
    .Y(net281));
 INVx1_ASAP7_75t_R _12182_ (.A(_02576_),
    .Y(net282));
 INVx1_ASAP7_75t_R _12183_ (.A(_02577_),
    .Y(net283));
 INVx2_ASAP7_75t_R _12184_ (.A(_02578_),
    .Y(net284));
 INVx2_ASAP7_75t_R _12185_ (.A(_02579_),
    .Y(net285));
 INVx1_ASAP7_75t_R _12186_ (.A(_02580_),
    .Y(net288));
 INVx1_ASAP7_75t_R _12187_ (.A(_02581_),
    .Y(net289));
 INVx1_ASAP7_75t_R _12188_ (.A(_02582_),
    .Y(net290));
 INVx2_ASAP7_75t_R _12189_ (.A(_02583_),
    .Y(net291));
 INVx1_ASAP7_75t_R _12190_ (.A(_02584_),
    .Y(net292));
 INVx1_ASAP7_75t_R _12191_ (.A(_02585_),
    .Y(net293));
 INVx1_ASAP7_75t_R _12192_ (.A(_02586_),
    .Y(net294));
 INVx1_ASAP7_75t_R _12193_ (.A(_02587_),
    .Y(net295));
 INVx2_ASAP7_75t_R _12194_ (.A(_02588_),
    .Y(net298));
 INVx1_ASAP7_75t_R _12195_ (.A(_02589_),
    .Y(net299));
 INVx1_ASAP7_75t_R _12196_ (.A(_02590_),
    .Y(net300));
 INVx1_ASAP7_75t_R _12197_ (.A(_02591_),
    .Y(net301));
 INVx1_ASAP7_75t_R _12198_ (.A(_02592_),
    .Y(net302));
 INVx1_ASAP7_75t_R _12199_ (.A(_02593_),
    .Y(net303));
 INVx1_ASAP7_75t_R _12200_ (.A(_02594_),
    .Y(net304));
 INVx2_ASAP7_75t_R _12201_ (.A(_02595_),
    .Y(net305));
 INVx1_ASAP7_75t_R _12202_ (.A(_02596_),
    .Y(net306));
 INVx2_ASAP7_75t_R _12203_ (.A(_02597_),
    .Y(net310));
 INVx2_ASAP7_75t_R _12204_ (.A(_02598_),
    .Y(net311));
 INVx2_ASAP7_75t_R _12205_ (.A(_02599_),
    .Y(net312));
 INVx2_ASAP7_75t_R _12206_ (.A(_02600_),
    .Y(net313));
 INVx2_ASAP7_75t_R _12207_ (.A(_02601_),
    .Y(net314));
 INVx2_ASAP7_75t_R _12208_ (.A(_02602_),
    .Y(net315));
 INVx1_ASAP7_75t_R _12209_ (.A(_02603_),
    .Y(net316));
 INVx2_ASAP7_75t_R _12210_ (.A(_02604_),
    .Y(net317));
 INVx2_ASAP7_75t_R _12211_ (.A(_02605_),
    .Y(net319));
 INVx2_ASAP7_75t_R _12212_ (.A(_02606_),
    .Y(net320));
 INVx2_ASAP7_75t_R _12213_ (.A(_02607_),
    .Y(net321));
 INVx2_ASAP7_75t_R _12214_ (.A(_02608_),
    .Y(net322));
 INVx2_ASAP7_75t_R _12215_ (.A(_02609_),
    .Y(net323));
 INVx2_ASAP7_75t_R _12216_ (.A(_02610_),
    .Y(net324));
 INVx8_ASAP7_75t_R _12217_ (.A(net21),
    .Y(_08526_));
 BUFx12f_ASAP7_75t_R _12218_ (.A(_08526_),
    .Y(_08527_));
 BUFx12f_ASAP7_75t_R _12219_ (.A(_08527_),
    .Y(_08528_));
 BUFx12f_ASAP7_75t_R _12220_ (.A(_08528_),
    .Y(_08529_));
 AND2x2_ASAP7_75t_R _12221_ (.A(_08529_),
    .B(_00000_),
    .Y(_02675_));
 BUFx6f_ASAP7_75t_R _12222_ (.A(_01994_),
    .Y(_08530_));
 BUFx6f_ASAP7_75t_R _12223_ (.A(_01995_),
    .Y(_08531_));
 INVx1_ASAP7_75t_R _12224_ (.A(_08531_),
    .Y(_08532_));
 INVx2_ASAP7_75t_R _12225_ (.A(_02000_),
    .Y(_08533_));
 INVx1_ASAP7_75t_R _12226_ (.A(_00897_),
    .Y(_08534_));
 AND4x1_ASAP7_75t_R _12227_ (.A(_00899_),
    .B(_00900_),
    .C(_00901_),
    .D(_00902_),
    .Y(_08535_));
 AND3x4_ASAP7_75t_R _12228_ (.A(_08534_),
    .B(_00903_),
    .C(_08535_),
    .Y(_08536_));
 AND4x1_ASAP7_75t_R _12229_ (.A(_01627_),
    .B(_01628_),
    .C(_01629_),
    .D(_01630_),
    .Y(_08537_));
 BUFx6f_ASAP7_75t_R _12230_ (.A(_08537_),
    .Y(_08538_));
 BUFx6f_ASAP7_75t_R _12231_ (.A(_01625_),
    .Y(_08539_));
 NOR2x1_ASAP7_75t_R _12232_ (.A(_08539_),
    .B(_01631_),
    .Y(_08540_));
 NOR2x1_ASAP7_75t_R _12233_ (.A(_08539_),
    .B(_01626_),
    .Y(_08541_));
 AO21x1_ASAP7_75t_R _12234_ (.A1(_08538_),
    .A2(_08540_),
    .B(_08541_),
    .Y(_08542_));
 OR2x6_ASAP7_75t_R _12235_ (.A(_08539_),
    .B(_01626_),
    .Y(_08543_));
 OR3x1_ASAP7_75t_R _12236_ (.A(_00897_),
    .B(_00898_),
    .C(_02000_),
    .Y(_08544_));
 OAI21x1_ASAP7_75t_R _12237_ (.A1(_08533_),
    .A2(_08543_),
    .B(_08544_),
    .Y(_08545_));
 AO21x1_ASAP7_75t_R _12238_ (.A1(_08536_),
    .A2(_08542_),
    .B(_08545_),
    .Y(_08546_));
 INVx1_ASAP7_75t_R _12239_ (.A(_00898_),
    .Y(_08547_));
 AND2x2_ASAP7_75t_R _12240_ (.A(_08538_),
    .B(_08540_),
    .Y(_08548_));
 OR2x6_ASAP7_75t_R _12241_ (.A(_08539_),
    .B(_08538_),
    .Y(_08549_));
 AO32x1_ASAP7_75t_R _12242_ (.A1(_08534_),
    .A2(_08547_),
    .A3(_08548_),
    .B1(_08536_),
    .B2(_08549_),
    .Y(_08550_));
 OR5x1_ASAP7_75t_R _12243_ (.A(_08530_),
    .B(_08532_),
    .C(_08533_),
    .D(_08546_),
    .E(_08550_),
    .Y(_08551_));
 NOR2x1_ASAP7_75t_R _12244_ (.A(_00897_),
    .B(_00898_),
    .Y(_08552_));
 AO21x1_ASAP7_75t_R _12245_ (.A1(_08531_),
    .A2(_08533_),
    .B(_08530_),
    .Y(_08553_));
 OA21x2_ASAP7_75t_R _12246_ (.A1(_08549_),
    .A2(_08553_),
    .B(_08543_),
    .Y(_08554_));
 OA21x2_ASAP7_75t_R _12247_ (.A1(_08552_),
    .A2(_08554_),
    .B(_08536_),
    .Y(_08555_));
 NOR2x1_ASAP7_75t_R _12248_ (.A(_08551_),
    .B(_08555_),
    .Y(_08556_));
 BUFx6f_ASAP7_75t_R _12249_ (.A(_08556_),
    .Y(_08557_));
 INVx1_ASAP7_75t_R _12250_ (.A(_08530_),
    .Y(_08558_));
 AO221x1_ASAP7_75t_R _12251_ (.A1(_08558_),
    .A2(_02000_),
    .B1(_08535_),
    .B2(_00898_),
    .C(_00897_),
    .Y(_08559_));
 OR3x1_ASAP7_75t_R _12252_ (.A(_00897_),
    .B(_00000_),
    .C(_08535_),
    .Y(_08560_));
 AO22x2_ASAP7_75t_R _12253_ (.A1(_08531_),
    .A2(_08559_),
    .B1(_08560_),
    .B2(_08530_),
    .Y(_08561_));
 OR2x6_ASAP7_75t_R _12254_ (.A(_00897_),
    .B(_08535_),
    .Y(_08562_));
 AO21x1_ASAP7_75t_R _12255_ (.A1(_08531_),
    .A2(_02000_),
    .B(_08530_),
    .Y(_08563_));
 OR2x2_ASAP7_75t_R _12256_ (.A(_00897_),
    .B(_00898_),
    .Y(_08564_));
 OA21x2_ASAP7_75t_R _12257_ (.A1(_08562_),
    .A2(_08563_),
    .B(_08564_),
    .Y(_08565_));
 NAND2x1_ASAP7_75t_R _12258_ (.A(_08538_),
    .B(_08540_),
    .Y(_08566_));
 OA22x2_ASAP7_75t_R _12259_ (.A1(_08549_),
    .A2(_08561_),
    .B1(_08565_),
    .B2(_08566_),
    .Y(_08567_));
 AND3x4_ASAP7_75t_R _12260_ (.A(_08543_),
    .B(_08567_),
    .C(_08555_),
    .Y(_08568_));
 NOR2x1_ASAP7_75t_R _12261_ (.A(_08556_),
    .B(_08568_),
    .Y(_08569_));
 BUFx6f_ASAP7_75t_R _12262_ (.A(_08569_),
    .Y(_08570_));
 BUFx12f_ASAP7_75t_R _12263_ (.A(net21),
    .Y(_08571_));
 BUFx12f_ASAP7_75t_R _12264_ (.A(_08571_),
    .Y(_08572_));
 BUFx12f_ASAP7_75t_R _12265_ (.A(_08572_),
    .Y(_08573_));
 AO21x1_ASAP7_75t_R _12266_ (.A1(_00908_),
    .A2(_08568_),
    .B(_08573_),
    .Y(_08574_));
 AOI221x1_ASAP7_75t_R _12267_ (.A1(_02005_),
    .A2(_08557_),
    .B1(_08570_),
    .B2(_01636_),
    .C(_08574_),
    .Y(_02676_));
 AO21x1_ASAP7_75t_R _12268_ (.A1(_00907_),
    .A2(_08568_),
    .B(_08573_),
    .Y(_08575_));
 AOI221x1_ASAP7_75t_R _12269_ (.A1(_02004_),
    .A2(_08557_),
    .B1(_08570_),
    .B2(_01635_),
    .C(_08575_),
    .Y(_02677_));
 AO21x1_ASAP7_75t_R _12270_ (.A1(_00906_),
    .A2(_08568_),
    .B(_08573_),
    .Y(_08576_));
 AOI221x1_ASAP7_75t_R _12271_ (.A1(_02003_),
    .A2(_08557_),
    .B1(_08570_),
    .B2(_01634_),
    .C(_08576_),
    .Y(_02678_));
 AO21x1_ASAP7_75t_R _12272_ (.A1(_00905_),
    .A2(_08568_),
    .B(_08573_),
    .Y(_08577_));
 AOI221x1_ASAP7_75t_R _12273_ (.A1(_02002_),
    .A2(_08557_),
    .B1(_08570_),
    .B2(_01633_),
    .C(_08577_),
    .Y(_02679_));
 BUFx12f_ASAP7_75t_R _12274_ (.A(_08571_),
    .Y(_08578_));
 BUFx6f_ASAP7_75t_R _12275_ (.A(_08578_),
    .Y(_08579_));
 AO21x1_ASAP7_75t_R _12276_ (.A1(_00904_),
    .A2(_08568_),
    .B(_08579_),
    .Y(_08580_));
 AOI221x1_ASAP7_75t_R _12277_ (.A1(_02001_),
    .A2(_08557_),
    .B1(_08570_),
    .B2(_01632_),
    .C(_08580_),
    .Y(_02680_));
 BUFx12f_ASAP7_75t_R _12278_ (.A(_08527_),
    .Y(_08581_));
 BUFx12f_ASAP7_75t_R _12279_ (.A(_08581_),
    .Y(_08582_));
 INVx2_ASAP7_75t_R _12280_ (.A(_01631_),
    .Y(_08583_));
 AND3x1_ASAP7_75t_R _12281_ (.A(_08582_),
    .B(_08583_),
    .C(_08570_),
    .Y(_02681_));
 BUFx12f_ASAP7_75t_R _12282_ (.A(_08527_),
    .Y(_08584_));
 BUFx12f_ASAP7_75t_R _12283_ (.A(_08584_),
    .Y(_08585_));
 INVx1_ASAP7_75t_R _12284_ (.A(_01630_),
    .Y(_08586_));
 BUFx12f_ASAP7_75t_R _12285_ (.A(_08578_),
    .Y(_08587_));
 NOR2x1_ASAP7_75t_R _12286_ (.A(_08587_),
    .B(_01999_),
    .Y(_08588_));
 AO32x1_ASAP7_75t_R _12287_ (.A1(_08585_),
    .A2(_08586_),
    .A3(_08570_),
    .B1(_08588_),
    .B2(_08557_),
    .Y(_02682_));
 INVx1_ASAP7_75t_R _12288_ (.A(_01629_),
    .Y(_08589_));
 NOR2x1_ASAP7_75t_R _12289_ (.A(_08587_),
    .B(_01998_),
    .Y(_08590_));
 AO32x1_ASAP7_75t_R _12290_ (.A1(_08585_),
    .A2(_08589_),
    .A3(_08570_),
    .B1(_08590_),
    .B2(_08557_),
    .Y(_02683_));
 INVx1_ASAP7_75t_R _12291_ (.A(_01628_),
    .Y(_08591_));
 NOR2x1_ASAP7_75t_R _12292_ (.A(_08587_),
    .B(_01997_),
    .Y(_08592_));
 AO32x1_ASAP7_75t_R _12293_ (.A1(_08585_),
    .A2(_08591_),
    .A3(_08569_),
    .B1(_08592_),
    .B2(_08557_),
    .Y(_02684_));
 INVx1_ASAP7_75t_R _12294_ (.A(_01627_),
    .Y(_08593_));
 NOR2x1_ASAP7_75t_R _12295_ (.A(_08587_),
    .B(_01996_),
    .Y(_08594_));
 AO32x1_ASAP7_75t_R _12296_ (.A1(_08585_),
    .A2(_08593_),
    .A3(_08569_),
    .B1(_08594_),
    .B2(_08556_),
    .Y(_02685_));
 OAI22x1_ASAP7_75t_R _12297_ (.A1(_08549_),
    .A2(_08561_),
    .B1(_08565_),
    .B2(_08566_),
    .Y(_08595_));
 AND3x1_ASAP7_75t_R _12298_ (.A(_08582_),
    .B(_08543_),
    .C(_08595_),
    .Y(_02686_));
 INVx1_ASAP7_75t_R _12299_ (.A(_08551_),
    .Y(_08596_));
 OR3x1_ASAP7_75t_R _12300_ (.A(_08541_),
    .B(_08595_),
    .C(_08555_),
    .Y(_08597_));
 BUFx12f_ASAP7_75t_R _12301_ (.A(_08526_),
    .Y(_08598_));
 BUFx12f_ASAP7_75t_R _12302_ (.A(_08598_),
    .Y(_08599_));
 BUFx6f_ASAP7_75t_R _12303_ (.A(_08599_),
    .Y(_08600_));
 OA21x2_ASAP7_75t_R _12304_ (.A1(_08596_),
    .A2(_08597_),
    .B(_08600_),
    .Y(_02687_));
 AO21x1_ASAP7_75t_R _12305_ (.A1(_00896_),
    .A2(_08568_),
    .B(_08579_),
    .Y(_08601_));
 AOI221x1_ASAP7_75t_R _12306_ (.A1(_01993_),
    .A2(_08557_),
    .B1(_08570_),
    .B2(_01624_),
    .C(_08601_),
    .Y(_02688_));
 AO21x1_ASAP7_75t_R _12307_ (.A1(_00895_),
    .A2(_08568_),
    .B(_08579_),
    .Y(_08602_));
 AOI221x1_ASAP7_75t_R _12308_ (.A1(_01992_),
    .A2(_08557_),
    .B1(_08570_),
    .B2(_01623_),
    .C(_08602_),
    .Y(_02689_));
 OAI21x1_ASAP7_75t_R _12309_ (.A1(_08549_),
    .A2(_08553_),
    .B(_08543_),
    .Y(_08603_));
 AO221x1_ASAP7_75t_R _12310_ (.A1(_08558_),
    .A2(_08533_),
    .B1(_08538_),
    .B2(_01626_),
    .C(_08539_),
    .Y(_08604_));
 INVx1_ASAP7_75t_R _12311_ (.A(_00000_),
    .Y(_08605_));
 OA31x2_ASAP7_75t_R _12312_ (.A1(_08539_),
    .A2(_08605_),
    .A3(_08538_),
    .B1(_08530_),
    .Y(_08606_));
 AOI211x1_ASAP7_75t_R _12313_ (.A1(_08531_),
    .A2(_08604_),
    .B(_08606_),
    .C(_08562_),
    .Y(_08607_));
 AO221x1_ASAP7_75t_R _12314_ (.A1(_08534_),
    .A2(_08547_),
    .B1(_08536_),
    .B2(_08603_),
    .C(_08607_),
    .Y(_08608_));
 BUFx6f_ASAP7_75t_R _12315_ (.A(_08608_),
    .Y(_08609_));
 OA21x2_ASAP7_75t_R _12316_ (.A1(_08541_),
    .A2(_08565_),
    .B(_08548_),
    .Y(_08610_));
 AND3x1_ASAP7_75t_R _12317_ (.A(_08533_),
    .B(_08548_),
    .C(_08562_),
    .Y(_08611_));
 AO211x2_ASAP7_75t_R _12318_ (.A1(_08536_),
    .A2(_08542_),
    .B(_08545_),
    .C(_08532_),
    .Y(_08612_));
 OR4x1_ASAP7_75t_R _12319_ (.A(_08530_),
    .B(_02000_),
    .C(_08611_),
    .D(_08612_),
    .Y(_08613_));
 OR3x2_ASAP7_75t_R _12320_ (.A(_08609_),
    .B(_08610_),
    .C(_08613_),
    .Y(_08614_));
 BUFx12f_ASAP7_75t_R _12321_ (.A(_08614_),
    .Y(_08615_));
 NOR2x1_ASAP7_75t_R _12322_ (.A(_02005_),
    .B(_08615_),
    .Y(_08616_));
 INVx1_ASAP7_75t_R _12323_ (.A(_01636_),
    .Y(_08617_));
 BUFx6f_ASAP7_75t_R _12324_ (.A(_08609_),
    .Y(_08618_));
 BUFx6f_ASAP7_75t_R _12325_ (.A(_08614_),
    .Y(_08619_));
 BUFx6f_ASAP7_75t_R _12326_ (.A(_08609_),
    .Y(_08620_));
 NAND2x1_ASAP7_75t_R _12327_ (.A(_00908_),
    .B(_08620_),
    .Y(_08621_));
 OA211x2_ASAP7_75t_R _12328_ (.A1(_08617_),
    .A2(_08618_),
    .B(_08619_),
    .C(_08621_),
    .Y(_08622_));
 OA21x2_ASAP7_75t_R _12329_ (.A1(_08616_),
    .A2(_08622_),
    .B(_08600_),
    .Y(_02690_));
 NOR2x1_ASAP7_75t_R _12330_ (.A(_02004_),
    .B(_08615_),
    .Y(_08623_));
 INVx1_ASAP7_75t_R _12331_ (.A(_01635_),
    .Y(_08624_));
 NAND2x1_ASAP7_75t_R _12332_ (.A(_00907_),
    .B(_08620_),
    .Y(_08625_));
 OA211x2_ASAP7_75t_R _12333_ (.A1(_08624_),
    .A2(_08618_),
    .B(_08619_),
    .C(_08625_),
    .Y(_08626_));
 OA21x2_ASAP7_75t_R _12334_ (.A1(_08623_),
    .A2(_08626_),
    .B(_08600_),
    .Y(_02691_));
 NOR2x1_ASAP7_75t_R _12335_ (.A(_02003_),
    .B(_08615_),
    .Y(_08627_));
 INVx1_ASAP7_75t_R _12336_ (.A(_01634_),
    .Y(_08628_));
 NAND2x1_ASAP7_75t_R _12337_ (.A(_00906_),
    .B(_08620_),
    .Y(_08629_));
 OA211x2_ASAP7_75t_R _12338_ (.A1(_08628_),
    .A2(_08618_),
    .B(_08619_),
    .C(_08629_),
    .Y(_08630_));
 OA21x2_ASAP7_75t_R _12339_ (.A1(_08627_),
    .A2(_08630_),
    .B(_08600_),
    .Y(_02692_));
 NOR2x1_ASAP7_75t_R _12340_ (.A(_02002_),
    .B(_08615_),
    .Y(_08631_));
 INVx1_ASAP7_75t_R _12341_ (.A(_01633_),
    .Y(_08632_));
 NAND2x1_ASAP7_75t_R _12342_ (.A(_00905_),
    .B(_08620_),
    .Y(_08633_));
 OA211x2_ASAP7_75t_R _12343_ (.A1(_08632_),
    .A2(_08618_),
    .B(_08619_),
    .C(_08633_),
    .Y(_08634_));
 OA21x2_ASAP7_75t_R _12344_ (.A1(_08631_),
    .A2(_08634_),
    .B(_08600_),
    .Y(_02693_));
 NOR2x1_ASAP7_75t_R _12345_ (.A(_02001_),
    .B(_08615_),
    .Y(_08635_));
 INVx1_ASAP7_75t_R _12346_ (.A(_01632_),
    .Y(_08636_));
 NAND2x1_ASAP7_75t_R _12347_ (.A(_00904_),
    .B(_08620_),
    .Y(_08637_));
 OA211x2_ASAP7_75t_R _12348_ (.A1(_08636_),
    .A2(_08618_),
    .B(_08619_),
    .C(_08637_),
    .Y(_08638_));
 OA21x2_ASAP7_75t_R _12349_ (.A1(_08635_),
    .A2(_08638_),
    .B(_08600_),
    .Y(_02694_));
 NOR2x1_ASAP7_75t_R _12350_ (.A(_08583_),
    .B(_08618_),
    .Y(_08639_));
 AO21x1_ASAP7_75t_R _12351_ (.A1(_00903_),
    .A2(_08618_),
    .B(_08639_),
    .Y(_08640_));
 BUFx12f_ASAP7_75t_R _12352_ (.A(_08571_),
    .Y(_08641_));
 BUFx12f_ASAP7_75t_R _12353_ (.A(_08641_),
    .Y(_08642_));
 BUFx12f_ASAP7_75t_R _12354_ (.A(_08642_),
    .Y(_08643_));
 AOI21x1_ASAP7_75t_R _12355_ (.A1(_08615_),
    .A2(_08640_),
    .B(_08643_),
    .Y(_02695_));
 NOR2x1_ASAP7_75t_R _12356_ (.A(_01999_),
    .B(_08615_),
    .Y(_08644_));
 NAND2x1_ASAP7_75t_R _12357_ (.A(_00902_),
    .B(_08620_),
    .Y(_08645_));
 OA211x2_ASAP7_75t_R _12358_ (.A1(_08586_),
    .A2(_08618_),
    .B(_08619_),
    .C(_08645_),
    .Y(_08646_));
 OA21x2_ASAP7_75t_R _12359_ (.A1(_08644_),
    .A2(_08646_),
    .B(_08600_),
    .Y(_02696_));
 NOR2x1_ASAP7_75t_R _12360_ (.A(_01998_),
    .B(_08615_),
    .Y(_08647_));
 NAND2x1_ASAP7_75t_R _12361_ (.A(_00901_),
    .B(_08609_),
    .Y(_08648_));
 OA211x2_ASAP7_75t_R _12362_ (.A1(_08589_),
    .A2(_08618_),
    .B(_08619_),
    .C(_08648_),
    .Y(_08649_));
 OA21x2_ASAP7_75t_R _12363_ (.A1(_08647_),
    .A2(_08649_),
    .B(_08600_),
    .Y(_02697_));
 NOR2x1_ASAP7_75t_R _12364_ (.A(_01997_),
    .B(_08615_),
    .Y(_08650_));
 NAND2x1_ASAP7_75t_R _12365_ (.A(_00900_),
    .B(_08609_),
    .Y(_08651_));
 OA211x2_ASAP7_75t_R _12366_ (.A1(_08591_),
    .A2(_08620_),
    .B(_08619_),
    .C(_08651_),
    .Y(_08652_));
 OA21x2_ASAP7_75t_R _12367_ (.A1(_08650_),
    .A2(_08652_),
    .B(_08600_),
    .Y(_02698_));
 NOR2x1_ASAP7_75t_R _12368_ (.A(_01996_),
    .B(_08615_),
    .Y(_08653_));
 NAND2x1_ASAP7_75t_R _12369_ (.A(_00899_),
    .B(_08609_),
    .Y(_08654_));
 OA211x2_ASAP7_75t_R _12370_ (.A1(_08593_),
    .A2(_08620_),
    .B(_08614_),
    .C(_08654_),
    .Y(_08655_));
 OA21x2_ASAP7_75t_R _12371_ (.A1(_08653_),
    .A2(_08655_),
    .B(_08600_),
    .Y(_02699_));
 BUFx12f_ASAP7_75t_R _12372_ (.A(_08571_),
    .Y(_08656_));
 BUFx12f_ASAP7_75t_R _12373_ (.A(_08656_),
    .Y(_08657_));
 AOI21x1_ASAP7_75t_R _12374_ (.A1(_08536_),
    .A2(_08603_),
    .B(_08607_),
    .Y(_08658_));
 OR3x1_ASAP7_75t_R _12375_ (.A(_08657_),
    .B(_08552_),
    .C(_08658_),
    .Y(_08659_));
 INVx1_ASAP7_75t_R _12376_ (.A(_08659_),
    .Y(_02700_));
 NOR2x1_ASAP7_75t_R _12377_ (.A(_08618_),
    .B(_08610_),
    .Y(_08660_));
 AOI21x1_ASAP7_75t_R _12378_ (.A1(_08660_),
    .A2(_08613_),
    .B(_08643_),
    .Y(_02701_));
 NOR2x1_ASAP7_75t_R _12379_ (.A(_01993_),
    .B(_08619_),
    .Y(_08661_));
 INVx1_ASAP7_75t_R _12380_ (.A(_01624_),
    .Y(_08662_));
 NAND2x1_ASAP7_75t_R _12381_ (.A(_00896_),
    .B(_08609_),
    .Y(_08663_));
 OA211x2_ASAP7_75t_R _12382_ (.A1(_08662_),
    .A2(_08620_),
    .B(_08614_),
    .C(_08663_),
    .Y(_08664_));
 BUFx12f_ASAP7_75t_R _12383_ (.A(_08598_),
    .Y(_08665_));
 BUFx6f_ASAP7_75t_R _12384_ (.A(_08665_),
    .Y(_08666_));
 OA21x2_ASAP7_75t_R _12385_ (.A1(_08661_),
    .A2(_08664_),
    .B(_08666_),
    .Y(_02702_));
 NOR2x1_ASAP7_75t_R _12386_ (.A(_01992_),
    .B(_08619_),
    .Y(_08667_));
 INVx1_ASAP7_75t_R _12387_ (.A(_01623_),
    .Y(_08668_));
 NAND2x1_ASAP7_75t_R _12388_ (.A(_00895_),
    .B(_08609_),
    .Y(_08669_));
 OA211x2_ASAP7_75t_R _12389_ (.A1(_08668_),
    .A2(_08620_),
    .B(_08614_),
    .C(_08669_),
    .Y(_08670_));
 OA21x2_ASAP7_75t_R _12390_ (.A1(_08667_),
    .A2(_08670_),
    .B(_08666_),
    .Y(_02703_));
 NOR2x1_ASAP7_75t_R _12391_ (.A(_08539_),
    .B(_08538_),
    .Y(_08671_));
 OR2x6_ASAP7_75t_R _12392_ (.A(_08541_),
    .B(_08561_),
    .Y(_08672_));
 AOI21x1_ASAP7_75t_R _12393_ (.A1(_08531_),
    .A2(_08604_),
    .B(_08606_),
    .Y(_08673_));
 AO21x1_ASAP7_75t_R _12394_ (.A1(_08564_),
    .A2(_08673_),
    .B(_08562_),
    .Y(_08674_));
 AOI21x1_ASAP7_75t_R _12395_ (.A1(_08671_),
    .A2(_08672_),
    .B(_08674_),
    .Y(_08675_));
 BUFx6f_ASAP7_75t_R _12396_ (.A(_08675_),
    .Y(_08676_));
 NAND2x1_ASAP7_75t_R _12397_ (.A(_00908_),
    .B(_08676_),
    .Y(_08677_));
 BUFx6f_ASAP7_75t_R _12398_ (.A(_08675_),
    .Y(_08678_));
 OR2x2_ASAP7_75t_R _12399_ (.A(_08617_),
    .B(_08678_),
    .Y(_08679_));
 AOI211x1_ASAP7_75t_R _12400_ (.A1(_02000_),
    .A2(_08550_),
    .B(_08611_),
    .C(_08546_),
    .Y(_08680_));
 AOI21x1_ASAP7_75t_R _12401_ (.A1(_08531_),
    .A2(_08680_),
    .B(_08530_),
    .Y(_08681_));
 NOR2x1_ASAP7_75t_R _12402_ (.A(_08572_),
    .B(_08681_),
    .Y(_08682_));
 BUFx12f_ASAP7_75t_R _12403_ (.A(net21),
    .Y(_08683_));
 BUFx12f_ASAP7_75t_R _12404_ (.A(_08683_),
    .Y(_08684_));
 NOR2x1_ASAP7_75t_R _12405_ (.A(_08684_),
    .B(_02005_),
    .Y(_08685_));
 BUFx3_ASAP7_75t_R _12406_ (.A(_08681_),
    .Y(_08686_));
 AO32x1_ASAP7_75t_R _12407_ (.A1(_08677_),
    .A2(_08679_),
    .A3(_08682_),
    .B1(_08685_),
    .B2(_08686_),
    .Y(_02704_));
 BUFx6f_ASAP7_75t_R _12408_ (.A(_08682_),
    .Y(_08687_));
 NAND2x1_ASAP7_75t_R _12409_ (.A(_00907_),
    .B(_08676_),
    .Y(_08688_));
 OR2x2_ASAP7_75t_R _12410_ (.A(_08624_),
    .B(_08678_),
    .Y(_08689_));
 NOR2x1_ASAP7_75t_R _12411_ (.A(_08684_),
    .B(_02004_),
    .Y(_08690_));
 AO32x1_ASAP7_75t_R _12412_ (.A1(_08687_),
    .A2(_08688_),
    .A3(_08689_),
    .B1(_08690_),
    .B2(_08686_),
    .Y(_02705_));
 NAND2x1_ASAP7_75t_R _12413_ (.A(_00906_),
    .B(_08676_),
    .Y(_08691_));
 OR2x2_ASAP7_75t_R _12414_ (.A(_08628_),
    .B(_08678_),
    .Y(_08692_));
 NOR2x1_ASAP7_75t_R _12415_ (.A(_08684_),
    .B(_02003_),
    .Y(_08693_));
 AO32x1_ASAP7_75t_R _12416_ (.A1(_08687_),
    .A2(_08691_),
    .A3(_08692_),
    .B1(_08693_),
    .B2(_08686_),
    .Y(_02706_));
 NAND2x1_ASAP7_75t_R _12417_ (.A(_00905_),
    .B(_08676_),
    .Y(_08694_));
 OR2x2_ASAP7_75t_R _12418_ (.A(_08632_),
    .B(_08678_),
    .Y(_08695_));
 BUFx12f_ASAP7_75t_R _12419_ (.A(_08656_),
    .Y(_08696_));
 NOR2x1_ASAP7_75t_R _12420_ (.A(_08696_),
    .B(_02002_),
    .Y(_08697_));
 AO32x1_ASAP7_75t_R _12421_ (.A1(_08687_),
    .A2(_08694_),
    .A3(_08695_),
    .B1(_08697_),
    .B2(_08686_),
    .Y(_02707_));
 NAND2x1_ASAP7_75t_R _12422_ (.A(_00904_),
    .B(_08676_),
    .Y(_08698_));
 OR2x2_ASAP7_75t_R _12423_ (.A(_08636_),
    .B(_08678_),
    .Y(_08699_));
 NOR2x1_ASAP7_75t_R _12424_ (.A(_08696_),
    .B(_02001_),
    .Y(_08700_));
 AO32x1_ASAP7_75t_R _12425_ (.A1(_08687_),
    .A2(_08698_),
    .A3(_08699_),
    .B1(_08700_),
    .B2(_08686_),
    .Y(_02708_));
 NAND2x1_ASAP7_75t_R _12426_ (.A(_00903_),
    .B(_08676_),
    .Y(_08701_));
 OR2x2_ASAP7_75t_R _12427_ (.A(_08583_),
    .B(_08678_),
    .Y(_08702_));
 NOR2x1_ASAP7_75t_R _12428_ (.A(_08696_),
    .B(_02000_),
    .Y(_08703_));
 AO32x1_ASAP7_75t_R _12429_ (.A1(_08687_),
    .A2(_08701_),
    .A3(_08702_),
    .B1(_08703_),
    .B2(_08686_),
    .Y(_02709_));
 NAND2x1_ASAP7_75t_R _12430_ (.A(_00902_),
    .B(_08676_),
    .Y(_08704_));
 OR2x2_ASAP7_75t_R _12431_ (.A(_08586_),
    .B(_08678_),
    .Y(_08705_));
 AO32x1_ASAP7_75t_R _12432_ (.A1(_08687_),
    .A2(_08704_),
    .A3(_08705_),
    .B1(_08686_),
    .B2(_08588_),
    .Y(_02710_));
 NAND2x1_ASAP7_75t_R _12433_ (.A(_00901_),
    .B(_08676_),
    .Y(_08706_));
 OR2x2_ASAP7_75t_R _12434_ (.A(_08589_),
    .B(_08678_),
    .Y(_08707_));
 AO32x1_ASAP7_75t_R _12435_ (.A1(_08687_),
    .A2(_08706_),
    .A3(_08707_),
    .B1(_08681_),
    .B2(_08590_),
    .Y(_02711_));
 NAND2x1_ASAP7_75t_R _12436_ (.A(_00900_),
    .B(_08676_),
    .Y(_08708_));
 OR2x2_ASAP7_75t_R _12437_ (.A(_08591_),
    .B(_08675_),
    .Y(_08709_));
 AO32x1_ASAP7_75t_R _12438_ (.A1(_08687_),
    .A2(_08708_),
    .A3(_08709_),
    .B1(_08681_),
    .B2(_08592_),
    .Y(_02712_));
 NAND2x1_ASAP7_75t_R _12439_ (.A(_00899_),
    .B(_08676_),
    .Y(_08710_));
 OR2x2_ASAP7_75t_R _12440_ (.A(_08593_),
    .B(_08675_),
    .Y(_08711_));
 AO32x1_ASAP7_75t_R _12441_ (.A1(_08687_),
    .A2(_08710_),
    .A3(_08711_),
    .B1(_08681_),
    .B2(_08594_),
    .Y(_02713_));
 BUFx12f_ASAP7_75t_R _12442_ (.A(_08572_),
    .Y(_08712_));
 OR4x1_ASAP7_75t_R _12443_ (.A(_08712_),
    .B(_08530_),
    .C(_08532_),
    .D(_08680_),
    .Y(_08713_));
 INVx1_ASAP7_75t_R _12444_ (.A(_08713_),
    .Y(_02714_));
 NAND2x1_ASAP7_75t_R _12445_ (.A(_08671_),
    .B(_08672_),
    .Y(_08714_));
 NAND2x1_ASAP7_75t_R _12446_ (.A(_08674_),
    .B(_08714_),
    .Y(_08715_));
 OA21x2_ASAP7_75t_R _12447_ (.A1(_08686_),
    .A2(_08715_),
    .B(_08666_),
    .Y(_02715_));
 NAND2x1_ASAP7_75t_R _12448_ (.A(_00896_),
    .B(_08678_),
    .Y(_08716_));
 OR2x2_ASAP7_75t_R _12449_ (.A(_08662_),
    .B(_08675_),
    .Y(_08717_));
 NOR2x1_ASAP7_75t_R _12450_ (.A(_08696_),
    .B(_01993_),
    .Y(_08718_));
 AO32x1_ASAP7_75t_R _12451_ (.A1(_08687_),
    .A2(_08716_),
    .A3(_08717_),
    .B1(_08718_),
    .B2(_08686_),
    .Y(_02716_));
 NAND2x1_ASAP7_75t_R _12452_ (.A(_00895_),
    .B(_08678_),
    .Y(_08719_));
 OR2x2_ASAP7_75t_R _12453_ (.A(_08668_),
    .B(_08675_),
    .Y(_08720_));
 NOR2x1_ASAP7_75t_R _12454_ (.A(_08696_),
    .B(_01992_),
    .Y(_08721_));
 AO32x1_ASAP7_75t_R _12455_ (.A1(_08682_),
    .A2(_08719_),
    .A3(_08720_),
    .B1(_08721_),
    .B2(_08686_),
    .Y(_02717_));
 BUFx12f_ASAP7_75t_R _12456_ (.A(_08527_),
    .Y(_08722_));
 BUFx12f_ASAP7_75t_R _12457_ (.A(_08722_),
    .Y(_08723_));
 AND2x2_ASAP7_75t_R _12458_ (.A(_08723_),
    .B(_00001_),
    .Y(_02718_));
 INVx1_ASAP7_75t_R _12459_ (.A(_00793_),
    .Y(_08724_));
 INVx2_ASAP7_75t_R _12460_ (.A(_00797_),
    .Y(_08725_));
 NAND2x1_ASAP7_75t_R _12461_ (.A(_00795_),
    .B(_00796_),
    .Y(_08726_));
 OR3x2_ASAP7_75t_R _12462_ (.A(_08725_),
    .B(_00798_),
    .C(_08726_),
    .Y(_08727_));
 NAND2x1_ASAP7_75t_R _12463_ (.A(_08724_),
    .B(_08727_),
    .Y(_08728_));
 INVx2_ASAP7_75t_R _12464_ (.A(_00693_),
    .Y(_08729_));
 NAND2x1_ASAP7_75t_R _12465_ (.A(_00691_),
    .B(_00692_),
    .Y(_08730_));
 OR3x1_ASAP7_75t_R _12466_ (.A(_08729_),
    .B(_00694_),
    .C(_08730_),
    .Y(_08731_));
 BUFx6f_ASAP7_75t_R _12467_ (.A(_01980_),
    .Y(_08732_));
 BUFx6f_ASAP7_75t_R _12468_ (.A(_01986_),
    .Y(_08733_));
 INVx2_ASAP7_75t_R _12469_ (.A(_08733_),
    .Y(_08734_));
 INVx1_ASAP7_75t_R _12470_ (.A(_00689_),
    .Y(_08735_));
 OA21x2_ASAP7_75t_R _12471_ (.A1(_08732_),
    .A2(_08734_),
    .B(_08735_),
    .Y(_08736_));
 NOR2x1_ASAP7_75t_R _12472_ (.A(_00689_),
    .B(_00690_),
    .Y(_08737_));
 OA21x2_ASAP7_75t_R _12473_ (.A1(_08732_),
    .A2(_08734_),
    .B(_08737_),
    .Y(_08738_));
 BUFx6f_ASAP7_75t_R _12474_ (.A(_01981_),
    .Y(_08739_));
 INVx2_ASAP7_75t_R _12475_ (.A(_08739_),
    .Y(_08740_));
 AOI211x1_ASAP7_75t_R _12476_ (.A1(_08731_),
    .A2(_08736_),
    .B(_08738_),
    .C(_08740_),
    .Y(_08741_));
 INVx1_ASAP7_75t_R _12477_ (.A(_00694_),
    .Y(_08742_));
 AND2x2_ASAP7_75t_R _12478_ (.A(_00691_),
    .B(_00692_),
    .Y(_08743_));
 AO31x2_ASAP7_75t_R _12479_ (.A1(_00693_),
    .A2(_08742_),
    .A3(_08743_),
    .B(_00689_),
    .Y(_08744_));
 OA21x2_ASAP7_75t_R _12480_ (.A1(_00001_),
    .A2(_08744_),
    .B(_08732_),
    .Y(_08745_));
 OR2x2_ASAP7_75t_R _12481_ (.A(_00793_),
    .B(_00799_),
    .Y(_08746_));
 AO21x1_ASAP7_75t_R _12482_ (.A1(_08739_),
    .A2(_08733_),
    .B(_08732_),
    .Y(_08747_));
 OR2x2_ASAP7_75t_R _12483_ (.A(_00689_),
    .B(_00690_),
    .Y(_08748_));
 BUFx6f_ASAP7_75t_R _12484_ (.A(_08748_),
    .Y(_08749_));
 OA21x2_ASAP7_75t_R _12485_ (.A1(_08744_),
    .A2(_08747_),
    .B(_08749_),
    .Y(_08750_));
 OA33x2_ASAP7_75t_R _12486_ (.A1(_08728_),
    .A2(_08741_),
    .A3(_08745_),
    .B1(_08746_),
    .B2(_08750_),
    .B3(_08727_),
    .Y(_08751_));
 NOR2x2_ASAP7_75t_R _12487_ (.A(_00793_),
    .B(_00794_),
    .Y(_08752_));
 INVx1_ASAP7_75t_R _12488_ (.A(_00695_),
    .Y(_08753_));
 OR5x2_ASAP7_75t_R _12489_ (.A(_00689_),
    .B(_08729_),
    .C(_00694_),
    .D(_08753_),
    .E(_08730_),
    .Y(_08754_));
 INVx2_ASAP7_75t_R _12490_ (.A(_08732_),
    .Y(_08755_));
 OA31x2_ASAP7_75t_R _12491_ (.A1(_08725_),
    .A2(_00798_),
    .A3(_08726_),
    .B1(_08724_),
    .Y(_08756_));
 OA21x2_ASAP7_75t_R _12492_ (.A1(_08740_),
    .A2(_08733_),
    .B(_08749_),
    .Y(_08757_));
 AND3x1_ASAP7_75t_R _12493_ (.A(_08755_),
    .B(_08756_),
    .C(_08757_),
    .Y(_08758_));
 NOR3x1_ASAP7_75t_R _12494_ (.A(_08752_),
    .B(_08754_),
    .C(_08758_),
    .Y(_08759_));
 AND2x4_ASAP7_75t_R _12495_ (.A(_08751_),
    .B(_08759_),
    .Y(_08760_));
 BUFx6f_ASAP7_75t_R _12496_ (.A(_08760_),
    .Y(_08761_));
 NAND2x1_ASAP7_75t_R _12497_ (.A(_00700_),
    .B(_08761_),
    .Y(_08762_));
 NAND2x2_ASAP7_75t_R _12498_ (.A(_08751_),
    .B(_08759_),
    .Y(_08763_));
 NAND2x1_ASAP7_75t_R _12499_ (.A(_00804_),
    .B(_08763_),
    .Y(_08764_));
 BUFx12f_ASAP7_75t_R _12500_ (.A(_08571_),
    .Y(_08765_));
 OR2x6_ASAP7_75t_R _12501_ (.A(_00793_),
    .B(_00794_),
    .Y(_08766_));
 OA21x2_ASAP7_75t_R _12502_ (.A1(_08754_),
    .A2(_08758_),
    .B(_08766_),
    .Y(_08767_));
 OA31x2_ASAP7_75t_R _12503_ (.A1(_08729_),
    .A2(_00694_),
    .A3(_08730_),
    .B1(_08735_),
    .Y(_08768_));
 OR4x1_ASAP7_75t_R _12504_ (.A(_08725_),
    .B(_00798_),
    .C(_08726_),
    .D(_08746_),
    .Y(_08769_));
 OA21x2_ASAP7_75t_R _12505_ (.A1(_08768_),
    .A2(_08769_),
    .B(_08734_),
    .Y(_08770_));
 OA211x2_ASAP7_75t_R _12506_ (.A1(_08756_),
    .A2(_08754_),
    .B(_08766_),
    .C(_08733_),
    .Y(_08771_));
 AO21x1_ASAP7_75t_R _12507_ (.A1(_08733_),
    .A2(_08769_),
    .B(_08749_),
    .Y(_08772_));
 AO21x1_ASAP7_75t_R _12508_ (.A1(_08769_),
    .A2(_08766_),
    .B(_08754_),
    .Y(_08773_));
 OA211x2_ASAP7_75t_R _12509_ (.A1(_08770_),
    .A2(_08771_),
    .B(_08772_),
    .C(_08773_),
    .Y(_08774_));
 AND3x1_ASAP7_75t_R _12510_ (.A(_08755_),
    .B(_08739_),
    .C(_08733_),
    .Y(_08775_));
 AND4x1_ASAP7_75t_R _12511_ (.A(_08751_),
    .B(_08767_),
    .C(_08774_),
    .D(_08775_),
    .Y(_08776_));
 BUFx6f_ASAP7_75t_R _12512_ (.A(_08776_),
    .Y(_08777_));
 NOR2x2_ASAP7_75t_R _12513_ (.A(_08765_),
    .B(_08777_),
    .Y(_08778_));
 NOR2x1_ASAP7_75t_R _12514_ (.A(_08696_),
    .B(_01991_),
    .Y(_08779_));
 BUFx6f_ASAP7_75t_R _12515_ (.A(_08777_),
    .Y(_08780_));
 AO32x1_ASAP7_75t_R _12516_ (.A1(_08762_),
    .A2(_08764_),
    .A3(_08778_),
    .B1(_08779_),
    .B2(_08780_),
    .Y(_02719_));
 NAND2x1_ASAP7_75t_R _12517_ (.A(_00699_),
    .B(_08761_),
    .Y(_08781_));
 NAND2x1_ASAP7_75t_R _12518_ (.A(_00803_),
    .B(_08763_),
    .Y(_08782_));
 NOR2x1_ASAP7_75t_R _12519_ (.A(_08696_),
    .B(_01990_),
    .Y(_08783_));
 AO32x1_ASAP7_75t_R _12520_ (.A1(_08778_),
    .A2(_08781_),
    .A3(_08782_),
    .B1(_08783_),
    .B2(_08780_),
    .Y(_02720_));
 NAND2x1_ASAP7_75t_R _12521_ (.A(_00698_),
    .B(_08761_),
    .Y(_08784_));
 NAND2x1_ASAP7_75t_R _12522_ (.A(_00802_),
    .B(_08763_),
    .Y(_08785_));
 NOR2x1_ASAP7_75t_R _12523_ (.A(_08696_),
    .B(_01989_),
    .Y(_08786_));
 AO32x1_ASAP7_75t_R _12524_ (.A1(_08778_),
    .A2(_08784_),
    .A3(_08785_),
    .B1(_08786_),
    .B2(_08780_),
    .Y(_02721_));
 NAND2x1_ASAP7_75t_R _12525_ (.A(_00697_),
    .B(_08761_),
    .Y(_08787_));
 NAND2x1_ASAP7_75t_R _12526_ (.A(_00801_),
    .B(_08763_),
    .Y(_08788_));
 NOR2x1_ASAP7_75t_R _12527_ (.A(_08696_),
    .B(_01988_),
    .Y(_08789_));
 AO32x1_ASAP7_75t_R _12528_ (.A1(_08778_),
    .A2(_08787_),
    .A3(_08788_),
    .B1(_08789_),
    .B2(_08780_),
    .Y(_02722_));
 NAND2x1_ASAP7_75t_R _12529_ (.A(_00696_),
    .B(_08761_),
    .Y(_08790_));
 NAND2x1_ASAP7_75t_R _12530_ (.A(_00800_),
    .B(_08763_),
    .Y(_08791_));
 NOR2x1_ASAP7_75t_R _12531_ (.A(_08696_),
    .B(_01987_),
    .Y(_08792_));
 AO32x1_ASAP7_75t_R _12532_ (.A1(_08778_),
    .A2(_08790_),
    .A3(_08791_),
    .B1(_08792_),
    .B2(_08780_),
    .Y(_02723_));
 OR4x1_ASAP7_75t_R _12533_ (.A(_08712_),
    .B(_00799_),
    .C(_08760_),
    .D(_08777_),
    .Y(_08793_));
 INVx1_ASAP7_75t_R _12534_ (.A(_08793_),
    .Y(_02724_));
 NAND2x1_ASAP7_75t_R _12535_ (.A(_01985_),
    .B(_08777_),
    .Y(_08794_));
 INVx1_ASAP7_75t_R _12536_ (.A(_00798_),
    .Y(_08795_));
 OR3x1_ASAP7_75t_R _12537_ (.A(_08795_),
    .B(_08760_),
    .C(_08777_),
    .Y(_08796_));
 AND3x1_ASAP7_75t_R _12538_ (.A(_08582_),
    .B(_08794_),
    .C(_08796_),
    .Y(_02725_));
 INVx2_ASAP7_75t_R _12539_ (.A(_01984_),
    .Y(_08797_));
 NAND2x1_ASAP7_75t_R _12540_ (.A(_08797_),
    .B(_08780_),
    .Y(_08798_));
 OR3x1_ASAP7_75t_R _12541_ (.A(_00797_),
    .B(_08761_),
    .C(_08777_),
    .Y(_08799_));
 AOI21x1_ASAP7_75t_R _12542_ (.A1(_08798_),
    .A2(_08799_),
    .B(_08643_),
    .Y(_02726_));
 INVx2_ASAP7_75t_R _12543_ (.A(_01983_),
    .Y(_08800_));
 NAND2x1_ASAP7_75t_R _12544_ (.A(_08800_),
    .B(_08780_),
    .Y(_08801_));
 OR3x1_ASAP7_75t_R _12545_ (.A(_00796_),
    .B(_08761_),
    .C(_08777_),
    .Y(_08802_));
 AOI21x1_ASAP7_75t_R _12546_ (.A1(_08801_),
    .A2(_08802_),
    .B(_08643_),
    .Y(_02727_));
 INVx2_ASAP7_75t_R _12547_ (.A(_01982_),
    .Y(_08803_));
 NAND2x1_ASAP7_75t_R _12548_ (.A(_08803_),
    .B(_08780_),
    .Y(_08804_));
 OR3x1_ASAP7_75t_R _12549_ (.A(_00795_),
    .B(_08761_),
    .C(_08777_),
    .Y(_08805_));
 AOI21x1_ASAP7_75t_R _12550_ (.A1(_08804_),
    .A2(_08805_),
    .B(_08643_),
    .Y(_02728_));
 OR3x1_ASAP7_75t_R _12551_ (.A(_08657_),
    .B(_08751_),
    .C(_08752_),
    .Y(_08806_));
 INVx1_ASAP7_75t_R _12552_ (.A(_08806_),
    .Y(_02729_));
 NAND2x1_ASAP7_75t_R _12553_ (.A(_08751_),
    .B(_08767_),
    .Y(_08807_));
 AND2x2_ASAP7_75t_R _12554_ (.A(_08774_),
    .B(_08775_),
    .Y(_08808_));
 OA21x2_ASAP7_75t_R _12555_ (.A1(_08807_),
    .A2(_08808_),
    .B(_08666_),
    .Y(_02730_));
 NAND2x1_ASAP7_75t_R _12556_ (.A(_00688_),
    .B(_08761_),
    .Y(_08809_));
 NAND2x1_ASAP7_75t_R _12557_ (.A(_00792_),
    .B(_08763_),
    .Y(_08810_));
 BUFx12f_ASAP7_75t_R _12558_ (.A(_08656_),
    .Y(_08811_));
 NOR2x1_ASAP7_75t_R _12559_ (.A(_08811_),
    .B(_01979_),
    .Y(_08812_));
 AO32x1_ASAP7_75t_R _12560_ (.A1(_08778_),
    .A2(_08809_),
    .A3(_08810_),
    .B1(_08812_),
    .B2(_08780_),
    .Y(_02731_));
 NAND2x1_ASAP7_75t_R _12561_ (.A(_00687_),
    .B(_08761_),
    .Y(_08813_));
 NAND2x1_ASAP7_75t_R _12562_ (.A(_00791_),
    .B(_08763_),
    .Y(_08814_));
 NOR2x1_ASAP7_75t_R _12563_ (.A(_08811_),
    .B(_01978_),
    .Y(_08815_));
 AO32x1_ASAP7_75t_R _12564_ (.A1(_08778_),
    .A2(_08813_),
    .A3(_08814_),
    .B1(_08815_),
    .B2(_08780_),
    .Y(_02732_));
 INVx1_ASAP7_75t_R _12565_ (.A(_01991_),
    .Y(_08816_));
 AO211x2_ASAP7_75t_R _12566_ (.A1(_08731_),
    .A2(_08736_),
    .B(_08738_),
    .C(_08740_),
    .Y(_08817_));
 INVx1_ASAP7_75t_R _12567_ (.A(_00001_),
    .Y(_08818_));
 AO21x1_ASAP7_75t_R _12568_ (.A1(_08818_),
    .A2(_08768_),
    .B(_08755_),
    .Y(_08819_));
 AND2x2_ASAP7_75t_R _12569_ (.A(_08756_),
    .B(_08766_),
    .Y(_08820_));
 OAI21x1_ASAP7_75t_R _12570_ (.A1(_08744_),
    .A2(_08747_),
    .B(_08749_),
    .Y(_08821_));
 AO32x1_ASAP7_75t_R _12571_ (.A1(_08817_),
    .A2(_08819_),
    .A3(_08820_),
    .B1(_08766_),
    .B2(_08821_),
    .Y(_08822_));
 AND3x1_ASAP7_75t_R _12572_ (.A(_08755_),
    .B(_08739_),
    .C(_08734_),
    .Y(_08823_));
 OA211x2_ASAP7_75t_R _12573_ (.A1(_08769_),
    .A2(_08822_),
    .B(_08823_),
    .C(_08774_),
    .Y(_08824_));
 BUFx6f_ASAP7_75t_R _12574_ (.A(_08824_),
    .Y(_08825_));
 NAND2x1_ASAP7_75t_R _12575_ (.A(_08816_),
    .B(_08825_),
    .Y(_08826_));
 AND5x1_ASAP7_75t_R _12576_ (.A(_08735_),
    .B(_00693_),
    .C(_08742_),
    .D(_00695_),
    .E(_08743_),
    .Y(_08827_));
 OA21x2_ASAP7_75t_R _12577_ (.A1(_08740_),
    .A2(_08733_),
    .B(_08755_),
    .Y(_08828_));
 AO21x1_ASAP7_75t_R _12578_ (.A1(_08756_),
    .A2(_08828_),
    .B(_08752_),
    .Y(_08829_));
 AO21x1_ASAP7_75t_R _12579_ (.A1(_08733_),
    .A2(_08752_),
    .B(_08740_),
    .Y(_08830_));
 AO21x1_ASAP7_75t_R _12580_ (.A1(_08755_),
    .A2(_08830_),
    .B(_08756_),
    .Y(_08831_));
 AOI211x1_ASAP7_75t_R _12581_ (.A1(_08732_),
    .A2(_08818_),
    .B(_08744_),
    .C(_08823_),
    .Y(_08832_));
 AOI22x1_ASAP7_75t_R _12582_ (.A1(_08827_),
    .A2(_08829_),
    .B1(_08831_),
    .B2(_08832_),
    .Y(_08833_));
 NAND2x1_ASAP7_75t_R _12583_ (.A(_08749_),
    .B(_08833_),
    .Y(_08834_));
 BUFx6f_ASAP7_75t_R _12584_ (.A(_08834_),
    .Y(_08835_));
 BUFx6f_ASAP7_75t_R _12585_ (.A(_08749_),
    .Y(_08836_));
 AND2x2_ASAP7_75t_R _12586_ (.A(_00804_),
    .B(_08836_),
    .Y(_08837_));
 BUFx6f_ASAP7_75t_R _12587_ (.A(_08833_),
    .Y(_08838_));
 BUFx6f_ASAP7_75t_R _12588_ (.A(_08824_),
    .Y(_08839_));
 AO221x1_ASAP7_75t_R _12589_ (.A1(_00700_),
    .A2(_08835_),
    .B1(_08837_),
    .B2(_08838_),
    .C(_08839_),
    .Y(_08840_));
 AOI21x1_ASAP7_75t_R _12590_ (.A1(_08826_),
    .A2(_08840_),
    .B(_08643_),
    .Y(_02733_));
 INVx1_ASAP7_75t_R _12591_ (.A(_01990_),
    .Y(_08841_));
 NAND2x1_ASAP7_75t_R _12592_ (.A(_08841_),
    .B(_08825_),
    .Y(_08842_));
 AND2x2_ASAP7_75t_R _12593_ (.A(_00803_),
    .B(_08836_),
    .Y(_08843_));
 AO221x1_ASAP7_75t_R _12594_ (.A1(_00699_),
    .A2(_08835_),
    .B1(_08843_),
    .B2(_08838_),
    .C(_08839_),
    .Y(_08844_));
 AOI21x1_ASAP7_75t_R _12595_ (.A1(_08842_),
    .A2(_08844_),
    .B(_08643_),
    .Y(_02734_));
 INVx1_ASAP7_75t_R _12596_ (.A(_01989_),
    .Y(_08845_));
 NAND2x1_ASAP7_75t_R _12597_ (.A(_08845_),
    .B(_08825_),
    .Y(_08846_));
 AND2x2_ASAP7_75t_R _12598_ (.A(_00802_),
    .B(_08836_),
    .Y(_08847_));
 AO221x1_ASAP7_75t_R _12599_ (.A1(_00698_),
    .A2(_08835_),
    .B1(_08847_),
    .B2(_08838_),
    .C(_08839_),
    .Y(_08848_));
 AOI21x1_ASAP7_75t_R _12600_ (.A1(_08846_),
    .A2(_08848_),
    .B(_08643_),
    .Y(_02735_));
 INVx1_ASAP7_75t_R _12601_ (.A(_01988_),
    .Y(_08849_));
 NAND2x1_ASAP7_75t_R _12602_ (.A(_08849_),
    .B(_08825_),
    .Y(_08850_));
 AND2x2_ASAP7_75t_R _12603_ (.A(_00801_),
    .B(_08836_),
    .Y(_08851_));
 AO221x1_ASAP7_75t_R _12604_ (.A1(_00697_),
    .A2(_08835_),
    .B1(_08851_),
    .B2(_08838_),
    .C(_08839_),
    .Y(_08852_));
 AOI21x1_ASAP7_75t_R _12605_ (.A1(_08850_),
    .A2(_08852_),
    .B(_08643_),
    .Y(_02736_));
 INVx1_ASAP7_75t_R _12606_ (.A(_01987_),
    .Y(_08853_));
 NAND2x1_ASAP7_75t_R _12607_ (.A(_08853_),
    .B(_08825_),
    .Y(_08854_));
 AND2x2_ASAP7_75t_R _12608_ (.A(_00800_),
    .B(_08836_),
    .Y(_08855_));
 AO221x1_ASAP7_75t_R _12609_ (.A1(_00696_),
    .A2(_08835_),
    .B1(_08855_),
    .B2(_08838_),
    .C(_08839_),
    .Y(_08856_));
 AOI21x1_ASAP7_75t_R _12610_ (.A1(_08854_),
    .A2(_08856_),
    .B(_08643_),
    .Y(_02737_));
 AND3x1_ASAP7_75t_R _12611_ (.A(_00799_),
    .B(_08836_),
    .C(_08833_),
    .Y(_08857_));
 AOI21x1_ASAP7_75t_R _12612_ (.A1(_00695_),
    .A2(_08835_),
    .B(_08857_),
    .Y(_08858_));
 OA21x2_ASAP7_75t_R _12613_ (.A1(_08825_),
    .A2(_08858_),
    .B(_08666_),
    .Y(_02738_));
 INVx1_ASAP7_75t_R _12614_ (.A(_01985_),
    .Y(_08859_));
 NAND2x1_ASAP7_75t_R _12615_ (.A(_08859_),
    .B(_08825_),
    .Y(_08860_));
 AND2x2_ASAP7_75t_R _12616_ (.A(_00798_),
    .B(_08836_),
    .Y(_08861_));
 AO221x1_ASAP7_75t_R _12617_ (.A1(_00694_),
    .A2(_08835_),
    .B1(_08861_),
    .B2(_08838_),
    .C(_08839_),
    .Y(_08862_));
 BUFx12f_ASAP7_75t_R _12618_ (.A(_08642_),
    .Y(_08863_));
 AOI21x1_ASAP7_75t_R _12619_ (.A1(_08860_),
    .A2(_08862_),
    .B(_08863_),
    .Y(_02739_));
 NAND2x1_ASAP7_75t_R _12620_ (.A(_08797_),
    .B(_08825_),
    .Y(_08864_));
 AND2x2_ASAP7_75t_R _12621_ (.A(_00797_),
    .B(_08836_),
    .Y(_08865_));
 AO221x1_ASAP7_75t_R _12622_ (.A1(_00693_),
    .A2(_08835_),
    .B1(_08865_),
    .B2(_08838_),
    .C(_08839_),
    .Y(_08866_));
 AOI21x1_ASAP7_75t_R _12623_ (.A1(_08864_),
    .A2(_08866_),
    .B(_08863_),
    .Y(_02740_));
 NAND2x1_ASAP7_75t_R _12624_ (.A(_08800_),
    .B(_08825_),
    .Y(_08867_));
 AND2x2_ASAP7_75t_R _12625_ (.A(_00796_),
    .B(_08836_),
    .Y(_08868_));
 AO221x1_ASAP7_75t_R _12626_ (.A1(_00692_),
    .A2(_08835_),
    .B1(_08868_),
    .B2(_08838_),
    .C(_08839_),
    .Y(_08869_));
 AOI21x1_ASAP7_75t_R _12627_ (.A1(_08867_),
    .A2(_08869_),
    .B(_08863_),
    .Y(_02741_));
 NAND2x1_ASAP7_75t_R _12628_ (.A(_08803_),
    .B(_08825_),
    .Y(_08870_));
 AND2x2_ASAP7_75t_R _12629_ (.A(_00795_),
    .B(_08836_),
    .Y(_08871_));
 AO221x1_ASAP7_75t_R _12630_ (.A1(_00691_),
    .A2(_08834_),
    .B1(_08871_),
    .B2(_08838_),
    .C(_08824_),
    .Y(_08872_));
 AOI21x1_ASAP7_75t_R _12631_ (.A1(_08870_),
    .A2(_08872_),
    .B(_08863_),
    .Y(_02742_));
 OR3x1_ASAP7_75t_R _12632_ (.A(_08657_),
    .B(_08737_),
    .C(_08838_),
    .Y(_08873_));
 INVx1_ASAP7_75t_R _12633_ (.A(_08873_),
    .Y(_02743_));
 NOR2x1_ASAP7_75t_R _12634_ (.A(_08769_),
    .B(_08822_),
    .Y(_08874_));
 AND2x2_ASAP7_75t_R _12635_ (.A(_08774_),
    .B(_08823_),
    .Y(_08875_));
 BUFx12f_ASAP7_75t_R _12636_ (.A(_08526_),
    .Y(_08876_));
 BUFx12f_ASAP7_75t_R _12637_ (.A(_08876_),
    .Y(_08877_));
 OA31x2_ASAP7_75t_R _12638_ (.A1(_08874_),
    .A2(_08875_),
    .A3(_08835_),
    .B1(_08877_),
    .Y(_02744_));
 INVx2_ASAP7_75t_R _12639_ (.A(_01979_),
    .Y(_08878_));
 NAND2x1_ASAP7_75t_R _12640_ (.A(_08878_),
    .B(_08839_),
    .Y(_08879_));
 AND2x2_ASAP7_75t_R _12641_ (.A(_00792_),
    .B(_08749_),
    .Y(_08880_));
 AO221x1_ASAP7_75t_R _12642_ (.A1(_00688_),
    .A2(_08834_),
    .B1(_08880_),
    .B2(_08833_),
    .C(_08824_),
    .Y(_08881_));
 AOI21x1_ASAP7_75t_R _12643_ (.A1(_08879_),
    .A2(_08881_),
    .B(_08863_),
    .Y(_02745_));
 INVx1_ASAP7_75t_R _12644_ (.A(_01978_),
    .Y(_08882_));
 NAND2x1_ASAP7_75t_R _12645_ (.A(_08882_),
    .B(_08839_),
    .Y(_08883_));
 AND2x2_ASAP7_75t_R _12646_ (.A(_00791_),
    .B(_08749_),
    .Y(_08884_));
 AO221x1_ASAP7_75t_R _12647_ (.A1(_00687_),
    .A2(_08834_),
    .B1(_08884_),
    .B2(_08833_),
    .C(_08824_),
    .Y(_08885_));
 AOI21x1_ASAP7_75t_R _12648_ (.A1(_08883_),
    .A2(_08885_),
    .B(_08863_),
    .Y(_02746_));
 AOI21x1_ASAP7_75t_R _12649_ (.A1(_08739_),
    .A2(_08774_),
    .B(_08732_),
    .Y(_08886_));
 BUFx6f_ASAP7_75t_R _12650_ (.A(_08886_),
    .Y(_08887_));
 AND2x2_ASAP7_75t_R _12651_ (.A(_08816_),
    .B(_08887_),
    .Y(_08888_));
 AO21x1_ASAP7_75t_R _12652_ (.A1(_00001_),
    .A2(_08756_),
    .B(_08755_),
    .Y(_08889_));
 NOR2x1_ASAP7_75t_R _12653_ (.A(_08732_),
    .B(_08733_),
    .Y(_08890_));
 NOR2x1_ASAP7_75t_R _12654_ (.A(_00793_),
    .B(_08890_),
    .Y(_08891_));
 OAI21x1_ASAP7_75t_R _12655_ (.A1(_08766_),
    .A2(_08890_),
    .B(_08739_),
    .Y(_08892_));
 AO21x1_ASAP7_75t_R _12656_ (.A1(_08727_),
    .A2(_08891_),
    .B(_08892_),
    .Y(_08893_));
 AO31x2_ASAP7_75t_R _12657_ (.A1(_08749_),
    .A2(_08889_),
    .A3(_08893_),
    .B(_08744_),
    .Y(_08894_));
 OA31x2_ASAP7_75t_R _12658_ (.A1(_08741_),
    .A2(_08745_),
    .A3(_08752_),
    .B1(_08756_),
    .Y(_08895_));
 NOR2x1_ASAP7_75t_R _12659_ (.A(_08894_),
    .B(_08895_),
    .Y(_08896_));
 BUFx6f_ASAP7_75t_R _12660_ (.A(_08896_),
    .Y(_08897_));
 BUFx6f_ASAP7_75t_R _12661_ (.A(_08894_),
    .Y(_08898_));
 BUFx6f_ASAP7_75t_R _12662_ (.A(_08895_),
    .Y(_08899_));
 OA21x2_ASAP7_75t_R _12663_ (.A1(_08898_),
    .A2(_08899_),
    .B(_00804_),
    .Y(_08900_));
 BUFx12f_ASAP7_75t_R _12664_ (.A(_08886_),
    .Y(_08901_));
 AOI211x1_ASAP7_75t_R _12665_ (.A1(_00700_),
    .A2(_08897_),
    .B(_08900_),
    .C(_08901_),
    .Y(_08902_));
 OA21x2_ASAP7_75t_R _12666_ (.A1(_08888_),
    .A2(_08902_),
    .B(_08666_),
    .Y(_02747_));
 AND2x2_ASAP7_75t_R _12667_ (.A(_08841_),
    .B(_08887_),
    .Y(_08903_));
 OA21x2_ASAP7_75t_R _12668_ (.A1(_08898_),
    .A2(_08899_),
    .B(_00803_),
    .Y(_08904_));
 AOI211x1_ASAP7_75t_R _12669_ (.A1(_00699_),
    .A2(_08897_),
    .B(_08904_),
    .C(_08901_),
    .Y(_08905_));
 OA21x2_ASAP7_75t_R _12670_ (.A1(_08903_),
    .A2(_08905_),
    .B(_08666_),
    .Y(_02748_));
 AND2x2_ASAP7_75t_R _12671_ (.A(_08845_),
    .B(_08887_),
    .Y(_08906_));
 OA21x2_ASAP7_75t_R _12672_ (.A1(_08898_),
    .A2(_08899_),
    .B(_00802_),
    .Y(_08907_));
 AOI211x1_ASAP7_75t_R _12673_ (.A1(_00698_),
    .A2(_08897_),
    .B(_08907_),
    .C(_08901_),
    .Y(_08908_));
 OA21x2_ASAP7_75t_R _12674_ (.A1(_08906_),
    .A2(_08908_),
    .B(_08666_),
    .Y(_02749_));
 AND2x2_ASAP7_75t_R _12675_ (.A(_08849_),
    .B(_08887_),
    .Y(_08909_));
 OA21x2_ASAP7_75t_R _12676_ (.A1(_08898_),
    .A2(_08899_),
    .B(_00801_),
    .Y(_08910_));
 AOI211x1_ASAP7_75t_R _12677_ (.A1(_00697_),
    .A2(_08897_),
    .B(_08910_),
    .C(_08901_),
    .Y(_08911_));
 OA21x2_ASAP7_75t_R _12678_ (.A1(_08909_),
    .A2(_08911_),
    .B(_08666_),
    .Y(_02750_));
 AND2x2_ASAP7_75t_R _12679_ (.A(_08853_),
    .B(_08887_),
    .Y(_08912_));
 OA21x2_ASAP7_75t_R _12680_ (.A1(_08898_),
    .A2(_08899_),
    .B(_00800_),
    .Y(_08913_));
 AOI211x1_ASAP7_75t_R _12681_ (.A1(_00696_),
    .A2(_08897_),
    .B(_08913_),
    .C(_08901_),
    .Y(_08914_));
 OA21x2_ASAP7_75t_R _12682_ (.A1(_08912_),
    .A2(_08914_),
    .B(_08666_),
    .Y(_02751_));
 NAND2x1_ASAP7_75t_R _12683_ (.A(_08734_),
    .B(_08901_),
    .Y(_08915_));
 OA21x2_ASAP7_75t_R _12684_ (.A1(_08894_),
    .A2(_08895_),
    .B(_00799_),
    .Y(_08916_));
 AO211x2_ASAP7_75t_R _12685_ (.A1(_00695_),
    .A2(_08897_),
    .B(_08916_),
    .C(_08887_),
    .Y(_08917_));
 AOI21x1_ASAP7_75t_R _12686_ (.A1(_08915_),
    .A2(_08917_),
    .B(_08863_),
    .Y(_02752_));
 AND2x2_ASAP7_75t_R _12687_ (.A(_08859_),
    .B(_08887_),
    .Y(_08918_));
 OR3x1_ASAP7_75t_R _12688_ (.A(_08742_),
    .B(_08894_),
    .C(_08895_),
    .Y(_08919_));
 AO21x1_ASAP7_75t_R _12689_ (.A1(_08739_),
    .A2(_08774_),
    .B(_08732_),
    .Y(_08920_));
 OA211x2_ASAP7_75t_R _12690_ (.A1(_08795_),
    .A2(_08896_),
    .B(_08919_),
    .C(_08920_),
    .Y(_08921_));
 BUFx6f_ASAP7_75t_R _12691_ (.A(_08665_),
    .Y(_08922_));
 OA21x2_ASAP7_75t_R _12692_ (.A1(_08918_),
    .A2(_08921_),
    .B(_08922_),
    .Y(_02753_));
 AND2x2_ASAP7_75t_R _12693_ (.A(_08797_),
    .B(_08887_),
    .Y(_08923_));
 OR3x1_ASAP7_75t_R _12694_ (.A(_08729_),
    .B(_08894_),
    .C(_08895_),
    .Y(_08924_));
 OA211x2_ASAP7_75t_R _12695_ (.A1(_08725_),
    .A2(_08896_),
    .B(_08924_),
    .C(_08920_),
    .Y(_08925_));
 OA21x2_ASAP7_75t_R _12696_ (.A1(_08923_),
    .A2(_08925_),
    .B(_08922_),
    .Y(_02754_));
 AND2x2_ASAP7_75t_R _12697_ (.A(_08800_),
    .B(_08887_),
    .Y(_08926_));
 OA21x2_ASAP7_75t_R _12698_ (.A1(_08898_),
    .A2(_08899_),
    .B(_00796_),
    .Y(_08927_));
 AOI211x1_ASAP7_75t_R _12699_ (.A1(_00692_),
    .A2(_08897_),
    .B(_08927_),
    .C(_08901_),
    .Y(_08928_));
 OA21x2_ASAP7_75t_R _12700_ (.A1(_08926_),
    .A2(_08928_),
    .B(_08922_),
    .Y(_02755_));
 AND2x2_ASAP7_75t_R _12701_ (.A(_08803_),
    .B(_08887_),
    .Y(_08929_));
 OA21x2_ASAP7_75t_R _12702_ (.A1(_08898_),
    .A2(_08899_),
    .B(_00795_),
    .Y(_08930_));
 AOI211x1_ASAP7_75t_R _12703_ (.A1(_00691_),
    .A2(_08897_),
    .B(_08930_),
    .C(_08901_),
    .Y(_08931_));
 OA21x2_ASAP7_75t_R _12704_ (.A1(_08929_),
    .A2(_08931_),
    .B(_08922_),
    .Y(_02756_));
 OR4x1_ASAP7_75t_R _12705_ (.A(_08712_),
    .B(_08732_),
    .C(_08740_),
    .D(_08774_),
    .Y(_08932_));
 INVx1_ASAP7_75t_R _12706_ (.A(_08932_),
    .Y(_02757_));
 INVx1_ASAP7_75t_R _12707_ (.A(_08898_),
    .Y(_08933_));
 OR3x1_ASAP7_75t_R _12708_ (.A(_08886_),
    .B(_08933_),
    .C(_08899_),
    .Y(_08934_));
 AND2x2_ASAP7_75t_R _12709_ (.A(_08723_),
    .B(_08934_),
    .Y(_02758_));
 AND2x2_ASAP7_75t_R _12710_ (.A(_08878_),
    .B(_08886_),
    .Y(_08935_));
 OA21x2_ASAP7_75t_R _12711_ (.A1(_08898_),
    .A2(_08899_),
    .B(_00792_),
    .Y(_08936_));
 AOI211x1_ASAP7_75t_R _12712_ (.A1(_00688_),
    .A2(_08897_),
    .B(_08936_),
    .C(_08901_),
    .Y(_08937_));
 OA21x2_ASAP7_75t_R _12713_ (.A1(_08935_),
    .A2(_08937_),
    .B(_08922_),
    .Y(_02759_));
 AND2x2_ASAP7_75t_R _12714_ (.A(_08882_),
    .B(_08886_),
    .Y(_08938_));
 OA21x2_ASAP7_75t_R _12715_ (.A1(_08898_),
    .A2(_08899_),
    .B(_00791_),
    .Y(_08939_));
 AOI211x1_ASAP7_75t_R _12716_ (.A1(_00687_),
    .A2(_08897_),
    .B(_08939_),
    .C(_08901_),
    .Y(_08940_));
 OA21x2_ASAP7_75t_R _12717_ (.A1(_08938_),
    .A2(_08940_),
    .B(_08922_),
    .Y(_02760_));
 AND2x2_ASAP7_75t_R _12718_ (.A(_08723_),
    .B(_00002_),
    .Y(_02761_));
 BUFx12f_ASAP7_75t_R _12719_ (.A(_08578_),
    .Y(_08941_));
 BUFx12f_ASAP7_75t_R _12720_ (.A(_08941_),
    .Y(_08942_));
 OR2x2_ASAP7_75t_R _12721_ (.A(_00481_),
    .B(_00482_),
    .Y(_08943_));
 BUFx6f_ASAP7_75t_R _12722_ (.A(_08943_),
    .Y(_08944_));
 INVx3_ASAP7_75t_R _12723_ (.A(_00590_),
    .Y(_08945_));
 NAND2x1_ASAP7_75t_R _12724_ (.A(_00587_),
    .B(_00588_),
    .Y(_08946_));
 INVx2_ASAP7_75t_R _12725_ (.A(_00585_),
    .Y(_08947_));
 OA31x2_ASAP7_75t_R _12726_ (.A1(_00589_),
    .A2(_08945_),
    .A3(_08946_),
    .B1(_08947_),
    .Y(_08948_));
 BUFx6f_ASAP7_75t_R _12727_ (.A(_01958_),
    .Y(_08949_));
 INVx2_ASAP7_75t_R _12728_ (.A(_08949_),
    .Y(_08950_));
 BUFx6f_ASAP7_75t_R _12729_ (.A(_01952_),
    .Y(_08951_));
 AOI21x1_ASAP7_75t_R _12730_ (.A1(_01953_),
    .A2(_08950_),
    .B(_08951_),
    .Y(_08952_));
 NOR2x1_ASAP7_75t_R _12731_ (.A(_00585_),
    .B(_00586_),
    .Y(_08953_));
 AO21x2_ASAP7_75t_R _12732_ (.A1(_08948_),
    .A2(_08952_),
    .B(_08953_),
    .Y(_08954_));
 INVx1_ASAP7_75t_R _12733_ (.A(_00486_),
    .Y(_08955_));
 INVx1_ASAP7_75t_R _12734_ (.A(_00487_),
    .Y(_08956_));
 NAND2x1_ASAP7_75t_R _12735_ (.A(_00483_),
    .B(_00484_),
    .Y(_08957_));
 OR5x2_ASAP7_75t_R _12736_ (.A(_00481_),
    .B(_00485_),
    .C(_08955_),
    .D(_08956_),
    .E(_08957_),
    .Y(_08958_));
 AOI21x1_ASAP7_75t_R _12737_ (.A1(_08944_),
    .A2(_08954_),
    .B(_08958_),
    .Y(_08959_));
 INVx3_ASAP7_75t_R _12738_ (.A(_00589_),
    .Y(_08960_));
 INVx2_ASAP7_75t_R _12739_ (.A(_00591_),
    .Y(_08961_));
 AND2x4_ASAP7_75t_R _12740_ (.A(_00587_),
    .B(_00588_),
    .Y(_08962_));
 AND5x2_ASAP7_75t_R _12741_ (.A(_08947_),
    .B(_08960_),
    .C(_00590_),
    .D(_08961_),
    .E(_08962_),
    .Y(_08963_));
 INVx2_ASAP7_75t_R _12742_ (.A(_00485_),
    .Y(_08964_));
 AND2x4_ASAP7_75t_R _12743_ (.A(_00483_),
    .B(_00484_),
    .Y(_08965_));
 AO31x2_ASAP7_75t_R _12744_ (.A1(_08964_),
    .A2(_00486_),
    .A3(_08965_),
    .B(_00481_),
    .Y(_08966_));
 AO21x1_ASAP7_75t_R _12745_ (.A1(_01953_),
    .A2(_08949_),
    .B(_08951_),
    .Y(_08967_));
 OAI21x1_ASAP7_75t_R _12746_ (.A1(_08966_),
    .A2(_08967_),
    .B(_08944_),
    .Y(_08968_));
 OR4x1_ASAP7_75t_R _12747_ (.A(_08951_),
    .B(_00481_),
    .C(_00482_),
    .D(_08949_),
    .Y(_08969_));
 OA21x2_ASAP7_75t_R _12748_ (.A1(_08951_),
    .A2(_01953_),
    .B(_08969_),
    .Y(_08970_));
 INVx3_ASAP7_75t_R _12749_ (.A(_08951_),
    .Y(_08971_));
 AND2x2_ASAP7_75t_R _12750_ (.A(_01953_),
    .B(_08949_),
    .Y(_08972_));
 AND2x2_ASAP7_75t_R _12751_ (.A(_08951_),
    .B(_00002_),
    .Y(_08973_));
 AO21x1_ASAP7_75t_R _12752_ (.A1(_08971_),
    .A2(_08972_),
    .B(_08973_),
    .Y(_08974_));
 AO31x2_ASAP7_75t_R _12753_ (.A1(_08960_),
    .A2(_00590_),
    .A3(_08962_),
    .B(_00585_),
    .Y(_08975_));
 AOI211x1_ASAP7_75t_R _12754_ (.A1(_08966_),
    .A2(_08970_),
    .B(_08974_),
    .C(_08975_),
    .Y(_08976_));
 AOI211x1_ASAP7_75t_R _12755_ (.A1(_08963_),
    .A2(_08968_),
    .B(_08976_),
    .C(_08953_),
    .Y(_08977_));
 NAND2x1_ASAP7_75t_R _12756_ (.A(_08959_),
    .B(_08977_),
    .Y(_08978_));
 BUFx6f_ASAP7_75t_R _12757_ (.A(_08978_),
    .Y(_08979_));
 OR2x2_ASAP7_75t_R _12758_ (.A(_00585_),
    .B(_00586_),
    .Y(_08980_));
 AND2x2_ASAP7_75t_R _12759_ (.A(_08947_),
    .B(_00586_),
    .Y(_08981_));
 OR3x1_ASAP7_75t_R _12760_ (.A(_00589_),
    .B(_08945_),
    .C(_08946_),
    .Y(_08982_));
 AO221x1_ASAP7_75t_R _12761_ (.A1(_08958_),
    .A2(_08980_),
    .B1(_08981_),
    .B2(_08982_),
    .C(_08950_),
    .Y(_08983_));
 OR5x2_ASAP7_75t_R _12762_ (.A(_00585_),
    .B(_00589_),
    .C(_08945_),
    .D(_00591_),
    .E(_08946_),
    .Y(_08984_));
 OR3x1_ASAP7_75t_R _12763_ (.A(_00481_),
    .B(_00482_),
    .C(_08949_),
    .Y(_08985_));
 OA21x2_ASAP7_75t_R _12764_ (.A1(_08958_),
    .A2(_08984_),
    .B(_08985_),
    .Y(_08986_));
 OA211x2_ASAP7_75t_R _12765_ (.A1(_08984_),
    .A2(_08944_),
    .B(_08972_),
    .C(_08971_),
    .Y(_08987_));
 AND3x4_ASAP7_75t_R _12766_ (.A(_08983_),
    .B(_08986_),
    .C(_08987_),
    .Y(_08988_));
 OA21x2_ASAP7_75t_R _12767_ (.A1(_08988_),
    .A2(_08959_),
    .B(_08977_),
    .Y(_08989_));
 AO21x2_ASAP7_75t_R _12768_ (.A1(_08944_),
    .A2(_08954_),
    .B(_08958_),
    .Y(_08990_));
 NAND3x1_ASAP7_75t_R _12769_ (.A(_08988_),
    .B(_08990_),
    .C(_08977_),
    .Y(_08991_));
 BUFx6f_ASAP7_75t_R _12770_ (.A(_08991_),
    .Y(_08992_));
 OA222x2_ASAP7_75t_R _12771_ (.A1(_00492_),
    .A2(_08979_),
    .B1(_08989_),
    .B2(_00596_),
    .C1(_01963_),
    .C2(_08992_),
    .Y(_08993_));
 NOR2x1_ASAP7_75t_R _12772_ (.A(_08942_),
    .B(_08993_),
    .Y(_02762_));
 OA222x2_ASAP7_75t_R _12773_ (.A1(_00491_),
    .A2(_08979_),
    .B1(_08989_),
    .B2(_00595_),
    .C1(_01962_),
    .C2(_08992_),
    .Y(_08994_));
 NOR2x1_ASAP7_75t_R _12774_ (.A(_08942_),
    .B(_08994_),
    .Y(_02763_));
 OA222x2_ASAP7_75t_R _12775_ (.A1(_00490_),
    .A2(_08979_),
    .B1(_08989_),
    .B2(_00594_),
    .C1(_01961_),
    .C2(_08992_),
    .Y(_08995_));
 NOR2x1_ASAP7_75t_R _12776_ (.A(_08942_),
    .B(_08995_),
    .Y(_02764_));
 OA222x2_ASAP7_75t_R _12777_ (.A1(_00489_),
    .A2(_08979_),
    .B1(_08989_),
    .B2(_00593_),
    .C1(_01960_),
    .C2(_08992_),
    .Y(_08996_));
 NOR2x1_ASAP7_75t_R _12778_ (.A(_08942_),
    .B(_08996_),
    .Y(_02765_));
 OA222x2_ASAP7_75t_R _12779_ (.A1(_00488_),
    .A2(_08979_),
    .B1(_08989_),
    .B2(_00592_),
    .C1(_01959_),
    .C2(_08992_),
    .Y(_08997_));
 NOR2x1_ASAP7_75t_R _12780_ (.A(_08942_),
    .B(_08997_),
    .Y(_02766_));
 BUFx12f_ASAP7_75t_R _12781_ (.A(_08527_),
    .Y(_08998_));
 BUFx12f_ASAP7_75t_R _12782_ (.A(_08998_),
    .Y(_08999_));
 AND4x1_ASAP7_75t_R _12783_ (.A(_08999_),
    .B(_08961_),
    .C(_08992_),
    .D(_08979_),
    .Y(_02767_));
 AND3x1_ASAP7_75t_R _12784_ (.A(_08988_),
    .B(_08990_),
    .C(_08977_),
    .Y(_09000_));
 NOR2x1_ASAP7_75t_R _12785_ (.A(_08641_),
    .B(_01957_),
    .Y(_09001_));
 AND4x1_ASAP7_75t_R _12786_ (.A(_08528_),
    .B(_08945_),
    .C(_08992_),
    .D(_08979_),
    .Y(_09002_));
 AO21x1_ASAP7_75t_R _12787_ (.A1(_09000_),
    .A2(_09001_),
    .B(_09002_),
    .Y(_02768_));
 INVx1_ASAP7_75t_R _12788_ (.A(_01956_),
    .Y(_09003_));
 OA21x2_ASAP7_75t_R _12789_ (.A1(_08960_),
    .A2(_08989_),
    .B(_08599_),
    .Y(_09004_));
 OA21x2_ASAP7_75t_R _12790_ (.A1(_09003_),
    .A2(_08992_),
    .B(_09004_),
    .Y(_02769_));
 NOR2x1_ASAP7_75t_R _12791_ (.A(_08641_),
    .B(_01955_),
    .Y(_09005_));
 INVx2_ASAP7_75t_R _12792_ (.A(_00588_),
    .Y(_09006_));
 AND4x1_ASAP7_75t_R _12793_ (.A(_08528_),
    .B(_09006_),
    .C(_08991_),
    .D(_08979_),
    .Y(_09007_));
 AO21x1_ASAP7_75t_R _12794_ (.A1(_09000_),
    .A2(_09005_),
    .B(_09007_),
    .Y(_02770_));
 NOR2x1_ASAP7_75t_R _12795_ (.A(_08641_),
    .B(_01954_),
    .Y(_09008_));
 INVx2_ASAP7_75t_R _12796_ (.A(_00587_),
    .Y(_09009_));
 AND4x1_ASAP7_75t_R _12797_ (.A(_08528_),
    .B(_09009_),
    .C(_08991_),
    .D(_08978_),
    .Y(_09010_));
 AO21x1_ASAP7_75t_R _12798_ (.A1(_09000_),
    .A2(_09008_),
    .B(_09010_),
    .Y(_02771_));
 AO21x1_ASAP7_75t_R _12799_ (.A1(_08963_),
    .A2(_08968_),
    .B(_08976_),
    .Y(_09011_));
 AND3x1_ASAP7_75t_R _12800_ (.A(_08582_),
    .B(_08980_),
    .C(_09011_),
    .Y(_02772_));
 NAND2x1_ASAP7_75t_R _12801_ (.A(_08990_),
    .B(_08977_),
    .Y(_09012_));
 OA21x2_ASAP7_75t_R _12802_ (.A1(_08988_),
    .A2(_09012_),
    .B(_08922_),
    .Y(_02773_));
 OA222x2_ASAP7_75t_R _12803_ (.A1(_00480_),
    .A2(_08979_),
    .B1(_08989_),
    .B2(_00584_),
    .C1(_01951_),
    .C2(_08992_),
    .Y(_09013_));
 NOR2x1_ASAP7_75t_R _12804_ (.A(_08942_),
    .B(_09013_),
    .Y(_02774_));
 OA222x2_ASAP7_75t_R _12805_ (.A1(_00479_),
    .A2(_08979_),
    .B1(_08989_),
    .B2(_00583_),
    .C1(_01950_),
    .C2(_08992_),
    .Y(_09014_));
 NOR2x1_ASAP7_75t_R _12806_ (.A(_08942_),
    .B(_09014_),
    .Y(_02775_));
 INVx1_ASAP7_75t_R _12807_ (.A(_00596_),
    .Y(_09015_));
 INVx1_ASAP7_75t_R _12808_ (.A(_00481_),
    .Y(_09016_));
 AND5x2_ASAP7_75t_R _12809_ (.A(_09016_),
    .B(_08964_),
    .C(_00486_),
    .D(_00487_),
    .E(_08965_),
    .Y(_09017_));
 INVx1_ASAP7_75t_R _12810_ (.A(_08966_),
    .Y(_09018_));
 AO21x1_ASAP7_75t_R _12811_ (.A1(_08971_),
    .A2(_08949_),
    .B(_08973_),
    .Y(_09019_));
 NOR2x1_ASAP7_75t_R _12812_ (.A(_08951_),
    .B(_01953_),
    .Y(_09020_));
 AO31x2_ASAP7_75t_R _12813_ (.A1(_08971_),
    .A2(_08949_),
    .A3(_08953_),
    .B(_09020_),
    .Y(_09021_));
 AO21x2_ASAP7_75t_R _12814_ (.A1(_08948_),
    .A2(_09019_),
    .B(_09021_),
    .Y(_09022_));
 NOR2x1_ASAP7_75t_R _12815_ (.A(_00481_),
    .B(_00482_),
    .Y(_09023_));
 AO221x1_ASAP7_75t_R _12816_ (.A1(_09017_),
    .A2(_08954_),
    .B1(_09018_),
    .B2(_09022_),
    .C(_09023_),
    .Y(_09024_));
 BUFx6f_ASAP7_75t_R _12817_ (.A(_09024_),
    .Y(_09025_));
 BUFx6f_ASAP7_75t_R _12818_ (.A(_09025_),
    .Y(_09026_));
 BUFx6f_ASAP7_75t_R _12819_ (.A(_09025_),
    .Y(_09027_));
 NAND2x1_ASAP7_75t_R _12820_ (.A(_00492_),
    .B(_09027_),
    .Y(_09028_));
 BUFx12f_ASAP7_75t_R _12821_ (.A(_08527_),
    .Y(_09029_));
 OA211x2_ASAP7_75t_R _12822_ (.A1(_09015_),
    .A2(_09026_),
    .B(_09028_),
    .C(_09029_),
    .Y(_09030_));
 OA21x2_ASAP7_75t_R _12823_ (.A1(_08976_),
    .A2(_08968_),
    .B(_08980_),
    .Y(_09031_));
 AOI22x1_ASAP7_75t_R _12824_ (.A1(_09017_),
    .A2(_08954_),
    .B1(_09018_),
    .B2(_09022_),
    .Y(_09032_));
 OA211x2_ASAP7_75t_R _12825_ (.A1(_08984_),
    .A2(_09031_),
    .B(_09032_),
    .C(_08944_),
    .Y(_09033_));
 OA211x2_ASAP7_75t_R _12826_ (.A1(_08958_),
    .A2(_08984_),
    .B(_08985_),
    .C(_01953_),
    .Y(_09034_));
 AO21x2_ASAP7_75t_R _12827_ (.A1(_08983_),
    .A2(_09034_),
    .B(_08951_),
    .Y(_09035_));
 AO21x2_ASAP7_75t_R _12828_ (.A1(_08963_),
    .A2(_09023_),
    .B(_08950_),
    .Y(_09036_));
 AO221x1_ASAP7_75t_R _12829_ (.A1(_09017_),
    .A2(_08953_),
    .B1(_08966_),
    .B2(_08963_),
    .C(_08949_),
    .Y(_09037_));
 NAND3x2_ASAP7_75t_R _12830_ (.B(_09036_),
    .C(_09037_),
    .Y(_09038_),
    .A(_08971_));
 AND4x1_ASAP7_75t_R _12831_ (.A(_08971_),
    .B(_08950_),
    .C(_09035_),
    .D(_09038_),
    .Y(_09039_));
 NAND2x1_ASAP7_75t_R _12832_ (.A(_09033_),
    .B(_09039_),
    .Y(_09040_));
 INVx1_ASAP7_75t_R _12833_ (.A(_01963_),
    .Y(_09041_));
 BUFx6f_ASAP7_75t_R _12834_ (.A(_09033_),
    .Y(_09042_));
 BUFx6f_ASAP7_75t_R _12835_ (.A(_09039_),
    .Y(_09043_));
 AND4x1_ASAP7_75t_R _12836_ (.A(_08528_),
    .B(_09041_),
    .C(_09042_),
    .D(_09043_),
    .Y(_09044_));
 AO21x1_ASAP7_75t_R _12837_ (.A1(_09030_),
    .A2(_09040_),
    .B(_09044_),
    .Y(_02776_));
 BUFx6f_ASAP7_75t_R _12838_ (.A(_09040_),
    .Y(_09045_));
 INVx1_ASAP7_75t_R _12839_ (.A(_00595_),
    .Y(_09046_));
 NAND2x1_ASAP7_75t_R _12840_ (.A(_00491_),
    .B(_09027_),
    .Y(_09047_));
 OA211x2_ASAP7_75t_R _12841_ (.A1(_09046_),
    .A2(_09026_),
    .B(_09047_),
    .C(_09029_),
    .Y(_09048_));
 INVx1_ASAP7_75t_R _12842_ (.A(_01962_),
    .Y(_09049_));
 AND4x1_ASAP7_75t_R _12843_ (.A(_08528_),
    .B(_09049_),
    .C(_09042_),
    .D(_09043_),
    .Y(_09050_));
 AO21x1_ASAP7_75t_R _12844_ (.A1(_09045_),
    .A2(_09048_),
    .B(_09050_),
    .Y(_02777_));
 INVx1_ASAP7_75t_R _12845_ (.A(_00594_),
    .Y(_09051_));
 NAND2x1_ASAP7_75t_R _12846_ (.A(_00490_),
    .B(_09027_),
    .Y(_09052_));
 OA211x2_ASAP7_75t_R _12847_ (.A1(_09051_),
    .A2(_09026_),
    .B(_09052_),
    .C(_09029_),
    .Y(_09053_));
 INVx1_ASAP7_75t_R _12848_ (.A(_01961_),
    .Y(_09054_));
 AND4x1_ASAP7_75t_R _12849_ (.A(_08722_),
    .B(_09054_),
    .C(_09042_),
    .D(_09043_),
    .Y(_09055_));
 AO21x1_ASAP7_75t_R _12850_ (.A1(_09045_),
    .A2(_09053_),
    .B(_09055_),
    .Y(_02778_));
 INVx1_ASAP7_75t_R _12851_ (.A(_00593_),
    .Y(_09056_));
 NAND2x1_ASAP7_75t_R _12852_ (.A(_00489_),
    .B(_09027_),
    .Y(_09057_));
 BUFx6f_ASAP7_75t_R _12853_ (.A(_08527_),
    .Y(_09058_));
 OA211x2_ASAP7_75t_R _12854_ (.A1(_09056_),
    .A2(_09026_),
    .B(_09057_),
    .C(_09058_),
    .Y(_09059_));
 INVx1_ASAP7_75t_R _12855_ (.A(_01960_),
    .Y(_09060_));
 AND4x1_ASAP7_75t_R _12856_ (.A(_08722_),
    .B(_09060_),
    .C(_09042_),
    .D(_09043_),
    .Y(_09061_));
 AO21x1_ASAP7_75t_R _12857_ (.A1(_09045_),
    .A2(_09059_),
    .B(_09061_),
    .Y(_02779_));
 INVx1_ASAP7_75t_R _12858_ (.A(_00592_),
    .Y(_09062_));
 NAND2x1_ASAP7_75t_R _12859_ (.A(_00488_),
    .B(_09027_),
    .Y(_09063_));
 OA211x2_ASAP7_75t_R _12860_ (.A1(_09062_),
    .A2(_09026_),
    .B(_09063_),
    .C(_09058_),
    .Y(_09064_));
 INVx1_ASAP7_75t_R _12861_ (.A(_01959_),
    .Y(_09065_));
 AND4x1_ASAP7_75t_R _12862_ (.A(_08722_),
    .B(_09065_),
    .C(_09042_),
    .D(_09043_),
    .Y(_09066_));
 AO21x1_ASAP7_75t_R _12863_ (.A1(_09045_),
    .A2(_09064_),
    .B(_09066_),
    .Y(_02780_));
 NAND2x1_ASAP7_75t_R _12864_ (.A(_00487_),
    .B(_09026_),
    .Y(_09067_));
 OAI21x1_ASAP7_75t_R _12865_ (.A1(_08961_),
    .A2(_09026_),
    .B(_09067_),
    .Y(_09068_));
 AOI21x1_ASAP7_75t_R _12866_ (.A1(_09045_),
    .A2(_09068_),
    .B(_08863_),
    .Y(_02781_));
 NAND2x1_ASAP7_75t_R _12867_ (.A(_00486_),
    .B(_09027_),
    .Y(_09069_));
 OA211x2_ASAP7_75t_R _12868_ (.A1(_08945_),
    .A2(_09026_),
    .B(_09069_),
    .C(_09058_),
    .Y(_09070_));
 AND3x1_ASAP7_75t_R _12869_ (.A(_09001_),
    .B(_09042_),
    .C(_09043_),
    .Y(_09071_));
 AO21x1_ASAP7_75t_R _12870_ (.A1(_09045_),
    .A2(_09070_),
    .B(_09071_),
    .Y(_02782_));
 NAND2x1_ASAP7_75t_R _12871_ (.A(_00485_),
    .B(_09027_),
    .Y(_09072_));
 OA211x2_ASAP7_75t_R _12872_ (.A1(_08960_),
    .A2(_09026_),
    .B(_09072_),
    .C(_09058_),
    .Y(_09073_));
 AND4x1_ASAP7_75t_R _12873_ (.A(_08722_),
    .B(_09003_),
    .C(_09042_),
    .D(_09043_),
    .Y(_09074_));
 AO21x1_ASAP7_75t_R _12874_ (.A1(_09045_),
    .A2(_09073_),
    .B(_09074_),
    .Y(_02783_));
 NAND2x1_ASAP7_75t_R _12875_ (.A(_00484_),
    .B(_09025_),
    .Y(_09075_));
 OA211x2_ASAP7_75t_R _12876_ (.A1(_09006_),
    .A2(_09026_),
    .B(_09075_),
    .C(_09058_),
    .Y(_09076_));
 AND3x1_ASAP7_75t_R _12877_ (.A(_09005_),
    .B(_09042_),
    .C(_09043_),
    .Y(_09077_));
 AO21x1_ASAP7_75t_R _12878_ (.A1(_09045_),
    .A2(_09076_),
    .B(_09077_),
    .Y(_02784_));
 NAND2x1_ASAP7_75t_R _12879_ (.A(_00483_),
    .B(_09025_),
    .Y(_09078_));
 OA211x2_ASAP7_75t_R _12880_ (.A1(_09009_),
    .A2(_09027_),
    .B(_09078_),
    .C(_09058_),
    .Y(_09079_));
 AND3x1_ASAP7_75t_R _12881_ (.A(_09008_),
    .B(_09042_),
    .C(_09043_),
    .Y(_09080_));
 AO21x1_ASAP7_75t_R _12882_ (.A1(_09045_),
    .A2(_09079_),
    .B(_09080_),
    .Y(_02785_));
 BUFx12f_ASAP7_75t_R _12883_ (.A(_08573_),
    .Y(_09081_));
 NOR3x1_ASAP7_75t_R _12884_ (.A(_09081_),
    .B(_09023_),
    .C(_09032_),
    .Y(_02786_));
 INVx1_ASAP7_75t_R _12885_ (.A(_09042_),
    .Y(_09082_));
 OA21x2_ASAP7_75t_R _12886_ (.A1(_09082_),
    .A2(_09043_),
    .B(_08922_),
    .Y(_02787_));
 INVx1_ASAP7_75t_R _12887_ (.A(_00584_),
    .Y(_09083_));
 NAND2x1_ASAP7_75t_R _12888_ (.A(_00480_),
    .B(_09025_),
    .Y(_09084_));
 OA211x2_ASAP7_75t_R _12889_ (.A1(_09083_),
    .A2(_09027_),
    .B(_09084_),
    .C(_09058_),
    .Y(_09085_));
 INVx1_ASAP7_75t_R _12890_ (.A(_01951_),
    .Y(_09086_));
 AND4x1_ASAP7_75t_R _12891_ (.A(_08722_),
    .B(_09086_),
    .C(_09033_),
    .D(_09039_),
    .Y(_09087_));
 AO21x1_ASAP7_75t_R _12892_ (.A1(_09045_),
    .A2(_09085_),
    .B(_09087_),
    .Y(_02788_));
 INVx1_ASAP7_75t_R _12893_ (.A(_00583_),
    .Y(_09088_));
 NAND2x1_ASAP7_75t_R _12894_ (.A(_00479_),
    .B(_09025_),
    .Y(_09089_));
 OA211x2_ASAP7_75t_R _12895_ (.A1(_09088_),
    .A2(_09027_),
    .B(_09089_),
    .C(_09058_),
    .Y(_09090_));
 INVx1_ASAP7_75t_R _12896_ (.A(_01950_),
    .Y(_09091_));
 AND4x1_ASAP7_75t_R _12897_ (.A(_08722_),
    .B(_09091_),
    .C(_09033_),
    .D(_09039_),
    .Y(_09092_));
 AO21x1_ASAP7_75t_R _12898_ (.A1(_09040_),
    .A2(_09090_),
    .B(_09092_),
    .Y(_02789_));
 NAND2x2_ASAP7_75t_R _12899_ (.A(_09035_),
    .B(_09038_),
    .Y(_09093_));
 AND2x2_ASAP7_75t_R _12900_ (.A(_09041_),
    .B(_09093_),
    .Y(_09094_));
 INVx1_ASAP7_75t_R _12901_ (.A(_00586_),
    .Y(_09095_));
 AO221x1_ASAP7_75t_R _12902_ (.A1(_08947_),
    .A2(_09095_),
    .B1(_08966_),
    .B2(_08970_),
    .C(_08974_),
    .Y(_09096_));
 AO221x1_ASAP7_75t_R _12903_ (.A1(_08944_),
    .A2(_09022_),
    .B1(_09096_),
    .B2(_08948_),
    .C(_08966_),
    .Y(_09097_));
 BUFx12f_ASAP7_75t_R _12904_ (.A(_09097_),
    .Y(_09098_));
 AOI221x1_ASAP7_75t_R _12905_ (.A1(_08944_),
    .A2(_09022_),
    .B1(_09096_),
    .B2(_08948_),
    .C(_08966_),
    .Y(_09099_));
 AND2x2_ASAP7_75t_R _12906_ (.A(_00492_),
    .B(_09099_),
    .Y(_09100_));
 AOI211x1_ASAP7_75t_R _12907_ (.A1(_00596_),
    .A2(_09098_),
    .B(_09100_),
    .C(_09093_),
    .Y(_09101_));
 OA21x2_ASAP7_75t_R _12908_ (.A1(_09094_),
    .A2(_09101_),
    .B(_08922_),
    .Y(_02790_));
 BUFx6f_ASAP7_75t_R _12909_ (.A(_09035_),
    .Y(_09102_));
 BUFx6f_ASAP7_75t_R _12910_ (.A(_09038_),
    .Y(_09103_));
 AO21x1_ASAP7_75t_R _12911_ (.A1(_09102_),
    .A2(_09103_),
    .B(_01962_),
    .Y(_09104_));
 BUFx6f_ASAP7_75t_R _12912_ (.A(_09097_),
    .Y(_09105_));
 OR2x2_ASAP7_75t_R _12913_ (.A(_00491_),
    .B(_09105_),
    .Y(_09106_));
 NAND2x1_ASAP7_75t_R _12914_ (.A(_09046_),
    .B(_09098_),
    .Y(_09107_));
 BUFx6f_ASAP7_75t_R _12915_ (.A(_09093_),
    .Y(_09108_));
 AO21x1_ASAP7_75t_R _12916_ (.A1(_09106_),
    .A2(_09107_),
    .B(_09108_),
    .Y(_09109_));
 AOI21x1_ASAP7_75t_R _12917_ (.A1(_09104_),
    .A2(_09109_),
    .B(_08863_),
    .Y(_02791_));
 AO21x1_ASAP7_75t_R _12918_ (.A1(_09102_),
    .A2(_09103_),
    .B(_01961_),
    .Y(_09110_));
 OR2x2_ASAP7_75t_R _12919_ (.A(_00490_),
    .B(_09105_),
    .Y(_09111_));
 NAND2x1_ASAP7_75t_R _12920_ (.A(_09051_),
    .B(_09098_),
    .Y(_09112_));
 AO21x1_ASAP7_75t_R _12921_ (.A1(_09111_),
    .A2(_09112_),
    .B(_09108_),
    .Y(_09113_));
 AOI21x1_ASAP7_75t_R _12922_ (.A1(_09110_),
    .A2(_09113_),
    .B(_08863_),
    .Y(_02792_));
 AO21x1_ASAP7_75t_R _12923_ (.A1(_09102_),
    .A2(_09103_),
    .B(_01960_),
    .Y(_09114_));
 OR2x2_ASAP7_75t_R _12924_ (.A(_00489_),
    .B(_09105_),
    .Y(_09115_));
 NAND2x1_ASAP7_75t_R _12925_ (.A(_09056_),
    .B(_09098_),
    .Y(_09116_));
 AO21x1_ASAP7_75t_R _12926_ (.A1(_09115_),
    .A2(_09116_),
    .B(_09108_),
    .Y(_09117_));
 BUFx12f_ASAP7_75t_R _12927_ (.A(_08641_),
    .Y(_09118_));
 BUFx12f_ASAP7_75t_R _12928_ (.A(_09118_),
    .Y(_09119_));
 AOI21x1_ASAP7_75t_R _12929_ (.A1(_09114_),
    .A2(_09117_),
    .B(_09119_),
    .Y(_02793_));
 AO21x1_ASAP7_75t_R _12930_ (.A1(_09102_),
    .A2(_09103_),
    .B(_01959_),
    .Y(_09120_));
 OR2x2_ASAP7_75t_R _12931_ (.A(_00488_),
    .B(_09105_),
    .Y(_09121_));
 NAND2x1_ASAP7_75t_R _12932_ (.A(_09062_),
    .B(_09098_),
    .Y(_09122_));
 AO21x1_ASAP7_75t_R _12933_ (.A1(_09121_),
    .A2(_09122_),
    .B(_09108_),
    .Y(_09123_));
 AOI21x1_ASAP7_75t_R _12934_ (.A1(_09120_),
    .A2(_09123_),
    .B(_09119_),
    .Y(_02794_));
 AO21x1_ASAP7_75t_R _12935_ (.A1(_09102_),
    .A2(_09103_),
    .B(_08949_),
    .Y(_09124_));
 NAND2x1_ASAP7_75t_R _12936_ (.A(_08956_),
    .B(_09099_),
    .Y(_09125_));
 NAND2x1_ASAP7_75t_R _12937_ (.A(_08961_),
    .B(_09098_),
    .Y(_09126_));
 AO21x1_ASAP7_75t_R _12938_ (.A1(_09125_),
    .A2(_09126_),
    .B(_09108_),
    .Y(_09127_));
 AOI21x1_ASAP7_75t_R _12939_ (.A1(_09124_),
    .A2(_09127_),
    .B(_09119_),
    .Y(_02795_));
 AO21x1_ASAP7_75t_R _12940_ (.A1(_09102_),
    .A2(_09103_),
    .B(_01957_),
    .Y(_09128_));
 NAND2x1_ASAP7_75t_R _12941_ (.A(_08955_),
    .B(_09099_),
    .Y(_09129_));
 NAND2x1_ASAP7_75t_R _12942_ (.A(_08945_),
    .B(_09098_),
    .Y(_09130_));
 AO21x1_ASAP7_75t_R _12943_ (.A1(_09129_),
    .A2(_09130_),
    .B(_09108_),
    .Y(_09131_));
 AOI21x1_ASAP7_75t_R _12944_ (.A1(_09128_),
    .A2(_09131_),
    .B(_09119_),
    .Y(_02796_));
 AO21x1_ASAP7_75t_R _12945_ (.A1(_09102_),
    .A2(_09103_),
    .B(_01956_),
    .Y(_09132_));
 NAND2x1_ASAP7_75t_R _12946_ (.A(_08964_),
    .B(_09099_),
    .Y(_09133_));
 NAND2x1_ASAP7_75t_R _12947_ (.A(_08960_),
    .B(_09098_),
    .Y(_09134_));
 AO21x1_ASAP7_75t_R _12948_ (.A1(_09133_),
    .A2(_09134_),
    .B(_09108_),
    .Y(_09135_));
 AOI21x1_ASAP7_75t_R _12949_ (.A1(_09132_),
    .A2(_09135_),
    .B(_09119_),
    .Y(_02797_));
 AO21x1_ASAP7_75t_R _12950_ (.A1(_09102_),
    .A2(_09103_),
    .B(_01955_),
    .Y(_09136_));
 OR2x2_ASAP7_75t_R _12951_ (.A(_00484_),
    .B(_09105_),
    .Y(_09137_));
 NAND2x1_ASAP7_75t_R _12952_ (.A(_09006_),
    .B(_09098_),
    .Y(_09138_));
 AO21x1_ASAP7_75t_R _12953_ (.A1(_09137_),
    .A2(_09138_),
    .B(_09108_),
    .Y(_09139_));
 AOI21x1_ASAP7_75t_R _12954_ (.A1(_09136_),
    .A2(_09139_),
    .B(_09119_),
    .Y(_02798_));
 AO21x1_ASAP7_75t_R _12955_ (.A1(_09102_),
    .A2(_09103_),
    .B(_01954_),
    .Y(_09140_));
 OR2x2_ASAP7_75t_R _12956_ (.A(_00483_),
    .B(_09105_),
    .Y(_09141_));
 NAND2x1_ASAP7_75t_R _12957_ (.A(_09009_),
    .B(_09098_),
    .Y(_09142_));
 AO21x1_ASAP7_75t_R _12958_ (.A1(_09141_),
    .A2(_09142_),
    .B(_09108_),
    .Y(_09143_));
 AOI21x1_ASAP7_75t_R _12959_ (.A1(_09140_),
    .A2(_09143_),
    .B(_09119_),
    .Y(_02799_));
 AO21x1_ASAP7_75t_R _12960_ (.A1(_08983_),
    .A2(_08986_),
    .B(_08951_),
    .Y(_09144_));
 BUFx12f_ASAP7_75t_R _12961_ (.A(_08587_),
    .Y(_09145_));
 AOI211x1_ASAP7_75t_R _12962_ (.A1(_09103_),
    .A2(_09144_),
    .B(_09145_),
    .C(_09020_),
    .Y(_02800_));
 AOI21x1_ASAP7_75t_R _12963_ (.A1(_08944_),
    .A2(_09022_),
    .B(_08966_),
    .Y(_09146_));
 AO21x1_ASAP7_75t_R _12964_ (.A1(_08948_),
    .A2(_09096_),
    .B(_09146_),
    .Y(_09147_));
 OA21x2_ASAP7_75t_R _12965_ (.A1(_09108_),
    .A2(_09147_),
    .B(_08922_),
    .Y(_02801_));
 AO21x1_ASAP7_75t_R _12966_ (.A1(_09102_),
    .A2(_09038_),
    .B(_01951_),
    .Y(_09148_));
 OR2x2_ASAP7_75t_R _12967_ (.A(_00480_),
    .B(_09105_),
    .Y(_09149_));
 NAND2x1_ASAP7_75t_R _12968_ (.A(_09083_),
    .B(_09105_),
    .Y(_09150_));
 AO21x1_ASAP7_75t_R _12969_ (.A1(_09149_),
    .A2(_09150_),
    .B(_09093_),
    .Y(_09151_));
 AOI21x1_ASAP7_75t_R _12970_ (.A1(_09148_),
    .A2(_09151_),
    .B(_09119_),
    .Y(_02802_));
 AO21x1_ASAP7_75t_R _12971_ (.A1(_09035_),
    .A2(_09038_),
    .B(_01950_),
    .Y(_09152_));
 OR2x2_ASAP7_75t_R _12972_ (.A(_00479_),
    .B(_09105_),
    .Y(_09153_));
 NAND2x1_ASAP7_75t_R _12973_ (.A(_09088_),
    .B(_09105_),
    .Y(_09154_));
 AO21x1_ASAP7_75t_R _12974_ (.A1(_09153_),
    .A2(_09154_),
    .B(_09093_),
    .Y(_09155_));
 AOI21x1_ASAP7_75t_R _12975_ (.A1(_09152_),
    .A2(_09155_),
    .B(_09119_),
    .Y(_02803_));
 AND2x2_ASAP7_75t_R _12976_ (.A(_08723_),
    .B(_00003_),
    .Y(_02804_));
 OR2x6_ASAP7_75t_R _12977_ (.A(_00377_),
    .B(_00378_),
    .Y(_09156_));
 NOR2x1_ASAP7_75t_R _12978_ (.A(_00381_),
    .B(_00382_),
    .Y(_09157_));
 AND2x2_ASAP7_75t_R _12979_ (.A(_00379_),
    .B(_00380_),
    .Y(_09158_));
 AO21x2_ASAP7_75t_R _12980_ (.A1(_09157_),
    .A2(_09158_),
    .B(_00377_),
    .Y(_09159_));
 NOR2x1_ASAP7_75t_R _12981_ (.A(_00277_),
    .B(_00278_),
    .Y(_09160_));
 AND2x4_ASAP7_75t_R _12982_ (.A(_00275_),
    .B(_00276_),
    .Y(_09161_));
 AND3x1_ASAP7_75t_R _12983_ (.A(_00274_),
    .B(_09160_),
    .C(_09161_),
    .Y(_09162_));
 INVx2_ASAP7_75t_R _12984_ (.A(_01938_),
    .Y(_09163_));
 BUFx3_ASAP7_75t_R _12985_ (.A(_01944_),
    .Y(_09164_));
 BUFx6f_ASAP7_75t_R _12986_ (.A(_00273_),
    .Y(_09165_));
 AO21x1_ASAP7_75t_R _12987_ (.A1(_09163_),
    .A2(_09164_),
    .B(_09165_),
    .Y(_09166_));
 BUFx6f_ASAP7_75t_R _12988_ (.A(_01939_),
    .Y(_09167_));
 OA21x2_ASAP7_75t_R _12989_ (.A1(_09162_),
    .A2(_09166_),
    .B(_09167_),
    .Y(_09168_));
 AO21x2_ASAP7_75t_R _12990_ (.A1(_09160_),
    .A2(_09161_),
    .B(_09165_),
    .Y(_09169_));
 OA21x2_ASAP7_75t_R _12991_ (.A1(_00003_),
    .A2(_09169_),
    .B(_01938_),
    .Y(_09170_));
 OR3x2_ASAP7_75t_R _12992_ (.A(_09159_),
    .B(_09168_),
    .C(_09170_),
    .Y(_09171_));
 OR2x2_ASAP7_75t_R _12993_ (.A(_00381_),
    .B(_00382_),
    .Y(_09172_));
 NAND2x1_ASAP7_75t_R _12994_ (.A(_00379_),
    .B(_00380_),
    .Y(_09173_));
 OR4x1_ASAP7_75t_R _12995_ (.A(_00377_),
    .B(_00383_),
    .C(_09172_),
    .D(_09173_),
    .Y(_09174_));
 AO21x1_ASAP7_75t_R _12996_ (.A1(_09167_),
    .A2(_09164_),
    .B(_01938_),
    .Y(_09175_));
 OR2x2_ASAP7_75t_R _12997_ (.A(_09165_),
    .B(_00274_),
    .Y(_09176_));
 BUFx3_ASAP7_75t_R _12998_ (.A(_09176_),
    .Y(_09177_));
 OA21x2_ASAP7_75t_R _12999_ (.A1(_09169_),
    .A2(_09175_),
    .B(_09177_),
    .Y(_09178_));
 OR2x6_ASAP7_75t_R _13000_ (.A(_09174_),
    .B(_09178_),
    .Y(_09179_));
 AND3x4_ASAP7_75t_R _13001_ (.A(_09156_),
    .B(_09171_),
    .C(_09179_),
    .Y(_09180_));
 INVx1_ASAP7_75t_R _13002_ (.A(_09164_),
    .Y(_09181_));
 AO21x1_ASAP7_75t_R _13003_ (.A1(_09167_),
    .A2(_09181_),
    .B(_01938_),
    .Y(_09182_));
 OAI21x1_ASAP7_75t_R _13004_ (.A1(_09159_),
    .A2(_09182_),
    .B(_09156_),
    .Y(_09183_));
 INVx1_ASAP7_75t_R _13005_ (.A(_00279_),
    .Y(_09184_));
 NAND2x1_ASAP7_75t_R _13006_ (.A(_00275_),
    .B(_00276_),
    .Y(_09185_));
 OR5x2_ASAP7_75t_R _13007_ (.A(_09165_),
    .B(_00277_),
    .C(_00278_),
    .D(_09184_),
    .E(_09185_),
    .Y(_09186_));
 AOI21x1_ASAP7_75t_R _13008_ (.A1(_09177_),
    .A2(_09183_),
    .B(_09186_),
    .Y(_09187_));
 INVx1_ASAP7_75t_R _13009_ (.A(_00377_),
    .Y(_09188_));
 INVx2_ASAP7_75t_R _13010_ (.A(_00383_),
    .Y(_09189_));
 AND4x1_ASAP7_75t_R _13011_ (.A(_09188_),
    .B(_09189_),
    .C(_09157_),
    .D(_09158_),
    .Y(_09190_));
 NOR2x1_ASAP7_75t_R _13012_ (.A(_09165_),
    .B(_00274_),
    .Y(_09191_));
 INVx1_ASAP7_75t_R _13013_ (.A(_09165_),
    .Y(_09192_));
 AND4x1_ASAP7_75t_R _13014_ (.A(_09192_),
    .B(_00279_),
    .C(_09160_),
    .D(_09161_),
    .Y(_09193_));
 AOI221x1_ASAP7_75t_R _13015_ (.A1(_09190_),
    .A2(_09191_),
    .B1(_09193_),
    .B2(_09159_),
    .C(_09181_),
    .Y(_09194_));
 OA21x2_ASAP7_75t_R _13016_ (.A1(_00377_),
    .A2(_00378_),
    .B(_09164_),
    .Y(_09195_));
 AO21x1_ASAP7_75t_R _13017_ (.A1(_09181_),
    .A2(_09177_),
    .B(_09195_),
    .Y(_09196_));
 OA21x2_ASAP7_75t_R _13018_ (.A1(_09174_),
    .A2(_09186_),
    .B(_09196_),
    .Y(_09197_));
 AND2x4_ASAP7_75t_R _13019_ (.A(_09163_),
    .B(_09167_),
    .Y(_09198_));
 AND3x4_ASAP7_75t_R _13020_ (.A(_09194_),
    .B(_09197_),
    .C(_09198_),
    .Y(_09199_));
 OR2x6_ASAP7_75t_R _13021_ (.A(_09187_),
    .B(_09199_),
    .Y(_09200_));
 NAND2x2_ASAP7_75t_R _13022_ (.A(_09180_),
    .B(_09200_),
    .Y(_09201_));
 AND4x1_ASAP7_75t_R _13023_ (.A(_09156_),
    .B(_09171_),
    .C(_09179_),
    .D(_09187_),
    .Y(_09202_));
 BUFx3_ASAP7_75t_R _13024_ (.A(_09202_),
    .Y(_09203_));
 AO21x1_ASAP7_75t_R _13025_ (.A1(_09177_),
    .A2(_09183_),
    .B(_09186_),
    .Y(_09204_));
 AND2x6_ASAP7_75t_R _13026_ (.A(_09204_),
    .B(_09199_),
    .Y(_09205_));
 BUFx6f_ASAP7_75t_R _13027_ (.A(_09205_),
    .Y(_09206_));
 BUFx12f_ASAP7_75t_R _13028_ (.A(_08572_),
    .Y(_09207_));
 AO221x1_ASAP7_75t_R _13029_ (.A1(_00284_),
    .A2(_09203_),
    .B1(_09206_),
    .B2(_01949_),
    .C(_09207_),
    .Y(_09208_));
 AOI21x1_ASAP7_75t_R _13030_ (.A1(_00388_),
    .A2(_09201_),
    .B(_09208_),
    .Y(_02805_));
 AO221x1_ASAP7_75t_R _13031_ (.A1(_00283_),
    .A2(_09203_),
    .B1(_09206_),
    .B2(_01948_),
    .C(_09207_),
    .Y(_09209_));
 AOI21x1_ASAP7_75t_R _13032_ (.A1(_00387_),
    .A2(_09201_),
    .B(_09209_),
    .Y(_02806_));
 AO221x1_ASAP7_75t_R _13033_ (.A1(_00282_),
    .A2(_09203_),
    .B1(_09206_),
    .B2(_01947_),
    .C(_09207_),
    .Y(_09210_));
 AOI21x1_ASAP7_75t_R _13034_ (.A1(_00386_),
    .A2(_09201_),
    .B(_09210_),
    .Y(_02807_));
 BUFx6f_ASAP7_75t_R _13035_ (.A(_08656_),
    .Y(_09211_));
 AO221x1_ASAP7_75t_R _13036_ (.A1(_00281_),
    .A2(_09203_),
    .B1(_09206_),
    .B2(_01946_),
    .C(_09211_),
    .Y(_09212_));
 AOI21x1_ASAP7_75t_R _13037_ (.A1(_00385_),
    .A2(_09201_),
    .B(_09212_),
    .Y(_02808_));
 AO221x1_ASAP7_75t_R _13038_ (.A1(_00280_),
    .A2(_09203_),
    .B1(_09206_),
    .B2(_01945_),
    .C(_09211_),
    .Y(_09213_));
 AOI21x1_ASAP7_75t_R _13039_ (.A1(_00384_),
    .A2(_09201_),
    .B(_09213_),
    .Y(_02809_));
 AND3x1_ASAP7_75t_R _13040_ (.A(_08582_),
    .B(_09189_),
    .C(_09201_),
    .Y(_02810_));
 INVx1_ASAP7_75t_R _13041_ (.A(_00382_),
    .Y(_09214_));
 OR3x1_ASAP7_75t_R _13042_ (.A(_09214_),
    .B(_09203_),
    .C(_09205_),
    .Y(_09215_));
 NAND2x1_ASAP7_75t_R _13043_ (.A(_01943_),
    .B(_09206_),
    .Y(_09216_));
 AND3x1_ASAP7_75t_R _13044_ (.A(_08582_),
    .B(_09215_),
    .C(_09216_),
    .Y(_02811_));
 INVx1_ASAP7_75t_R _13045_ (.A(_00381_),
    .Y(_09217_));
 OR3x1_ASAP7_75t_R _13046_ (.A(_09217_),
    .B(_09202_),
    .C(_09205_),
    .Y(_09218_));
 NAND2x1_ASAP7_75t_R _13047_ (.A(_01942_),
    .B(_09206_),
    .Y(_09219_));
 AND3x1_ASAP7_75t_R _13048_ (.A(_08582_),
    .B(_09218_),
    .C(_09219_),
    .Y(_02812_));
 BUFx12f_ASAP7_75t_R _13049_ (.A(net21),
    .Y(_09220_));
 BUFx12f_ASAP7_75t_R _13050_ (.A(_09220_),
    .Y(_09221_));
 OR4x1_ASAP7_75t_R _13051_ (.A(_09221_),
    .B(_00380_),
    .C(_09203_),
    .D(_09205_),
    .Y(_09222_));
 BUFx12f_ASAP7_75t_R _13052_ (.A(_08572_),
    .Y(_09223_));
 NOR2x1_ASAP7_75t_R _13053_ (.A(_09223_),
    .B(_01941_),
    .Y(_09224_));
 NAND2x1_ASAP7_75t_R _13054_ (.A(_09206_),
    .B(_09224_),
    .Y(_09225_));
 NAND2x1_ASAP7_75t_R _13055_ (.A(_09222_),
    .B(_09225_),
    .Y(_02813_));
 OR4x1_ASAP7_75t_R _13056_ (.A(_09221_),
    .B(_00379_),
    .C(_09203_),
    .D(_09205_),
    .Y(_09226_));
 NOR2x1_ASAP7_75t_R _13057_ (.A(_09223_),
    .B(_01940_),
    .Y(_09227_));
 NAND2x1_ASAP7_75t_R _13058_ (.A(_09206_),
    .B(_09227_),
    .Y(_09228_));
 NAND2x1_ASAP7_75t_R _13059_ (.A(_09226_),
    .B(_09228_),
    .Y(_02814_));
 BUFx12f_ASAP7_75t_R _13060_ (.A(_08598_),
    .Y(_09229_));
 NAND2x1_ASAP7_75t_R _13061_ (.A(_09229_),
    .B(_09156_),
    .Y(_09230_));
 AO21x1_ASAP7_75t_R _13062_ (.A1(_09171_),
    .A2(_09179_),
    .B(_09230_),
    .Y(_09231_));
 INVx1_ASAP7_75t_R _13063_ (.A(_09231_),
    .Y(_02815_));
 INVx1_ASAP7_75t_R _13064_ (.A(_09200_),
    .Y(_09232_));
 AOI21x1_ASAP7_75t_R _13065_ (.A1(_09180_),
    .A2(_09232_),
    .B(_09119_),
    .Y(_02816_));
 AO221x1_ASAP7_75t_R _13066_ (.A1(_00272_),
    .A2(_09203_),
    .B1(_09206_),
    .B2(_01937_),
    .C(_09211_),
    .Y(_09233_));
 AOI21x1_ASAP7_75t_R _13067_ (.A1(_00376_),
    .A2(_09201_),
    .B(_09233_),
    .Y(_02817_));
 AO221x1_ASAP7_75t_R _13068_ (.A1(_00271_),
    .A2(_09203_),
    .B1(_09205_),
    .B2(_01936_),
    .C(_09211_),
    .Y(_09234_));
 AOI21x1_ASAP7_75t_R _13069_ (.A1(_00375_),
    .A2(_09201_),
    .B(_09234_),
    .Y(_02818_));
 NAND2x1_ASAP7_75t_R _13070_ (.A(_09163_),
    .B(_09167_),
    .Y(_09235_));
 NAND2x1_ASAP7_75t_R _13071_ (.A(_09167_),
    .B(_09156_),
    .Y(_09236_));
 OA21x2_ASAP7_75t_R _13072_ (.A1(_09172_),
    .A2(_09173_),
    .B(_09188_),
    .Y(_09237_));
 OA211x2_ASAP7_75t_R _13073_ (.A1(_09172_),
    .A2(_09173_),
    .B(_09188_),
    .C(_00003_),
    .Y(_09238_));
 OA222x2_ASAP7_75t_R _13074_ (.A1(_09164_),
    .A2(_09235_),
    .B1(_09236_),
    .B2(_09237_),
    .C1(_09238_),
    .C2(_09163_),
    .Y(_09239_));
 AOI21x1_ASAP7_75t_R _13075_ (.A1(_09160_),
    .A2(_09161_),
    .B(_09165_),
    .Y(_09240_));
 AO221x1_ASAP7_75t_R _13076_ (.A1(_09193_),
    .A2(_09183_),
    .B1(_09239_),
    .B2(_09240_),
    .C(_09191_),
    .Y(_09241_));
 BUFx6f_ASAP7_75t_R _13077_ (.A(_09241_),
    .Y(_09242_));
 NOR2x1_ASAP7_75t_R _13078_ (.A(_00377_),
    .B(_00378_),
    .Y(_09243_));
 OA21x2_ASAP7_75t_R _13079_ (.A1(_09243_),
    .A2(_09178_),
    .B(_09190_),
    .Y(_09244_));
 AOI221x1_ASAP7_75t_R _13080_ (.A1(_09169_),
    .A2(_09190_),
    .B1(_09193_),
    .B2(_09243_),
    .C(_09164_),
    .Y(_09245_));
 NAND3x1_ASAP7_75t_R _13081_ (.A(_09197_),
    .B(_09198_),
    .C(_09245_),
    .Y(_09246_));
 OR3x2_ASAP7_75t_R _13082_ (.A(_09242_),
    .B(_09244_),
    .C(_09246_),
    .Y(_09247_));
 BUFx12f_ASAP7_75t_R _13083_ (.A(_09247_),
    .Y(_09248_));
 NOR2x1_ASAP7_75t_R _13084_ (.A(_01949_),
    .B(_09248_),
    .Y(_09249_));
 INVx1_ASAP7_75t_R _13085_ (.A(_00388_),
    .Y(_09250_));
 BUFx6f_ASAP7_75t_R _13086_ (.A(_09242_),
    .Y(_09251_));
 BUFx6f_ASAP7_75t_R _13087_ (.A(_09247_),
    .Y(_09252_));
 BUFx6f_ASAP7_75t_R _13088_ (.A(_09242_),
    .Y(_09253_));
 NAND2x1_ASAP7_75t_R _13089_ (.A(_00284_),
    .B(_09253_),
    .Y(_09254_));
 OA211x2_ASAP7_75t_R _13090_ (.A1(_09250_),
    .A2(_09251_),
    .B(_09252_),
    .C(_09254_),
    .Y(_09255_));
 BUFx6f_ASAP7_75t_R _13091_ (.A(_08665_),
    .Y(_09256_));
 OA21x2_ASAP7_75t_R _13092_ (.A1(_09249_),
    .A2(_09255_),
    .B(_09256_),
    .Y(_02819_));
 NOR2x1_ASAP7_75t_R _13093_ (.A(_01948_),
    .B(_09248_),
    .Y(_09257_));
 INVx1_ASAP7_75t_R _13094_ (.A(_00387_),
    .Y(_09258_));
 NAND2x1_ASAP7_75t_R _13095_ (.A(_00283_),
    .B(_09253_),
    .Y(_09259_));
 OA211x2_ASAP7_75t_R _13096_ (.A1(_09258_),
    .A2(_09251_),
    .B(_09252_),
    .C(_09259_),
    .Y(_09260_));
 OA21x2_ASAP7_75t_R _13097_ (.A1(_09257_),
    .A2(_09260_),
    .B(_09256_),
    .Y(_02820_));
 NOR2x1_ASAP7_75t_R _13098_ (.A(_01947_),
    .B(_09248_),
    .Y(_09261_));
 INVx1_ASAP7_75t_R _13099_ (.A(_00386_),
    .Y(_09262_));
 NAND2x1_ASAP7_75t_R _13100_ (.A(_00282_),
    .B(_09253_),
    .Y(_09263_));
 OA211x2_ASAP7_75t_R _13101_ (.A1(_09262_),
    .A2(_09251_),
    .B(_09252_),
    .C(_09263_),
    .Y(_09264_));
 OA21x2_ASAP7_75t_R _13102_ (.A1(_09261_),
    .A2(_09264_),
    .B(_09256_),
    .Y(_02821_));
 NOR2x1_ASAP7_75t_R _13103_ (.A(_01946_),
    .B(_09248_),
    .Y(_09265_));
 INVx1_ASAP7_75t_R _13104_ (.A(_00385_),
    .Y(_09266_));
 NAND2x1_ASAP7_75t_R _13105_ (.A(_00281_),
    .B(_09253_),
    .Y(_09267_));
 OA211x2_ASAP7_75t_R _13106_ (.A1(_09266_),
    .A2(_09251_),
    .B(_09252_),
    .C(_09267_),
    .Y(_09268_));
 OA21x2_ASAP7_75t_R _13107_ (.A1(_09265_),
    .A2(_09268_),
    .B(_09256_),
    .Y(_02822_));
 NOR2x1_ASAP7_75t_R _13108_ (.A(_01945_),
    .B(_09248_),
    .Y(_09269_));
 INVx1_ASAP7_75t_R _13109_ (.A(_00384_),
    .Y(_09270_));
 NAND2x1_ASAP7_75t_R _13110_ (.A(_00280_),
    .B(_09253_),
    .Y(_09271_));
 OA211x2_ASAP7_75t_R _13111_ (.A1(_09270_),
    .A2(_09251_),
    .B(_09252_),
    .C(_09271_),
    .Y(_09272_));
 OA21x2_ASAP7_75t_R _13112_ (.A1(_09269_),
    .A2(_09272_),
    .B(_09256_),
    .Y(_02823_));
 NOR2x1_ASAP7_75t_R _13113_ (.A(_09189_),
    .B(_09251_),
    .Y(_09273_));
 AO21x1_ASAP7_75t_R _13114_ (.A1(_00279_),
    .A2(_09251_),
    .B(_09273_),
    .Y(_09274_));
 BUFx12f_ASAP7_75t_R _13115_ (.A(_09118_),
    .Y(_09275_));
 AOI21x1_ASAP7_75t_R _13116_ (.A1(_09248_),
    .A2(_09274_),
    .B(_09275_),
    .Y(_02824_));
 NOR2x1_ASAP7_75t_R _13117_ (.A(_01943_),
    .B(_09248_),
    .Y(_09276_));
 NAND2x1_ASAP7_75t_R _13118_ (.A(_00278_),
    .B(_09253_),
    .Y(_09277_));
 OA211x2_ASAP7_75t_R _13119_ (.A1(_09214_),
    .A2(_09251_),
    .B(_09252_),
    .C(_09277_),
    .Y(_09278_));
 OA21x2_ASAP7_75t_R _13120_ (.A1(_09276_),
    .A2(_09278_),
    .B(_09256_),
    .Y(_02825_));
 NOR2x1_ASAP7_75t_R _13121_ (.A(_01942_),
    .B(_09248_),
    .Y(_09279_));
 NAND2x1_ASAP7_75t_R _13122_ (.A(_00277_),
    .B(_09242_),
    .Y(_09280_));
 OA211x2_ASAP7_75t_R _13123_ (.A1(_09217_),
    .A2(_09251_),
    .B(_09252_),
    .C(_09280_),
    .Y(_09281_));
 OA21x2_ASAP7_75t_R _13124_ (.A1(_09279_),
    .A2(_09281_),
    .B(_09256_),
    .Y(_02826_));
 NOR2x1_ASAP7_75t_R _13125_ (.A(_01941_),
    .B(_09248_),
    .Y(_09282_));
 INVx1_ASAP7_75t_R _13126_ (.A(_00380_),
    .Y(_09283_));
 NAND2x1_ASAP7_75t_R _13127_ (.A(_00276_),
    .B(_09242_),
    .Y(_09284_));
 OA211x2_ASAP7_75t_R _13128_ (.A1(_09283_),
    .A2(_09253_),
    .B(_09252_),
    .C(_09284_),
    .Y(_09285_));
 OA21x2_ASAP7_75t_R _13129_ (.A1(_09282_),
    .A2(_09285_),
    .B(_09256_),
    .Y(_02827_));
 NOR2x1_ASAP7_75t_R _13130_ (.A(_01940_),
    .B(_09248_),
    .Y(_09286_));
 INVx1_ASAP7_75t_R _13131_ (.A(_00379_),
    .Y(_09287_));
 NAND2x1_ASAP7_75t_R _13132_ (.A(_00275_),
    .B(_09242_),
    .Y(_09288_));
 OA211x2_ASAP7_75t_R _13133_ (.A1(_09287_),
    .A2(_09253_),
    .B(_09247_),
    .C(_09288_),
    .Y(_09289_));
 OA21x2_ASAP7_75t_R _13134_ (.A1(_09286_),
    .A2(_09289_),
    .B(_09256_),
    .Y(_02828_));
 AO22x1_ASAP7_75t_R _13135_ (.A1(_09193_),
    .A2(_09183_),
    .B1(_09239_),
    .B2(_09240_),
    .Y(_09290_));
 AND3x1_ASAP7_75t_R _13136_ (.A(_08582_),
    .B(_09177_),
    .C(_09290_),
    .Y(_02829_));
 NOR2x1_ASAP7_75t_R _13137_ (.A(_09251_),
    .B(_09244_),
    .Y(_09291_));
 AOI21x1_ASAP7_75t_R _13138_ (.A1(_09291_),
    .A2(_09246_),
    .B(_09275_),
    .Y(_02830_));
 NOR2x1_ASAP7_75t_R _13139_ (.A(_01937_),
    .B(_09252_),
    .Y(_09292_));
 INVx1_ASAP7_75t_R _13140_ (.A(_00376_),
    .Y(_09293_));
 NAND2x1_ASAP7_75t_R _13141_ (.A(_00272_),
    .B(_09242_),
    .Y(_09294_));
 OA211x2_ASAP7_75t_R _13142_ (.A1(_09293_),
    .A2(_09253_),
    .B(_09247_),
    .C(_09294_),
    .Y(_09295_));
 OA21x2_ASAP7_75t_R _13143_ (.A1(_09292_),
    .A2(_09295_),
    .B(_09256_),
    .Y(_02831_));
 NOR2x1_ASAP7_75t_R _13144_ (.A(_01936_),
    .B(_09252_),
    .Y(_09296_));
 INVx1_ASAP7_75t_R _13145_ (.A(_00375_),
    .Y(_09297_));
 NAND2x1_ASAP7_75t_R _13146_ (.A(_00271_),
    .B(_09242_),
    .Y(_09298_));
 OA211x2_ASAP7_75t_R _13147_ (.A1(_09297_),
    .A2(_09253_),
    .B(_09247_),
    .C(_09298_),
    .Y(_09299_));
 BUFx12f_ASAP7_75t_R _13148_ (.A(_08665_),
    .Y(_09300_));
 OA21x2_ASAP7_75t_R _13149_ (.A1(_09296_),
    .A2(_09299_),
    .B(_09300_),
    .Y(_02832_));
 OA21x2_ASAP7_75t_R _13150_ (.A1(_09194_),
    .A2(_09245_),
    .B(_09197_),
    .Y(_09301_));
 AOI21x1_ASAP7_75t_R _13151_ (.A1(_09167_),
    .A2(_09301_),
    .B(_01938_),
    .Y(_09302_));
 NOR2x1_ASAP7_75t_R _13152_ (.A(_08683_),
    .B(_09302_),
    .Y(_09303_));
 BUFx6f_ASAP7_75t_R _13153_ (.A(_09303_),
    .Y(_09304_));
 OA31x2_ASAP7_75t_R _13154_ (.A1(_09243_),
    .A2(_09168_),
    .A3(_09170_),
    .B1(_09237_),
    .Y(_09305_));
 AO21x2_ASAP7_75t_R _13155_ (.A1(_09177_),
    .A2(_09239_),
    .B(_09169_),
    .Y(_09306_));
 NOR2x1_ASAP7_75t_R _13156_ (.A(_09305_),
    .B(_09306_),
    .Y(_09307_));
 BUFx6f_ASAP7_75t_R _13157_ (.A(_09307_),
    .Y(_09308_));
 NAND2x1_ASAP7_75t_R _13158_ (.A(_00284_),
    .B(_09308_),
    .Y(_09309_));
 OR2x6_ASAP7_75t_R _13159_ (.A(_09305_),
    .B(_09306_),
    .Y(_09310_));
 BUFx6f_ASAP7_75t_R _13160_ (.A(_09310_),
    .Y(_09311_));
 NAND2x1_ASAP7_75t_R _13161_ (.A(_00388_),
    .B(_09311_),
    .Y(_09312_));
 BUFx3_ASAP7_75t_R _13162_ (.A(_09302_),
    .Y(_09313_));
 BUFx12f_ASAP7_75t_R _13163_ (.A(_08578_),
    .Y(_09314_));
 NOR2x1_ASAP7_75t_R _13164_ (.A(_09314_),
    .B(_01949_),
    .Y(_09315_));
 AO32x1_ASAP7_75t_R _13165_ (.A1(_09304_),
    .A2(_09309_),
    .A3(_09312_),
    .B1(_09313_),
    .B2(_09315_),
    .Y(_02833_));
 NAND2x1_ASAP7_75t_R _13166_ (.A(_00283_),
    .B(_09308_),
    .Y(_09316_));
 NAND2x1_ASAP7_75t_R _13167_ (.A(_00387_),
    .B(_09311_),
    .Y(_09317_));
 BUFx12f_ASAP7_75t_R _13168_ (.A(_08656_),
    .Y(_09318_));
 NOR2x1_ASAP7_75t_R _13169_ (.A(_09318_),
    .B(_01948_),
    .Y(_09319_));
 AO32x1_ASAP7_75t_R _13170_ (.A1(_09304_),
    .A2(_09316_),
    .A3(_09317_),
    .B1(_09313_),
    .B2(_09319_),
    .Y(_02834_));
 NAND2x1_ASAP7_75t_R _13171_ (.A(_00282_),
    .B(_09308_),
    .Y(_09320_));
 NAND2x1_ASAP7_75t_R _13172_ (.A(_00386_),
    .B(_09311_),
    .Y(_09321_));
 NOR2x1_ASAP7_75t_R _13173_ (.A(_09318_),
    .B(_01947_),
    .Y(_09322_));
 AO32x1_ASAP7_75t_R _13174_ (.A1(_09304_),
    .A2(_09320_),
    .A3(_09321_),
    .B1(_09313_),
    .B2(_09322_),
    .Y(_02835_));
 NAND2x1_ASAP7_75t_R _13175_ (.A(_00281_),
    .B(_09308_),
    .Y(_09323_));
 NAND2x1_ASAP7_75t_R _13176_ (.A(_00385_),
    .B(_09311_),
    .Y(_09324_));
 NOR2x1_ASAP7_75t_R _13177_ (.A(_09318_),
    .B(_01946_),
    .Y(_09325_));
 AO32x2_ASAP7_75t_R _13178_ (.A1(_09304_),
    .A2(_09323_),
    .A3(_09324_),
    .B1(_09313_),
    .B2(_09325_),
    .Y(_02836_));
 NAND2x1_ASAP7_75t_R _13179_ (.A(_00280_),
    .B(_09308_),
    .Y(_09326_));
 NAND2x1_ASAP7_75t_R _13180_ (.A(_00384_),
    .B(_09311_),
    .Y(_09327_));
 NOR2x1_ASAP7_75t_R _13181_ (.A(_09318_),
    .B(_01945_),
    .Y(_09328_));
 AO32x2_ASAP7_75t_R _13182_ (.A1(_09304_),
    .A2(_09326_),
    .A3(_09327_),
    .B1(_09313_),
    .B2(_09328_),
    .Y(_02837_));
 OR3x1_ASAP7_75t_R _13183_ (.A(_09184_),
    .B(_09305_),
    .C(_09306_),
    .Y(_09329_));
 NAND2x1_ASAP7_75t_R _13184_ (.A(_00383_),
    .B(_09311_),
    .Y(_09330_));
 NOR2x1_ASAP7_75t_R _13185_ (.A(_08811_),
    .B(_09164_),
    .Y(_09331_));
 AO32x1_ASAP7_75t_R _13186_ (.A1(_09304_),
    .A2(_09329_),
    .A3(_09330_),
    .B1(_09331_),
    .B2(_09313_),
    .Y(_02838_));
 NAND2x1_ASAP7_75t_R _13187_ (.A(_00278_),
    .B(_09308_),
    .Y(_09332_));
 NAND2x1_ASAP7_75t_R _13188_ (.A(_00382_),
    .B(_09311_),
    .Y(_09333_));
 NOR2x1_ASAP7_75t_R _13189_ (.A(_09318_),
    .B(_01943_),
    .Y(_09334_));
 AO32x1_ASAP7_75t_R _13190_ (.A1(_09304_),
    .A2(_09332_),
    .A3(_09333_),
    .B1(_09313_),
    .B2(_09334_),
    .Y(_02839_));
 NAND2x1_ASAP7_75t_R _13191_ (.A(_00277_),
    .B(_09308_),
    .Y(_09335_));
 NAND2x1_ASAP7_75t_R _13192_ (.A(_00381_),
    .B(_09311_),
    .Y(_09336_));
 NOR2x1_ASAP7_75t_R _13193_ (.A(_09318_),
    .B(_01942_),
    .Y(_09337_));
 AO32x1_ASAP7_75t_R _13194_ (.A1(_09304_),
    .A2(_09335_),
    .A3(_09336_),
    .B1(_09313_),
    .B2(_09337_),
    .Y(_02840_));
 NAND2x1_ASAP7_75t_R _13195_ (.A(_00276_),
    .B(_09308_),
    .Y(_09338_));
 NAND2x1_ASAP7_75t_R _13196_ (.A(_00380_),
    .B(_09311_),
    .Y(_09339_));
 AO32x1_ASAP7_75t_R _13197_ (.A1(_09304_),
    .A2(_09338_),
    .A3(_09339_),
    .B1(_09313_),
    .B2(_09224_),
    .Y(_02841_));
 NAND2x1_ASAP7_75t_R _13198_ (.A(_00275_),
    .B(_09308_),
    .Y(_09340_));
 NAND2x1_ASAP7_75t_R _13199_ (.A(_00379_),
    .B(_09311_),
    .Y(_09341_));
 AO32x1_ASAP7_75t_R _13200_ (.A1(_09304_),
    .A2(_09340_),
    .A3(_09341_),
    .B1(_09302_),
    .B2(_09227_),
    .Y(_02842_));
 OR3x1_ASAP7_75t_R _13201_ (.A(_08657_),
    .B(_09235_),
    .C(_09301_),
    .Y(_09342_));
 INVx1_ASAP7_75t_R _13202_ (.A(_09342_),
    .Y(_02843_));
 NAND2x1_ASAP7_75t_R _13203_ (.A(_09177_),
    .B(_09239_),
    .Y(_09343_));
 AO21x1_ASAP7_75t_R _13204_ (.A1(_09240_),
    .A2(_09343_),
    .B(_09305_),
    .Y(_09344_));
 OA21x2_ASAP7_75t_R _13205_ (.A1(_09313_),
    .A2(_09344_),
    .B(_09300_),
    .Y(_02844_));
 NAND2x1_ASAP7_75t_R _13206_ (.A(_00272_),
    .B(_09308_),
    .Y(_09345_));
 NAND2x1_ASAP7_75t_R _13207_ (.A(_00376_),
    .B(_09310_),
    .Y(_09346_));
 NOR2x1_ASAP7_75t_R _13208_ (.A(_09318_),
    .B(_01937_),
    .Y(_09347_));
 AO32x1_ASAP7_75t_R _13209_ (.A1(_09303_),
    .A2(_09345_),
    .A3(_09346_),
    .B1(_09302_),
    .B2(_09347_),
    .Y(_02845_));
 NAND2x1_ASAP7_75t_R _13210_ (.A(_00271_),
    .B(_09307_),
    .Y(_09348_));
 NAND2x1_ASAP7_75t_R _13211_ (.A(_00375_),
    .B(_09310_),
    .Y(_09349_));
 NOR2x1_ASAP7_75t_R _13212_ (.A(_09318_),
    .B(_01936_),
    .Y(_09350_));
 AO32x1_ASAP7_75t_R _13213_ (.A1(_09303_),
    .A2(_09348_),
    .A3(_09349_),
    .B1(_09302_),
    .B2(_09350_),
    .Y(_02846_));
 AND2x2_ASAP7_75t_R _13214_ (.A(_08723_),
    .B(_00004_),
    .Y(_02847_));
 BUFx6f_ASAP7_75t_R _13215_ (.A(_00065_),
    .Y(_09351_));
 NOR2x1_ASAP7_75t_R _13216_ (.A(_09351_),
    .B(_00066_),
    .Y(_09352_));
 INVx2_ASAP7_75t_R _13217_ (.A(_00171_),
    .Y(_09353_));
 NAND2x1_ASAP7_75t_R _13218_ (.A(_00173_),
    .B(_00174_),
    .Y(_09354_));
 INVx1_ASAP7_75t_R _13219_ (.A(_00169_),
    .Y(_09355_));
 OA31x2_ASAP7_75t_R _13220_ (.A1(_09353_),
    .A2(_00172_),
    .A3(_09354_),
    .B1(_09355_),
    .Y(_09356_));
 BUFx6f_ASAP7_75t_R _13221_ (.A(_09356_),
    .Y(_09357_));
 INVx2_ASAP7_75t_R _13222_ (.A(_00068_),
    .Y(_09358_));
 INVx2_ASAP7_75t_R _13223_ (.A(_01911_),
    .Y(_09359_));
 AND2x4_ASAP7_75t_R _13224_ (.A(_00069_),
    .B(_00070_),
    .Y(_09360_));
 AND4x1_ASAP7_75t_R _13225_ (.A(_00067_),
    .B(_09358_),
    .C(_09359_),
    .D(_09360_),
    .Y(_09361_));
 INVx2_ASAP7_75t_R _13226_ (.A(_00067_),
    .Y(_09362_));
 NAND2x1_ASAP7_75t_R _13227_ (.A(_00069_),
    .B(_00070_),
    .Y(_09363_));
 OR4x1_ASAP7_75t_R _13228_ (.A(_09362_),
    .B(_00068_),
    .C(_00071_),
    .D(_09363_),
    .Y(_09364_));
 BUFx6f_ASAP7_75t_R _13229_ (.A(_01910_),
    .Y(_09365_));
 NOR2x1_ASAP7_75t_R _13230_ (.A(_09365_),
    .B(_09351_),
    .Y(_09366_));
 OA211x2_ASAP7_75t_R _13231_ (.A1(_01916_),
    .A2(_09361_),
    .B(_09364_),
    .C(_09366_),
    .Y(_09367_));
 INVx1_ASAP7_75t_R _13232_ (.A(_09351_),
    .Y(_09368_));
 OA31x2_ASAP7_75t_R _13233_ (.A1(_09362_),
    .A2(_00068_),
    .A3(_09363_),
    .B1(_09368_),
    .Y(_09369_));
 AND4x1_ASAP7_75t_R _13234_ (.A(_09365_),
    .B(_00004_),
    .C(_09357_),
    .D(_09369_),
    .Y(_09370_));
 NOR2x2_ASAP7_75t_R _13235_ (.A(_00169_),
    .B(_00170_),
    .Y(_09371_));
 AND5x1_ASAP7_75t_R _13236_ (.A(_09368_),
    .B(_00067_),
    .C(_09358_),
    .D(_00071_),
    .E(_09360_),
    .Y(_09372_));
 AO21x1_ASAP7_75t_R _13237_ (.A1(_01916_),
    .A2(_09371_),
    .B(_09359_),
    .Y(_09373_));
 OA31x2_ASAP7_75t_R _13238_ (.A1(_09362_),
    .A2(_00068_),
    .A3(_09363_),
    .B1(_09366_),
    .Y(_09374_));
 AO22x2_ASAP7_75t_R _13239_ (.A1(_09371_),
    .A2(_09372_),
    .B1(_09373_),
    .B2(_09374_),
    .Y(_09375_));
 AOI211x1_ASAP7_75t_R _13240_ (.A1(_09357_),
    .A2(_09367_),
    .B(_09370_),
    .C(_09375_),
    .Y(_09376_));
 INVx2_ASAP7_75t_R _13241_ (.A(_09365_),
    .Y(_09377_));
 INVx1_ASAP7_75t_R _13242_ (.A(_00004_),
    .Y(_09378_));
 INVx3_ASAP7_75t_R _13243_ (.A(_01916_),
    .Y(_09379_));
 AO32x1_ASAP7_75t_R _13244_ (.A1(_09365_),
    .A2(_09378_),
    .A3(_09369_),
    .B1(_09374_),
    .B2(_09379_),
    .Y(_09380_));
 AO21x2_ASAP7_75t_R _13245_ (.A1(_09377_),
    .A2(_09359_),
    .B(_09380_),
    .Y(_09381_));
 OR5x2_ASAP7_75t_R _13246_ (.A(_00169_),
    .B(_09353_),
    .C(_00172_),
    .D(_00175_),
    .E(_09354_),
    .Y(_09382_));
 NAND3x1_ASAP7_75t_R _13247_ (.A(_09377_),
    .B(_09379_),
    .C(_09357_),
    .Y(_09383_));
 OR2x6_ASAP7_75t_R _13248_ (.A(_09351_),
    .B(_00066_),
    .Y(_09384_));
 BUFx6f_ASAP7_75t_R _13249_ (.A(_09384_),
    .Y(_09385_));
 AND3x1_ASAP7_75t_R _13250_ (.A(_00067_),
    .B(_09358_),
    .C(_09360_),
    .Y(_09386_));
 AND2x2_ASAP7_75t_R _13251_ (.A(_01911_),
    .B(_01916_),
    .Y(_09387_));
 OR5x1_ASAP7_75t_R _13252_ (.A(_09365_),
    .B(_09351_),
    .C(_09386_),
    .D(_09382_),
    .E(_09387_),
    .Y(_09388_));
 AOI22x1_ASAP7_75t_R _13253_ (.A1(_09382_),
    .A2(_09383_),
    .B1(_09385_),
    .B2(_09388_),
    .Y(_09389_));
 AOI211x1_ASAP7_75t_R _13254_ (.A1(_09357_),
    .A2(_09381_),
    .B(_09389_),
    .C(_09371_),
    .Y(_09390_));
 OA211x2_ASAP7_75t_R _13255_ (.A1(_09352_),
    .A2(_09376_),
    .B(_09372_),
    .C(_09390_),
    .Y(_09391_));
 BUFx6f_ASAP7_75t_R _13256_ (.A(_09391_),
    .Y(_09392_));
 INVx1_ASAP7_75t_R _13257_ (.A(_00170_),
    .Y(_09393_));
 AO211x2_ASAP7_75t_R _13258_ (.A1(_09357_),
    .A2(_09367_),
    .B(_09370_),
    .C(_09375_),
    .Y(_09394_));
 INVx2_ASAP7_75t_R _13259_ (.A(_00071_),
    .Y(_09395_));
 OR3x2_ASAP7_75t_R _13260_ (.A(_09362_),
    .B(_00068_),
    .C(_09363_),
    .Y(_09396_));
 OR3x1_ASAP7_75t_R _13261_ (.A(_09351_),
    .B(_09395_),
    .C(_09396_),
    .Y(_09397_));
 AO21x2_ASAP7_75t_R _13262_ (.A1(_09385_),
    .A2(_09394_),
    .B(_09397_),
    .Y(_09398_));
 OR4x1_ASAP7_75t_R _13263_ (.A(_09351_),
    .B(_09395_),
    .C(_00169_),
    .D(_00175_),
    .Y(_09399_));
 OA33x2_ASAP7_75t_R _13264_ (.A1(_00169_),
    .A2(_00170_),
    .A3(_09379_),
    .B1(_09356_),
    .B2(_09396_),
    .B3(_09399_),
    .Y(_09400_));
 OR3x1_ASAP7_75t_R _13265_ (.A(_09351_),
    .B(_09395_),
    .C(_09379_),
    .Y(_09401_));
 OR3x1_ASAP7_75t_R _13266_ (.A(_09357_),
    .B(_09396_),
    .C(_09401_),
    .Y(_09402_));
 AND2x4_ASAP7_75t_R _13267_ (.A(_09377_),
    .B(_01911_),
    .Y(_09403_));
 OA211x2_ASAP7_75t_R _13268_ (.A1(_09382_),
    .A2(_09384_),
    .B(_09403_),
    .C(_01916_),
    .Y(_09404_));
 AND3x4_ASAP7_75t_R _13269_ (.A(_09400_),
    .B(_09402_),
    .C(_09404_),
    .Y(_09405_));
 INVx1_ASAP7_75t_R _13270_ (.A(_09405_),
    .Y(_09406_));
 AO21x1_ASAP7_75t_R _13271_ (.A1(_09357_),
    .A2(_09381_),
    .B(_09389_),
    .Y(_09407_));
 AO221x1_ASAP7_75t_R _13272_ (.A1(_09355_),
    .A2(_09393_),
    .B1(_09398_),
    .B2(_09406_),
    .C(_09407_),
    .Y(_09408_));
 BUFx6f_ASAP7_75t_R _13273_ (.A(_09408_),
    .Y(_09409_));
 AND4x1_ASAP7_75t_R _13274_ (.A(_09397_),
    .B(_09400_),
    .C(_09402_),
    .D(_09404_),
    .Y(_09410_));
 AO31x2_ASAP7_75t_R _13275_ (.A1(_09385_),
    .A2(_09394_),
    .A3(_09405_),
    .B(_09410_),
    .Y(_09411_));
 AO21x1_ASAP7_75t_R _13276_ (.A1(_01921_),
    .A2(_09411_),
    .B(_08579_),
    .Y(_09412_));
 AOI221x1_ASAP7_75t_R _13277_ (.A1(_00076_),
    .A2(_09392_),
    .B1(_09409_),
    .B2(_00180_),
    .C(_09412_),
    .Y(_02848_));
 AO21x1_ASAP7_75t_R _13278_ (.A1(_01920_),
    .A2(_09411_),
    .B(_08579_),
    .Y(_09413_));
 AOI221x1_ASAP7_75t_R _13279_ (.A1(_00075_),
    .A2(_09392_),
    .B1(_09409_),
    .B2(_00179_),
    .C(_09413_),
    .Y(_02849_));
 AO21x1_ASAP7_75t_R _13280_ (.A1(_01919_),
    .A2(_09411_),
    .B(_08579_),
    .Y(_09414_));
 AOI221x1_ASAP7_75t_R _13281_ (.A1(_00074_),
    .A2(_09392_),
    .B1(_09409_),
    .B2(_00178_),
    .C(_09414_),
    .Y(_02850_));
 AO21x1_ASAP7_75t_R _13282_ (.A1(_01918_),
    .A2(_09411_),
    .B(_08579_),
    .Y(_09415_));
 AOI221x1_ASAP7_75t_R _13283_ (.A1(_00073_),
    .A2(_09392_),
    .B1(_09409_),
    .B2(_00177_),
    .C(_09415_),
    .Y(_02851_));
 AO21x1_ASAP7_75t_R _13284_ (.A1(_01917_),
    .A2(_09411_),
    .B(_08579_),
    .Y(_09416_));
 AOI221x1_ASAP7_75t_R _13285_ (.A1(_00072_),
    .A2(_09392_),
    .B1(_09409_),
    .B2(_00176_),
    .C(_09416_),
    .Y(_02852_));
 NOR2x1_ASAP7_75t_R _13286_ (.A(_08578_),
    .B(_00175_),
    .Y(_09417_));
 AND2x2_ASAP7_75t_R _13287_ (.A(_09409_),
    .B(_09417_),
    .Y(_02853_));
 INVx1_ASAP7_75t_R _13288_ (.A(_00174_),
    .Y(_09418_));
 INVx2_ASAP7_75t_R _13289_ (.A(_01915_),
    .Y(_09419_));
 AND3x1_ASAP7_75t_R _13290_ (.A(_08584_),
    .B(_09419_),
    .C(_09405_),
    .Y(_09420_));
 AO32x1_ASAP7_75t_R _13291_ (.A1(_08585_),
    .A2(_09418_),
    .A3(_09409_),
    .B1(_09420_),
    .B2(_09398_),
    .Y(_02854_));
 INVx1_ASAP7_75t_R _13292_ (.A(_00173_),
    .Y(_09421_));
 INVx2_ASAP7_75t_R _13293_ (.A(_01914_),
    .Y(_09422_));
 AND3x1_ASAP7_75t_R _13294_ (.A(_08584_),
    .B(_09422_),
    .C(_09405_),
    .Y(_09423_));
 AO32x1_ASAP7_75t_R _13295_ (.A1(_08585_),
    .A2(_09421_),
    .A3(_09408_),
    .B1(_09423_),
    .B2(_09398_),
    .Y(_02855_));
 AOI221x1_ASAP7_75t_R _13296_ (.A1(_00172_),
    .A2(_09409_),
    .B1(_09411_),
    .B2(_01913_),
    .C(_09145_),
    .Y(_02856_));
 INVx2_ASAP7_75t_R _13297_ (.A(_01912_),
    .Y(_09424_));
 AND3x1_ASAP7_75t_R _13298_ (.A(_08584_),
    .B(_09424_),
    .C(_09405_),
    .Y(_09425_));
 AO32x1_ASAP7_75t_R _13299_ (.A1(_08585_),
    .A2(_09353_),
    .A3(_09408_),
    .B1(_09425_),
    .B2(_09398_),
    .Y(_02857_));
 OR2x2_ASAP7_75t_R _13300_ (.A(_00169_),
    .B(_00170_),
    .Y(_09426_));
 AND3x1_ASAP7_75t_R _13301_ (.A(_08582_),
    .B(_09426_),
    .C(_09407_),
    .Y(_02858_));
 AND3x1_ASAP7_75t_R _13302_ (.A(_09390_),
    .B(_09398_),
    .C(_09406_),
    .Y(_09427_));
 NOR2x1_ASAP7_75t_R _13303_ (.A(_08942_),
    .B(_09427_),
    .Y(_02859_));
 AO21x1_ASAP7_75t_R _13304_ (.A1(_01909_),
    .A2(_09411_),
    .B(_08579_),
    .Y(_09428_));
 AOI221x1_ASAP7_75t_R _13305_ (.A1(_00064_),
    .A2(_09392_),
    .B1(_09409_),
    .B2(_00168_),
    .C(_09428_),
    .Y(_02860_));
 AO21x1_ASAP7_75t_R _13306_ (.A1(_01908_),
    .A2(_09411_),
    .B(_08579_),
    .Y(_09429_));
 AOI221x1_ASAP7_75t_R _13307_ (.A1(_00063_),
    .A2(_09392_),
    .B1(_09409_),
    .B2(_00167_),
    .C(_09429_),
    .Y(_02861_));
 INVx1_ASAP7_75t_R _13308_ (.A(_01921_),
    .Y(_09430_));
 OR3x1_ASAP7_75t_R _13309_ (.A(_09351_),
    .B(_09395_),
    .C(_09426_),
    .Y(_09431_));
 OA221x2_ASAP7_75t_R _13310_ (.A1(_09369_),
    .A2(_09382_),
    .B1(_09431_),
    .B2(_09396_),
    .C(_09384_),
    .Y(_09432_));
 NOR2x1_ASAP7_75t_R _13311_ (.A(_09371_),
    .B(_09387_),
    .Y(_09433_));
 AO221x1_ASAP7_75t_R _13312_ (.A1(_09426_),
    .A2(_09352_),
    .B1(_09433_),
    .B2(_09374_),
    .C(_09382_),
    .Y(_09434_));
 AND4x1_ASAP7_75t_R _13313_ (.A(_09379_),
    .B(_09403_),
    .C(_09432_),
    .D(_09434_),
    .Y(_09435_));
 BUFx6f_ASAP7_75t_R _13314_ (.A(_09435_),
    .Y(_09436_));
 NAND2x1_ASAP7_75t_R _13315_ (.A(_09430_),
    .B(_09436_),
    .Y(_09437_));
 NAND2x1_ASAP7_75t_R _13316_ (.A(_09385_),
    .B(_09376_),
    .Y(_09438_));
 BUFx6f_ASAP7_75t_R _13317_ (.A(_09438_),
    .Y(_09439_));
 BUFx6f_ASAP7_75t_R _13318_ (.A(_09385_),
    .Y(_09440_));
 AND2x2_ASAP7_75t_R _13319_ (.A(_00180_),
    .B(_09440_),
    .Y(_09441_));
 BUFx6f_ASAP7_75t_R _13320_ (.A(_09376_),
    .Y(_09442_));
 BUFx6f_ASAP7_75t_R _13321_ (.A(_09435_),
    .Y(_09443_));
 AO221x1_ASAP7_75t_R _13322_ (.A1(_00076_),
    .A2(_09439_),
    .B1(_09441_),
    .B2(_09442_),
    .C(_09443_),
    .Y(_09444_));
 AOI21x1_ASAP7_75t_R _13323_ (.A1(_09437_),
    .A2(_09444_),
    .B(_09275_),
    .Y(_02862_));
 INVx1_ASAP7_75t_R _13324_ (.A(_01920_),
    .Y(_09445_));
 NAND2x1_ASAP7_75t_R _13325_ (.A(_09445_),
    .B(_09436_),
    .Y(_09446_));
 AND2x2_ASAP7_75t_R _13326_ (.A(_00179_),
    .B(_09440_),
    .Y(_09447_));
 AO221x1_ASAP7_75t_R _13327_ (.A1(_00075_),
    .A2(_09439_),
    .B1(_09447_),
    .B2(_09442_),
    .C(_09443_),
    .Y(_09448_));
 AOI21x1_ASAP7_75t_R _13328_ (.A1(_09446_),
    .A2(_09448_),
    .B(_09275_),
    .Y(_02863_));
 INVx1_ASAP7_75t_R _13329_ (.A(_01919_),
    .Y(_09449_));
 NAND2x1_ASAP7_75t_R _13330_ (.A(_09449_),
    .B(_09436_),
    .Y(_09450_));
 AND2x2_ASAP7_75t_R _13331_ (.A(_00178_),
    .B(_09440_),
    .Y(_09451_));
 AO221x1_ASAP7_75t_R _13332_ (.A1(_00074_),
    .A2(_09439_),
    .B1(_09451_),
    .B2(_09442_),
    .C(_09443_),
    .Y(_09452_));
 AOI21x1_ASAP7_75t_R _13333_ (.A1(_09450_),
    .A2(_09452_),
    .B(_09275_),
    .Y(_02864_));
 INVx1_ASAP7_75t_R _13334_ (.A(_01918_),
    .Y(_09453_));
 NAND2x1_ASAP7_75t_R _13335_ (.A(_09453_),
    .B(_09436_),
    .Y(_09454_));
 AND2x2_ASAP7_75t_R _13336_ (.A(_00177_),
    .B(_09440_),
    .Y(_09455_));
 AO221x1_ASAP7_75t_R _13337_ (.A1(_00073_),
    .A2(_09439_),
    .B1(_09455_),
    .B2(_09442_),
    .C(_09443_),
    .Y(_09456_));
 AOI21x1_ASAP7_75t_R _13338_ (.A1(_09454_),
    .A2(_09456_),
    .B(_09275_),
    .Y(_02865_));
 INVx1_ASAP7_75t_R _13339_ (.A(_01917_),
    .Y(_09457_));
 NAND2x1_ASAP7_75t_R _13340_ (.A(_09457_),
    .B(_09436_),
    .Y(_09458_));
 AND2x2_ASAP7_75t_R _13341_ (.A(_00176_),
    .B(_09440_),
    .Y(_09459_));
 AO221x1_ASAP7_75t_R _13342_ (.A1(_00072_),
    .A2(_09439_),
    .B1(_09459_),
    .B2(_09442_),
    .C(_09443_),
    .Y(_09460_));
 AOI21x1_ASAP7_75t_R _13343_ (.A1(_09458_),
    .A2(_09460_),
    .B(_09275_),
    .Y(_02866_));
 AND3x1_ASAP7_75t_R _13344_ (.A(_00175_),
    .B(_09440_),
    .C(_09376_),
    .Y(_09461_));
 AOI21x1_ASAP7_75t_R _13345_ (.A1(_00071_),
    .A2(_09439_),
    .B(_09461_),
    .Y(_09462_));
 OA21x2_ASAP7_75t_R _13346_ (.A1(_09436_),
    .A2(_09462_),
    .B(_09300_),
    .Y(_02867_));
 NAND2x1_ASAP7_75t_R _13347_ (.A(_09419_),
    .B(_09436_),
    .Y(_09463_));
 AND2x2_ASAP7_75t_R _13348_ (.A(_00174_),
    .B(_09440_),
    .Y(_09464_));
 AO221x1_ASAP7_75t_R _13349_ (.A1(_00070_),
    .A2(_09439_),
    .B1(_09464_),
    .B2(_09442_),
    .C(_09443_),
    .Y(_09465_));
 AOI21x1_ASAP7_75t_R _13350_ (.A1(_09463_),
    .A2(_09465_),
    .B(_09275_),
    .Y(_02868_));
 NAND2x1_ASAP7_75t_R _13351_ (.A(_09422_),
    .B(_09436_),
    .Y(_09466_));
 AND2x2_ASAP7_75t_R _13352_ (.A(_00173_),
    .B(_09440_),
    .Y(_09467_));
 AO221x1_ASAP7_75t_R _13353_ (.A1(_00069_),
    .A2(_09439_),
    .B1(_09467_),
    .B2(_09442_),
    .C(_09443_),
    .Y(_09468_));
 AOI21x1_ASAP7_75t_R _13354_ (.A1(_09466_),
    .A2(_09468_),
    .B(_09275_),
    .Y(_02869_));
 INVx1_ASAP7_75t_R _13355_ (.A(_01913_),
    .Y(_09469_));
 NAND2x1_ASAP7_75t_R _13356_ (.A(_09469_),
    .B(_09436_),
    .Y(_09470_));
 AND2x2_ASAP7_75t_R _13357_ (.A(_00172_),
    .B(_09440_),
    .Y(_09471_));
 AO221x1_ASAP7_75t_R _13358_ (.A1(_00068_),
    .A2(_09439_),
    .B1(_09471_),
    .B2(_09442_),
    .C(_09443_),
    .Y(_09472_));
 AOI21x1_ASAP7_75t_R _13359_ (.A1(_09470_),
    .A2(_09472_),
    .B(_09275_),
    .Y(_02870_));
 NAND2x1_ASAP7_75t_R _13360_ (.A(_09424_),
    .B(_09436_),
    .Y(_09473_));
 AND2x2_ASAP7_75t_R _13361_ (.A(_00171_),
    .B(_09385_),
    .Y(_09474_));
 AO221x1_ASAP7_75t_R _13362_ (.A1(_00067_),
    .A2(_09439_),
    .B1(_09474_),
    .B2(_09442_),
    .C(_09435_),
    .Y(_09475_));
 BUFx12f_ASAP7_75t_R _13363_ (.A(_09118_),
    .Y(_09476_));
 AOI21x1_ASAP7_75t_R _13364_ (.A1(_09473_),
    .A2(_09475_),
    .B(_09476_),
    .Y(_02871_));
 OR3x1_ASAP7_75t_R _13365_ (.A(_08657_),
    .B(_09352_),
    .C(_09442_),
    .Y(_09477_));
 INVx1_ASAP7_75t_R _13366_ (.A(_09477_),
    .Y(_02872_));
 NAND3x1_ASAP7_75t_R _13367_ (.A(_09379_),
    .B(_09403_),
    .C(_09432_),
    .Y(_09478_));
 AND4x1_ASAP7_75t_R _13368_ (.A(_09440_),
    .B(_09376_),
    .C(_09478_),
    .D(_09434_),
    .Y(_09479_));
 NOR2x1_ASAP7_75t_R _13369_ (.A(_08942_),
    .B(_09479_),
    .Y(_02873_));
 INVx1_ASAP7_75t_R _13370_ (.A(_01909_),
    .Y(_09480_));
 NAND2x1_ASAP7_75t_R _13371_ (.A(_09480_),
    .B(_09443_),
    .Y(_09481_));
 AND2x2_ASAP7_75t_R _13372_ (.A(_00168_),
    .B(_09385_),
    .Y(_09482_));
 AO221x1_ASAP7_75t_R _13373_ (.A1(_00064_),
    .A2(_09438_),
    .B1(_09482_),
    .B2(_09376_),
    .C(_09435_),
    .Y(_09483_));
 AOI21x1_ASAP7_75t_R _13374_ (.A1(_09481_),
    .A2(_09483_),
    .B(_09476_),
    .Y(_02874_));
 INVx1_ASAP7_75t_R _13375_ (.A(_01908_),
    .Y(_09484_));
 NAND2x1_ASAP7_75t_R _13376_ (.A(_09484_),
    .B(_09443_),
    .Y(_09485_));
 AND2x2_ASAP7_75t_R _13377_ (.A(_00167_),
    .B(_09385_),
    .Y(_09486_));
 AO221x1_ASAP7_75t_R _13378_ (.A1(_00063_),
    .A2(_09438_),
    .B1(_09486_),
    .B2(_09376_),
    .C(_09435_),
    .Y(_09487_));
 AOI21x1_ASAP7_75t_R _13379_ (.A1(_09485_),
    .A2(_09487_),
    .B(_09476_),
    .Y(_02875_));
 OA21x2_ASAP7_75t_R _13380_ (.A1(_09382_),
    .A2(_09384_),
    .B(_01916_),
    .Y(_09488_));
 OA31x2_ASAP7_75t_R _13381_ (.A1(_09357_),
    .A2(_09396_),
    .A3(_09401_),
    .B1(_01911_),
    .Y(_09489_));
 OA211x2_ASAP7_75t_R _13382_ (.A1(_09488_),
    .A2(_09432_),
    .B(_09489_),
    .C(_09400_),
    .Y(_09490_));
 NOR2x1_ASAP7_75t_R _13383_ (.A(_09365_),
    .B(_09490_),
    .Y(_09491_));
 AND2x2_ASAP7_75t_R _13384_ (.A(_08526_),
    .B(_09491_),
    .Y(_09492_));
 BUFx3_ASAP7_75t_R _13385_ (.A(_09492_),
    .Y(_09493_));
 OR3x1_ASAP7_75t_R _13386_ (.A(_09353_),
    .B(_00172_),
    .C(_09354_),
    .Y(_09494_));
 NAND2x1_ASAP7_75t_R _13387_ (.A(_09355_),
    .B(_09494_),
    .Y(_09495_));
 NAND2x1_ASAP7_75t_R _13388_ (.A(_09371_),
    .B(_09357_),
    .Y(_09496_));
 OA31x2_ASAP7_75t_R _13389_ (.A1(_09495_),
    .A2(_09381_),
    .A3(_09389_),
    .B1(_09496_),
    .Y(_09497_));
 AND3x1_ASAP7_75t_R _13390_ (.A(_09365_),
    .B(_00004_),
    .C(_09369_),
    .Y(_09498_));
 OA211x2_ASAP7_75t_R _13391_ (.A1(_09367_),
    .A2(_09498_),
    .B(_09357_),
    .C(_09385_),
    .Y(_09499_));
 NAND2x1_ASAP7_75t_R _13392_ (.A(_09368_),
    .B(_09396_),
    .Y(_09500_));
 AOI211x1_ASAP7_75t_R _13393_ (.A1(_09385_),
    .A2(_09375_),
    .B(_09499_),
    .C(_09500_),
    .Y(_09501_));
 NAND2x1_ASAP7_75t_R _13394_ (.A(_09497_),
    .B(_09501_),
    .Y(_09502_));
 BUFx6f_ASAP7_75t_R _13395_ (.A(_09502_),
    .Y(_09503_));
 INVx1_ASAP7_75t_R _13396_ (.A(_00180_),
    .Y(_09504_));
 OA21x2_ASAP7_75t_R _13397_ (.A1(_09365_),
    .A2(_09490_),
    .B(_08526_),
    .Y(_09505_));
 BUFx6f_ASAP7_75t_R _13398_ (.A(_09505_),
    .Y(_09506_));
 AND2x2_ASAP7_75t_R _13399_ (.A(_09504_),
    .B(_09506_),
    .Y(_09507_));
 INVx1_ASAP7_75t_R _13400_ (.A(_00076_),
    .Y(_09508_));
 BUFx6f_ASAP7_75t_R _13401_ (.A(_09505_),
    .Y(_09509_));
 BUFx6f_ASAP7_75t_R _13402_ (.A(_09497_),
    .Y(_09510_));
 BUFx6f_ASAP7_75t_R _13403_ (.A(_09501_),
    .Y(_09511_));
 AND4x1_ASAP7_75t_R _13404_ (.A(_09508_),
    .B(_09509_),
    .C(_09510_),
    .D(_09511_),
    .Y(_09512_));
 AO221x1_ASAP7_75t_R _13405_ (.A1(_09430_),
    .A2(_09493_),
    .B1(_09503_),
    .B2(_09507_),
    .C(_09512_),
    .Y(_02876_));
 INVx1_ASAP7_75t_R _13406_ (.A(_00179_),
    .Y(_09513_));
 AND2x2_ASAP7_75t_R _13407_ (.A(_09513_),
    .B(_09506_),
    .Y(_09514_));
 INVx1_ASAP7_75t_R _13408_ (.A(_00075_),
    .Y(_09515_));
 AND4x1_ASAP7_75t_R _13409_ (.A(_09515_),
    .B(_09509_),
    .C(_09510_),
    .D(_09511_),
    .Y(_09516_));
 AO221x1_ASAP7_75t_R _13410_ (.A1(_09445_),
    .A2(_09493_),
    .B1(_09503_),
    .B2(_09514_),
    .C(_09516_),
    .Y(_02877_));
 INVx1_ASAP7_75t_R _13411_ (.A(_00178_),
    .Y(_09517_));
 AND2x2_ASAP7_75t_R _13412_ (.A(_09517_),
    .B(_09506_),
    .Y(_09518_));
 INVx1_ASAP7_75t_R _13413_ (.A(_00074_),
    .Y(_09519_));
 AND4x1_ASAP7_75t_R _13414_ (.A(_09519_),
    .B(_09509_),
    .C(_09510_),
    .D(_09511_),
    .Y(_09520_));
 AO221x1_ASAP7_75t_R _13415_ (.A1(_09449_),
    .A2(_09493_),
    .B1(_09503_),
    .B2(_09518_),
    .C(_09520_),
    .Y(_02878_));
 INVx1_ASAP7_75t_R _13416_ (.A(_00177_),
    .Y(_09521_));
 AND2x2_ASAP7_75t_R _13417_ (.A(_09521_),
    .B(_09506_),
    .Y(_09522_));
 INVx1_ASAP7_75t_R _13418_ (.A(_00073_),
    .Y(_09523_));
 AND4x1_ASAP7_75t_R _13419_ (.A(_09523_),
    .B(_09509_),
    .C(_09510_),
    .D(_09511_),
    .Y(_09524_));
 AO221x1_ASAP7_75t_R _13420_ (.A1(_09453_),
    .A2(_09493_),
    .B1(_09503_),
    .B2(_09522_),
    .C(_09524_),
    .Y(_02879_));
 INVx1_ASAP7_75t_R _13421_ (.A(_00176_),
    .Y(_09525_));
 AND2x2_ASAP7_75t_R _13422_ (.A(_09525_),
    .B(_09506_),
    .Y(_09526_));
 INVx1_ASAP7_75t_R _13423_ (.A(_00072_),
    .Y(_09527_));
 AND4x1_ASAP7_75t_R _13424_ (.A(_09527_),
    .B(_09509_),
    .C(_09510_),
    .D(_09511_),
    .Y(_09528_));
 AO221x1_ASAP7_75t_R _13425_ (.A1(_09457_),
    .A2(_09493_),
    .B1(_09503_),
    .B2(_09526_),
    .C(_09528_),
    .Y(_02880_));
 OR2x6_ASAP7_75t_R _13426_ (.A(_09365_),
    .B(_09490_),
    .Y(_09529_));
 AND2x2_ASAP7_75t_R _13427_ (.A(_09417_),
    .B(_09529_),
    .Y(_09530_));
 NOR2x1_ASAP7_75t_R _13428_ (.A(_09207_),
    .B(_01916_),
    .Y(_09531_));
 AND5x1_ASAP7_75t_R _13429_ (.A(_08876_),
    .B(_09395_),
    .C(_09529_),
    .D(_09497_),
    .E(_09501_),
    .Y(_09532_));
 AO221x1_ASAP7_75t_R _13430_ (.A1(_09502_),
    .A2(_09530_),
    .B1(_09531_),
    .B2(_09491_),
    .C(_09532_),
    .Y(_02881_));
 AND2x2_ASAP7_75t_R _13431_ (.A(_09418_),
    .B(_09506_),
    .Y(_09533_));
 INVx1_ASAP7_75t_R _13432_ (.A(_00070_),
    .Y(_09534_));
 AND4x1_ASAP7_75t_R _13433_ (.A(_09534_),
    .B(_09509_),
    .C(_09510_),
    .D(_09511_),
    .Y(_09535_));
 AO221x1_ASAP7_75t_R _13434_ (.A1(_09419_),
    .A2(_09493_),
    .B1(_09503_),
    .B2(_09533_),
    .C(_09535_),
    .Y(_02882_));
 AND2x2_ASAP7_75t_R _13435_ (.A(_09421_),
    .B(_09506_),
    .Y(_09536_));
 INVx1_ASAP7_75t_R _13436_ (.A(_00069_),
    .Y(_09537_));
 AND4x1_ASAP7_75t_R _13437_ (.A(_09537_),
    .B(_09509_),
    .C(_09510_),
    .D(_09511_),
    .Y(_09538_));
 AO221x1_ASAP7_75t_R _13438_ (.A1(_09422_),
    .A2(_09493_),
    .B1(_09503_),
    .B2(_09536_),
    .C(_09538_),
    .Y(_02883_));
 INVx1_ASAP7_75t_R _13439_ (.A(_00172_),
    .Y(_09539_));
 AND2x2_ASAP7_75t_R _13440_ (.A(_09539_),
    .B(_09506_),
    .Y(_09540_));
 AND4x1_ASAP7_75t_R _13441_ (.A(_09358_),
    .B(_09509_),
    .C(_09510_),
    .D(_09511_),
    .Y(_09541_));
 AO221x1_ASAP7_75t_R _13442_ (.A1(_09469_),
    .A2(_09493_),
    .B1(_09503_),
    .B2(_09540_),
    .C(_09541_),
    .Y(_02884_));
 AND2x2_ASAP7_75t_R _13443_ (.A(_09353_),
    .B(_09506_),
    .Y(_09542_));
 AND4x1_ASAP7_75t_R _13444_ (.A(_09362_),
    .B(_09509_),
    .C(_09510_),
    .D(_09511_),
    .Y(_09543_));
 AO221x1_ASAP7_75t_R _13445_ (.A1(_09424_),
    .A2(_09493_),
    .B1(_09503_),
    .B2(_09542_),
    .C(_09543_),
    .Y(_02885_));
 OA211x2_ASAP7_75t_R _13446_ (.A1(_09488_),
    .A2(_09432_),
    .B(_09402_),
    .C(_09400_),
    .Y(_09544_));
 OR3x1_ASAP7_75t_R _13447_ (.A(_09207_),
    .B(_09365_),
    .C(_09359_),
    .Y(_09545_));
 NOR2x1_ASAP7_75t_R _13448_ (.A(_09544_),
    .B(_09545_),
    .Y(_02886_));
 NAND2x1_ASAP7_75t_R _13449_ (.A(_09529_),
    .B(_09510_),
    .Y(_09546_));
 OA21x2_ASAP7_75t_R _13450_ (.A1(_09511_),
    .A2(_09546_),
    .B(_09300_),
    .Y(_02887_));
 INVx1_ASAP7_75t_R _13451_ (.A(_00168_),
    .Y(_09547_));
 AND2x2_ASAP7_75t_R _13452_ (.A(_09547_),
    .B(_09506_),
    .Y(_09548_));
 INVx1_ASAP7_75t_R _13453_ (.A(_00064_),
    .Y(_09549_));
 AND4x1_ASAP7_75t_R _13454_ (.A(_09549_),
    .B(_09505_),
    .C(_09497_),
    .D(_09501_),
    .Y(_09550_));
 AO221x1_ASAP7_75t_R _13455_ (.A1(_09480_),
    .A2(_09493_),
    .B1(_09503_),
    .B2(_09548_),
    .C(_09550_),
    .Y(_02888_));
 INVx1_ASAP7_75t_R _13456_ (.A(_00167_),
    .Y(_09551_));
 AND2x2_ASAP7_75t_R _13457_ (.A(_09551_),
    .B(_09509_),
    .Y(_09552_));
 INVx1_ASAP7_75t_R _13458_ (.A(_00063_),
    .Y(_09553_));
 AND4x1_ASAP7_75t_R _13459_ (.A(_09553_),
    .B(_09505_),
    .C(_09497_),
    .D(_09501_),
    .Y(_09554_));
 AO221x1_ASAP7_75t_R _13460_ (.A1(_09484_),
    .A2(_09492_),
    .B1(_09502_),
    .B2(_09552_),
    .C(_09554_),
    .Y(_02889_));
 AND2x2_ASAP7_75t_R _13461_ (.A(_08723_),
    .B(_00005_),
    .Y(_02890_));
 AND2x4_ASAP7_75t_R _13462_ (.A(_01523_),
    .B(_01525_),
    .Y(_09555_));
 NOR2x1_ASAP7_75t_R _13463_ (.A(_01524_),
    .B(_01526_),
    .Y(_09556_));
 BUFx6f_ASAP7_75t_R _13464_ (.A(_01521_),
    .Y(_09557_));
 AO21x2_ASAP7_75t_R _13465_ (.A1(_09555_),
    .A2(_09556_),
    .B(_09557_),
    .Y(_09558_));
 INVx1_ASAP7_75t_R _13466_ (.A(_01419_),
    .Y(_09559_));
 INVx1_ASAP7_75t_R _13467_ (.A(_01421_),
    .Y(_09560_));
 OR4x1_ASAP7_75t_R _13468_ (.A(_09559_),
    .B(_01420_),
    .C(_09560_),
    .D(_01422_),
    .Y(_09561_));
 BUFx6f_ASAP7_75t_R _13469_ (.A(_09561_),
    .Y(_09562_));
 INVx3_ASAP7_75t_R _13470_ (.A(_01902_),
    .Y(_09563_));
 INVx3_ASAP7_75t_R _13471_ (.A(_01417_),
    .Y(_09564_));
 OA21x2_ASAP7_75t_R _13472_ (.A1(_01896_),
    .A2(_09563_),
    .B(_09564_),
    .Y(_09565_));
 BUFx6f_ASAP7_75t_R _13473_ (.A(_01896_),
    .Y(_09566_));
 NOR2x1_ASAP7_75t_R _13474_ (.A(_01417_),
    .B(_01418_),
    .Y(_09567_));
 OA21x2_ASAP7_75t_R _13475_ (.A1(_09566_),
    .A2(_09563_),
    .B(_09567_),
    .Y(_09568_));
 BUFx6f_ASAP7_75t_R _13476_ (.A(_01897_),
    .Y(_09569_));
 INVx2_ASAP7_75t_R _13477_ (.A(_09569_),
    .Y(_09570_));
 AOI211x1_ASAP7_75t_R _13478_ (.A1(_09562_),
    .A2(_09565_),
    .B(_09568_),
    .C(_09570_),
    .Y(_09571_));
 INVx1_ASAP7_75t_R _13479_ (.A(_01420_),
    .Y(_09572_));
 INVx1_ASAP7_75t_R _13480_ (.A(_01422_),
    .Y(_09573_));
 AND4x1_ASAP7_75t_R _13481_ (.A(_01419_),
    .B(_09572_),
    .C(_01421_),
    .D(_09573_),
    .Y(_09574_));
 OR2x2_ASAP7_75t_R _13482_ (.A(_01417_),
    .B(_00005_),
    .Y(_09575_));
 OA21x2_ASAP7_75t_R _13483_ (.A1(_09574_),
    .A2(_09575_),
    .B(_09566_),
    .Y(_09576_));
 OR2x6_ASAP7_75t_R _13484_ (.A(_09557_),
    .B(_01527_),
    .Y(_09577_));
 AO21x1_ASAP7_75t_R _13485_ (.A1(_09569_),
    .A2(_01902_),
    .B(_09566_),
    .Y(_09578_));
 OR2x2_ASAP7_75t_R _13486_ (.A(_01417_),
    .B(_01418_),
    .Y(_09579_));
 BUFx6f_ASAP7_75t_R _13487_ (.A(_09579_),
    .Y(_09580_));
 OA31x2_ASAP7_75t_R _13488_ (.A1(_01417_),
    .A2(_09574_),
    .A3(_09578_),
    .B1(_09580_),
    .Y(_09581_));
 NAND2x1_ASAP7_75t_R _13489_ (.A(_09555_),
    .B(_09556_),
    .Y(_09582_));
 OA33x2_ASAP7_75t_R _13490_ (.A1(_09558_),
    .A2(_09571_),
    .A3(_09576_),
    .B1(_09577_),
    .B2(_09581_),
    .B3(_09582_),
    .Y(_09583_));
 AO21x1_ASAP7_75t_R _13491_ (.A1(_09569_),
    .A2(_09563_),
    .B(_09566_),
    .Y(_09584_));
 OR2x2_ASAP7_75t_R _13492_ (.A(_09557_),
    .B(_01522_),
    .Y(_09585_));
 BUFx6f_ASAP7_75t_R _13493_ (.A(_09585_),
    .Y(_09586_));
 OAI21x1_ASAP7_75t_R _13494_ (.A1(_09558_),
    .A2(_09584_),
    .B(_09586_),
    .Y(_09587_));
 NAND2x1_ASAP7_75t_R _13495_ (.A(_09564_),
    .B(_01423_),
    .Y(_09588_));
 OR2x6_ASAP7_75t_R _13496_ (.A(_09562_),
    .B(_09588_),
    .Y(_09589_));
 NOR2x1_ASAP7_75t_R _13497_ (.A(_09557_),
    .B(_01522_),
    .Y(_09590_));
 AOI211x1_ASAP7_75t_R _13498_ (.A1(_09580_),
    .A2(_09587_),
    .B(_09589_),
    .C(_09590_),
    .Y(_09591_));
 AND2x4_ASAP7_75t_R _13499_ (.A(_09583_),
    .B(_09591_),
    .Y(_09592_));
 BUFx6f_ASAP7_75t_R _13500_ (.A(_09592_),
    .Y(_09593_));
 NAND2x1_ASAP7_75t_R _13501_ (.A(_01428_),
    .B(_09593_),
    .Y(_09594_));
 NAND2x2_ASAP7_75t_R _13502_ (.A(_09583_),
    .B(_09591_),
    .Y(_09595_));
 NAND2x1_ASAP7_75t_R _13503_ (.A(_01532_),
    .B(_09595_),
    .Y(_09596_));
 AO21x1_ASAP7_75t_R _13504_ (.A1(_09580_),
    .A2(_09587_),
    .B(_09589_),
    .Y(_09597_));
 AOI21x1_ASAP7_75t_R _13505_ (.A1(_09555_),
    .A2(_09556_),
    .B(_09557_),
    .Y(_09598_));
 OA31x2_ASAP7_75t_R _13506_ (.A1(_09598_),
    .A2(_09562_),
    .A3(_09588_),
    .B1(_09586_),
    .Y(_09599_));
 NAND2x1_ASAP7_75t_R _13507_ (.A(_01523_),
    .B(_01525_),
    .Y(_09600_));
 OR2x6_ASAP7_75t_R _13508_ (.A(_01524_),
    .B(_01526_),
    .Y(_09601_));
 OA31x2_ASAP7_75t_R _13509_ (.A1(_09600_),
    .A2(_09601_),
    .A3(_09577_),
    .B1(_01902_),
    .Y(_09602_));
 OA31x2_ASAP7_75t_R _13510_ (.A1(_09600_),
    .A2(_09601_),
    .A3(_09577_),
    .B1(_09586_),
    .Y(_09603_));
 OA33x2_ASAP7_75t_R _13511_ (.A1(_01417_),
    .A2(_01418_),
    .A3(_09602_),
    .B1(_09603_),
    .B2(_09562_),
    .B3(_09588_),
    .Y(_09604_));
 INVx3_ASAP7_75t_R _13512_ (.A(_01896_),
    .Y(_09605_));
 AND2x2_ASAP7_75t_R _13513_ (.A(_09605_),
    .B(_09569_),
    .Y(_09606_));
 AND4x1_ASAP7_75t_R _13514_ (.A(_01902_),
    .B(_09599_),
    .C(_09604_),
    .D(_09606_),
    .Y(_09607_));
 AND4x1_ASAP7_75t_R _13515_ (.A(_09583_),
    .B(_09586_),
    .C(_09597_),
    .D(_09607_),
    .Y(_09608_));
 BUFx6f_ASAP7_75t_R _13516_ (.A(_09608_),
    .Y(_09609_));
 NOR2x2_ASAP7_75t_R _13517_ (.A(_08765_),
    .B(_09609_),
    .Y(_09610_));
 NOR2x1_ASAP7_75t_R _13518_ (.A(_08811_),
    .B(_01907_),
    .Y(_09611_));
 BUFx6f_ASAP7_75t_R _13519_ (.A(_09609_),
    .Y(_09612_));
 AO32x1_ASAP7_75t_R _13520_ (.A1(_09594_),
    .A2(_09596_),
    .A3(_09610_),
    .B1(_09611_),
    .B2(_09612_),
    .Y(_02891_));
 NAND2x1_ASAP7_75t_R _13521_ (.A(_01427_),
    .B(_09593_),
    .Y(_09613_));
 NAND2x1_ASAP7_75t_R _13522_ (.A(_01531_),
    .B(_09595_),
    .Y(_09614_));
 NOR2x1_ASAP7_75t_R _13523_ (.A(_08811_),
    .B(_01906_),
    .Y(_09615_));
 AO32x1_ASAP7_75t_R _13524_ (.A1(_09610_),
    .A2(_09613_),
    .A3(_09614_),
    .B1(_09615_),
    .B2(_09612_),
    .Y(_02892_));
 NAND2x1_ASAP7_75t_R _13525_ (.A(_01426_),
    .B(_09593_),
    .Y(_09616_));
 NAND2x1_ASAP7_75t_R _13526_ (.A(_01530_),
    .B(_09595_),
    .Y(_09617_));
 NOR2x1_ASAP7_75t_R _13527_ (.A(_08811_),
    .B(_01905_),
    .Y(_09618_));
 AO32x1_ASAP7_75t_R _13528_ (.A1(_09610_),
    .A2(_09616_),
    .A3(_09617_),
    .B1(_09618_),
    .B2(_09612_),
    .Y(_02893_));
 NAND2x1_ASAP7_75t_R _13529_ (.A(_01425_),
    .B(_09593_),
    .Y(_09619_));
 NAND2x1_ASAP7_75t_R _13530_ (.A(_01529_),
    .B(_09595_),
    .Y(_09620_));
 NOR2x1_ASAP7_75t_R _13531_ (.A(_08811_),
    .B(_01904_),
    .Y(_09621_));
 AO32x1_ASAP7_75t_R _13532_ (.A1(_09610_),
    .A2(_09619_),
    .A3(_09620_),
    .B1(_09621_),
    .B2(_09612_),
    .Y(_02894_));
 NAND2x1_ASAP7_75t_R _13533_ (.A(_01424_),
    .B(_09593_),
    .Y(_09622_));
 NAND2x1_ASAP7_75t_R _13534_ (.A(_01528_),
    .B(_09595_),
    .Y(_09623_));
 NOR2x1_ASAP7_75t_R _13535_ (.A(_08811_),
    .B(_01903_),
    .Y(_09624_));
 AO32x1_ASAP7_75t_R _13536_ (.A1(_09610_),
    .A2(_09622_),
    .A3(_09623_),
    .B1(_09624_),
    .B2(_09612_),
    .Y(_02895_));
 OR4x1_ASAP7_75t_R _13537_ (.A(_08712_),
    .B(_01527_),
    .C(_09593_),
    .D(_09609_),
    .Y(_09625_));
 INVx1_ASAP7_75t_R _13538_ (.A(_09625_),
    .Y(_02896_));
 NAND2x1_ASAP7_75t_R _13539_ (.A(_01901_),
    .B(_09612_),
    .Y(_09626_));
 INVx1_ASAP7_75t_R _13540_ (.A(_01526_),
    .Y(_09627_));
 OR3x1_ASAP7_75t_R _13541_ (.A(_09627_),
    .B(_09592_),
    .C(_09609_),
    .Y(_09628_));
 AND3x1_ASAP7_75t_R _13542_ (.A(_08582_),
    .B(_09626_),
    .C(_09628_),
    .Y(_02897_));
 INVx2_ASAP7_75t_R _13543_ (.A(_01900_),
    .Y(_09629_));
 NAND2x1_ASAP7_75t_R _13544_ (.A(_09629_),
    .B(_09612_),
    .Y(_09630_));
 OR3x1_ASAP7_75t_R _13545_ (.A(_01525_),
    .B(_09593_),
    .C(_09609_),
    .Y(_09631_));
 AOI21x1_ASAP7_75t_R _13546_ (.A1(_09630_),
    .A2(_09631_),
    .B(_09476_),
    .Y(_02898_));
 BUFx12f_ASAP7_75t_R _13547_ (.A(_08581_),
    .Y(_09632_));
 NAND2x1_ASAP7_75t_R _13548_ (.A(_01899_),
    .B(_09609_),
    .Y(_09633_));
 INVx1_ASAP7_75t_R _13549_ (.A(_01524_),
    .Y(_09634_));
 OR3x1_ASAP7_75t_R _13550_ (.A(_09634_),
    .B(_09592_),
    .C(_09609_),
    .Y(_09635_));
 AND3x1_ASAP7_75t_R _13551_ (.A(_09632_),
    .B(_09633_),
    .C(_09635_),
    .Y(_02899_));
 INVx2_ASAP7_75t_R _13552_ (.A(_01898_),
    .Y(_09636_));
 NAND2x1_ASAP7_75t_R _13553_ (.A(_09636_),
    .B(_09612_),
    .Y(_09637_));
 OR3x1_ASAP7_75t_R _13554_ (.A(_01523_),
    .B(_09593_),
    .C(_09609_),
    .Y(_09638_));
 AOI21x1_ASAP7_75t_R _13555_ (.A1(_09637_),
    .A2(_09638_),
    .B(_09476_),
    .Y(_02900_));
 OR3x1_ASAP7_75t_R _13556_ (.A(_08657_),
    .B(_09583_),
    .C(_09590_),
    .Y(_09639_));
 INVx1_ASAP7_75t_R _13557_ (.A(_09639_),
    .Y(_02901_));
 NAND3x1_ASAP7_75t_R _13558_ (.A(_09583_),
    .B(_09586_),
    .C(_09597_),
    .Y(_09640_));
 OA21x2_ASAP7_75t_R _13559_ (.A1(_09640_),
    .A2(_09607_),
    .B(_09300_),
    .Y(_02902_));
 NAND2x1_ASAP7_75t_R _13560_ (.A(_01416_),
    .B(_09593_),
    .Y(_09641_));
 NAND2x1_ASAP7_75t_R _13561_ (.A(_01520_),
    .B(_09595_),
    .Y(_09642_));
 NOR2x1_ASAP7_75t_R _13562_ (.A(_08811_),
    .B(_01895_),
    .Y(_09643_));
 AO32x1_ASAP7_75t_R _13563_ (.A1(_09610_),
    .A2(_09641_),
    .A3(_09642_),
    .B1(_09643_),
    .B2(_09612_),
    .Y(_02903_));
 NAND2x1_ASAP7_75t_R _13564_ (.A(_01415_),
    .B(_09593_),
    .Y(_09644_));
 NAND2x1_ASAP7_75t_R _13565_ (.A(_01519_),
    .B(_09595_),
    .Y(_09645_));
 NOR2x1_ASAP7_75t_R _13566_ (.A(_08811_),
    .B(_01894_),
    .Y(_09646_));
 AO32x1_ASAP7_75t_R _13567_ (.A1(_09610_),
    .A2(_09644_),
    .A3(_09645_),
    .B1(_09646_),
    .B2(_09612_),
    .Y(_02904_));
 OR3x2_ASAP7_75t_R _13568_ (.A(_09600_),
    .B(_09601_),
    .C(_09577_),
    .Y(_09647_));
 AO211x2_ASAP7_75t_R _13569_ (.A1(_09562_),
    .A2(_09565_),
    .B(_09568_),
    .C(_09570_),
    .Y(_09648_));
 OAI21x1_ASAP7_75t_R _13570_ (.A1(_09574_),
    .A2(_09575_),
    .B(_09566_),
    .Y(_09649_));
 AND2x2_ASAP7_75t_R _13571_ (.A(_09598_),
    .B(_09586_),
    .Y(_09650_));
 OA21x2_ASAP7_75t_R _13572_ (.A1(_09570_),
    .A2(_09563_),
    .B(_09605_),
    .Y(_09651_));
 AO31x2_ASAP7_75t_R _13573_ (.A1(_09564_),
    .A2(_09562_),
    .A3(_09651_),
    .B(_09567_),
    .Y(_09652_));
 AO32x2_ASAP7_75t_R _13574_ (.A1(_09648_),
    .A2(_09649_),
    .A3(_09650_),
    .B1(_09586_),
    .B2(_09652_),
    .Y(_09653_));
 AO211x2_ASAP7_75t_R _13575_ (.A1(_09564_),
    .A2(_09562_),
    .B(_09647_),
    .C(_01902_),
    .Y(_09654_));
 AND4x1_ASAP7_75t_R _13576_ (.A(_09563_),
    .B(_09654_),
    .C(_09604_),
    .D(_09606_),
    .Y(_09655_));
 OAI21x1_ASAP7_75t_R _13577_ (.A1(_09647_),
    .A2(_09653_),
    .B(_09655_),
    .Y(_09656_));
 OR2x2_ASAP7_75t_R _13578_ (.A(_01907_),
    .B(_09656_),
    .Y(_09657_));
 OA21x2_ASAP7_75t_R _13579_ (.A1(_09558_),
    .A2(_09584_),
    .B(_09586_),
    .Y(_09658_));
 OA21x2_ASAP7_75t_R _13580_ (.A1(_09563_),
    .A2(_09586_),
    .B(_09569_),
    .Y(_09659_));
 OA21x2_ASAP7_75t_R _13581_ (.A1(_09566_),
    .A2(_09659_),
    .B(_09558_),
    .Y(_09660_));
 AND3x1_ASAP7_75t_R _13582_ (.A(_09605_),
    .B(_09569_),
    .C(_09563_),
    .Y(_09661_));
 NOR2x1_ASAP7_75t_R _13583_ (.A(_09605_),
    .B(_00005_),
    .Y(_09662_));
 OR4x1_ASAP7_75t_R _13584_ (.A(_01417_),
    .B(_09574_),
    .C(_09661_),
    .D(_09662_),
    .Y(_09663_));
 OA22x2_ASAP7_75t_R _13585_ (.A1(_09589_),
    .A2(_09658_),
    .B1(_09660_),
    .B2(_09663_),
    .Y(_09664_));
 NAND2x1_ASAP7_75t_R _13586_ (.A(_09580_),
    .B(_09664_),
    .Y(_09665_));
 BUFx3_ASAP7_75t_R _13587_ (.A(_09665_),
    .Y(_09666_));
 BUFx6f_ASAP7_75t_R _13588_ (.A(_09580_),
    .Y(_09667_));
 AND2x2_ASAP7_75t_R _13589_ (.A(_01532_),
    .B(_09667_),
    .Y(_09668_));
 BUFx6f_ASAP7_75t_R _13590_ (.A(_09664_),
    .Y(_09669_));
 OA21x2_ASAP7_75t_R _13591_ (.A1(_09647_),
    .A2(_09653_),
    .B(_09655_),
    .Y(_09670_));
 BUFx6f_ASAP7_75t_R _13592_ (.A(_09670_),
    .Y(_09671_));
 AO221x1_ASAP7_75t_R _13593_ (.A1(_01428_),
    .A2(_09666_),
    .B1(_09668_),
    .B2(_09669_),
    .C(_09671_),
    .Y(_09672_));
 AOI21x1_ASAP7_75t_R _13594_ (.A1(_09657_),
    .A2(_09672_),
    .B(_09476_),
    .Y(_02905_));
 OR2x2_ASAP7_75t_R _13595_ (.A(_01906_),
    .B(_09656_),
    .Y(_09673_));
 AND2x2_ASAP7_75t_R _13596_ (.A(_01531_),
    .B(_09667_),
    .Y(_09674_));
 AO221x1_ASAP7_75t_R _13597_ (.A1(_01427_),
    .A2(_09666_),
    .B1(_09674_),
    .B2(_09669_),
    .C(_09671_),
    .Y(_09675_));
 AOI21x1_ASAP7_75t_R _13598_ (.A1(_09673_),
    .A2(_09675_),
    .B(_09476_),
    .Y(_02906_));
 OR2x2_ASAP7_75t_R _13599_ (.A(_01905_),
    .B(_09656_),
    .Y(_09676_));
 AND2x2_ASAP7_75t_R _13600_ (.A(_01530_),
    .B(_09667_),
    .Y(_09677_));
 AO221x1_ASAP7_75t_R _13601_ (.A1(_01426_),
    .A2(_09666_),
    .B1(_09677_),
    .B2(_09669_),
    .C(_09671_),
    .Y(_09678_));
 AOI21x1_ASAP7_75t_R _13602_ (.A1(_09676_),
    .A2(_09678_),
    .B(_09476_),
    .Y(_02907_));
 OR2x2_ASAP7_75t_R _13603_ (.A(_01904_),
    .B(_09656_),
    .Y(_09679_));
 AND2x2_ASAP7_75t_R _13604_ (.A(_01529_),
    .B(_09667_),
    .Y(_09680_));
 AO221x1_ASAP7_75t_R _13605_ (.A1(_01425_),
    .A2(_09666_),
    .B1(_09680_),
    .B2(_09669_),
    .C(_09671_),
    .Y(_09681_));
 AOI21x1_ASAP7_75t_R _13606_ (.A1(_09679_),
    .A2(_09681_),
    .B(_09476_),
    .Y(_02908_));
 OR2x2_ASAP7_75t_R _13607_ (.A(_01903_),
    .B(_09656_),
    .Y(_09682_));
 AND2x2_ASAP7_75t_R _13608_ (.A(_01528_),
    .B(_09667_),
    .Y(_09683_));
 AO221x1_ASAP7_75t_R _13609_ (.A1(_01424_),
    .A2(_09666_),
    .B1(_09683_),
    .B2(_09669_),
    .C(_09671_),
    .Y(_09684_));
 AOI21x1_ASAP7_75t_R _13610_ (.A1(_09682_),
    .A2(_09684_),
    .B(_09476_),
    .Y(_02909_));
 AND3x1_ASAP7_75t_R _13611_ (.A(_01527_),
    .B(_09667_),
    .C(_09664_),
    .Y(_09685_));
 AO21x1_ASAP7_75t_R _13612_ (.A1(_01423_),
    .A2(_09666_),
    .B(_09685_),
    .Y(_09686_));
 BUFx12f_ASAP7_75t_R _13613_ (.A(_09118_),
    .Y(_09687_));
 AOI21x1_ASAP7_75t_R _13614_ (.A1(_09656_),
    .A2(_09686_),
    .B(_09687_),
    .Y(_02910_));
 OR2x2_ASAP7_75t_R _13615_ (.A(_01901_),
    .B(_09656_),
    .Y(_09688_));
 AND2x2_ASAP7_75t_R _13616_ (.A(_01526_),
    .B(_09667_),
    .Y(_09689_));
 AO221x1_ASAP7_75t_R _13617_ (.A1(_01422_),
    .A2(_09666_),
    .B1(_09689_),
    .B2(_09669_),
    .C(_09671_),
    .Y(_09690_));
 AOI21x1_ASAP7_75t_R _13618_ (.A1(_09688_),
    .A2(_09690_),
    .B(_09687_),
    .Y(_02911_));
 NAND2x1_ASAP7_75t_R _13619_ (.A(_09629_),
    .B(_09671_),
    .Y(_09691_));
 AND2x2_ASAP7_75t_R _13620_ (.A(_01525_),
    .B(_09667_),
    .Y(_09692_));
 AO221x1_ASAP7_75t_R _13621_ (.A1(_01421_),
    .A2(_09666_),
    .B1(_09692_),
    .B2(_09669_),
    .C(_09671_),
    .Y(_09693_));
 AOI21x1_ASAP7_75t_R _13622_ (.A1(_09691_),
    .A2(_09693_),
    .B(_09687_),
    .Y(_02912_));
 OR2x2_ASAP7_75t_R _13623_ (.A(_01899_),
    .B(_09656_),
    .Y(_09694_));
 AND2x2_ASAP7_75t_R _13624_ (.A(_01524_),
    .B(_09667_),
    .Y(_09695_));
 AO221x1_ASAP7_75t_R _13625_ (.A1(_01420_),
    .A2(_09666_),
    .B1(_09695_),
    .B2(_09669_),
    .C(_09671_),
    .Y(_09696_));
 AOI21x1_ASAP7_75t_R _13626_ (.A1(_09694_),
    .A2(_09696_),
    .B(_09687_),
    .Y(_02913_));
 NAND2x1_ASAP7_75t_R _13627_ (.A(_09636_),
    .B(_09671_),
    .Y(_09697_));
 AND2x2_ASAP7_75t_R _13628_ (.A(_01523_),
    .B(_09667_),
    .Y(_09698_));
 AO221x1_ASAP7_75t_R _13629_ (.A1(_01419_),
    .A2(_09666_),
    .B1(_09698_),
    .B2(_09669_),
    .C(_09670_),
    .Y(_09699_));
 AOI21x1_ASAP7_75t_R _13630_ (.A1(_09697_),
    .A2(_09699_),
    .B(_09687_),
    .Y(_02914_));
 OR3x1_ASAP7_75t_R _13631_ (.A(_08657_),
    .B(_09567_),
    .C(_09669_),
    .Y(_09700_));
 INVx1_ASAP7_75t_R _13632_ (.A(_09700_),
    .Y(_02915_));
 NOR2x1_ASAP7_75t_R _13633_ (.A(_09647_),
    .B(_09653_),
    .Y(_09701_));
 OR3x1_ASAP7_75t_R _13634_ (.A(_09701_),
    .B(_09655_),
    .C(_09665_),
    .Y(_09702_));
 AND2x2_ASAP7_75t_R _13635_ (.A(_08723_),
    .B(_09702_),
    .Y(_02916_));
 OR2x2_ASAP7_75t_R _13636_ (.A(_01895_),
    .B(_09656_),
    .Y(_09703_));
 AND2x2_ASAP7_75t_R _13637_ (.A(_01520_),
    .B(_09580_),
    .Y(_09704_));
 AO221x1_ASAP7_75t_R _13638_ (.A1(_01416_),
    .A2(_09665_),
    .B1(_09704_),
    .B2(_09664_),
    .C(_09670_),
    .Y(_09705_));
 AOI21x1_ASAP7_75t_R _13639_ (.A1(_09703_),
    .A2(_09705_),
    .B(_09687_),
    .Y(_02917_));
 OR2x2_ASAP7_75t_R _13640_ (.A(_01894_),
    .B(_09656_),
    .Y(_09706_));
 AND2x2_ASAP7_75t_R _13641_ (.A(_01519_),
    .B(_09580_),
    .Y(_09707_));
 AO221x1_ASAP7_75t_R _13642_ (.A1(_01415_),
    .A2(_09665_),
    .B1(_09707_),
    .B2(_09664_),
    .C(_09670_),
    .Y(_09708_));
 AOI21x1_ASAP7_75t_R _13643_ (.A1(_09706_),
    .A2(_09708_),
    .B(_09687_),
    .Y(_02918_));
 OA211x2_ASAP7_75t_R _13644_ (.A1(_09563_),
    .A2(_09599_),
    .B(_09604_),
    .C(_09654_),
    .Y(_09709_));
 AO21x2_ASAP7_75t_R _13645_ (.A1(_09569_),
    .A2(_09709_),
    .B(_09566_),
    .Y(_09710_));
 BUFx6f_ASAP7_75t_R _13646_ (.A(_09710_),
    .Y(_09711_));
 NOR2x1_ASAP7_75t_R _13647_ (.A(_01907_),
    .B(_09711_),
    .Y(_09712_));
 AO21x1_ASAP7_75t_R _13648_ (.A1(_00005_),
    .A2(_09598_),
    .B(_09605_),
    .Y(_09713_));
 OR2x2_ASAP7_75t_R _13649_ (.A(_09566_),
    .B(_01902_),
    .Y(_09714_));
 AOI21x1_ASAP7_75t_R _13650_ (.A1(_09605_),
    .A2(_09563_),
    .B(_09557_),
    .Y(_09715_));
 AO221x1_ASAP7_75t_R _13651_ (.A1(_09590_),
    .A2(_09714_),
    .B1(_09715_),
    .B2(_09582_),
    .C(_09570_),
    .Y(_09716_));
 NAND2x1_ASAP7_75t_R _13652_ (.A(_09564_),
    .B(_09562_),
    .Y(_09717_));
 AO31x2_ASAP7_75t_R _13653_ (.A1(_09580_),
    .A2(_09713_),
    .A3(_09716_),
    .B(_09717_),
    .Y(_09718_));
 OA31x2_ASAP7_75t_R _13654_ (.A1(_09571_),
    .A2(_09576_),
    .A3(_09590_),
    .B1(_09598_),
    .Y(_09719_));
 NOR2x1_ASAP7_75t_R _13655_ (.A(_09718_),
    .B(_09719_),
    .Y(_09720_));
 BUFx6f_ASAP7_75t_R _13656_ (.A(_09720_),
    .Y(_09721_));
 BUFx6f_ASAP7_75t_R _13657_ (.A(_09718_),
    .Y(_09722_));
 BUFx6f_ASAP7_75t_R _13658_ (.A(_09719_),
    .Y(_09723_));
 OA21x2_ASAP7_75t_R _13659_ (.A1(_09722_),
    .A2(_09723_),
    .B(_01532_),
    .Y(_09724_));
 AOI21x1_ASAP7_75t_R _13660_ (.A1(_09569_),
    .A2(_09709_),
    .B(_09566_),
    .Y(_09725_));
 BUFx6f_ASAP7_75t_R _13661_ (.A(_09725_),
    .Y(_09726_));
 AOI211x1_ASAP7_75t_R _13662_ (.A1(_01428_),
    .A2(_09721_),
    .B(_09724_),
    .C(_09726_),
    .Y(_09727_));
 OA21x2_ASAP7_75t_R _13663_ (.A1(_09712_),
    .A2(_09727_),
    .B(_09300_),
    .Y(_02919_));
 NOR2x1_ASAP7_75t_R _13664_ (.A(_01906_),
    .B(_09711_),
    .Y(_09728_));
 OA21x2_ASAP7_75t_R _13665_ (.A1(_09722_),
    .A2(_09723_),
    .B(_01531_),
    .Y(_09729_));
 AOI211x1_ASAP7_75t_R _13666_ (.A1(_01427_),
    .A2(_09721_),
    .B(_09729_),
    .C(_09726_),
    .Y(_09730_));
 OA21x2_ASAP7_75t_R _13667_ (.A1(_09728_),
    .A2(_09730_),
    .B(_09300_),
    .Y(_02920_));
 NOR2x1_ASAP7_75t_R _13668_ (.A(_01905_),
    .B(_09711_),
    .Y(_09731_));
 OA21x2_ASAP7_75t_R _13669_ (.A1(_09722_),
    .A2(_09723_),
    .B(_01530_),
    .Y(_09732_));
 AOI211x1_ASAP7_75t_R _13670_ (.A1(_01426_),
    .A2(_09721_),
    .B(_09732_),
    .C(_09726_),
    .Y(_09733_));
 OA21x2_ASAP7_75t_R _13671_ (.A1(_09731_),
    .A2(_09733_),
    .B(_09300_),
    .Y(_02921_));
 NOR2x1_ASAP7_75t_R _13672_ (.A(_01904_),
    .B(_09711_),
    .Y(_09734_));
 OA21x2_ASAP7_75t_R _13673_ (.A1(_09722_),
    .A2(_09723_),
    .B(_01529_),
    .Y(_09735_));
 AOI211x1_ASAP7_75t_R _13674_ (.A1(_01425_),
    .A2(_09721_),
    .B(_09735_),
    .C(_09726_),
    .Y(_09736_));
 OA21x2_ASAP7_75t_R _13675_ (.A1(_09734_),
    .A2(_09736_),
    .B(_09300_),
    .Y(_02922_));
 NOR2x1_ASAP7_75t_R _13676_ (.A(_01903_),
    .B(_09711_),
    .Y(_09737_));
 OA21x2_ASAP7_75t_R _13677_ (.A1(_09722_),
    .A2(_09723_),
    .B(_01528_),
    .Y(_09738_));
 AOI211x1_ASAP7_75t_R _13678_ (.A1(_01424_),
    .A2(_09721_),
    .B(_09738_),
    .C(_09726_),
    .Y(_09739_));
 OA21x2_ASAP7_75t_R _13679_ (.A1(_09737_),
    .A2(_09739_),
    .B(_09300_),
    .Y(_02923_));
 AND2x2_ASAP7_75t_R _13680_ (.A(_09563_),
    .B(_09726_),
    .Y(_09740_));
 OA21x2_ASAP7_75t_R _13681_ (.A1(_09722_),
    .A2(_09723_),
    .B(_01527_),
    .Y(_09741_));
 AOI211x1_ASAP7_75t_R _13682_ (.A1(_01423_),
    .A2(_09721_),
    .B(_09741_),
    .C(_09726_),
    .Y(_09742_));
 BUFx6f_ASAP7_75t_R _13683_ (.A(_08665_),
    .Y(_09743_));
 OA21x2_ASAP7_75t_R _13684_ (.A1(_09740_),
    .A2(_09742_),
    .B(_09743_),
    .Y(_02924_));
 NOR2x1_ASAP7_75t_R _13685_ (.A(_01901_),
    .B(_09711_),
    .Y(_09744_));
 OR3x1_ASAP7_75t_R _13686_ (.A(_09573_),
    .B(_09722_),
    .C(_09723_),
    .Y(_09745_));
 OA211x2_ASAP7_75t_R _13687_ (.A1(_09627_),
    .A2(_09721_),
    .B(_09745_),
    .C(_09711_),
    .Y(_09746_));
 OA21x2_ASAP7_75t_R _13688_ (.A1(_09744_),
    .A2(_09746_),
    .B(_09743_),
    .Y(_02925_));
 AND2x2_ASAP7_75t_R _13689_ (.A(_09629_),
    .B(_09726_),
    .Y(_09747_));
 INVx1_ASAP7_75t_R _13690_ (.A(_01525_),
    .Y(_09748_));
 OR3x1_ASAP7_75t_R _13691_ (.A(_09560_),
    .B(_09718_),
    .C(_09719_),
    .Y(_09749_));
 OA211x2_ASAP7_75t_R _13692_ (.A1(_09748_),
    .A2(_09721_),
    .B(_09749_),
    .C(_09710_),
    .Y(_09750_));
 OA21x2_ASAP7_75t_R _13693_ (.A1(_09747_),
    .A2(_09750_),
    .B(_09743_),
    .Y(_02926_));
 NOR2x1_ASAP7_75t_R _13694_ (.A(_01899_),
    .B(_09711_),
    .Y(_09751_));
 OR3x1_ASAP7_75t_R _13695_ (.A(_09572_),
    .B(_09718_),
    .C(_09719_),
    .Y(_09752_));
 OA211x2_ASAP7_75t_R _13696_ (.A1(_09634_),
    .A2(_09720_),
    .B(_09752_),
    .C(_09710_),
    .Y(_09753_));
 OA21x2_ASAP7_75t_R _13697_ (.A1(_09751_),
    .A2(_09753_),
    .B(_09743_),
    .Y(_02927_));
 AND2x2_ASAP7_75t_R _13698_ (.A(_09636_),
    .B(_09725_),
    .Y(_09754_));
 INVx1_ASAP7_75t_R _13699_ (.A(_01523_),
    .Y(_09755_));
 OR3x1_ASAP7_75t_R _13700_ (.A(_09559_),
    .B(_09718_),
    .C(_09719_),
    .Y(_09756_));
 OA211x2_ASAP7_75t_R _13701_ (.A1(_09755_),
    .A2(_09720_),
    .B(_09756_),
    .C(_09710_),
    .Y(_09757_));
 OA21x2_ASAP7_75t_R _13702_ (.A1(_09754_),
    .A2(_09757_),
    .B(_09743_),
    .Y(_02928_));
 OR4x1_ASAP7_75t_R _13703_ (.A(_08712_),
    .B(_09566_),
    .C(_09570_),
    .D(_09709_),
    .Y(_09758_));
 INVx1_ASAP7_75t_R _13704_ (.A(_09758_),
    .Y(_02929_));
 INVx1_ASAP7_75t_R _13705_ (.A(_09722_),
    .Y(_09759_));
 OR3x1_ASAP7_75t_R _13706_ (.A(_09725_),
    .B(_09759_),
    .C(_09723_),
    .Y(_09760_));
 AND2x2_ASAP7_75t_R _13707_ (.A(_08723_),
    .B(_09760_),
    .Y(_02930_));
 NOR2x1_ASAP7_75t_R _13708_ (.A(_01895_),
    .B(_09711_),
    .Y(_09761_));
 OA21x2_ASAP7_75t_R _13709_ (.A1(_09722_),
    .A2(_09723_),
    .B(_01520_),
    .Y(_09762_));
 AOI211x1_ASAP7_75t_R _13710_ (.A1(_01416_),
    .A2(_09721_),
    .B(_09762_),
    .C(_09726_),
    .Y(_09763_));
 OA21x2_ASAP7_75t_R _13711_ (.A1(_09761_),
    .A2(_09763_),
    .B(_09743_),
    .Y(_02931_));
 NOR2x1_ASAP7_75t_R _13712_ (.A(_01894_),
    .B(_09711_),
    .Y(_09764_));
 OA21x2_ASAP7_75t_R _13713_ (.A1(_09722_),
    .A2(_09723_),
    .B(_01519_),
    .Y(_09765_));
 AOI211x1_ASAP7_75t_R _13714_ (.A1(_01415_),
    .A2(_09721_),
    .B(_09765_),
    .C(_09726_),
    .Y(_09766_));
 OA21x2_ASAP7_75t_R _13715_ (.A1(_09764_),
    .A2(_09766_),
    .B(_09743_),
    .Y(_02932_));
 AND2x2_ASAP7_75t_R _13716_ (.A(_08723_),
    .B(_00006_),
    .Y(_02933_));
 NOR2x2_ASAP7_75t_R _13717_ (.A(_01209_),
    .B(_01210_),
    .Y(_09767_));
 BUFx6f_ASAP7_75t_R _13718_ (.A(_01313_),
    .Y(_09768_));
 INVx2_ASAP7_75t_R _13719_ (.A(_01316_),
    .Y(_09769_));
 INVx2_ASAP7_75t_R _13720_ (.A(_01317_),
    .Y(_09770_));
 AND4x1_ASAP7_75t_R _13721_ (.A(_01315_),
    .B(_09769_),
    .C(_09770_),
    .D(_01318_),
    .Y(_09771_));
 INVx2_ASAP7_75t_R _13722_ (.A(_01874_),
    .Y(_09772_));
 BUFx6f_ASAP7_75t_R _13723_ (.A(_01868_),
    .Y(_09773_));
 AO21x1_ASAP7_75t_R _13724_ (.A1(_01869_),
    .A2(_09772_),
    .B(_09773_),
    .Y(_09774_));
 OR2x2_ASAP7_75t_R _13725_ (.A(_09768_),
    .B(_01314_),
    .Y(_09775_));
 OA31x2_ASAP7_75t_R _13726_ (.A1(_09768_),
    .A2(_09771_),
    .A3(_09774_),
    .B1(_09775_),
    .Y(_09776_));
 INVx1_ASAP7_75t_R _13727_ (.A(_01209_),
    .Y(_09777_));
 NOR2x1_ASAP7_75t_R _13728_ (.A(_01212_),
    .B(_01213_),
    .Y(_09778_));
 AND2x2_ASAP7_75t_R _13729_ (.A(_01211_),
    .B(_01214_),
    .Y(_09779_));
 AND4x1_ASAP7_75t_R _13730_ (.A(_09777_),
    .B(_01215_),
    .C(_09778_),
    .D(_09779_),
    .Y(_09780_));
 OA21x2_ASAP7_75t_R _13731_ (.A1(_09767_),
    .A2(_09776_),
    .B(_09780_),
    .Y(_09781_));
 NOR2x2_ASAP7_75t_R _13732_ (.A(_09768_),
    .B(_01314_),
    .Y(_09782_));
 INVx1_ASAP7_75t_R _13733_ (.A(_09768_),
    .Y(_09783_));
 INVx1_ASAP7_75t_R _13734_ (.A(_01315_),
    .Y(_09784_));
 INVx1_ASAP7_75t_R _13735_ (.A(_01318_),
    .Y(_09785_));
 OR4x1_ASAP7_75t_R _13736_ (.A(_09784_),
    .B(_01316_),
    .C(_01317_),
    .D(_09785_),
    .Y(_09786_));
 AND2x2_ASAP7_75t_R _13737_ (.A(_09783_),
    .B(_09786_),
    .Y(_09787_));
 AND3x1_ASAP7_75t_R _13738_ (.A(_01210_),
    .B(_09778_),
    .C(_09779_),
    .Y(_09788_));
 INVx2_ASAP7_75t_R _13739_ (.A(_09773_),
    .Y(_09789_));
 AO21x1_ASAP7_75t_R _13740_ (.A1(_09789_),
    .A2(_01874_),
    .B(_01209_),
    .Y(_09790_));
 OAI21x1_ASAP7_75t_R _13741_ (.A1(_09788_),
    .A2(_09790_),
    .B(_01869_),
    .Y(_09791_));
 AO21x1_ASAP7_75t_R _13742_ (.A1(_09778_),
    .A2(_09779_),
    .B(_01209_),
    .Y(_09792_));
 BUFx6f_ASAP7_75t_R _13743_ (.A(_09792_),
    .Y(_09793_));
 OAI21x1_ASAP7_75t_R _13744_ (.A1(_00006_),
    .A2(_09793_),
    .B(_09773_),
    .Y(_09794_));
 NOR2x1_ASAP7_75t_R _13745_ (.A(_09768_),
    .B(_01319_),
    .Y(_09795_));
 AND5x2_ASAP7_75t_R _13746_ (.A(_01315_),
    .B(_09769_),
    .C(_09770_),
    .D(_01318_),
    .E(_09795_),
    .Y(_09796_));
 AO21x1_ASAP7_75t_R _13747_ (.A1(_01869_),
    .A2(_01874_),
    .B(_09773_),
    .Y(_09797_));
 OR2x6_ASAP7_75t_R _13748_ (.A(_01209_),
    .B(_01210_),
    .Y(_09798_));
 OAI21x1_ASAP7_75t_R _13749_ (.A1(_09793_),
    .A2(_09797_),
    .B(_09798_),
    .Y(_09799_));
 AO32x2_ASAP7_75t_R _13750_ (.A1(_09787_),
    .A2(_09791_),
    .A3(_09794_),
    .B1(_09796_),
    .B2(_09799_),
    .Y(_09800_));
 NOR2x1_ASAP7_75t_R _13751_ (.A(_09782_),
    .B(_09800_),
    .Y(_09801_));
 AND2x2_ASAP7_75t_R _13752_ (.A(_09781_),
    .B(_09801_),
    .Y(_09802_));
 BUFx6f_ASAP7_75t_R _13753_ (.A(_09802_),
    .Y(_09803_));
 INVx1_ASAP7_75t_R _13754_ (.A(_01215_),
    .Y(_09804_));
 NAND2x1_ASAP7_75t_R _13755_ (.A(_01211_),
    .B(_01214_),
    .Y(_09805_));
 OR5x2_ASAP7_75t_R _13756_ (.A(_01209_),
    .B(_01212_),
    .C(_01213_),
    .D(_09804_),
    .E(_09805_),
    .Y(_09806_));
 AO21x1_ASAP7_75t_R _13757_ (.A1(_09783_),
    .A2(_09786_),
    .B(_09806_),
    .Y(_09807_));
 AOI21x1_ASAP7_75t_R _13758_ (.A1(_09767_),
    .A2(_09796_),
    .B(_09772_),
    .Y(_09808_));
 AND2x2_ASAP7_75t_R _13759_ (.A(_01874_),
    .B(_09782_),
    .Y(_09809_));
 AOI221x1_ASAP7_75t_R _13760_ (.A1(_09772_),
    .A2(_09767_),
    .B1(_09796_),
    .B2(_09780_),
    .C(_09809_),
    .Y(_09810_));
 AND2x4_ASAP7_75t_R _13761_ (.A(_09789_),
    .B(_01869_),
    .Y(_09811_));
 AND4x1_ASAP7_75t_R _13762_ (.A(_09807_),
    .B(_09808_),
    .C(_09810_),
    .D(_09811_),
    .Y(_09812_));
 OR2x6_ASAP7_75t_R _13763_ (.A(_09781_),
    .B(_09812_),
    .Y(_09813_));
 NAND2x2_ASAP7_75t_R _13764_ (.A(_09801_),
    .B(_09813_),
    .Y(_09814_));
 OAI21x1_ASAP7_75t_R _13765_ (.A1(_09767_),
    .A2(_09776_),
    .B(_09780_),
    .Y(_09815_));
 AND2x2_ASAP7_75t_R _13766_ (.A(_09815_),
    .B(_09812_),
    .Y(_09816_));
 BUFx6f_ASAP7_75t_R _13767_ (.A(_09816_),
    .Y(_09817_));
 BUFx12f_ASAP7_75t_R _13768_ (.A(_08572_),
    .Y(_09818_));
 AO21x1_ASAP7_75t_R _13769_ (.A1(_01879_),
    .A2(_09817_),
    .B(_09818_),
    .Y(_09819_));
 AOI221x1_ASAP7_75t_R _13770_ (.A1(_01220_),
    .A2(_09803_),
    .B1(_09814_),
    .B2(_01324_),
    .C(_09819_),
    .Y(_02934_));
 AO21x1_ASAP7_75t_R _13771_ (.A1(_01878_),
    .A2(_09817_),
    .B(_09818_),
    .Y(_09820_));
 AOI221x1_ASAP7_75t_R _13772_ (.A1(_01219_),
    .A2(_09803_),
    .B1(_09814_),
    .B2(_01323_),
    .C(_09820_),
    .Y(_02935_));
 AO21x1_ASAP7_75t_R _13773_ (.A1(_01877_),
    .A2(_09817_),
    .B(_09818_),
    .Y(_09821_));
 AOI221x1_ASAP7_75t_R _13774_ (.A1(_01218_),
    .A2(_09803_),
    .B1(_09814_),
    .B2(_01322_),
    .C(_09821_),
    .Y(_02936_));
 AO21x1_ASAP7_75t_R _13775_ (.A1(_01876_),
    .A2(_09817_),
    .B(_09818_),
    .Y(_09822_));
 AOI221x1_ASAP7_75t_R _13776_ (.A1(_01217_),
    .A2(_09803_),
    .B1(_09814_),
    .B2(_01321_),
    .C(_09822_),
    .Y(_02937_));
 AO21x1_ASAP7_75t_R _13777_ (.A1(_01875_),
    .A2(_09817_),
    .B(_09818_),
    .Y(_09823_));
 AOI221x1_ASAP7_75t_R _13778_ (.A1(_01216_),
    .A2(_09803_),
    .B1(_09814_),
    .B2(_01320_),
    .C(_09823_),
    .Y(_02938_));
 INVx1_ASAP7_75t_R _13779_ (.A(_01319_),
    .Y(_09824_));
 AND3x1_ASAP7_75t_R _13780_ (.A(_09632_),
    .B(_09824_),
    .C(_09814_),
    .Y(_02939_));
 OR3x1_ASAP7_75t_R _13781_ (.A(_09207_),
    .B(_01318_),
    .C(_09817_),
    .Y(_09825_));
 OR2x2_ASAP7_75t_R _13782_ (.A(_08683_),
    .B(_01873_),
    .Y(_09826_));
 NAND2x1_ASAP7_75t_R _13783_ (.A(_09815_),
    .B(_09812_),
    .Y(_09827_));
 OAI22x1_ASAP7_75t_R _13784_ (.A1(_09803_),
    .A2(_09825_),
    .B1(_09826_),
    .B2(_09827_),
    .Y(_02940_));
 AO21x1_ASAP7_75t_R _13785_ (.A1(_09815_),
    .A2(_09812_),
    .B(_09770_),
    .Y(_09828_));
 NAND2x1_ASAP7_75t_R _13786_ (.A(_01872_),
    .B(_09817_),
    .Y(_09829_));
 BUFx12f_ASAP7_75t_R _13787_ (.A(_08876_),
    .Y(_09830_));
 OA211x2_ASAP7_75t_R _13788_ (.A1(_09803_),
    .A2(_09828_),
    .B(_09829_),
    .C(_09830_),
    .Y(_02941_));
 AO21x1_ASAP7_75t_R _13789_ (.A1(_09815_),
    .A2(_09812_),
    .B(_09769_),
    .Y(_09831_));
 NAND2x1_ASAP7_75t_R _13790_ (.A(_01871_),
    .B(_09817_),
    .Y(_09832_));
 OA211x2_ASAP7_75t_R _13791_ (.A1(_09802_),
    .A2(_09831_),
    .B(_09832_),
    .C(_09830_),
    .Y(_02942_));
 OR3x1_ASAP7_75t_R _13792_ (.A(_09207_),
    .B(_01315_),
    .C(_09816_),
    .Y(_09833_));
 OR2x2_ASAP7_75t_R _13793_ (.A(_08683_),
    .B(_01870_),
    .Y(_09834_));
 OAI22x1_ASAP7_75t_R _13794_ (.A1(_09803_),
    .A2(_09833_),
    .B1(_09834_),
    .B2(_09827_),
    .Y(_02943_));
 AND3x1_ASAP7_75t_R _13795_ (.A(_09632_),
    .B(_09775_),
    .C(_09800_),
    .Y(_02944_));
 INVx1_ASAP7_75t_R _13796_ (.A(_09813_),
    .Y(_09835_));
 AOI21x1_ASAP7_75t_R _13797_ (.A1(_09801_),
    .A2(_09835_),
    .B(_09687_),
    .Y(_02945_));
 AO21x1_ASAP7_75t_R _13798_ (.A1(_01867_),
    .A2(_09817_),
    .B(_09818_),
    .Y(_09836_));
 AOI221x1_ASAP7_75t_R _13799_ (.A1(_01208_),
    .A2(_09803_),
    .B1(_09814_),
    .B2(_01312_),
    .C(_09836_),
    .Y(_02946_));
 AO21x1_ASAP7_75t_R _13800_ (.A1(_01866_),
    .A2(_09817_),
    .B(_09818_),
    .Y(_09837_));
 AOI221x1_ASAP7_75t_R _13801_ (.A1(_01207_),
    .A2(_09803_),
    .B1(_09814_),
    .B2(_01311_),
    .C(_09837_),
    .Y(_02947_));
 INVx1_ASAP7_75t_R _13802_ (.A(_01869_),
    .Y(_09838_));
 AOI221x1_ASAP7_75t_R _13803_ (.A1(_09789_),
    .A2(_09772_),
    .B1(_09771_),
    .B2(_01314_),
    .C(_09768_),
    .Y(_09839_));
 AO31x2_ASAP7_75t_R _13804_ (.A1(_09783_),
    .A2(_00006_),
    .A3(_09786_),
    .B(_09789_),
    .Y(_09840_));
 INVx1_ASAP7_75t_R _13805_ (.A(_09793_),
    .Y(_09841_));
 OA211x2_ASAP7_75t_R _13806_ (.A1(_09838_),
    .A2(_09839_),
    .B(_09840_),
    .C(_09841_),
    .Y(_09842_));
 BUFx6f_ASAP7_75t_R _13807_ (.A(_09842_),
    .Y(_09843_));
 OAI21x1_ASAP7_75t_R _13808_ (.A1(_09806_),
    .A2(_09776_),
    .B(_09798_),
    .Y(_09844_));
 OA21x2_ASAP7_75t_R _13809_ (.A1(_09793_),
    .A2(_09797_),
    .B(_09798_),
    .Y(_09845_));
 OA21x2_ASAP7_75t_R _13810_ (.A1(_09782_),
    .A2(_09845_),
    .B(_09796_),
    .Y(_09846_));
 AOI221x1_ASAP7_75t_R _13811_ (.A1(_09780_),
    .A2(_09782_),
    .B1(_09796_),
    .B2(_09793_),
    .C(_01874_),
    .Y(_09847_));
 NAND3x1_ASAP7_75t_R _13812_ (.A(_09810_),
    .B(_09811_),
    .C(_09847_),
    .Y(_09848_));
 OR4x1_ASAP7_75t_R _13813_ (.A(_09843_),
    .B(_09844_),
    .C(_09846_),
    .D(_09848_),
    .Y(_09849_));
 BUFx12f_ASAP7_75t_R _13814_ (.A(_09849_),
    .Y(_09850_));
 NOR2x1_ASAP7_75t_R _13815_ (.A(_01879_),
    .B(_09850_),
    .Y(_09851_));
 INVx1_ASAP7_75t_R _13816_ (.A(_01324_),
    .Y(_09852_));
 OR2x6_ASAP7_75t_R _13817_ (.A(_09843_),
    .B(_09844_),
    .Y(_09853_));
 BUFx6f_ASAP7_75t_R _13818_ (.A(_09853_),
    .Y(_09854_));
 BUFx6f_ASAP7_75t_R _13819_ (.A(_09849_),
    .Y(_09855_));
 BUFx12f_ASAP7_75t_R _13820_ (.A(_09843_),
    .Y(_09856_));
 BUFx6f_ASAP7_75t_R _13821_ (.A(_09844_),
    .Y(_09857_));
 OAI21x1_ASAP7_75t_R _13822_ (.A1(_09856_),
    .A2(_09857_),
    .B(_01220_),
    .Y(_09858_));
 OA211x2_ASAP7_75t_R _13823_ (.A1(_09852_),
    .A2(_09854_),
    .B(_09855_),
    .C(_09858_),
    .Y(_09859_));
 OA21x2_ASAP7_75t_R _13824_ (.A1(_09851_),
    .A2(_09859_),
    .B(_09743_),
    .Y(_02948_));
 NOR2x1_ASAP7_75t_R _13825_ (.A(_01878_),
    .B(_09850_),
    .Y(_09860_));
 INVx1_ASAP7_75t_R _13826_ (.A(_01323_),
    .Y(_09861_));
 OAI21x1_ASAP7_75t_R _13827_ (.A1(_09856_),
    .A2(_09857_),
    .B(_01219_),
    .Y(_09862_));
 OA211x2_ASAP7_75t_R _13828_ (.A1(_09861_),
    .A2(_09854_),
    .B(_09855_),
    .C(_09862_),
    .Y(_09863_));
 OA21x2_ASAP7_75t_R _13829_ (.A1(_09860_),
    .A2(_09863_),
    .B(_09743_),
    .Y(_02949_));
 NOR2x1_ASAP7_75t_R _13830_ (.A(_01877_),
    .B(_09850_),
    .Y(_09864_));
 INVx1_ASAP7_75t_R _13831_ (.A(_01322_),
    .Y(_09865_));
 OAI21x1_ASAP7_75t_R _13832_ (.A1(_09856_),
    .A2(_09857_),
    .B(_01218_),
    .Y(_09866_));
 OA211x2_ASAP7_75t_R _13833_ (.A1(_09865_),
    .A2(_09854_),
    .B(_09855_),
    .C(_09866_),
    .Y(_09867_));
 OA21x2_ASAP7_75t_R _13834_ (.A1(_09864_),
    .A2(_09867_),
    .B(_09743_),
    .Y(_02950_));
 NOR2x1_ASAP7_75t_R _13835_ (.A(_01876_),
    .B(_09850_),
    .Y(_09868_));
 INVx1_ASAP7_75t_R _13836_ (.A(_01321_),
    .Y(_09869_));
 OAI21x1_ASAP7_75t_R _13837_ (.A1(_09856_),
    .A2(_09857_),
    .B(_01217_),
    .Y(_09870_));
 OA211x2_ASAP7_75t_R _13838_ (.A1(_09869_),
    .A2(_09854_),
    .B(_09855_),
    .C(_09870_),
    .Y(_09871_));
 BUFx6f_ASAP7_75t_R _13839_ (.A(_08665_),
    .Y(_09872_));
 OA21x2_ASAP7_75t_R _13840_ (.A1(_09868_),
    .A2(_09871_),
    .B(_09872_),
    .Y(_02951_));
 NOR2x1_ASAP7_75t_R _13841_ (.A(_01875_),
    .B(_09850_),
    .Y(_09873_));
 INVx1_ASAP7_75t_R _13842_ (.A(_01320_),
    .Y(_09874_));
 OAI21x1_ASAP7_75t_R _13843_ (.A1(_09856_),
    .A2(_09857_),
    .B(_01216_),
    .Y(_09875_));
 OA211x2_ASAP7_75t_R _13844_ (.A1(_09874_),
    .A2(_09854_),
    .B(_09855_),
    .C(_09875_),
    .Y(_09876_));
 OA21x2_ASAP7_75t_R _13845_ (.A1(_09873_),
    .A2(_09876_),
    .B(_09872_),
    .Y(_02952_));
 OAI21x1_ASAP7_75t_R _13846_ (.A1(_09856_),
    .A2(_09857_),
    .B(_01215_),
    .Y(_09877_));
 OAI21x1_ASAP7_75t_R _13847_ (.A1(_09824_),
    .A2(_09854_),
    .B(_09877_),
    .Y(_09878_));
 AOI21x1_ASAP7_75t_R _13848_ (.A1(_09850_),
    .A2(_09878_),
    .B(_09687_),
    .Y(_02953_));
 NOR2x1_ASAP7_75t_R _13849_ (.A(_01873_),
    .B(_09850_),
    .Y(_09879_));
 OAI21x1_ASAP7_75t_R _13850_ (.A1(_09856_),
    .A2(_09857_),
    .B(_01214_),
    .Y(_09880_));
 OA211x2_ASAP7_75t_R _13851_ (.A1(_09785_),
    .A2(_09854_),
    .B(_09855_),
    .C(_09880_),
    .Y(_09881_));
 OA21x2_ASAP7_75t_R _13852_ (.A1(_09879_),
    .A2(_09881_),
    .B(_09872_),
    .Y(_02954_));
 NOR2x1_ASAP7_75t_R _13853_ (.A(_01872_),
    .B(_09850_),
    .Y(_09882_));
 OAI21x1_ASAP7_75t_R _13854_ (.A1(_09856_),
    .A2(_09857_),
    .B(_01213_),
    .Y(_09883_));
 OA211x2_ASAP7_75t_R _13855_ (.A1(_09770_),
    .A2(_09854_),
    .B(_09855_),
    .C(_09883_),
    .Y(_09884_));
 OA21x2_ASAP7_75t_R _13856_ (.A1(_09882_),
    .A2(_09884_),
    .B(_09872_),
    .Y(_02955_));
 NOR2x1_ASAP7_75t_R _13857_ (.A(_01871_),
    .B(_09850_),
    .Y(_09885_));
 OAI21x1_ASAP7_75t_R _13858_ (.A1(_09843_),
    .A2(_09857_),
    .B(_01212_),
    .Y(_09886_));
 OA211x2_ASAP7_75t_R _13859_ (.A1(_09769_),
    .A2(_09854_),
    .B(_09855_),
    .C(_09886_),
    .Y(_09887_));
 OA21x2_ASAP7_75t_R _13860_ (.A1(_09885_),
    .A2(_09887_),
    .B(_09872_),
    .Y(_02956_));
 NOR2x1_ASAP7_75t_R _13861_ (.A(_01870_),
    .B(_09850_),
    .Y(_09888_));
 OAI21x1_ASAP7_75t_R _13862_ (.A1(_09843_),
    .A2(_09844_),
    .B(_01211_),
    .Y(_09889_));
 OA211x2_ASAP7_75t_R _13863_ (.A1(_09784_),
    .A2(_09854_),
    .B(_09849_),
    .C(_09889_),
    .Y(_09890_));
 OA21x2_ASAP7_75t_R _13864_ (.A1(_09888_),
    .A2(_09890_),
    .B(_09872_),
    .Y(_02957_));
 NOR2x1_ASAP7_75t_R _13865_ (.A(_09806_),
    .B(_09776_),
    .Y(_09891_));
 OA211x2_ASAP7_75t_R _13866_ (.A1(_09856_),
    .A2(_09891_),
    .B(_09830_),
    .C(_09798_),
    .Y(_02958_));
 OR3x1_ASAP7_75t_R _13867_ (.A(_09856_),
    .B(_09857_),
    .C(_09846_),
    .Y(_09892_));
 INVx1_ASAP7_75t_R _13868_ (.A(_09892_),
    .Y(_09893_));
 AOI21x1_ASAP7_75t_R _13869_ (.A1(_09893_),
    .A2(_09848_),
    .B(_09687_),
    .Y(_02959_));
 NOR2x1_ASAP7_75t_R _13870_ (.A(_01867_),
    .B(_09855_),
    .Y(_09894_));
 INVx1_ASAP7_75t_R _13871_ (.A(_01312_),
    .Y(_09895_));
 OAI21x1_ASAP7_75t_R _13872_ (.A1(_09843_),
    .A2(_09844_),
    .B(_01208_),
    .Y(_09896_));
 OA211x2_ASAP7_75t_R _13873_ (.A1(_09895_),
    .A2(_09853_),
    .B(_09849_),
    .C(_09896_),
    .Y(_09897_));
 OA21x2_ASAP7_75t_R _13874_ (.A1(_09894_),
    .A2(_09897_),
    .B(_09872_),
    .Y(_02960_));
 NOR2x1_ASAP7_75t_R _13875_ (.A(_01866_),
    .B(_09855_),
    .Y(_09898_));
 INVx1_ASAP7_75t_R _13876_ (.A(_01311_),
    .Y(_09899_));
 OAI21x1_ASAP7_75t_R _13877_ (.A1(_09843_),
    .A2(_09844_),
    .B(_01207_),
    .Y(_09900_));
 OA211x2_ASAP7_75t_R _13878_ (.A1(_09899_),
    .A2(_09853_),
    .B(_09849_),
    .C(_09900_),
    .Y(_09901_));
 OA21x2_ASAP7_75t_R _13879_ (.A1(_09898_),
    .A2(_09901_),
    .B(_09872_),
    .Y(_02961_));
 OA21x2_ASAP7_75t_R _13880_ (.A1(_09788_),
    .A2(_09790_),
    .B(_01869_),
    .Y(_09902_));
 OA21x2_ASAP7_75t_R _13881_ (.A1(_00006_),
    .A2(_09793_),
    .B(_09773_),
    .Y(_09903_));
 OA31x2_ASAP7_75t_R _13882_ (.A1(_09782_),
    .A2(_09902_),
    .A3(_09903_),
    .B1(_09787_),
    .Y(_09904_));
 OA211x2_ASAP7_75t_R _13883_ (.A1(_09838_),
    .A2(_09839_),
    .B(_09840_),
    .C(_09798_),
    .Y(_09905_));
 NOR3x1_ASAP7_75t_R _13884_ (.A(_09793_),
    .B(_09904_),
    .C(_09905_),
    .Y(_09906_));
 BUFx6f_ASAP7_75t_R _13885_ (.A(_09906_),
    .Y(_09907_));
 NAND2x1_ASAP7_75t_R _13886_ (.A(_01220_),
    .B(_09907_),
    .Y(_09908_));
 OR3x2_ASAP7_75t_R _13887_ (.A(_09793_),
    .B(_09904_),
    .C(_09905_),
    .Y(_09909_));
 BUFx6f_ASAP7_75t_R _13888_ (.A(_09909_),
    .Y(_09910_));
 NAND2x1_ASAP7_75t_R _13889_ (.A(_01324_),
    .B(_09910_),
    .Y(_09911_));
 AO21x1_ASAP7_75t_R _13890_ (.A1(_09807_),
    .A2(_09808_),
    .B(_09847_),
    .Y(_09912_));
 AND2x2_ASAP7_75t_R _13891_ (.A(_01869_),
    .B(_09810_),
    .Y(_09913_));
 AOI21x1_ASAP7_75t_R _13892_ (.A1(_09912_),
    .A2(_09913_),
    .B(_09773_),
    .Y(_09914_));
 NOR2x1_ASAP7_75t_R _13893_ (.A(_08572_),
    .B(_09914_),
    .Y(_09915_));
 BUFx3_ASAP7_75t_R _13894_ (.A(_09914_),
    .Y(_09916_));
 NOR2x1_ASAP7_75t_R _13895_ (.A(_09318_),
    .B(_01879_),
    .Y(_09917_));
 AO32x1_ASAP7_75t_R _13896_ (.A1(_09908_),
    .A2(_09911_),
    .A3(_09915_),
    .B1(_09916_),
    .B2(_09917_),
    .Y(_02962_));
 BUFx6f_ASAP7_75t_R _13897_ (.A(_09915_),
    .Y(_09918_));
 NAND2x1_ASAP7_75t_R _13898_ (.A(_01219_),
    .B(_09907_),
    .Y(_09919_));
 NAND2x1_ASAP7_75t_R _13899_ (.A(_01323_),
    .B(_09910_),
    .Y(_09920_));
 NOR2x1_ASAP7_75t_R _13900_ (.A(_09318_),
    .B(_01878_),
    .Y(_09921_));
 AO32x1_ASAP7_75t_R _13901_ (.A1(_09918_),
    .A2(_09919_),
    .A3(_09920_),
    .B1(_09916_),
    .B2(_09921_),
    .Y(_02963_));
 NAND2x1_ASAP7_75t_R _13902_ (.A(_01218_),
    .B(_09907_),
    .Y(_09922_));
 NAND2x1_ASAP7_75t_R _13903_ (.A(_01322_),
    .B(_09910_),
    .Y(_09923_));
 BUFx12f_ASAP7_75t_R _13904_ (.A(_08656_),
    .Y(_09924_));
 NOR2x1_ASAP7_75t_R _13905_ (.A(_09924_),
    .B(_01877_),
    .Y(_09925_));
 AO32x1_ASAP7_75t_R _13906_ (.A1(_09918_),
    .A2(_09922_),
    .A3(_09923_),
    .B1(_09916_),
    .B2(_09925_),
    .Y(_02964_));
 NAND2x1_ASAP7_75t_R _13907_ (.A(_01217_),
    .B(_09907_),
    .Y(_09926_));
 NAND2x1_ASAP7_75t_R _13908_ (.A(_01321_),
    .B(_09910_),
    .Y(_09927_));
 NOR2x1_ASAP7_75t_R _13909_ (.A(_09924_),
    .B(_01876_),
    .Y(_09928_));
 AO32x1_ASAP7_75t_R _13910_ (.A1(_09918_),
    .A2(_09926_),
    .A3(_09927_),
    .B1(_09916_),
    .B2(_09928_),
    .Y(_02965_));
 NAND2x1_ASAP7_75t_R _13911_ (.A(_01216_),
    .B(_09907_),
    .Y(_09929_));
 NAND2x1_ASAP7_75t_R _13912_ (.A(_01320_),
    .B(_09910_),
    .Y(_09930_));
 NOR2x1_ASAP7_75t_R _13913_ (.A(_09924_),
    .B(_01875_),
    .Y(_09931_));
 AO32x1_ASAP7_75t_R _13914_ (.A1(_09918_),
    .A2(_09929_),
    .A3(_09930_),
    .B1(_09916_),
    .B2(_09931_),
    .Y(_02966_));
 NAND2x1_ASAP7_75t_R _13915_ (.A(_01215_),
    .B(_09907_),
    .Y(_09932_));
 NAND2x1_ASAP7_75t_R _13916_ (.A(_01319_),
    .B(_09910_),
    .Y(_09933_));
 BUFx12f_ASAP7_75t_R _13917_ (.A(_08656_),
    .Y(_09934_));
 NOR2x1_ASAP7_75t_R _13918_ (.A(_09934_),
    .B(_01874_),
    .Y(_09935_));
 AO32x1_ASAP7_75t_R _13919_ (.A1(_09918_),
    .A2(_09932_),
    .A3(_09933_),
    .B1(_09935_),
    .B2(_09916_),
    .Y(_02967_));
 NAND2x1_ASAP7_75t_R _13920_ (.A(_01214_),
    .B(_09907_),
    .Y(_09936_));
 NAND2x1_ASAP7_75t_R _13921_ (.A(_01318_),
    .B(_09910_),
    .Y(_09937_));
 INVx1_ASAP7_75t_R _13922_ (.A(_09826_),
    .Y(_09938_));
 AO32x1_ASAP7_75t_R _13923_ (.A1(_09918_),
    .A2(_09936_),
    .A3(_09937_),
    .B1(_09916_),
    .B2(_09938_),
    .Y(_02968_));
 NAND2x1_ASAP7_75t_R _13924_ (.A(_01213_),
    .B(_09907_),
    .Y(_09939_));
 NAND2x1_ASAP7_75t_R _13925_ (.A(_01317_),
    .B(_09910_),
    .Y(_09940_));
 NOR2x1_ASAP7_75t_R _13926_ (.A(_09924_),
    .B(_01872_),
    .Y(_09941_));
 AO32x1_ASAP7_75t_R _13927_ (.A1(_09918_),
    .A2(_09939_),
    .A3(_09940_),
    .B1(_09916_),
    .B2(_09941_),
    .Y(_02969_));
 NAND2x1_ASAP7_75t_R _13928_ (.A(_01212_),
    .B(_09907_),
    .Y(_09942_));
 NAND2x1_ASAP7_75t_R _13929_ (.A(_01316_),
    .B(_09910_),
    .Y(_09943_));
 NOR2x1_ASAP7_75t_R _13930_ (.A(_09924_),
    .B(_01871_),
    .Y(_09944_));
 AO32x1_ASAP7_75t_R _13931_ (.A1(_09918_),
    .A2(_09942_),
    .A3(_09943_),
    .B1(_09916_),
    .B2(_09944_),
    .Y(_02970_));
 NAND2x1_ASAP7_75t_R _13932_ (.A(_01211_),
    .B(_09907_),
    .Y(_09945_));
 NAND2x1_ASAP7_75t_R _13933_ (.A(_01315_),
    .B(_09910_),
    .Y(_09946_));
 INVx1_ASAP7_75t_R _13934_ (.A(_09834_),
    .Y(_09947_));
 AO32x1_ASAP7_75t_R _13935_ (.A1(_09918_),
    .A2(_09945_),
    .A3(_09946_),
    .B1(_09916_),
    .B2(_09947_),
    .Y(_02971_));
 NAND2x1_ASAP7_75t_R _13936_ (.A(_09810_),
    .B(_09912_),
    .Y(_09948_));
 AND3x1_ASAP7_75t_R _13937_ (.A(_09632_),
    .B(_09811_),
    .C(_09948_),
    .Y(_02972_));
 NOR2x1_ASAP7_75t_R _13938_ (.A(_09793_),
    .B(_09905_),
    .Y(_09949_));
 OR3x1_ASAP7_75t_R _13939_ (.A(_09914_),
    .B(_09904_),
    .C(_09949_),
    .Y(_09950_));
 AND2x2_ASAP7_75t_R _13940_ (.A(_08723_),
    .B(_09950_),
    .Y(_02973_));
 NAND2x1_ASAP7_75t_R _13941_ (.A(_01208_),
    .B(_09906_),
    .Y(_09951_));
 NAND2x1_ASAP7_75t_R _13942_ (.A(_01312_),
    .B(_09909_),
    .Y(_09952_));
 NOR2x1_ASAP7_75t_R _13943_ (.A(_09924_),
    .B(_01867_),
    .Y(_09953_));
 AO32x1_ASAP7_75t_R _13944_ (.A1(_09918_),
    .A2(_09951_),
    .A3(_09952_),
    .B1(_09914_),
    .B2(_09953_),
    .Y(_02974_));
 NAND2x1_ASAP7_75t_R _13945_ (.A(_01207_),
    .B(_09906_),
    .Y(_09954_));
 NAND2x1_ASAP7_75t_R _13946_ (.A(_01311_),
    .B(_09909_),
    .Y(_09955_));
 NOR2x1_ASAP7_75t_R _13947_ (.A(_09924_),
    .B(_01866_),
    .Y(_09956_));
 AO32x1_ASAP7_75t_R _13948_ (.A1(_09915_),
    .A2(_09954_),
    .A3(_09955_),
    .B1(_09914_),
    .B2(_09956_),
    .Y(_02975_));
 BUFx6f_ASAP7_75t_R _13949_ (.A(_08722_),
    .Y(_09957_));
 AND2x2_ASAP7_75t_R _13950_ (.A(_09957_),
    .B(_00007_),
    .Y(_02976_));
 OR2x2_ASAP7_75t_R _13951_ (.A(_01001_),
    .B(_01002_),
    .Y(_09958_));
 BUFx6f_ASAP7_75t_R _13952_ (.A(_09958_),
    .Y(_09959_));
 BUFx6f_ASAP7_75t_R _13953_ (.A(_01854_),
    .Y(_09960_));
 INVx2_ASAP7_75t_R _13954_ (.A(_09960_),
    .Y(_09961_));
 INVx2_ASAP7_75t_R _13955_ (.A(_01107_),
    .Y(_09962_));
 OR2x6_ASAP7_75t_R _13956_ (.A(_01109_),
    .B(_01110_),
    .Y(_09963_));
 INVx1_ASAP7_75t_R _13957_ (.A(_01105_),
    .Y(_09964_));
 OA31x2_ASAP7_75t_R _13958_ (.A1(_09962_),
    .A2(_01108_),
    .A3(_09963_),
    .B1(_09964_),
    .Y(_09965_));
 BUFx6f_ASAP7_75t_R _13959_ (.A(_01855_),
    .Y(_09966_));
 BUFx6f_ASAP7_75t_R _13960_ (.A(_01860_),
    .Y(_09967_));
 INVx2_ASAP7_75t_R _13961_ (.A(_09967_),
    .Y(_09968_));
 NAND2x1_ASAP7_75t_R _13962_ (.A(_09966_),
    .B(_09968_),
    .Y(_09969_));
 INVx1_ASAP7_75t_R _13963_ (.A(_01106_),
    .Y(_09970_));
 AO32x2_ASAP7_75t_R _13964_ (.A1(_09961_),
    .A2(_09965_),
    .A3(_09969_),
    .B1(_09964_),
    .B2(_09970_),
    .Y(_09971_));
 INVx1_ASAP7_75t_R _13965_ (.A(_01003_),
    .Y(_09972_));
 INVx1_ASAP7_75t_R _13966_ (.A(_01007_),
    .Y(_09973_));
 OR2x2_ASAP7_75t_R _13967_ (.A(_01005_),
    .B(_01006_),
    .Y(_09974_));
 OR5x2_ASAP7_75t_R _13968_ (.A(_01001_),
    .B(_09972_),
    .C(_01004_),
    .D(_09973_),
    .E(_09974_),
    .Y(_09975_));
 AOI21x1_ASAP7_75t_R _13969_ (.A1(_09959_),
    .A2(_09971_),
    .B(_09975_),
    .Y(_09976_));
 OR2x2_ASAP7_75t_R _13970_ (.A(_01105_),
    .B(_01106_),
    .Y(_09977_));
 AND2x2_ASAP7_75t_R _13971_ (.A(_09964_),
    .B(_01106_),
    .Y(_09978_));
 OR3x1_ASAP7_75t_R _13972_ (.A(_09962_),
    .B(_01108_),
    .C(_09963_),
    .Y(_09979_));
 AO221x1_ASAP7_75t_R _13973_ (.A1(_09977_),
    .A2(_09975_),
    .B1(_09978_),
    .B2(_09979_),
    .C(_09968_),
    .Y(_09980_));
 NOR2x1_ASAP7_75t_R _13974_ (.A(_01001_),
    .B(_01002_),
    .Y(_09981_));
 INVx1_ASAP7_75t_R _13975_ (.A(_01108_),
    .Y(_09982_));
 NOR2x1_ASAP7_75t_R _13976_ (.A(_01109_),
    .B(_01110_),
    .Y(_09983_));
 NOR2x1_ASAP7_75t_R _13977_ (.A(_01105_),
    .B(_01111_),
    .Y(_09984_));
 AND4x1_ASAP7_75t_R _13978_ (.A(_01107_),
    .B(_09982_),
    .C(_09983_),
    .D(_09984_),
    .Y(_09985_));
 INVx1_ASAP7_75t_R _13979_ (.A(_01001_),
    .Y(_09986_));
 INVx2_ASAP7_75t_R _13980_ (.A(_01004_),
    .Y(_09987_));
 NOR2x1_ASAP7_75t_R _13981_ (.A(_01005_),
    .B(_01006_),
    .Y(_09988_));
 AND5x2_ASAP7_75t_R _13982_ (.A(_09986_),
    .B(_01003_),
    .C(_09987_),
    .D(_01007_),
    .E(_09988_),
    .Y(_09989_));
 AOI22x1_ASAP7_75t_R _13983_ (.A1(_09968_),
    .A2(_09981_),
    .B1(_09985_),
    .B2(_09989_),
    .Y(_09990_));
 OR5x2_ASAP7_75t_R _13984_ (.A(_01105_),
    .B(_09962_),
    .C(_01108_),
    .D(_01111_),
    .E(_09963_),
    .Y(_09991_));
 AND2x2_ASAP7_75t_R _13985_ (.A(_09961_),
    .B(_09967_),
    .Y(_09992_));
 OA211x2_ASAP7_75t_R _13986_ (.A1(_09959_),
    .A2(_09991_),
    .B(_09966_),
    .C(_09992_),
    .Y(_09993_));
 AND3x4_ASAP7_75t_R _13987_ (.A(_09980_),
    .B(_09990_),
    .C(_09993_),
    .Y(_09994_));
 AO31x2_ASAP7_75t_R _13988_ (.A1(_01003_),
    .A2(_09987_),
    .A3(_09988_),
    .B(_01001_),
    .Y(_09995_));
 OR2x6_ASAP7_75t_R _13989_ (.A(_09960_),
    .B(_09967_),
    .Y(_09996_));
 OA22x2_ASAP7_75t_R _13990_ (.A1(_09960_),
    .A2(_09966_),
    .B1(_09959_),
    .B2(_09996_),
    .Y(_09997_));
 AND2x2_ASAP7_75t_R _13991_ (.A(_09995_),
    .B(_09997_),
    .Y(_09998_));
 AND3x1_ASAP7_75t_R _13992_ (.A(_01107_),
    .B(_09982_),
    .C(_09983_),
    .Y(_09999_));
 AND2x2_ASAP7_75t_R _13993_ (.A(_09960_),
    .B(_00007_),
    .Y(_10000_));
 AO31x2_ASAP7_75t_R _13994_ (.A1(_09961_),
    .A2(_09966_),
    .A3(_09967_),
    .B(_10000_),
    .Y(_10001_));
 OR3x1_ASAP7_75t_R _13995_ (.A(_01105_),
    .B(_09999_),
    .C(_10001_),
    .Y(_10002_));
 AO21x1_ASAP7_75t_R _13996_ (.A1(_09966_),
    .A2(_09967_),
    .B(_09960_),
    .Y(_10003_));
 OA21x2_ASAP7_75t_R _13997_ (.A1(_09995_),
    .A2(_10003_),
    .B(_09959_),
    .Y(_10004_));
 OA222x2_ASAP7_75t_R _13998_ (.A1(_01105_),
    .A2(_01106_),
    .B1(_09998_),
    .B2(_10002_),
    .C1(_09991_),
    .C2(_10004_),
    .Y(_10005_));
 OA21x2_ASAP7_75t_R _13999_ (.A1(_09976_),
    .A2(_09994_),
    .B(_10005_),
    .Y(_10006_));
 BUFx6f_ASAP7_75t_R _14000_ (.A(_10006_),
    .Y(_10007_));
 AO21x2_ASAP7_75t_R _14001_ (.A1(_09959_),
    .A2(_09971_),
    .B(_09975_),
    .Y(_10008_));
 NAND2x2_ASAP7_75t_R _14002_ (.A(_10008_),
    .B(_09994_),
    .Y(_10009_));
 NAND2x2_ASAP7_75t_R _14003_ (.A(_10005_),
    .B(_09976_),
    .Y(_10010_));
 OA222x2_ASAP7_75t_R _14004_ (.A1(_01116_),
    .A2(_10007_),
    .B1(_10009_),
    .B2(_01865_),
    .C1(_10010_),
    .C2(_01012_),
    .Y(_10011_));
 NOR2x1_ASAP7_75t_R _14005_ (.A(_08942_),
    .B(_10011_),
    .Y(_02977_));
 BUFx12f_ASAP7_75t_R _14006_ (.A(_08656_),
    .Y(_10012_));
 BUFx12f_ASAP7_75t_R _14007_ (.A(_10012_),
    .Y(_10013_));
 OA222x2_ASAP7_75t_R _14008_ (.A1(_01115_),
    .A2(_10007_),
    .B1(_10009_),
    .B2(_01864_),
    .C1(_10010_),
    .C2(_01011_),
    .Y(_10014_));
 NOR2x1_ASAP7_75t_R _14009_ (.A(_10013_),
    .B(_10014_),
    .Y(_02978_));
 OA222x2_ASAP7_75t_R _14010_ (.A1(_01114_),
    .A2(_10007_),
    .B1(_10009_),
    .B2(_01863_),
    .C1(_10010_),
    .C2(_01010_),
    .Y(_10015_));
 NOR2x1_ASAP7_75t_R _14011_ (.A(_10013_),
    .B(_10015_),
    .Y(_02979_));
 OA222x2_ASAP7_75t_R _14012_ (.A1(_01113_),
    .A2(_10007_),
    .B1(_10009_),
    .B2(_01862_),
    .C1(_10010_),
    .C2(_01009_),
    .Y(_10016_));
 NOR2x1_ASAP7_75t_R _14013_ (.A(_10013_),
    .B(_10016_),
    .Y(_02980_));
 OA222x2_ASAP7_75t_R _14014_ (.A1(_01112_),
    .A2(_10007_),
    .B1(_10009_),
    .B2(_01861_),
    .C1(_10010_),
    .C2(_01008_),
    .Y(_10017_));
 NOR2x1_ASAP7_75t_R _14015_ (.A(_10013_),
    .B(_10017_),
    .Y(_02981_));
 OR3x1_ASAP7_75t_R _14016_ (.A(_08657_),
    .B(_01111_),
    .C(_10007_),
    .Y(_10018_));
 INVx1_ASAP7_75t_R _14017_ (.A(_10018_),
    .Y(_02982_));
 INVx2_ASAP7_75t_R _14018_ (.A(_10007_),
    .Y(_10019_));
 INVx2_ASAP7_75t_R _14019_ (.A(_10009_),
    .Y(_10020_));
 AOI221x1_ASAP7_75t_R _14020_ (.A1(_01110_),
    .A2(_10019_),
    .B1(_10020_),
    .B2(_01859_),
    .C(_09145_),
    .Y(_02983_));
 AOI221x1_ASAP7_75t_R _14021_ (.A1(_01109_),
    .A2(_10019_),
    .B1(_10020_),
    .B2(_01858_),
    .C(_09145_),
    .Y(_02984_));
 BUFx12f_ASAP7_75t_R _14022_ (.A(_08641_),
    .Y(_10021_));
 AOI221x1_ASAP7_75t_R _14023_ (.A1(_01108_),
    .A2(_10019_),
    .B1(_10020_),
    .B2(_01857_),
    .C(_10021_),
    .Y(_02985_));
 OAI22x1_ASAP7_75t_R _14024_ (.A1(_01107_),
    .A2(_10007_),
    .B1(_10009_),
    .B2(_01856_),
    .Y(_10022_));
 AND2x2_ASAP7_75t_R _14025_ (.A(_09957_),
    .B(_10022_),
    .Y(_02986_));
 OAI22x1_ASAP7_75t_R _14026_ (.A1(_09998_),
    .A2(_10002_),
    .B1(_09991_),
    .B2(_10004_),
    .Y(_10023_));
 AND3x1_ASAP7_75t_R _14027_ (.A(_09632_),
    .B(_09977_),
    .C(_10023_),
    .Y(_02987_));
 NAND2x1_ASAP7_75t_R _14028_ (.A(_10005_),
    .B(_10008_),
    .Y(_10024_));
 OA21x2_ASAP7_75t_R _14029_ (.A1(_09994_),
    .A2(_10024_),
    .B(_09872_),
    .Y(_02988_));
 OA222x2_ASAP7_75t_R _14030_ (.A1(_01104_),
    .A2(_10007_),
    .B1(_10009_),
    .B2(_01853_),
    .C1(_10010_),
    .C2(_01000_),
    .Y(_10025_));
 NOR2x1_ASAP7_75t_R _14031_ (.A(_10013_),
    .B(_10025_),
    .Y(_02989_));
 OA222x2_ASAP7_75t_R _14032_ (.A1(_01103_),
    .A2(_10007_),
    .B1(_10009_),
    .B2(_01852_),
    .C1(_10010_),
    .C2(_00999_),
    .Y(_10026_));
 NOR2x1_ASAP7_75t_R _14033_ (.A(_10013_),
    .B(_10026_),
    .Y(_02990_));
 AO21x1_ASAP7_75t_R _14034_ (.A1(_09961_),
    .A2(_09967_),
    .B(_10000_),
    .Y(_10027_));
 NOR2x1_ASAP7_75t_R _14035_ (.A(_01105_),
    .B(_01106_),
    .Y(_10028_));
 NOR2x1_ASAP7_75t_R _14036_ (.A(_09960_),
    .B(_09966_),
    .Y(_10029_));
 AO31x2_ASAP7_75t_R _14037_ (.A1(_09961_),
    .A2(_09967_),
    .A3(_10028_),
    .B(_10029_),
    .Y(_10030_));
 AO21x2_ASAP7_75t_R _14038_ (.A1(_09965_),
    .A2(_10027_),
    .B(_10030_),
    .Y(_10031_));
 AND3x1_ASAP7_75t_R _14039_ (.A(_01003_),
    .B(_09987_),
    .C(_09988_),
    .Y(_10032_));
 NOR2x1_ASAP7_75t_R _14040_ (.A(_01001_),
    .B(_10032_),
    .Y(_10033_));
 AO221x1_ASAP7_75t_R _14041_ (.A1(_09989_),
    .A2(_09971_),
    .B1(_10031_),
    .B2(_10033_),
    .C(_09981_),
    .Y(_10034_));
 AND2x2_ASAP7_75t_R _14042_ (.A(_01116_),
    .B(_09959_),
    .Y(_10035_));
 AOI22x1_ASAP7_75t_R _14043_ (.A1(_09989_),
    .A2(_09971_),
    .B1(_10031_),
    .B2(_10033_),
    .Y(_10036_));
 AO221x1_ASAP7_75t_R _14044_ (.A1(_01012_),
    .A2(_10034_),
    .B1(_10035_),
    .B2(_10036_),
    .C(_09207_),
    .Y(_10037_));
 OA211x2_ASAP7_75t_R _14045_ (.A1(_10028_),
    .A2(_10004_),
    .B(_09984_),
    .C(_09999_),
    .Y(_10038_));
 OR2x6_ASAP7_75t_R _14046_ (.A(_10034_),
    .B(_10038_),
    .Y(_10039_));
 AND3x1_ASAP7_75t_R _14047_ (.A(_09966_),
    .B(_09980_),
    .C(_09990_),
    .Y(_10040_));
 AO21x1_ASAP7_75t_R _14048_ (.A1(_09981_),
    .A2(_09985_),
    .B(_09968_),
    .Y(_10041_));
 AO221x1_ASAP7_75t_R _14049_ (.A1(_09995_),
    .A2(_09985_),
    .B1(_09989_),
    .B2(_10028_),
    .C(_09967_),
    .Y(_10042_));
 NAND2x1_ASAP7_75t_R _14050_ (.A(_10041_),
    .B(_10042_),
    .Y(_10043_));
 AOI21x1_ASAP7_75t_R _14051_ (.A1(_10040_),
    .A2(_10043_),
    .B(_09960_),
    .Y(_10044_));
 NOR3x1_ASAP7_75t_R _14052_ (.A(_09996_),
    .B(_10039_),
    .C(_10044_),
    .Y(_10045_));
 BUFx12f_ASAP7_75t_R _14053_ (.A(_10045_),
    .Y(_10046_));
 BUFx6f_ASAP7_75t_R _14054_ (.A(_08572_),
    .Y(_10047_));
 BUFx6f_ASAP7_75t_R _14055_ (.A(_09996_),
    .Y(_10048_));
 BUFx3_ASAP7_75t_R _14056_ (.A(_10039_),
    .Y(_10049_));
 BUFx6f_ASAP7_75t_R _14057_ (.A(_10044_),
    .Y(_10050_));
 OR5x1_ASAP7_75t_R _14058_ (.A(_10047_),
    .B(_01865_),
    .C(_10048_),
    .D(_10049_),
    .E(_10050_),
    .Y(_10051_));
 OAI21x1_ASAP7_75t_R _14059_ (.A1(_10037_),
    .A2(_10046_),
    .B(_10051_),
    .Y(_02991_));
 BUFx3_ASAP7_75t_R _14060_ (.A(_10034_),
    .Y(_10052_));
 BUFx6f_ASAP7_75t_R _14061_ (.A(_09959_),
    .Y(_10053_));
 AND2x2_ASAP7_75t_R _14062_ (.A(_01115_),
    .B(_10053_),
    .Y(_10054_));
 BUFx3_ASAP7_75t_R _14063_ (.A(_10036_),
    .Y(_10055_));
 AO221x1_ASAP7_75t_R _14064_ (.A1(_01011_),
    .A2(_10052_),
    .B1(_10054_),
    .B2(_10055_),
    .C(_10012_),
    .Y(_10056_));
 OR5x1_ASAP7_75t_R _14065_ (.A(_10047_),
    .B(_01864_),
    .C(_10048_),
    .D(_10049_),
    .E(_10050_),
    .Y(_10057_));
 OAI21x1_ASAP7_75t_R _14066_ (.A1(_10046_),
    .A2(_10056_),
    .B(_10057_),
    .Y(_02992_));
 AND2x2_ASAP7_75t_R _14067_ (.A(_01114_),
    .B(_10053_),
    .Y(_10058_));
 AO221x1_ASAP7_75t_R _14068_ (.A1(_01010_),
    .A2(_10052_),
    .B1(_10058_),
    .B2(_10055_),
    .C(_10012_),
    .Y(_10059_));
 OR5x1_ASAP7_75t_R _14069_ (.A(_10047_),
    .B(_01863_),
    .C(_10048_),
    .D(_10049_),
    .E(_10050_),
    .Y(_10060_));
 OAI21x1_ASAP7_75t_R _14070_ (.A1(_10046_),
    .A2(_10059_),
    .B(_10060_),
    .Y(_02993_));
 AND2x2_ASAP7_75t_R _14071_ (.A(_01113_),
    .B(_10053_),
    .Y(_10061_));
 AO221x1_ASAP7_75t_R _14072_ (.A1(_01009_),
    .A2(_10052_),
    .B1(_10061_),
    .B2(_10055_),
    .C(_10012_),
    .Y(_10062_));
 OR5x1_ASAP7_75t_R _14073_ (.A(_10047_),
    .B(_01862_),
    .C(_10048_),
    .D(_10049_),
    .E(_10050_),
    .Y(_10063_));
 OAI21x1_ASAP7_75t_R _14074_ (.A1(_10046_),
    .A2(_10062_),
    .B(_10063_),
    .Y(_02994_));
 AND2x2_ASAP7_75t_R _14075_ (.A(_01112_),
    .B(_10053_),
    .Y(_10064_));
 AO221x1_ASAP7_75t_R _14076_ (.A1(_01008_),
    .A2(_10052_),
    .B1(_10064_),
    .B2(_10055_),
    .C(_10012_),
    .Y(_10065_));
 OR5x1_ASAP7_75t_R _14077_ (.A(_10047_),
    .B(_01861_),
    .C(_10048_),
    .D(_10049_),
    .E(_10050_),
    .Y(_10066_));
 OAI21x1_ASAP7_75t_R _14078_ (.A1(_10046_),
    .A2(_10065_),
    .B(_10066_),
    .Y(_02995_));
 INVx1_ASAP7_75t_R _14079_ (.A(_01111_),
    .Y(_10067_));
 NAND2x1_ASAP7_75t_R _14080_ (.A(_01007_),
    .B(_10034_),
    .Y(_10068_));
 OA21x2_ASAP7_75t_R _14081_ (.A1(_10067_),
    .A2(_10052_),
    .B(_10068_),
    .Y(_10069_));
 OA21x2_ASAP7_75t_R _14082_ (.A1(_10045_),
    .A2(_10069_),
    .B(_09872_),
    .Y(_02996_));
 AND2x2_ASAP7_75t_R _14083_ (.A(_01110_),
    .B(_10053_),
    .Y(_10070_));
 AO221x1_ASAP7_75t_R _14084_ (.A1(_01006_),
    .A2(_10052_),
    .B1(_10070_),
    .B2(_10055_),
    .C(_10012_),
    .Y(_10071_));
 OR5x1_ASAP7_75t_R _14085_ (.A(_10047_),
    .B(_01859_),
    .C(_10048_),
    .D(_10049_),
    .E(_10050_),
    .Y(_10072_));
 OAI21x1_ASAP7_75t_R _14086_ (.A1(_10046_),
    .A2(_10071_),
    .B(_10072_),
    .Y(_02997_));
 AND2x2_ASAP7_75t_R _14087_ (.A(_01109_),
    .B(_10053_),
    .Y(_10073_));
 AO221x1_ASAP7_75t_R _14088_ (.A1(_01005_),
    .A2(_10052_),
    .B1(_10073_),
    .B2(_10055_),
    .C(_08573_),
    .Y(_10074_));
 OR5x1_ASAP7_75t_R _14089_ (.A(_10047_),
    .B(_01858_),
    .C(_10048_),
    .D(_10049_),
    .E(_10050_),
    .Y(_10075_));
 OAI21x1_ASAP7_75t_R _14090_ (.A1(_10046_),
    .A2(_10074_),
    .B(_10075_),
    .Y(_02998_));
 AND2x2_ASAP7_75t_R _14091_ (.A(_01108_),
    .B(_10053_),
    .Y(_10076_));
 AO221x1_ASAP7_75t_R _14092_ (.A1(_01004_),
    .A2(_10052_),
    .B1(_10076_),
    .B2(_10055_),
    .C(_08573_),
    .Y(_10077_));
 OR5x1_ASAP7_75t_R _14093_ (.A(_10047_),
    .B(_01857_),
    .C(_10048_),
    .D(_10049_),
    .E(_10044_),
    .Y(_10078_));
 OAI21x1_ASAP7_75t_R _14094_ (.A1(_10046_),
    .A2(_10077_),
    .B(_10078_),
    .Y(_02999_));
 AND2x2_ASAP7_75t_R _14095_ (.A(_01107_),
    .B(_10053_),
    .Y(_10079_));
 AO221x1_ASAP7_75t_R _14096_ (.A1(_01003_),
    .A2(_10052_),
    .B1(_10079_),
    .B2(_10055_),
    .C(_08573_),
    .Y(_10080_));
 OR5x1_ASAP7_75t_R _14097_ (.A(_10047_),
    .B(_01856_),
    .C(_10048_),
    .D(_10049_),
    .E(_10044_),
    .Y(_10081_));
 OAI21x1_ASAP7_75t_R _14098_ (.A1(_10046_),
    .A2(_10080_),
    .B(_10081_),
    .Y(_03000_));
 OR3x1_ASAP7_75t_R _14099_ (.A(_08657_),
    .B(_09981_),
    .C(_10055_),
    .Y(_10082_));
 INVx1_ASAP7_75t_R _14100_ (.A(_10082_),
    .Y(_03001_));
 NOR2x1_ASAP7_75t_R _14101_ (.A(_10048_),
    .B(_10050_),
    .Y(_10083_));
 BUFx6f_ASAP7_75t_R _14102_ (.A(_08665_),
    .Y(_10084_));
 OA21x2_ASAP7_75t_R _14103_ (.A1(_10049_),
    .A2(_10083_),
    .B(_10084_),
    .Y(_03002_));
 AND2x2_ASAP7_75t_R _14104_ (.A(_01104_),
    .B(_10053_),
    .Y(_10085_));
 AO221x1_ASAP7_75t_R _14105_ (.A1(_01000_),
    .A2(_10052_),
    .B1(_10085_),
    .B2(_10055_),
    .C(_08573_),
    .Y(_10086_));
 OR5x1_ASAP7_75t_R _14106_ (.A(_08587_),
    .B(_01853_),
    .C(_09996_),
    .D(_10039_),
    .E(_10044_),
    .Y(_10087_));
 OAI21x1_ASAP7_75t_R _14107_ (.A1(_10046_),
    .A2(_10086_),
    .B(_10087_),
    .Y(_03003_));
 AND2x2_ASAP7_75t_R _14108_ (.A(_01103_),
    .B(_09959_),
    .Y(_10088_));
 AO221x1_ASAP7_75t_R _14109_ (.A1(_00999_),
    .A2(_10034_),
    .B1(_10088_),
    .B2(_10036_),
    .C(_08573_),
    .Y(_10089_));
 OR5x1_ASAP7_75t_R _14110_ (.A(_08587_),
    .B(_01852_),
    .C(_09996_),
    .D(_10039_),
    .E(_10044_),
    .Y(_10090_));
 OAI21x1_ASAP7_75t_R _14111_ (.A1(_10045_),
    .A2(_10089_),
    .B(_10090_),
    .Y(_03004_));
 AO21x2_ASAP7_75t_R _14112_ (.A1(_10040_),
    .A2(_10043_),
    .B(_09960_),
    .Y(_10091_));
 BUFx6f_ASAP7_75t_R _14113_ (.A(_10091_),
    .Y(_10092_));
 NOR2x1_ASAP7_75t_R _14114_ (.A(_01865_),
    .B(_10092_),
    .Y(_10093_));
 INVx1_ASAP7_75t_R _14115_ (.A(_01116_),
    .Y(_10094_));
 AO221x1_ASAP7_75t_R _14116_ (.A1(_09964_),
    .A2(_09970_),
    .B1(_09995_),
    .B2(_09997_),
    .C(_10001_),
    .Y(_10095_));
 AOI221x1_ASAP7_75t_R _14117_ (.A1(_09959_),
    .A2(_10031_),
    .B1(_10095_),
    .B2(_09965_),
    .C(_09995_),
    .Y(_10096_));
 BUFx6f_ASAP7_75t_R _14118_ (.A(_10096_),
    .Y(_10097_));
 BUFx6f_ASAP7_75t_R _14119_ (.A(_10096_),
    .Y(_10098_));
 NAND2x1_ASAP7_75t_R _14120_ (.A(_01012_),
    .B(_10098_),
    .Y(_10099_));
 BUFx6f_ASAP7_75t_R _14121_ (.A(_10091_),
    .Y(_10100_));
 OA211x2_ASAP7_75t_R _14122_ (.A1(_10094_),
    .A2(_10097_),
    .B(_10099_),
    .C(_10100_),
    .Y(_10101_));
 OA21x2_ASAP7_75t_R _14123_ (.A1(_10093_),
    .A2(_10101_),
    .B(_10084_),
    .Y(_03005_));
 NOR2x1_ASAP7_75t_R _14124_ (.A(_01864_),
    .B(_10092_),
    .Y(_10102_));
 INVx1_ASAP7_75t_R _14125_ (.A(_01115_),
    .Y(_10103_));
 NAND2x1_ASAP7_75t_R _14126_ (.A(_01011_),
    .B(_10098_),
    .Y(_10104_));
 OA211x2_ASAP7_75t_R _14127_ (.A1(_10103_),
    .A2(_10097_),
    .B(_10104_),
    .C(_10100_),
    .Y(_10105_));
 OA21x2_ASAP7_75t_R _14128_ (.A1(_10102_),
    .A2(_10105_),
    .B(_10084_),
    .Y(_03006_));
 NOR2x1_ASAP7_75t_R _14129_ (.A(_01863_),
    .B(_10092_),
    .Y(_10106_));
 INVx1_ASAP7_75t_R _14130_ (.A(_01114_),
    .Y(_10107_));
 NAND2x1_ASAP7_75t_R _14131_ (.A(_01010_),
    .B(_10098_),
    .Y(_10108_));
 OA211x2_ASAP7_75t_R _14132_ (.A1(_10107_),
    .A2(_10097_),
    .B(_10108_),
    .C(_10100_),
    .Y(_10109_));
 OA21x2_ASAP7_75t_R _14133_ (.A1(_10106_),
    .A2(_10109_),
    .B(_10084_),
    .Y(_03007_));
 NOR2x1_ASAP7_75t_R _14134_ (.A(_01862_),
    .B(_10092_),
    .Y(_10110_));
 INVx1_ASAP7_75t_R _14135_ (.A(_01113_),
    .Y(_10111_));
 NAND2x1_ASAP7_75t_R _14136_ (.A(_01009_),
    .B(_10098_),
    .Y(_10112_));
 OA211x2_ASAP7_75t_R _14137_ (.A1(_10111_),
    .A2(_10097_),
    .B(_10112_),
    .C(_10100_),
    .Y(_10113_));
 OA21x2_ASAP7_75t_R _14138_ (.A1(_10110_),
    .A2(_10113_),
    .B(_10084_),
    .Y(_03008_));
 NOR2x1_ASAP7_75t_R _14139_ (.A(_01861_),
    .B(_10092_),
    .Y(_10114_));
 INVx1_ASAP7_75t_R _14140_ (.A(_01112_),
    .Y(_10115_));
 NAND2x1_ASAP7_75t_R _14141_ (.A(_01008_),
    .B(_10098_),
    .Y(_10116_));
 OA211x2_ASAP7_75t_R _14142_ (.A1(_10115_),
    .A2(_10097_),
    .B(_10116_),
    .C(_10100_),
    .Y(_10117_));
 OA21x2_ASAP7_75t_R _14143_ (.A1(_10114_),
    .A2(_10117_),
    .B(_10084_),
    .Y(_03009_));
 AND2x2_ASAP7_75t_R _14144_ (.A(_09968_),
    .B(_10050_),
    .Y(_10118_));
 NAND2x1_ASAP7_75t_R _14145_ (.A(_01007_),
    .B(_10098_),
    .Y(_10119_));
 OA211x2_ASAP7_75t_R _14146_ (.A1(_10067_),
    .A2(_10097_),
    .B(_10119_),
    .C(_10100_),
    .Y(_10120_));
 OA21x2_ASAP7_75t_R _14147_ (.A1(_10118_),
    .A2(_10120_),
    .B(_10084_),
    .Y(_03010_));
 NOR2x1_ASAP7_75t_R _14148_ (.A(_01859_),
    .B(_10092_),
    .Y(_10121_));
 INVx1_ASAP7_75t_R _14149_ (.A(_01110_),
    .Y(_10122_));
 NAND2x1_ASAP7_75t_R _14150_ (.A(_01006_),
    .B(_10098_),
    .Y(_10123_));
 OA211x2_ASAP7_75t_R _14151_ (.A1(_10122_),
    .A2(_10097_),
    .B(_10123_),
    .C(_10100_),
    .Y(_10124_));
 OA21x2_ASAP7_75t_R _14152_ (.A1(_10121_),
    .A2(_10124_),
    .B(_10084_),
    .Y(_03011_));
 NOR2x1_ASAP7_75t_R _14153_ (.A(_01858_),
    .B(_10092_),
    .Y(_10125_));
 INVx1_ASAP7_75t_R _14154_ (.A(_01109_),
    .Y(_10126_));
 NAND2x1_ASAP7_75t_R _14155_ (.A(_01005_),
    .B(_10098_),
    .Y(_10127_));
 OA211x2_ASAP7_75t_R _14156_ (.A1(_10126_),
    .A2(_10097_),
    .B(_10127_),
    .C(_10100_),
    .Y(_10128_));
 OA21x2_ASAP7_75t_R _14157_ (.A1(_10125_),
    .A2(_10128_),
    .B(_10084_),
    .Y(_03012_));
 NOR2x1_ASAP7_75t_R _14158_ (.A(_01857_),
    .B(_10092_),
    .Y(_10129_));
 NAND2x1_ASAP7_75t_R _14159_ (.A(_01004_),
    .B(_10096_),
    .Y(_10130_));
 OA211x2_ASAP7_75t_R _14160_ (.A1(_09982_),
    .A2(_10097_),
    .B(_10130_),
    .C(_10100_),
    .Y(_10131_));
 OA21x2_ASAP7_75t_R _14161_ (.A1(_10129_),
    .A2(_10131_),
    .B(_10084_),
    .Y(_03013_));
 NOR2x1_ASAP7_75t_R _14162_ (.A(_01856_),
    .B(_10092_),
    .Y(_10132_));
 NAND2x1_ASAP7_75t_R _14163_ (.A(_01003_),
    .B(_10096_),
    .Y(_10133_));
 OA211x2_ASAP7_75t_R _14164_ (.A1(_09962_),
    .A2(_10097_),
    .B(_10133_),
    .C(_10091_),
    .Y(_10134_));
 BUFx6f_ASAP7_75t_R _14165_ (.A(_08665_),
    .Y(_10135_));
 OA21x2_ASAP7_75t_R _14166_ (.A1(_10132_),
    .A2(_10134_),
    .B(_10135_),
    .Y(_03014_));
 NAND3x1_ASAP7_75t_R _14167_ (.A(_09980_),
    .B(_09990_),
    .C(_10043_),
    .Y(_10136_));
 AND4x1_ASAP7_75t_R _14168_ (.A(_08999_),
    .B(_09961_),
    .C(_09966_),
    .D(_10136_),
    .Y(_03015_));
 AOI21x1_ASAP7_75t_R _14169_ (.A1(_10053_),
    .A2(_10031_),
    .B(_09995_),
    .Y(_10137_));
 AO21x1_ASAP7_75t_R _14170_ (.A1(_09965_),
    .A2(_10095_),
    .B(_10137_),
    .Y(_10138_));
 OA21x2_ASAP7_75t_R _14171_ (.A1(_10050_),
    .A2(_10138_),
    .B(_10135_),
    .Y(_03016_));
 NOR2x1_ASAP7_75t_R _14172_ (.A(_01853_),
    .B(_10092_),
    .Y(_10139_));
 INVx1_ASAP7_75t_R _14173_ (.A(_01104_),
    .Y(_10140_));
 NAND2x1_ASAP7_75t_R _14174_ (.A(_01000_),
    .B(_10096_),
    .Y(_10141_));
 OA211x2_ASAP7_75t_R _14175_ (.A1(_10140_),
    .A2(_10098_),
    .B(_10141_),
    .C(_10091_),
    .Y(_10142_));
 OA21x2_ASAP7_75t_R _14176_ (.A1(_10139_),
    .A2(_10142_),
    .B(_10135_),
    .Y(_03017_));
 NOR2x1_ASAP7_75t_R _14177_ (.A(_01852_),
    .B(_10100_),
    .Y(_10143_));
 INVx1_ASAP7_75t_R _14178_ (.A(_01103_),
    .Y(_10144_));
 NAND2x1_ASAP7_75t_R _14179_ (.A(_00999_),
    .B(_10096_),
    .Y(_10145_));
 OA211x2_ASAP7_75t_R _14180_ (.A1(_10144_),
    .A2(_10098_),
    .B(_10145_),
    .C(_10091_),
    .Y(_10146_));
 OA21x2_ASAP7_75t_R _14181_ (.A1(_10143_),
    .A2(_10146_),
    .B(_10135_),
    .Y(_03018_));
 AND2x2_ASAP7_75t_R _14182_ (.A(_09957_),
    .B(_00008_),
    .Y(_03019_));
 OR2x6_ASAP7_75t_R _14183_ (.A(_02260_),
    .B(_02261_),
    .Y(_10147_));
 BUFx6f_ASAP7_75t_R _14184_ (.A(_10147_),
    .Y(_10148_));
 BUFx6f_ASAP7_75t_R _14185_ (.A(_02302_),
    .Y(_10149_));
 NOR2x2_ASAP7_75t_R _14186_ (.A(_10149_),
    .B(_02303_),
    .Y(_10150_));
 AND3x4_ASAP7_75t_R _14187_ (.A(_02304_),
    .B(_02305_),
    .C(_02306_),
    .Y(_10151_));
 NOR2x2_ASAP7_75t_R _14188_ (.A(_10149_),
    .B(_10151_),
    .Y(_10152_));
 INVx1_ASAP7_75t_R _14189_ (.A(_01827_),
    .Y(_10153_));
 BUFx6f_ASAP7_75t_R _14190_ (.A(_01831_),
    .Y(_10154_));
 INVx2_ASAP7_75t_R _14191_ (.A(_01826_),
    .Y(_10155_));
 OA211x2_ASAP7_75t_R _14192_ (.A1(_10153_),
    .A2(_10154_),
    .B(_10147_),
    .C(_10155_),
    .Y(_10156_));
 INVx2_ASAP7_75t_R _14193_ (.A(_02260_),
    .Y(_10157_));
 AND3x4_ASAP7_75t_R _14194_ (.A(_02262_),
    .B(_02263_),
    .C(_02264_),
    .Y(_10158_));
 NAND3x1_ASAP7_75t_R _14195_ (.A(_10157_),
    .B(_02265_),
    .C(_10158_),
    .Y(_10159_));
 AO221x1_ASAP7_75t_R _14196_ (.A1(_10148_),
    .A2(_10150_),
    .B1(_10152_),
    .B2(_10156_),
    .C(_10159_),
    .Y(_10160_));
 AND2x4_ASAP7_75t_R _14197_ (.A(_10155_),
    .B(_01827_),
    .Y(_10161_));
 OR2x2_ASAP7_75t_R _14198_ (.A(_10149_),
    .B(_10151_),
    .Y(_10162_));
 AND3x4_ASAP7_75t_R _14199_ (.A(_10157_),
    .B(_02265_),
    .C(_10158_),
    .Y(_10163_));
 NOR2x1_ASAP7_75t_R _14200_ (.A(_02260_),
    .B(_02261_),
    .Y(_10164_));
 AO31x2_ASAP7_75t_R _14201_ (.A1(_10157_),
    .A2(_02265_),
    .A3(_10158_),
    .B(_10164_),
    .Y(_10165_));
 INVx1_ASAP7_75t_R _14202_ (.A(_10149_),
    .Y(_10166_));
 INVx1_ASAP7_75t_R _14203_ (.A(_02307_),
    .Y(_10167_));
 AND3x4_ASAP7_75t_R _14204_ (.A(_10166_),
    .B(_10167_),
    .C(_10151_),
    .Y(_10168_));
 OR2x2_ASAP7_75t_R _14205_ (.A(_10149_),
    .B(_02303_),
    .Y(_10169_));
 NAND2x1_ASAP7_75t_R _14206_ (.A(_10154_),
    .B(_10169_),
    .Y(_10170_));
 AOI221x1_ASAP7_75t_R _14207_ (.A1(_10162_),
    .A2(_10163_),
    .B1(_10165_),
    .B2(_10168_),
    .C(_10170_),
    .Y(_10171_));
 AND2x4_ASAP7_75t_R _14208_ (.A(_10161_),
    .B(_10171_),
    .Y(_10172_));
 NAND2x1_ASAP7_75t_R _14209_ (.A(_10160_),
    .B(_10172_),
    .Y(_10173_));
 BUFx6f_ASAP7_75t_R _14210_ (.A(_10173_),
    .Y(_10174_));
 OR2x2_ASAP7_75t_R _14211_ (.A(_01837_),
    .B(_10174_),
    .Y(_10175_));
 AO31x2_ASAP7_75t_R _14212_ (.A1(_02262_),
    .A2(_02263_),
    .A3(_02264_),
    .B(_02260_),
    .Y(_10176_));
 OR2x2_ASAP7_75t_R _14213_ (.A(_01826_),
    .B(_01827_),
    .Y(_10177_));
 OA31x2_ASAP7_75t_R _14214_ (.A1(_10155_),
    .A2(_00008_),
    .A3(_10176_),
    .B1(_10177_),
    .Y(_10178_));
 OR3x1_ASAP7_75t_R _14215_ (.A(_01826_),
    .B(_10154_),
    .C(_02260_),
    .Y(_10179_));
 AO21x1_ASAP7_75t_R _14216_ (.A1(_02261_),
    .A2(_10158_),
    .B(_10179_),
    .Y(_10180_));
 AO21x2_ASAP7_75t_R _14217_ (.A1(_10178_),
    .A2(_10180_),
    .B(_10162_),
    .Y(_10181_));
 AO21x1_ASAP7_75t_R _14218_ (.A1(_01827_),
    .A2(_10154_),
    .B(_01826_),
    .Y(_10182_));
 OA21x2_ASAP7_75t_R _14219_ (.A1(_10176_),
    .A2(_10182_),
    .B(_10147_),
    .Y(_10183_));
 INVx1_ASAP7_75t_R _14220_ (.A(_02304_),
    .Y(_10184_));
 INVx1_ASAP7_75t_R _14221_ (.A(_02305_),
    .Y(_10185_));
 INVx1_ASAP7_75t_R _14222_ (.A(_02306_),
    .Y(_10186_));
 OR5x1_ASAP7_75t_R _14223_ (.A(_10149_),
    .B(_10184_),
    .C(_10185_),
    .D(_10186_),
    .E(_02307_),
    .Y(_10187_));
 OA21x2_ASAP7_75t_R _14224_ (.A1(_10183_),
    .A2(_10187_),
    .B(_10169_),
    .Y(_10188_));
 NAND2x1_ASAP7_75t_R _14225_ (.A(_10181_),
    .B(_10188_),
    .Y(_10189_));
 OR2x2_ASAP7_75t_R _14226_ (.A(_10189_),
    .B(_10160_),
    .Y(_10190_));
 BUFx3_ASAP7_75t_R _14227_ (.A(_10190_),
    .Y(_10191_));
 AOI221x1_ASAP7_75t_R _14228_ (.A1(_10148_),
    .A2(_10150_),
    .B1(_10152_),
    .B2(_10156_),
    .C(_10159_),
    .Y(_10192_));
 AND3x1_ASAP7_75t_R _14229_ (.A(_10181_),
    .B(_10188_),
    .C(_10192_),
    .Y(_10193_));
 BUFx6f_ASAP7_75t_R _14230_ (.A(_10193_),
    .Y(_10194_));
 AND3x1_ASAP7_75t_R _14231_ (.A(_10161_),
    .B(_10160_),
    .C(_10171_),
    .Y(_10195_));
 BUFx6f_ASAP7_75t_R _14232_ (.A(_10195_),
    .Y(_10196_));
 AO21x1_ASAP7_75t_R _14233_ (.A1(_02271_),
    .A2(_10194_),
    .B(_10196_),
    .Y(_10197_));
 AO21x1_ASAP7_75t_R _14234_ (.A1(_02313_),
    .A2(_10191_),
    .B(_10197_),
    .Y(_10198_));
 BUFx12f_ASAP7_75t_R _14235_ (.A(_09118_),
    .Y(_10199_));
 AOI21x1_ASAP7_75t_R _14236_ (.A1(_10175_),
    .A2(_10198_),
    .B(_10199_),
    .Y(_03020_));
 OR2x2_ASAP7_75t_R _14237_ (.A(_01836_),
    .B(_10174_),
    .Y(_10200_));
 AO21x1_ASAP7_75t_R _14238_ (.A1(_02270_),
    .A2(_10194_),
    .B(_10196_),
    .Y(_10201_));
 AO21x1_ASAP7_75t_R _14239_ (.A1(_02312_),
    .A2(_10191_),
    .B(_10201_),
    .Y(_10202_));
 AOI21x1_ASAP7_75t_R _14240_ (.A1(_10200_),
    .A2(_10202_),
    .B(_10199_),
    .Y(_03021_));
 OR2x2_ASAP7_75t_R _14241_ (.A(_01835_),
    .B(_10174_),
    .Y(_10203_));
 AO21x1_ASAP7_75t_R _14242_ (.A1(_02269_),
    .A2(_10194_),
    .B(_10196_),
    .Y(_10204_));
 AO21x1_ASAP7_75t_R _14243_ (.A1(_02311_),
    .A2(_10191_),
    .B(_10204_),
    .Y(_10205_));
 AOI21x1_ASAP7_75t_R _14244_ (.A1(_10203_),
    .A2(_10205_),
    .B(_10199_),
    .Y(_03022_));
 OR2x2_ASAP7_75t_R _14245_ (.A(_01834_),
    .B(_10174_),
    .Y(_10206_));
 AO21x1_ASAP7_75t_R _14246_ (.A1(_02268_),
    .A2(_10194_),
    .B(_10196_),
    .Y(_10207_));
 AO21x1_ASAP7_75t_R _14247_ (.A1(_02310_),
    .A2(_10191_),
    .B(_10207_),
    .Y(_10208_));
 AOI21x1_ASAP7_75t_R _14248_ (.A1(_10206_),
    .A2(_10208_),
    .B(_10199_),
    .Y(_03023_));
 OR2x2_ASAP7_75t_R _14249_ (.A(_01833_),
    .B(_10174_),
    .Y(_10209_));
 AO21x1_ASAP7_75t_R _14250_ (.A1(_02267_),
    .A2(_10194_),
    .B(_10196_),
    .Y(_10210_));
 AO21x1_ASAP7_75t_R _14251_ (.A1(_02309_),
    .A2(_10191_),
    .B(_10210_),
    .Y(_10211_));
 AOI21x1_ASAP7_75t_R _14252_ (.A1(_10209_),
    .A2(_10211_),
    .B(_10199_),
    .Y(_03024_));
 OR2x2_ASAP7_75t_R _14253_ (.A(_01832_),
    .B(_10174_),
    .Y(_10212_));
 AO21x1_ASAP7_75t_R _14254_ (.A1(_02266_),
    .A2(_10194_),
    .B(_10196_),
    .Y(_10213_));
 AO21x1_ASAP7_75t_R _14255_ (.A1(_02308_),
    .A2(_10191_),
    .B(_10213_),
    .Y(_10214_));
 AOI21x1_ASAP7_75t_R _14256_ (.A1(_10212_),
    .A2(_10214_),
    .B(_10199_),
    .Y(_03025_));
 OR2x6_ASAP7_75t_R _14257_ (.A(_10194_),
    .B(_10196_),
    .Y(_10215_));
 OR3x1_ASAP7_75t_R _14258_ (.A(_08657_),
    .B(_02307_),
    .C(_10215_),
    .Y(_10216_));
 INVx1_ASAP7_75t_R _14259_ (.A(_10216_),
    .Y(_03026_));
 OAI22x1_ASAP7_75t_R _14260_ (.A1(_01830_),
    .A2(_10174_),
    .B1(_10215_),
    .B2(_02306_),
    .Y(_10217_));
 AND2x2_ASAP7_75t_R _14261_ (.A(_09957_),
    .B(_10217_),
    .Y(_03027_));
 OAI22x1_ASAP7_75t_R _14262_ (.A1(_01829_),
    .A2(_10174_),
    .B1(_10215_),
    .B2(_02305_),
    .Y(_10218_));
 AND2x2_ASAP7_75t_R _14263_ (.A(_09957_),
    .B(_10218_),
    .Y(_03028_));
 OAI22x1_ASAP7_75t_R _14264_ (.A1(_01828_),
    .A2(_10174_),
    .B1(_10215_),
    .B2(_02304_),
    .Y(_10219_));
 AND2x2_ASAP7_75t_R _14265_ (.A(_09957_),
    .B(_10219_),
    .Y(_03029_));
 OA21x2_ASAP7_75t_R _14266_ (.A1(_10183_),
    .A2(_10187_),
    .B(_10181_),
    .Y(_10220_));
 OR3x1_ASAP7_75t_R _14267_ (.A(_08642_),
    .B(_10150_),
    .C(_10220_),
    .Y(_10221_));
 INVx1_ASAP7_75t_R _14268_ (.A(_10221_),
    .Y(_03030_));
 OA31x2_ASAP7_75t_R _14269_ (.A1(_10189_),
    .A2(_10192_),
    .A3(_10172_),
    .B1(_08877_),
    .Y(_03031_));
 OR2x2_ASAP7_75t_R _14270_ (.A(_01825_),
    .B(_10174_),
    .Y(_10222_));
 AO21x1_ASAP7_75t_R _14271_ (.A1(_02259_),
    .A2(_10194_),
    .B(_10196_),
    .Y(_10223_));
 AO21x1_ASAP7_75t_R _14272_ (.A1(_02301_),
    .A2(_10191_),
    .B(_10223_),
    .Y(_10224_));
 AOI21x1_ASAP7_75t_R _14273_ (.A1(_10222_),
    .A2(_10224_),
    .B(_10199_),
    .Y(_03032_));
 OR2x2_ASAP7_75t_R _14274_ (.A(_01824_),
    .B(_10173_),
    .Y(_10225_));
 AO21x1_ASAP7_75t_R _14275_ (.A1(_02258_),
    .A2(_10194_),
    .B(_10196_),
    .Y(_10226_));
 AO21x1_ASAP7_75t_R _14276_ (.A1(_02300_),
    .A2(_10191_),
    .B(_10226_),
    .Y(_10227_));
 AOI21x1_ASAP7_75t_R _14277_ (.A1(_10225_),
    .A2(_10227_),
    .B(_10199_),
    .Y(_03033_));
 AOI22x1_ASAP7_75t_R _14278_ (.A1(_10176_),
    .A2(_10168_),
    .B1(_10163_),
    .B2(_10150_),
    .Y(_10228_));
 INVx2_ASAP7_75t_R _14279_ (.A(_10154_),
    .Y(_10229_));
 AND2x2_ASAP7_75t_R _14280_ (.A(_10229_),
    .B(_10148_),
    .Y(_10230_));
 AO21x2_ASAP7_75t_R _14281_ (.A1(_10228_),
    .A2(_10230_),
    .B(_10171_),
    .Y(_10231_));
 OAI21x1_ASAP7_75t_R _14282_ (.A1(_10183_),
    .A2(_10150_),
    .B(_10168_),
    .Y(_10232_));
 AND3x1_ASAP7_75t_R _14283_ (.A(_10229_),
    .B(_10161_),
    .C(_10232_),
    .Y(_10233_));
 NAND2x1_ASAP7_75t_R _14284_ (.A(_10231_),
    .B(_10233_),
    .Y(_10234_));
 BUFx6f_ASAP7_75t_R _14285_ (.A(_10234_),
    .Y(_10235_));
 OR2x2_ASAP7_75t_R _14286_ (.A(_01837_),
    .B(_10235_),
    .Y(_10236_));
 OA21x2_ASAP7_75t_R _14287_ (.A1(_10153_),
    .A2(_10154_),
    .B(_10155_),
    .Y(_10237_));
 AO21x1_ASAP7_75t_R _14288_ (.A1(_10152_),
    .A2(_10237_),
    .B(_10150_),
    .Y(_10238_));
 AO221x1_ASAP7_75t_R _14289_ (.A1(_10155_),
    .A2(_10229_),
    .B1(_02303_),
    .B2(_10151_),
    .C(_10149_),
    .Y(_10239_));
 INVx1_ASAP7_75t_R _14290_ (.A(_00008_),
    .Y(_10240_));
 OR3x1_ASAP7_75t_R _14291_ (.A(_10240_),
    .B(_10149_),
    .C(_10151_),
    .Y(_10241_));
 AOI22x1_ASAP7_75t_R _14292_ (.A1(_01827_),
    .A2(_10239_),
    .B1(_10241_),
    .B2(_01826_),
    .Y(_10242_));
 NOR2x1_ASAP7_75t_R _14293_ (.A(_02260_),
    .B(_10158_),
    .Y(_10243_));
 AOI22x1_ASAP7_75t_R _14294_ (.A1(_10163_),
    .A2(_10238_),
    .B1(_10242_),
    .B2(_10243_),
    .Y(_10244_));
 NAND2x1_ASAP7_75t_R _14295_ (.A(_10148_),
    .B(_10244_),
    .Y(_10245_));
 BUFx3_ASAP7_75t_R _14296_ (.A(_10245_),
    .Y(_10246_));
 BUFx6f_ASAP7_75t_R _14297_ (.A(_10148_),
    .Y(_10247_));
 AND2x2_ASAP7_75t_R _14298_ (.A(_02313_),
    .B(_10247_),
    .Y(_10248_));
 BUFx6f_ASAP7_75t_R _14299_ (.A(_10244_),
    .Y(_10249_));
 AND2x2_ASAP7_75t_R _14300_ (.A(_10231_),
    .B(_10233_),
    .Y(_10250_));
 BUFx6f_ASAP7_75t_R _14301_ (.A(_10250_),
    .Y(_10251_));
 AO221x1_ASAP7_75t_R _14302_ (.A1(_02271_),
    .A2(_10246_),
    .B1(_10248_),
    .B2(_10249_),
    .C(_10251_),
    .Y(_10252_));
 AOI21x1_ASAP7_75t_R _14303_ (.A1(_10236_),
    .A2(_10252_),
    .B(_10199_),
    .Y(_03034_));
 OR2x2_ASAP7_75t_R _14304_ (.A(_01836_),
    .B(_10235_),
    .Y(_10253_));
 AND2x2_ASAP7_75t_R _14305_ (.A(_02312_),
    .B(_10247_),
    .Y(_10254_));
 AO221x1_ASAP7_75t_R _14306_ (.A1(_02270_),
    .A2(_10246_),
    .B1(_10254_),
    .B2(_10249_),
    .C(_10251_),
    .Y(_10255_));
 AOI21x1_ASAP7_75t_R _14307_ (.A1(_10253_),
    .A2(_10255_),
    .B(_10199_),
    .Y(_03035_));
 OR2x2_ASAP7_75t_R _14308_ (.A(_01835_),
    .B(_10235_),
    .Y(_10256_));
 AND2x2_ASAP7_75t_R _14309_ (.A(_02311_),
    .B(_10247_),
    .Y(_10257_));
 AO221x1_ASAP7_75t_R _14310_ (.A1(_02269_),
    .A2(_10246_),
    .B1(_10257_),
    .B2(_10249_),
    .C(_10251_),
    .Y(_10258_));
 BUFx12f_ASAP7_75t_R _14311_ (.A(_09118_),
    .Y(_10259_));
 AOI21x1_ASAP7_75t_R _14312_ (.A1(_10256_),
    .A2(_10258_),
    .B(_10259_),
    .Y(_03036_));
 OR2x2_ASAP7_75t_R _14313_ (.A(_01834_),
    .B(_10235_),
    .Y(_10260_));
 AND2x2_ASAP7_75t_R _14314_ (.A(_02310_),
    .B(_10247_),
    .Y(_10261_));
 AO221x1_ASAP7_75t_R _14315_ (.A1(_02268_),
    .A2(_10246_),
    .B1(_10261_),
    .B2(_10249_),
    .C(_10251_),
    .Y(_10262_));
 AOI21x1_ASAP7_75t_R _14316_ (.A1(_10260_),
    .A2(_10262_),
    .B(_10259_),
    .Y(_03037_));
 OR2x2_ASAP7_75t_R _14317_ (.A(_01833_),
    .B(_10235_),
    .Y(_10263_));
 AND2x2_ASAP7_75t_R _14318_ (.A(_02309_),
    .B(_10247_),
    .Y(_10264_));
 AO221x1_ASAP7_75t_R _14319_ (.A1(_02267_),
    .A2(_10246_),
    .B1(_10264_),
    .B2(_10249_),
    .C(_10251_),
    .Y(_10265_));
 AOI21x1_ASAP7_75t_R _14320_ (.A1(_10263_),
    .A2(_10265_),
    .B(_10259_),
    .Y(_03038_));
 OR2x2_ASAP7_75t_R _14321_ (.A(_01832_),
    .B(_10235_),
    .Y(_10266_));
 AND2x2_ASAP7_75t_R _14322_ (.A(_02308_),
    .B(_10247_),
    .Y(_10267_));
 AO221x1_ASAP7_75t_R _14323_ (.A1(_02266_),
    .A2(_10246_),
    .B1(_10267_),
    .B2(_10249_),
    .C(_10251_),
    .Y(_10268_));
 AOI21x1_ASAP7_75t_R _14324_ (.A1(_10266_),
    .A2(_10268_),
    .B(_10259_),
    .Y(_03039_));
 AND3x1_ASAP7_75t_R _14325_ (.A(_02307_),
    .B(_10247_),
    .C(_10244_),
    .Y(_10269_));
 AO21x1_ASAP7_75t_R _14326_ (.A1(_02265_),
    .A2(_10246_),
    .B(_10269_),
    .Y(_10270_));
 AOI21x1_ASAP7_75t_R _14327_ (.A1(_10235_),
    .A2(_10270_),
    .B(_10259_),
    .Y(_03040_));
 OR2x2_ASAP7_75t_R _14328_ (.A(_01830_),
    .B(_10235_),
    .Y(_10271_));
 AND2x2_ASAP7_75t_R _14329_ (.A(_02306_),
    .B(_10247_),
    .Y(_10272_));
 AO221x1_ASAP7_75t_R _14330_ (.A1(_02264_),
    .A2(_10246_),
    .B1(_10272_),
    .B2(_10249_),
    .C(_10251_),
    .Y(_10273_));
 AOI21x1_ASAP7_75t_R _14331_ (.A1(_10271_),
    .A2(_10273_),
    .B(_10259_),
    .Y(_03041_));
 OR2x2_ASAP7_75t_R _14332_ (.A(_01829_),
    .B(_10235_),
    .Y(_10274_));
 AND2x2_ASAP7_75t_R _14333_ (.A(_02305_),
    .B(_10148_),
    .Y(_10275_));
 AO221x1_ASAP7_75t_R _14334_ (.A1(_02263_),
    .A2(_10246_),
    .B1(_10275_),
    .B2(_10249_),
    .C(_10251_),
    .Y(_10276_));
 AOI21x1_ASAP7_75t_R _14335_ (.A1(_10274_),
    .A2(_10276_),
    .B(_10259_),
    .Y(_03042_));
 OR2x2_ASAP7_75t_R _14336_ (.A(_01828_),
    .B(_10235_),
    .Y(_10277_));
 AND2x2_ASAP7_75t_R _14337_ (.A(_02304_),
    .B(_10148_),
    .Y(_10278_));
 AO221x1_ASAP7_75t_R _14338_ (.A1(_02262_),
    .A2(_10246_),
    .B1(_10278_),
    .B2(_10244_),
    .C(_10251_),
    .Y(_10279_));
 AOI21x1_ASAP7_75t_R _14339_ (.A1(_10277_),
    .A2(_10279_),
    .B(_10259_),
    .Y(_03043_));
 OR3x1_ASAP7_75t_R _14340_ (.A(_08642_),
    .B(_10164_),
    .C(_10249_),
    .Y(_10280_));
 INVx1_ASAP7_75t_R _14341_ (.A(_10280_),
    .Y(_03044_));
 AND3x1_ASAP7_75t_R _14342_ (.A(_10247_),
    .B(_10232_),
    .C(_10249_),
    .Y(_10281_));
 NAND3x1_ASAP7_75t_R _14343_ (.A(_10229_),
    .B(_10161_),
    .C(_10231_),
    .Y(_10282_));
 AOI21x1_ASAP7_75t_R _14344_ (.A1(_10281_),
    .A2(_10282_),
    .B(_10259_),
    .Y(_03045_));
 OR2x2_ASAP7_75t_R _14345_ (.A(_01825_),
    .B(_10234_),
    .Y(_10283_));
 AND2x2_ASAP7_75t_R _14346_ (.A(_02301_),
    .B(_10148_),
    .Y(_10284_));
 AO221x1_ASAP7_75t_R _14347_ (.A1(_02259_),
    .A2(_10245_),
    .B1(_10284_),
    .B2(_10244_),
    .C(_10251_),
    .Y(_10285_));
 AOI21x1_ASAP7_75t_R _14348_ (.A1(_10283_),
    .A2(_10285_),
    .B(_10259_),
    .Y(_03046_));
 OR2x2_ASAP7_75t_R _14349_ (.A(_01824_),
    .B(_10234_),
    .Y(_10286_));
 AND2x2_ASAP7_75t_R _14350_ (.A(_02300_),
    .B(_10148_),
    .Y(_10287_));
 AO221x1_ASAP7_75t_R _14351_ (.A1(_02258_),
    .A2(_10245_),
    .B1(_10287_),
    .B2(_10244_),
    .C(_10250_),
    .Y(_10288_));
 BUFx12f_ASAP7_75t_R _14352_ (.A(_09118_),
    .Y(_10289_));
 AOI21x1_ASAP7_75t_R _14353_ (.A1(_10286_),
    .A2(_10288_),
    .B(_10289_),
    .Y(_03047_));
 AO21x2_ASAP7_75t_R _14354_ (.A1(_01827_),
    .A2(_10231_),
    .B(_01826_),
    .Y(_10290_));
 BUFx6f_ASAP7_75t_R _14355_ (.A(_10290_),
    .Y(_10291_));
 NOR2x1_ASAP7_75t_R _14356_ (.A(_01837_),
    .B(_10291_),
    .Y(_10292_));
 INVx1_ASAP7_75t_R _14357_ (.A(_02313_),
    .Y(_10293_));
 INVx1_ASAP7_75t_R _14358_ (.A(_02303_),
    .Y(_10294_));
 AO21x1_ASAP7_75t_R _14359_ (.A1(_10178_),
    .A2(_10180_),
    .B(_10294_),
    .Y(_10295_));
 AOI221x1_ASAP7_75t_R _14360_ (.A1(_10148_),
    .A2(_10242_),
    .B1(_10295_),
    .B2(_10152_),
    .C(_10176_),
    .Y(_10296_));
 BUFx6f_ASAP7_75t_R _14361_ (.A(_10296_),
    .Y(_10297_));
 BUFx6f_ASAP7_75t_R _14362_ (.A(_10296_),
    .Y(_10298_));
 NAND2x1_ASAP7_75t_R _14363_ (.A(_02271_),
    .B(_10298_),
    .Y(_10299_));
 BUFx6f_ASAP7_75t_R _14364_ (.A(_10290_),
    .Y(_10300_));
 OA211x2_ASAP7_75t_R _14365_ (.A1(_10293_),
    .A2(_10297_),
    .B(_10299_),
    .C(_10300_),
    .Y(_10301_));
 OA21x2_ASAP7_75t_R _14366_ (.A1(_10292_),
    .A2(_10301_),
    .B(_10135_),
    .Y(_03048_));
 NOR2x1_ASAP7_75t_R _14367_ (.A(_01836_),
    .B(_10291_),
    .Y(_10302_));
 INVx1_ASAP7_75t_R _14368_ (.A(_02312_),
    .Y(_10303_));
 NAND2x1_ASAP7_75t_R _14369_ (.A(_02270_),
    .B(_10298_),
    .Y(_10304_));
 OA211x2_ASAP7_75t_R _14370_ (.A1(_10303_),
    .A2(_10297_),
    .B(_10304_),
    .C(_10300_),
    .Y(_10305_));
 OA21x2_ASAP7_75t_R _14371_ (.A1(_10302_),
    .A2(_10305_),
    .B(_10135_),
    .Y(_03049_));
 NOR2x1_ASAP7_75t_R _14372_ (.A(_01835_),
    .B(_10291_),
    .Y(_10306_));
 INVx1_ASAP7_75t_R _14373_ (.A(_02311_),
    .Y(_10307_));
 NAND2x1_ASAP7_75t_R _14374_ (.A(_02269_),
    .B(_10298_),
    .Y(_10308_));
 OA211x2_ASAP7_75t_R _14375_ (.A1(_10307_),
    .A2(_10297_),
    .B(_10308_),
    .C(_10300_),
    .Y(_10309_));
 OA21x2_ASAP7_75t_R _14376_ (.A1(_10306_),
    .A2(_10309_),
    .B(_10135_),
    .Y(_03050_));
 NOR2x1_ASAP7_75t_R _14377_ (.A(_01834_),
    .B(_10291_),
    .Y(_10310_));
 INVx1_ASAP7_75t_R _14378_ (.A(_02310_),
    .Y(_10311_));
 NAND2x1_ASAP7_75t_R _14379_ (.A(_02268_),
    .B(_10298_),
    .Y(_10312_));
 OA211x2_ASAP7_75t_R _14380_ (.A1(_10311_),
    .A2(_10297_),
    .B(_10312_),
    .C(_10300_),
    .Y(_10313_));
 OA21x2_ASAP7_75t_R _14381_ (.A1(_10310_),
    .A2(_10313_),
    .B(_10135_),
    .Y(_03051_));
 NOR2x1_ASAP7_75t_R _14382_ (.A(_01833_),
    .B(_10291_),
    .Y(_10314_));
 INVx1_ASAP7_75t_R _14383_ (.A(_02309_),
    .Y(_10315_));
 NAND2x1_ASAP7_75t_R _14384_ (.A(_02267_),
    .B(_10298_),
    .Y(_10316_));
 OA211x2_ASAP7_75t_R _14385_ (.A1(_10315_),
    .A2(_10297_),
    .B(_10316_),
    .C(_10300_),
    .Y(_10317_));
 OA21x2_ASAP7_75t_R _14386_ (.A1(_10314_),
    .A2(_10317_),
    .B(_10135_),
    .Y(_03052_));
 NOR2x1_ASAP7_75t_R _14387_ (.A(_01832_),
    .B(_10291_),
    .Y(_10318_));
 INVx1_ASAP7_75t_R _14388_ (.A(_02308_),
    .Y(_10319_));
 NAND2x1_ASAP7_75t_R _14389_ (.A(_02266_),
    .B(_10298_),
    .Y(_10320_));
 OA211x2_ASAP7_75t_R _14390_ (.A1(_10319_),
    .A2(_10297_),
    .B(_10320_),
    .C(_10300_),
    .Y(_10321_));
 OA21x2_ASAP7_75t_R _14391_ (.A1(_10318_),
    .A2(_10321_),
    .B(_10135_),
    .Y(_03053_));
 NOR2x1_ASAP7_75t_R _14392_ (.A(_10154_),
    .B(_10291_),
    .Y(_10322_));
 NAND2x1_ASAP7_75t_R _14393_ (.A(_02265_),
    .B(_10298_),
    .Y(_10323_));
 OA211x2_ASAP7_75t_R _14394_ (.A1(_10167_),
    .A2(_10297_),
    .B(_10323_),
    .C(_10300_),
    .Y(_10324_));
 BUFx6f_ASAP7_75t_R _14395_ (.A(_08665_),
    .Y(_10325_));
 OA21x2_ASAP7_75t_R _14396_ (.A1(_10322_),
    .A2(_10324_),
    .B(_10325_),
    .Y(_03054_));
 NOR2x1_ASAP7_75t_R _14397_ (.A(_01830_),
    .B(_10291_),
    .Y(_10326_));
 NAND2x1_ASAP7_75t_R _14398_ (.A(_02264_),
    .B(_10298_),
    .Y(_10327_));
 OA211x2_ASAP7_75t_R _14399_ (.A1(_10186_),
    .A2(_10297_),
    .B(_10327_),
    .C(_10290_),
    .Y(_10328_));
 OA21x2_ASAP7_75t_R _14400_ (.A1(_10326_),
    .A2(_10328_),
    .B(_10325_),
    .Y(_03055_));
 NOR2x1_ASAP7_75t_R _14401_ (.A(_01829_),
    .B(_10291_),
    .Y(_10329_));
 NAND2x1_ASAP7_75t_R _14402_ (.A(_02263_),
    .B(_10296_),
    .Y(_10330_));
 OA211x2_ASAP7_75t_R _14403_ (.A1(_10185_),
    .A2(_10297_),
    .B(_10330_),
    .C(_10290_),
    .Y(_10331_));
 OA21x2_ASAP7_75t_R _14404_ (.A1(_10329_),
    .A2(_10331_),
    .B(_10325_),
    .Y(_03056_));
 NOR2x1_ASAP7_75t_R _14405_ (.A(_01828_),
    .B(_10291_),
    .Y(_10332_));
 NAND2x1_ASAP7_75t_R _14406_ (.A(_02262_),
    .B(_10296_),
    .Y(_10333_));
 OA211x2_ASAP7_75t_R _14407_ (.A1(_10184_),
    .A2(_10297_),
    .B(_10333_),
    .C(_10290_),
    .Y(_10334_));
 OA21x2_ASAP7_75t_R _14408_ (.A1(_10332_),
    .A2(_10334_),
    .B(_10325_),
    .Y(_03057_));
 OR4x1_ASAP7_75t_R _14409_ (.A(_08712_),
    .B(_01826_),
    .C(_10153_),
    .D(_10231_),
    .Y(_10335_));
 INVx1_ASAP7_75t_R _14410_ (.A(_10335_),
    .Y(_03058_));
 NAND2x1_ASAP7_75t_R _14411_ (.A(_10152_),
    .B(_10295_),
    .Y(_10336_));
 AO21x1_ASAP7_75t_R _14412_ (.A1(_10247_),
    .A2(_10242_),
    .B(_10176_),
    .Y(_10337_));
 AND3x1_ASAP7_75t_R _14413_ (.A(_10300_),
    .B(_10336_),
    .C(_10337_),
    .Y(_10338_));
 NOR2x1_ASAP7_75t_R _14414_ (.A(_10013_),
    .B(_10338_),
    .Y(_03059_));
 NOR2x1_ASAP7_75t_R _14415_ (.A(_01825_),
    .B(_10300_),
    .Y(_10339_));
 INVx1_ASAP7_75t_R _14416_ (.A(_02301_),
    .Y(_10340_));
 NAND2x1_ASAP7_75t_R _14417_ (.A(_02259_),
    .B(_10296_),
    .Y(_10341_));
 OA211x2_ASAP7_75t_R _14418_ (.A1(_10340_),
    .A2(_10298_),
    .B(_10341_),
    .C(_10290_),
    .Y(_10342_));
 OA21x2_ASAP7_75t_R _14419_ (.A1(_10339_),
    .A2(_10342_),
    .B(_10325_),
    .Y(_03060_));
 NOR2x1_ASAP7_75t_R _14420_ (.A(_01824_),
    .B(_10300_),
    .Y(_10343_));
 INVx1_ASAP7_75t_R _14421_ (.A(_02300_),
    .Y(_10344_));
 NAND2x1_ASAP7_75t_R _14422_ (.A(_02258_),
    .B(_10296_),
    .Y(_10345_));
 OA211x2_ASAP7_75t_R _14423_ (.A1(_10344_),
    .A2(_10298_),
    .B(_10345_),
    .C(_10290_),
    .Y(_10346_));
 OA21x2_ASAP7_75t_R _14424_ (.A1(_10343_),
    .A2(_10346_),
    .B(_10325_),
    .Y(_03061_));
 AND2x2_ASAP7_75t_R _14425_ (.A(_09957_),
    .B(_00009_),
    .Y(_03062_));
 BUFx6f_ASAP7_75t_R _14426_ (.A(_02218_),
    .Y(_10347_));
 NOR2x2_ASAP7_75t_R _14427_ (.A(_10347_),
    .B(_02219_),
    .Y(_10348_));
 BUFx6f_ASAP7_75t_R _14428_ (.A(_02176_),
    .Y(_10349_));
 OR2x6_ASAP7_75t_R _14429_ (.A(_10349_),
    .B(_02177_),
    .Y(_10350_));
 BUFx6f_ASAP7_75t_R _14430_ (.A(_01812_),
    .Y(_10351_));
 INVx3_ASAP7_75t_R _14431_ (.A(_10351_),
    .Y(_10352_));
 BUFx6f_ASAP7_75t_R _14432_ (.A(_01817_),
    .Y(_10353_));
 AND2x2_ASAP7_75t_R _14433_ (.A(_10351_),
    .B(_00009_),
    .Y(_10354_));
 AO21x1_ASAP7_75t_R _14434_ (.A1(_10352_),
    .A2(_10353_),
    .B(_10354_),
    .Y(_10355_));
 INVx1_ASAP7_75t_R _14435_ (.A(_02178_),
    .Y(_10356_));
 INVx1_ASAP7_75t_R _14436_ (.A(_02179_),
    .Y(_10357_));
 INVx1_ASAP7_75t_R _14437_ (.A(_02220_),
    .Y(_10358_));
 INVx1_ASAP7_75t_R _14438_ (.A(_02221_),
    .Y(_10359_));
 BUFx6f_ASAP7_75t_R _14439_ (.A(_02222_),
    .Y(_10360_));
 OA33x2_ASAP7_75t_R _14440_ (.A1(_10356_),
    .A2(_10357_),
    .A3(_02180_),
    .B1(_10358_),
    .B2(_10359_),
    .B3(_10360_),
    .Y(_10361_));
 NOR2x1_ASAP7_75t_R _14441_ (.A(_10349_),
    .B(_10347_),
    .Y(_10362_));
 INVx1_ASAP7_75t_R _14442_ (.A(_10349_),
    .Y(_10363_));
 INVx2_ASAP7_75t_R _14443_ (.A(_02180_),
    .Y(_10364_));
 AND2x4_ASAP7_75t_R _14444_ (.A(_02178_),
    .B(_02179_),
    .Y(_10365_));
 AND4x1_ASAP7_75t_R _14445_ (.A(_10363_),
    .B(_10364_),
    .C(_02181_),
    .D(_10365_),
    .Y(_10366_));
 AO32x2_ASAP7_75t_R _14446_ (.A1(_10355_),
    .A2(_10361_),
    .A3(_10362_),
    .B1(_10348_),
    .B2(_10366_),
    .Y(_10367_));
 BUFx6f_ASAP7_75t_R _14447_ (.A(_01813_),
    .Y(_10368_));
 INVx2_ASAP7_75t_R _14448_ (.A(_01817_),
    .Y(_10369_));
 NAND2x1_ASAP7_75t_R _14449_ (.A(_10368_),
    .B(_10369_),
    .Y(_10370_));
 INVx2_ASAP7_75t_R _14450_ (.A(_10360_),
    .Y(_10371_));
 AND2x4_ASAP7_75t_R _14451_ (.A(_02220_),
    .B(_02221_),
    .Y(_10372_));
 AOI21x1_ASAP7_75t_R _14452_ (.A1(_10371_),
    .A2(_10372_),
    .B(_10347_),
    .Y(_10373_));
 INVx1_ASAP7_75t_R _14453_ (.A(_10368_),
    .Y(_10374_));
 AO21x1_ASAP7_75t_R _14454_ (.A1(_10353_),
    .A2(_10348_),
    .B(_10374_),
    .Y(_10375_));
 NAND2x1_ASAP7_75t_R _14455_ (.A(_02178_),
    .B(_02179_),
    .Y(_10376_));
 OA21x2_ASAP7_75t_R _14456_ (.A1(_02180_),
    .A2(_10376_),
    .B(_10363_),
    .Y(_10377_));
 AO32x2_ASAP7_75t_R _14457_ (.A1(_10366_),
    .A2(_10370_),
    .A3(_10373_),
    .B1(_10375_),
    .B2(_10377_),
    .Y(_10378_));
 AND2x2_ASAP7_75t_R _14458_ (.A(_10352_),
    .B(_10350_),
    .Y(_10379_));
 INVx2_ASAP7_75t_R _14459_ (.A(_02181_),
    .Y(_10380_));
 OR4x1_ASAP7_75t_R _14460_ (.A(_10349_),
    .B(_02180_),
    .C(_10380_),
    .D(_10376_),
    .Y(_10381_));
 AO221x1_ASAP7_75t_R _14461_ (.A1(_10350_),
    .A2(_10367_),
    .B1(_10378_),
    .B2(_10379_),
    .C(_10381_),
    .Y(_10382_));
 AOI221x1_ASAP7_75t_R _14462_ (.A1(_10368_),
    .A2(_10353_),
    .B1(_10364_),
    .B2(_10365_),
    .C(_10351_),
    .Y(_10383_));
 INVx1_ASAP7_75t_R _14463_ (.A(_02177_),
    .Y(_10384_));
 NAND2x1_ASAP7_75t_R _14464_ (.A(_02220_),
    .B(_02221_),
    .Y(_10385_));
 OR3x1_ASAP7_75t_R _14465_ (.A(_10384_),
    .B(_10360_),
    .C(_10385_),
    .Y(_10386_));
 OR4x1_ASAP7_75t_R _14466_ (.A(_10351_),
    .B(_01817_),
    .C(_02177_),
    .D(_10347_),
    .Y(_10387_));
 OAI21x1_ASAP7_75t_R _14467_ (.A1(_10360_),
    .A2(_10385_),
    .B(_10387_),
    .Y(_10388_));
 NOR2x1_ASAP7_75t_R _14468_ (.A(_10347_),
    .B(_02223_),
    .Y(_10389_));
 OR3x1_ASAP7_75t_R _14469_ (.A(_10360_),
    .B(_10385_),
    .C(_10389_),
    .Y(_10390_));
 OA211x2_ASAP7_75t_R _14470_ (.A1(_10383_),
    .A2(_10386_),
    .B(_10388_),
    .C(_10390_),
    .Y(_10391_));
 INVx1_ASAP7_75t_R _14471_ (.A(_00009_),
    .Y(_10392_));
 OA211x2_ASAP7_75t_R _14472_ (.A1(_02180_),
    .A2(_10376_),
    .B(_10392_),
    .C(_10363_),
    .Y(_10393_));
 OR3x1_ASAP7_75t_R _14473_ (.A(_10351_),
    .B(_10353_),
    .C(_10349_),
    .Y(_10394_));
 AOI21x1_ASAP7_75t_R _14474_ (.A1(_10364_),
    .A2(_10365_),
    .B(_10394_),
    .Y(_10395_));
 NOR2x1_ASAP7_75t_R _14475_ (.A(_10351_),
    .B(_10368_),
    .Y(_10396_));
 AO211x2_ASAP7_75t_R _14476_ (.A1(_10351_),
    .A2(_10393_),
    .B(_10395_),
    .C(_10396_),
    .Y(_10397_));
 AO22x2_ASAP7_75t_R _14477_ (.A1(_10363_),
    .A2(_10391_),
    .B1(_10397_),
    .B2(_10373_),
    .Y(_10398_));
 NOR3x2_ASAP7_75t_R _14478_ (.B(_10382_),
    .C(_10398_),
    .Y(_10399_),
    .A(_10348_));
 AO21x2_ASAP7_75t_R _14479_ (.A1(_10371_),
    .A2(_10372_),
    .B(_10347_),
    .Y(_10400_));
 OR2x2_ASAP7_75t_R _14480_ (.A(_10353_),
    .B(_10389_),
    .Y(_10401_));
 AO31x2_ASAP7_75t_R _14481_ (.A1(_10371_),
    .A2(_10372_),
    .A3(_10389_),
    .B(_10369_),
    .Y(_10402_));
 NOR2x1_ASAP7_75t_R _14482_ (.A(_10349_),
    .B(_02177_),
    .Y(_10403_));
 AO32x2_ASAP7_75t_R _14483_ (.A1(_10366_),
    .A2(_10400_),
    .A3(_10401_),
    .B1(_10402_),
    .B2(_10403_),
    .Y(_10404_));
 AOI21x1_ASAP7_75t_R _14484_ (.A1(_10353_),
    .A2(_10348_),
    .B(_10404_),
    .Y(_10405_));
 AND5x2_ASAP7_75t_R _14485_ (.A(_10352_),
    .B(_10368_),
    .C(_10353_),
    .D(_10382_),
    .E(_10405_),
    .Y(_10406_));
 NOR2x1_ASAP7_75t_R _14486_ (.A(_10399_),
    .B(_10406_),
    .Y(_10407_));
 BUFx6f_ASAP7_75t_R _14487_ (.A(_10407_),
    .Y(_10408_));
 BUFx6f_ASAP7_75t_R _14488_ (.A(_10406_),
    .Y(_10409_));
 AO221x1_ASAP7_75t_R _14489_ (.A1(_02187_),
    .A2(_10399_),
    .B1(_10409_),
    .B2(_01823_),
    .C(_09211_),
    .Y(_10410_));
 AOI21x1_ASAP7_75t_R _14490_ (.A1(_02229_),
    .A2(_10408_),
    .B(_10410_),
    .Y(_03063_));
 AO221x1_ASAP7_75t_R _14491_ (.A1(_02186_),
    .A2(_10399_),
    .B1(_10409_),
    .B2(_01822_),
    .C(_09211_),
    .Y(_10411_));
 AOI21x1_ASAP7_75t_R _14492_ (.A1(_02228_),
    .A2(_10408_),
    .B(_10411_),
    .Y(_03064_));
 AO221x1_ASAP7_75t_R _14493_ (.A1(_02185_),
    .A2(_10399_),
    .B1(_10409_),
    .B2(_01821_),
    .C(_09211_),
    .Y(_10412_));
 AOI21x1_ASAP7_75t_R _14494_ (.A1(_02227_),
    .A2(_10408_),
    .B(_10412_),
    .Y(_03065_));
 AO221x1_ASAP7_75t_R _14495_ (.A1(_02184_),
    .A2(_10399_),
    .B1(_10409_),
    .B2(_01820_),
    .C(_09211_),
    .Y(_10413_));
 AOI21x1_ASAP7_75t_R _14496_ (.A1(_02226_),
    .A2(_10408_),
    .B(_10413_),
    .Y(_03066_));
 AO221x1_ASAP7_75t_R _14497_ (.A1(_02183_),
    .A2(_10399_),
    .B1(_10409_),
    .B2(_01819_),
    .C(_09211_),
    .Y(_10414_));
 AOI21x1_ASAP7_75t_R _14498_ (.A1(_02225_),
    .A2(_10408_),
    .B(_10414_),
    .Y(_03067_));
 AO221x1_ASAP7_75t_R _14499_ (.A1(_02182_),
    .A2(_10399_),
    .B1(_10409_),
    .B2(_01818_),
    .C(_09211_),
    .Y(_10415_));
 AOI21x1_ASAP7_75t_R _14500_ (.A1(_02224_),
    .A2(_10408_),
    .B(_10415_),
    .Y(_03068_));
 INVx1_ASAP7_75t_R _14501_ (.A(_02223_),
    .Y(_10416_));
 AND3x1_ASAP7_75t_R _14502_ (.A(_09632_),
    .B(_10416_),
    .C(_10408_),
    .Y(_03069_));
 AOI221x1_ASAP7_75t_R _14503_ (.A1(_01816_),
    .A2(_10409_),
    .B1(_10408_),
    .B2(_10360_),
    .C(_10021_),
    .Y(_03070_));
 INVx1_ASAP7_75t_R _14504_ (.A(_01815_),
    .Y(_10417_));
 NOR2x1_ASAP7_75t_R _14505_ (.A(_09924_),
    .B(_02221_),
    .Y(_10418_));
 AO32x1_ASAP7_75t_R _14506_ (.A1(_09830_),
    .A2(_10417_),
    .A3(_10409_),
    .B1(_10407_),
    .B2(_10418_),
    .Y(_03071_));
 INVx1_ASAP7_75t_R _14507_ (.A(_01814_),
    .Y(_10419_));
 NOR2x1_ASAP7_75t_R _14508_ (.A(_09924_),
    .B(_02220_),
    .Y(_10420_));
 AO32x1_ASAP7_75t_R _14509_ (.A1(_09830_),
    .A2(_10419_),
    .A3(_10409_),
    .B1(_10407_),
    .B2(_10420_),
    .Y(_03072_));
 NOR2x1_ASAP7_75t_R _14510_ (.A(_10348_),
    .B(_10400_),
    .Y(_10421_));
 NOR2x1_ASAP7_75t_R _14511_ (.A(_10349_),
    .B(_10348_),
    .Y(_10422_));
 AOI22x1_ASAP7_75t_R _14512_ (.A1(_10397_),
    .A2(_10421_),
    .B1(_10422_),
    .B2(_10391_),
    .Y(_10423_));
 NOR2x1_ASAP7_75t_R _14513_ (.A(_10013_),
    .B(_10423_),
    .Y(_03073_));
 NOR2x1_ASAP7_75t_R _14514_ (.A(_10348_),
    .B(_10398_),
    .Y(_10424_));
 NAND2x1_ASAP7_75t_R _14515_ (.A(_10352_),
    .B(_10368_),
    .Y(_10425_));
 OR4x1_ASAP7_75t_R _14516_ (.A(_10369_),
    .B(_10348_),
    .C(_10425_),
    .D(_10404_),
    .Y(_10426_));
 AND3x1_ASAP7_75t_R _14517_ (.A(_10382_),
    .B(_10424_),
    .C(_10426_),
    .Y(_10427_));
 NOR2x1_ASAP7_75t_R _14518_ (.A(_10013_),
    .B(_10427_),
    .Y(_03074_));
 AO221x1_ASAP7_75t_R _14519_ (.A1(_02175_),
    .A2(_10399_),
    .B1(_10409_),
    .B2(_01811_),
    .C(_09314_),
    .Y(_10428_));
 AOI21x1_ASAP7_75t_R _14520_ (.A1(_02217_),
    .A2(_10408_),
    .B(_10428_),
    .Y(_03075_));
 AO221x1_ASAP7_75t_R _14521_ (.A1(_02174_),
    .A2(_10399_),
    .B1(_10406_),
    .B2(_01810_),
    .C(_09314_),
    .Y(_10429_));
 AOI21x1_ASAP7_75t_R _14522_ (.A1(_02216_),
    .A2(_10408_),
    .B(_10429_),
    .Y(_03076_));
 AND3x4_ASAP7_75t_R _14523_ (.A(_10371_),
    .B(_10372_),
    .C(_10389_),
    .Y(_10430_));
 AO21x2_ASAP7_75t_R _14524_ (.A1(_10364_),
    .A2(_10365_),
    .B(_10349_),
    .Y(_10431_));
 AO22x1_ASAP7_75t_R _14525_ (.A1(_10366_),
    .A2(_10348_),
    .B1(_10430_),
    .B2(_10431_),
    .Y(_10432_));
 OR4x1_ASAP7_75t_R _14526_ (.A(_10353_),
    .B(_10425_),
    .C(_10404_),
    .D(_10432_),
    .Y(_10433_));
 AO21x2_ASAP7_75t_R _14527_ (.A1(_10430_),
    .A2(_10423_),
    .B(_10433_),
    .Y(_10434_));
 BUFx12f_ASAP7_75t_R _14528_ (.A(_10434_),
    .Y(_10435_));
 NOR2x1_ASAP7_75t_R _14529_ (.A(_01823_),
    .B(_10435_),
    .Y(_10436_));
 INVx1_ASAP7_75t_R _14530_ (.A(_02187_),
    .Y(_10437_));
 AOI211x1_ASAP7_75t_R _14531_ (.A1(_10352_),
    .A2(_10378_),
    .B(_10367_),
    .C(_10403_),
    .Y(_10438_));
 BUFx6f_ASAP7_75t_R _14532_ (.A(_10438_),
    .Y(_10439_));
 BUFx6f_ASAP7_75t_R _14533_ (.A(_10438_),
    .Y(_10440_));
 NAND2x1_ASAP7_75t_R _14534_ (.A(_02229_),
    .B(_10440_),
    .Y(_10441_));
 BUFx6f_ASAP7_75t_R _14535_ (.A(_10434_),
    .Y(_10442_));
 OA211x2_ASAP7_75t_R _14536_ (.A1(_10437_),
    .A2(_10439_),
    .B(_10441_),
    .C(_10442_),
    .Y(_10443_));
 OA21x2_ASAP7_75t_R _14537_ (.A1(_10436_),
    .A2(_10443_),
    .B(_10325_),
    .Y(_03077_));
 NOR2x1_ASAP7_75t_R _14538_ (.A(_01822_),
    .B(_10435_),
    .Y(_10444_));
 INVx1_ASAP7_75t_R _14539_ (.A(_02186_),
    .Y(_10445_));
 NAND2x1_ASAP7_75t_R _14540_ (.A(_02228_),
    .B(_10440_),
    .Y(_10446_));
 OA211x2_ASAP7_75t_R _14541_ (.A1(_10445_),
    .A2(_10439_),
    .B(_10446_),
    .C(_10442_),
    .Y(_10447_));
 OA21x2_ASAP7_75t_R _14542_ (.A1(_10444_),
    .A2(_10447_),
    .B(_10325_),
    .Y(_03078_));
 NOR2x1_ASAP7_75t_R _14543_ (.A(_01821_),
    .B(_10435_),
    .Y(_10448_));
 INVx1_ASAP7_75t_R _14544_ (.A(_02185_),
    .Y(_10449_));
 NAND2x1_ASAP7_75t_R _14545_ (.A(_02227_),
    .B(_10440_),
    .Y(_10450_));
 OA211x2_ASAP7_75t_R _14546_ (.A1(_10449_),
    .A2(_10439_),
    .B(_10450_),
    .C(_10442_),
    .Y(_10451_));
 OA21x2_ASAP7_75t_R _14547_ (.A1(_10448_),
    .A2(_10451_),
    .B(_10325_),
    .Y(_03079_));
 NOR2x1_ASAP7_75t_R _14548_ (.A(_01820_),
    .B(_10435_),
    .Y(_10452_));
 INVx1_ASAP7_75t_R _14549_ (.A(_02184_),
    .Y(_10453_));
 NAND2x1_ASAP7_75t_R _14550_ (.A(_02226_),
    .B(_10440_),
    .Y(_10454_));
 OA211x2_ASAP7_75t_R _14551_ (.A1(_10453_),
    .A2(_10439_),
    .B(_10454_),
    .C(_10442_),
    .Y(_10455_));
 OA21x2_ASAP7_75t_R _14552_ (.A1(_10452_),
    .A2(_10455_),
    .B(_10325_),
    .Y(_03080_));
 NOR2x1_ASAP7_75t_R _14553_ (.A(_01819_),
    .B(_10435_),
    .Y(_10456_));
 INVx1_ASAP7_75t_R _14554_ (.A(_02183_),
    .Y(_10457_));
 NAND2x1_ASAP7_75t_R _14555_ (.A(_02225_),
    .B(_10440_),
    .Y(_10458_));
 OA211x2_ASAP7_75t_R _14556_ (.A1(_10457_),
    .A2(_10439_),
    .B(_10458_),
    .C(_10442_),
    .Y(_10459_));
 BUFx6f_ASAP7_75t_R _14557_ (.A(_08665_),
    .Y(_10460_));
 OA21x2_ASAP7_75t_R _14558_ (.A1(_10456_),
    .A2(_10459_),
    .B(_10460_),
    .Y(_03081_));
 NOR2x1_ASAP7_75t_R _14559_ (.A(_01818_),
    .B(_10435_),
    .Y(_10461_));
 INVx1_ASAP7_75t_R _14560_ (.A(_02182_),
    .Y(_10462_));
 NAND2x1_ASAP7_75t_R _14561_ (.A(_02224_),
    .B(_10440_),
    .Y(_10463_));
 OA211x2_ASAP7_75t_R _14562_ (.A1(_10462_),
    .A2(_10439_),
    .B(_10463_),
    .C(_10442_),
    .Y(_10464_));
 OA21x2_ASAP7_75t_R _14563_ (.A1(_10461_),
    .A2(_10464_),
    .B(_10460_),
    .Y(_03082_));
 NOR2x1_ASAP7_75t_R _14564_ (.A(_10380_),
    .B(_10439_),
    .Y(_10465_));
 AO21x1_ASAP7_75t_R _14565_ (.A1(_02223_),
    .A2(_10439_),
    .B(_10465_),
    .Y(_10466_));
 AOI21x1_ASAP7_75t_R _14566_ (.A1(_10435_),
    .A2(_10466_),
    .B(_10289_),
    .Y(_03083_));
 NOR2x1_ASAP7_75t_R _14567_ (.A(_01816_),
    .B(_10435_),
    .Y(_10467_));
 NAND2x1_ASAP7_75t_R _14568_ (.A(_10360_),
    .B(_10438_),
    .Y(_10468_));
 OA211x2_ASAP7_75t_R _14569_ (.A1(_10364_),
    .A2(_10439_),
    .B(_10468_),
    .C(_10442_),
    .Y(_10469_));
 OA21x2_ASAP7_75t_R _14570_ (.A1(_10467_),
    .A2(_10469_),
    .B(_10460_),
    .Y(_03084_));
 NOR2x1_ASAP7_75t_R _14571_ (.A(_01815_),
    .B(_10435_),
    .Y(_10470_));
 NAND2x1_ASAP7_75t_R _14572_ (.A(_02221_),
    .B(_10438_),
    .Y(_10471_));
 OA211x2_ASAP7_75t_R _14573_ (.A1(_10357_),
    .A2(_10439_),
    .B(_10471_),
    .C(_10442_),
    .Y(_10472_));
 OA21x2_ASAP7_75t_R _14574_ (.A1(_10470_),
    .A2(_10472_),
    .B(_10460_),
    .Y(_03085_));
 NOR2x1_ASAP7_75t_R _14575_ (.A(_01814_),
    .B(_10435_),
    .Y(_10473_));
 NAND2x1_ASAP7_75t_R _14576_ (.A(_02220_),
    .B(_10438_),
    .Y(_10474_));
 OA211x2_ASAP7_75t_R _14577_ (.A1(_10356_),
    .A2(_10440_),
    .B(_10474_),
    .C(_10434_),
    .Y(_10475_));
 OA21x2_ASAP7_75t_R _14578_ (.A1(_10473_),
    .A2(_10475_),
    .B(_10460_),
    .Y(_03086_));
 AO21x1_ASAP7_75t_R _14579_ (.A1(_10352_),
    .A2(_10378_),
    .B(_10367_),
    .Y(_10476_));
 AND3x1_ASAP7_75t_R _14580_ (.A(_09632_),
    .B(_10350_),
    .C(_10476_),
    .Y(_03087_));
 NAND2x1_ASAP7_75t_R _14581_ (.A(_10433_),
    .B(_10440_),
    .Y(_10477_));
 AO21x1_ASAP7_75t_R _14582_ (.A1(_10430_),
    .A2(_10423_),
    .B(_10477_),
    .Y(_10478_));
 AND2x2_ASAP7_75t_R _14583_ (.A(_09957_),
    .B(_10478_),
    .Y(_03088_));
 NOR2x1_ASAP7_75t_R _14584_ (.A(_01811_),
    .B(_10442_),
    .Y(_10479_));
 INVx1_ASAP7_75t_R _14585_ (.A(_02175_),
    .Y(_10480_));
 NAND2x1_ASAP7_75t_R _14586_ (.A(_02217_),
    .B(_10438_),
    .Y(_10481_));
 OA211x2_ASAP7_75t_R _14587_ (.A1(_10480_),
    .A2(_10440_),
    .B(_10481_),
    .C(_10434_),
    .Y(_10482_));
 OA21x2_ASAP7_75t_R _14588_ (.A1(_10479_),
    .A2(_10482_),
    .B(_10460_),
    .Y(_03089_));
 NOR2x1_ASAP7_75t_R _14589_ (.A(_01810_),
    .B(_10442_),
    .Y(_10483_));
 INVx1_ASAP7_75t_R _14590_ (.A(_02174_),
    .Y(_10484_));
 NAND2x1_ASAP7_75t_R _14591_ (.A(_02216_),
    .B(_10438_),
    .Y(_10485_));
 OA211x2_ASAP7_75t_R _14592_ (.A1(_10484_),
    .A2(_10440_),
    .B(_10485_),
    .C(_10434_),
    .Y(_10486_));
 OA21x2_ASAP7_75t_R _14593_ (.A1(_10483_),
    .A2(_10486_),
    .B(_10460_),
    .Y(_03090_));
 AOI22x1_ASAP7_75t_R _14594_ (.A1(_10366_),
    .A2(_10348_),
    .B1(_10430_),
    .B2(_10431_),
    .Y(_10487_));
 OA21x2_ASAP7_75t_R _14595_ (.A1(_10353_),
    .A2(_10487_),
    .B(_10368_),
    .Y(_10488_));
 AO21x2_ASAP7_75t_R _14596_ (.A1(_10405_),
    .A2(_10488_),
    .B(_10351_),
    .Y(_10489_));
 BUFx6f_ASAP7_75t_R _14597_ (.A(_10489_),
    .Y(_10490_));
 NOR2x1_ASAP7_75t_R _14598_ (.A(_10349_),
    .B(_10387_),
    .Y(_10491_));
 OA21x2_ASAP7_75t_R _14599_ (.A1(_10397_),
    .A2(_10491_),
    .B(_02219_),
    .Y(_10492_));
 OR2x2_ASAP7_75t_R _14600_ (.A(_10431_),
    .B(_10375_),
    .Y(_10493_));
 OAI22x1_ASAP7_75t_R _14601_ (.A1(_10352_),
    .A2(_10431_),
    .B1(_10404_),
    .B2(_10493_),
    .Y(_10494_));
 OAI21x1_ASAP7_75t_R _14602_ (.A1(_10400_),
    .A2(_10492_),
    .B(_10494_),
    .Y(_10495_));
 BUFx6f_ASAP7_75t_R _14603_ (.A(_10495_),
    .Y(_10496_));
 OA22x2_ASAP7_75t_R _14604_ (.A1(_01823_),
    .A2(_10490_),
    .B1(_10496_),
    .B2(_02187_),
    .Y(_10497_));
 AOI21x1_ASAP7_75t_R _14605_ (.A1(_10405_),
    .A2(_10488_),
    .B(_10351_),
    .Y(_10498_));
 BUFx6f_ASAP7_75t_R _14606_ (.A(_10498_),
    .Y(_10499_));
 OA21x2_ASAP7_75t_R _14607_ (.A1(_10400_),
    .A2(_10492_),
    .B(_10494_),
    .Y(_10500_));
 OR3x1_ASAP7_75t_R _14608_ (.A(_02229_),
    .B(_10499_),
    .C(_10500_),
    .Y(_10501_));
 AOI21x1_ASAP7_75t_R _14609_ (.A1(_10497_),
    .A2(_10501_),
    .B(_10289_),
    .Y(_03091_));
 OA22x2_ASAP7_75t_R _14610_ (.A1(_01822_),
    .A2(_10490_),
    .B1(_10496_),
    .B2(_02186_),
    .Y(_10502_));
 OR3x1_ASAP7_75t_R _14611_ (.A(_02228_),
    .B(_10499_),
    .C(_10500_),
    .Y(_10503_));
 AOI21x1_ASAP7_75t_R _14612_ (.A1(_10502_),
    .A2(_10503_),
    .B(_10289_),
    .Y(_03092_));
 OA22x2_ASAP7_75t_R _14613_ (.A1(_01821_),
    .A2(_10490_),
    .B1(_10496_),
    .B2(_02185_),
    .Y(_10504_));
 OR3x1_ASAP7_75t_R _14614_ (.A(_02227_),
    .B(_10499_),
    .C(_10500_),
    .Y(_10505_));
 AOI21x1_ASAP7_75t_R _14615_ (.A1(_10504_),
    .A2(_10505_),
    .B(_10289_),
    .Y(_03093_));
 OA22x2_ASAP7_75t_R _14616_ (.A1(_01820_),
    .A2(_10490_),
    .B1(_10496_),
    .B2(_02184_),
    .Y(_10506_));
 OR3x1_ASAP7_75t_R _14617_ (.A(_02226_),
    .B(_10499_),
    .C(_10500_),
    .Y(_10507_));
 AOI21x1_ASAP7_75t_R _14618_ (.A1(_10506_),
    .A2(_10507_),
    .B(_10289_),
    .Y(_03094_));
 OA22x2_ASAP7_75t_R _14619_ (.A1(_01819_),
    .A2(_10490_),
    .B1(_10496_),
    .B2(_02183_),
    .Y(_10508_));
 OR3x1_ASAP7_75t_R _14620_ (.A(_02225_),
    .B(_10499_),
    .C(_10500_),
    .Y(_10509_));
 AOI21x1_ASAP7_75t_R _14621_ (.A1(_10508_),
    .A2(_10509_),
    .B(_10289_),
    .Y(_03095_));
 OA22x2_ASAP7_75t_R _14622_ (.A1(_01818_),
    .A2(_10490_),
    .B1(_10496_),
    .B2(_02182_),
    .Y(_10510_));
 OR3x1_ASAP7_75t_R _14623_ (.A(_02224_),
    .B(_10499_),
    .C(_10500_),
    .Y(_10511_));
 AOI21x1_ASAP7_75t_R _14624_ (.A1(_10510_),
    .A2(_10511_),
    .B(_10289_),
    .Y(_03096_));
 OR2x6_ASAP7_75t_R _14625_ (.A(_10400_),
    .B(_10492_),
    .Y(_10512_));
 AO32x1_ASAP7_75t_R _14626_ (.A1(_10380_),
    .A2(_10512_),
    .A3(_10494_),
    .B1(_10499_),
    .B2(_10369_),
    .Y(_10513_));
 AND3x1_ASAP7_75t_R _14627_ (.A(_10416_),
    .B(_10489_),
    .C(_10496_),
    .Y(_10514_));
 OA21x2_ASAP7_75t_R _14628_ (.A1(_10513_),
    .A2(_10514_),
    .B(_10460_),
    .Y(_03097_));
 OAI22x1_ASAP7_75t_R _14629_ (.A1(_01816_),
    .A2(_10490_),
    .B1(_10496_),
    .B2(_02180_),
    .Y(_10515_));
 AND3x1_ASAP7_75t_R _14630_ (.A(_10371_),
    .B(_10489_),
    .C(_10495_),
    .Y(_10516_));
 OA21x2_ASAP7_75t_R _14631_ (.A1(_10515_),
    .A2(_10516_),
    .B(_10460_),
    .Y(_03098_));
 AO32x1_ASAP7_75t_R _14632_ (.A1(_10357_),
    .A2(_10512_),
    .A3(_10494_),
    .B1(_10499_),
    .B2(_10417_),
    .Y(_10517_));
 AND3x1_ASAP7_75t_R _14633_ (.A(_10359_),
    .B(_10489_),
    .C(_10495_),
    .Y(_10518_));
 OA21x2_ASAP7_75t_R _14634_ (.A1(_10517_),
    .A2(_10518_),
    .B(_10460_),
    .Y(_03099_));
 AO32x1_ASAP7_75t_R _14635_ (.A1(_10356_),
    .A2(_10512_),
    .A3(_10494_),
    .B1(_10498_),
    .B2(_10419_),
    .Y(_10519_));
 AND3x1_ASAP7_75t_R _14636_ (.A(_10358_),
    .B(_10489_),
    .C(_10495_),
    .Y(_10520_));
 BUFx6f_ASAP7_75t_R _14637_ (.A(_09229_),
    .Y(_10521_));
 OA21x2_ASAP7_75t_R _14638_ (.A1(_10519_),
    .A2(_10520_),
    .B(_10521_),
    .Y(_03100_));
 OA21x2_ASAP7_75t_R _14639_ (.A1(_10353_),
    .A2(_10487_),
    .B(_10405_),
    .Y(_10522_));
 OR3x1_ASAP7_75t_R _14640_ (.A(_08642_),
    .B(_10425_),
    .C(_10522_),
    .Y(_10523_));
 INVx1_ASAP7_75t_R _14641_ (.A(_10523_),
    .Y(_03101_));
 AND2x2_ASAP7_75t_R _14642_ (.A(_10350_),
    .B(_10476_),
    .Y(_10524_));
 OA21x2_ASAP7_75t_R _14643_ (.A1(_10431_),
    .A2(_10524_),
    .B(_10490_),
    .Y(_10525_));
 AOI21x1_ASAP7_75t_R _14644_ (.A1(_10512_),
    .A2(_10525_),
    .B(_10289_),
    .Y(_03102_));
 OA22x2_ASAP7_75t_R _14645_ (.A1(_01811_),
    .A2(_10490_),
    .B1(_10496_),
    .B2(_02175_),
    .Y(_10526_));
 OR3x1_ASAP7_75t_R _14646_ (.A(_02217_),
    .B(_10499_),
    .C(_10500_),
    .Y(_10527_));
 AOI21x1_ASAP7_75t_R _14647_ (.A1(_10526_),
    .A2(_10527_),
    .B(_10289_),
    .Y(_03103_));
 OA22x2_ASAP7_75t_R _14648_ (.A1(_01810_),
    .A2(_10490_),
    .B1(_10496_),
    .B2(_02174_),
    .Y(_10528_));
 OR3x1_ASAP7_75t_R _14649_ (.A(_02216_),
    .B(_10499_),
    .C(_10500_),
    .Y(_10529_));
 BUFx12f_ASAP7_75t_R _14650_ (.A(_09118_),
    .Y(_10530_));
 AOI21x1_ASAP7_75t_R _14651_ (.A1(_10528_),
    .A2(_10529_),
    .B(_10530_),
    .Y(_03104_));
 AND2x2_ASAP7_75t_R _14652_ (.A(_09957_),
    .B(_00010_),
    .Y(_03105_));
 OR2x6_ASAP7_75t_R _14653_ (.A(_02092_),
    .B(_02093_),
    .Y(_10531_));
 INVx1_ASAP7_75t_R _14654_ (.A(_02136_),
    .Y(_10532_));
 INVx1_ASAP7_75t_R _14655_ (.A(_02138_),
    .Y(_10533_));
 INVx2_ASAP7_75t_R _14656_ (.A(_02134_),
    .Y(_10534_));
 OA31x2_ASAP7_75t_R _14657_ (.A1(_10532_),
    .A2(_02137_),
    .A3(_10533_),
    .B1(_10534_),
    .Y(_10535_));
 BUFx6f_ASAP7_75t_R _14658_ (.A(_01785_),
    .Y(_10536_));
 INVx1_ASAP7_75t_R _14659_ (.A(_10536_),
    .Y(_10537_));
 BUFx6f_ASAP7_75t_R _14660_ (.A(_01784_),
    .Y(_10538_));
 INVx1_ASAP7_75t_R _14661_ (.A(_10538_),
    .Y(_10539_));
 OA21x2_ASAP7_75t_R _14662_ (.A1(_10537_),
    .A2(_01789_),
    .B(_10539_),
    .Y(_10540_));
 OR2x6_ASAP7_75t_R _14663_ (.A(_02134_),
    .B(_02135_),
    .Y(_10541_));
 INVx1_ASAP7_75t_R _14664_ (.A(_10541_),
    .Y(_10542_));
 AO21x1_ASAP7_75t_R _14665_ (.A1(_10535_),
    .A2(_10540_),
    .B(_10542_),
    .Y(_10543_));
 INVx1_ASAP7_75t_R _14666_ (.A(_02097_),
    .Y(_10544_));
 NAND2x1_ASAP7_75t_R _14667_ (.A(_02094_),
    .B(_02096_),
    .Y(_10545_));
 OR4x1_ASAP7_75t_R _14668_ (.A(_02092_),
    .B(_02095_),
    .C(_10544_),
    .D(_10545_),
    .Y(_10546_));
 AO21x2_ASAP7_75t_R _14669_ (.A1(_10531_),
    .A2(_10543_),
    .B(_10546_),
    .Y(_10547_));
 OR5x2_ASAP7_75t_R _14670_ (.A(_02134_),
    .B(_10532_),
    .C(_02137_),
    .D(_10533_),
    .E(_02139_),
    .Y(_10548_));
 AO21x1_ASAP7_75t_R _14671_ (.A1(_10531_),
    .A2(_10546_),
    .B(_10548_),
    .Y(_10549_));
 OA211x2_ASAP7_75t_R _14672_ (.A1(_10535_),
    .A2(_10546_),
    .B(_01789_),
    .C(_10541_),
    .Y(_10550_));
 AND4x1_ASAP7_75t_R _14673_ (.A(_10539_),
    .B(_10536_),
    .C(_10549_),
    .D(_10550_),
    .Y(_10551_));
 NAND2x1_ASAP7_75t_R _14674_ (.A(_10547_),
    .B(_10551_),
    .Y(_10552_));
 BUFx6f_ASAP7_75t_R _14675_ (.A(_10552_),
    .Y(_10553_));
 NOR2x1_ASAP7_75t_R _14676_ (.A(_01795_),
    .B(_10553_),
    .Y(_10554_));
 INVx1_ASAP7_75t_R _14677_ (.A(_00010_),
    .Y(_10555_));
 INVx1_ASAP7_75t_R _14678_ (.A(_02092_),
    .Y(_10556_));
 OA211x2_ASAP7_75t_R _14679_ (.A1(_02095_),
    .A2(_10545_),
    .B(_10555_),
    .C(_10556_),
    .Y(_10557_));
 INVx1_ASAP7_75t_R _14680_ (.A(_02093_),
    .Y(_10558_));
 OR3x1_ASAP7_75t_R _14681_ (.A(_10558_),
    .B(_02095_),
    .C(_10545_),
    .Y(_10559_));
 OR3x1_ASAP7_75t_R _14682_ (.A(_10538_),
    .B(_01789_),
    .C(_02092_),
    .Y(_10560_));
 INVx1_ASAP7_75t_R _14683_ (.A(_10560_),
    .Y(_10561_));
 NOR2x1_ASAP7_75t_R _14684_ (.A(_10538_),
    .B(_10536_),
    .Y(_10562_));
 AO221x1_ASAP7_75t_R _14685_ (.A1(_10538_),
    .A2(_10557_),
    .B1(_10559_),
    .B2(_10561_),
    .C(_10562_),
    .Y(_10563_));
 INVx1_ASAP7_75t_R _14686_ (.A(_02139_),
    .Y(_10564_));
 INVx2_ASAP7_75t_R _14687_ (.A(_02137_),
    .Y(_10565_));
 AND3x4_ASAP7_75t_R _14688_ (.A(_02136_),
    .B(_10565_),
    .C(_02138_),
    .Y(_10566_));
 AND3x1_ASAP7_75t_R _14689_ (.A(_10534_),
    .B(_10564_),
    .C(_10566_),
    .Y(_10567_));
 OA21x2_ASAP7_75t_R _14690_ (.A1(_02095_),
    .A2(_10545_),
    .B(_10556_),
    .Y(_10568_));
 INVx1_ASAP7_75t_R _14691_ (.A(_01789_),
    .Y(_10569_));
 OA21x2_ASAP7_75t_R _14692_ (.A1(_10537_),
    .A2(_10569_),
    .B(_10539_),
    .Y(_10570_));
 NOR2x2_ASAP7_75t_R _14693_ (.A(_02092_),
    .B(_02093_),
    .Y(_10571_));
 AO21x1_ASAP7_75t_R _14694_ (.A1(_10568_),
    .A2(_10570_),
    .B(_10571_),
    .Y(_10572_));
 AO221x1_ASAP7_75t_R _14695_ (.A1(_10563_),
    .A2(_10535_),
    .B1(_10567_),
    .B2(_10572_),
    .C(_10542_),
    .Y(_10573_));
 BUFx6f_ASAP7_75t_R _14696_ (.A(_10573_),
    .Y(_10574_));
 BUFx6f_ASAP7_75t_R _14697_ (.A(_10547_),
    .Y(_10575_));
 NOR2x1_ASAP7_75t_R _14698_ (.A(_10574_),
    .B(_10575_),
    .Y(_10576_));
 BUFx6f_ASAP7_75t_R _14699_ (.A(_10576_),
    .Y(_10577_));
 AND2x4_ASAP7_75t_R _14700_ (.A(_10547_),
    .B(_10551_),
    .Y(_10578_));
 BUFx6f_ASAP7_75t_R _14701_ (.A(_10578_),
    .Y(_10579_));
 OA21x2_ASAP7_75t_R _14702_ (.A1(_10574_),
    .A2(_10575_),
    .B(_02145_),
    .Y(_10580_));
 AOI211x1_ASAP7_75t_R _14703_ (.A1(_02103_),
    .A2(_10577_),
    .B(_10579_),
    .C(_10580_),
    .Y(_10581_));
 OA21x2_ASAP7_75t_R _14704_ (.A1(_10554_),
    .A2(_10581_),
    .B(_10521_),
    .Y(_03106_));
 NOR2x1_ASAP7_75t_R _14705_ (.A(_01794_),
    .B(_10553_),
    .Y(_10582_));
 OA21x2_ASAP7_75t_R _14706_ (.A1(_10574_),
    .A2(_10575_),
    .B(_02144_),
    .Y(_10583_));
 AOI211x1_ASAP7_75t_R _14707_ (.A1(_02102_),
    .A2(_10577_),
    .B(_10579_),
    .C(_10583_),
    .Y(_10584_));
 OA21x2_ASAP7_75t_R _14708_ (.A1(_10582_),
    .A2(_10584_),
    .B(_10521_),
    .Y(_03107_));
 NOR2x1_ASAP7_75t_R _14709_ (.A(_01793_),
    .B(_10553_),
    .Y(_10585_));
 OA21x2_ASAP7_75t_R _14710_ (.A1(_10574_),
    .A2(_10575_),
    .B(_02143_),
    .Y(_10586_));
 AOI211x1_ASAP7_75t_R _14711_ (.A1(_02101_),
    .A2(_10577_),
    .B(_10579_),
    .C(_10586_),
    .Y(_10587_));
 OA21x2_ASAP7_75t_R _14712_ (.A1(_10585_),
    .A2(_10587_),
    .B(_10521_),
    .Y(_03108_));
 NOR2x1_ASAP7_75t_R _14713_ (.A(_01792_),
    .B(_10553_),
    .Y(_10588_));
 OA21x2_ASAP7_75t_R _14714_ (.A1(_10574_),
    .A2(_10575_),
    .B(_02142_),
    .Y(_10589_));
 AOI211x1_ASAP7_75t_R _14715_ (.A1(_02100_),
    .A2(_10577_),
    .B(_10579_),
    .C(_10589_),
    .Y(_10590_));
 OA21x2_ASAP7_75t_R _14716_ (.A1(_10588_),
    .A2(_10590_),
    .B(_10521_),
    .Y(_03109_));
 NOR2x1_ASAP7_75t_R _14717_ (.A(_01791_),
    .B(_10553_),
    .Y(_10591_));
 OA21x2_ASAP7_75t_R _14718_ (.A1(_10574_),
    .A2(_10575_),
    .B(_02141_),
    .Y(_10592_));
 AOI211x1_ASAP7_75t_R _14719_ (.A1(_02099_),
    .A2(_10577_),
    .B(_10579_),
    .C(_10592_),
    .Y(_10593_));
 OA21x2_ASAP7_75t_R _14720_ (.A1(_10591_),
    .A2(_10593_),
    .B(_10521_),
    .Y(_03110_));
 NOR2x1_ASAP7_75t_R _14721_ (.A(_01790_),
    .B(_10553_),
    .Y(_10594_));
 OA21x2_ASAP7_75t_R _14722_ (.A1(_10574_),
    .A2(_10575_),
    .B(_02140_),
    .Y(_10595_));
 AOI211x1_ASAP7_75t_R _14723_ (.A1(_02098_),
    .A2(_10577_),
    .B(_10579_),
    .C(_10595_),
    .Y(_10596_));
 OA21x2_ASAP7_75t_R _14724_ (.A1(_10594_),
    .A2(_10596_),
    .B(_10521_),
    .Y(_03111_));
 OR4x1_ASAP7_75t_R _14725_ (.A(_08712_),
    .B(_02139_),
    .C(_10576_),
    .D(_10578_),
    .Y(_10597_));
 INVx1_ASAP7_75t_R _14726_ (.A(_10597_),
    .Y(_03112_));
 OR3x1_ASAP7_75t_R _14727_ (.A(_02138_),
    .B(_10577_),
    .C(_10579_),
    .Y(_10598_));
 OR2x2_ASAP7_75t_R _14728_ (.A(_01788_),
    .B(_10553_),
    .Y(_10599_));
 AOI21x1_ASAP7_75t_R _14729_ (.A1(_10598_),
    .A2(_10599_),
    .B(_10530_),
    .Y(_03113_));
 INVx1_ASAP7_75t_R _14730_ (.A(_01787_),
    .Y(_10600_));
 OR3x1_ASAP7_75t_R _14731_ (.A(_10565_),
    .B(_10576_),
    .C(_10578_),
    .Y(_10601_));
 OA211x2_ASAP7_75t_R _14732_ (.A1(_10600_),
    .A2(_10553_),
    .B(_10601_),
    .C(_09830_),
    .Y(_03114_));
 OR3x1_ASAP7_75t_R _14733_ (.A(_02136_),
    .B(_10577_),
    .C(_10579_),
    .Y(_10602_));
 OR2x2_ASAP7_75t_R _14734_ (.A(_01786_),
    .B(_10552_),
    .Y(_10603_));
 AOI21x1_ASAP7_75t_R _14735_ (.A1(_10602_),
    .A2(_10603_),
    .B(_10530_),
    .Y(_03115_));
 AO22x1_ASAP7_75t_R _14736_ (.A1(_10563_),
    .A2(_10535_),
    .B1(_10567_),
    .B2(_10572_),
    .Y(_10604_));
 AND3x1_ASAP7_75t_R _14737_ (.A(_09632_),
    .B(_10541_),
    .C(_10604_),
    .Y(_03116_));
 NOR2x1_ASAP7_75t_R _14738_ (.A(_10574_),
    .B(_10551_),
    .Y(_10605_));
 AOI21x1_ASAP7_75t_R _14739_ (.A1(_10575_),
    .A2(_10605_),
    .B(_10530_),
    .Y(_03117_));
 NOR2x1_ASAP7_75t_R _14740_ (.A(_01783_),
    .B(_10553_),
    .Y(_10606_));
 OA21x2_ASAP7_75t_R _14741_ (.A1(_10574_),
    .A2(_10575_),
    .B(_02133_),
    .Y(_10607_));
 AOI211x1_ASAP7_75t_R _14742_ (.A1(_02091_),
    .A2(_10577_),
    .B(_10579_),
    .C(_10607_),
    .Y(_10608_));
 OA21x2_ASAP7_75t_R _14743_ (.A1(_10606_),
    .A2(_10608_),
    .B(_10521_),
    .Y(_03118_));
 NOR2x1_ASAP7_75t_R _14744_ (.A(_01782_),
    .B(_10553_),
    .Y(_10609_));
 OA21x2_ASAP7_75t_R _14745_ (.A1(_10574_),
    .A2(_10575_),
    .B(_02132_),
    .Y(_10610_));
 AOI211x1_ASAP7_75t_R _14746_ (.A1(_02090_),
    .A2(_10577_),
    .B(_10579_),
    .C(_10610_),
    .Y(_10611_));
 OA21x2_ASAP7_75t_R _14747_ (.A1(_10609_),
    .A2(_10611_),
    .B(_10521_),
    .Y(_03119_));
 OA22x2_ASAP7_75t_R _14748_ (.A1(_10568_),
    .A2(_10548_),
    .B1(_10546_),
    .B2(_10541_),
    .Y(_10612_));
 AO32x2_ASAP7_75t_R _14749_ (.A1(_10569_),
    .A2(_10531_),
    .A3(_10612_),
    .B1(_10550_),
    .B2(_10549_),
    .Y(_10613_));
 AO21x2_ASAP7_75t_R _14750_ (.A1(_10572_),
    .A2(_10541_),
    .B(_10548_),
    .Y(_10614_));
 AND3x1_ASAP7_75t_R _14751_ (.A(_10539_),
    .B(_10536_),
    .C(_10569_),
    .Y(_10615_));
 NAND3x1_ASAP7_75t_R _14752_ (.A(_10613_),
    .B(_10614_),
    .C(_10615_),
    .Y(_10616_));
 BUFx12f_ASAP7_75t_R _14753_ (.A(_10616_),
    .Y(_10617_));
 NOR2x1_ASAP7_75t_R _14754_ (.A(_01795_),
    .B(_10617_),
    .Y(_10618_));
 AND4x1_ASAP7_75t_R _14755_ (.A(_02135_),
    .B(_02136_),
    .C(_10565_),
    .D(_02138_),
    .Y(_10619_));
 OR2x2_ASAP7_75t_R _14756_ (.A(_10538_),
    .B(_01789_),
    .Y(_10620_));
 NAND2x1_ASAP7_75t_R _14757_ (.A(_10534_),
    .B(_10620_),
    .Y(_10621_));
 OAI21x1_ASAP7_75t_R _14758_ (.A1(_10619_),
    .A2(_10621_),
    .B(_10536_),
    .Y(_10622_));
 NAND2x1_ASAP7_75t_R _14759_ (.A(_00010_),
    .B(_10534_),
    .Y(_10623_));
 OAI21x1_ASAP7_75t_R _14760_ (.A1(_10566_),
    .A2(_10623_),
    .B(_10538_),
    .Y(_10624_));
 INVx1_ASAP7_75t_R _14761_ (.A(_10546_),
    .Y(_10625_));
 AO32x2_ASAP7_75t_R _14762_ (.A1(_10568_),
    .A2(_10622_),
    .A3(_10624_),
    .B1(_10625_),
    .B2(_10543_),
    .Y(_10626_));
 NOR2x1_ASAP7_75t_R _14763_ (.A(_10571_),
    .B(_10626_),
    .Y(_10627_));
 BUFx6f_ASAP7_75t_R _14764_ (.A(_10627_),
    .Y(_10628_));
 AND3x2_ASAP7_75t_R _14765_ (.A(_10613_),
    .B(_10614_),
    .C(_10615_),
    .Y(_10629_));
 BUFx6f_ASAP7_75t_R _14766_ (.A(_10629_),
    .Y(_10630_));
 BUFx6f_ASAP7_75t_R _14767_ (.A(_10571_),
    .Y(_10631_));
 BUFx6f_ASAP7_75t_R _14768_ (.A(_10626_),
    .Y(_10632_));
 OA21x2_ASAP7_75t_R _14769_ (.A1(_10631_),
    .A2(_10632_),
    .B(_02103_),
    .Y(_10633_));
 AOI211x1_ASAP7_75t_R _14770_ (.A1(_02145_),
    .A2(_10628_),
    .B(_10630_),
    .C(_10633_),
    .Y(_10634_));
 OA21x2_ASAP7_75t_R _14771_ (.A1(_10618_),
    .A2(_10634_),
    .B(_10521_),
    .Y(_03120_));
 NOR2x1_ASAP7_75t_R _14772_ (.A(_01794_),
    .B(_10617_),
    .Y(_10635_));
 OA21x2_ASAP7_75t_R _14773_ (.A1(_10631_),
    .A2(_10632_),
    .B(_02102_),
    .Y(_10636_));
 AOI211x1_ASAP7_75t_R _14774_ (.A1(_02144_),
    .A2(_10628_),
    .B(_10630_),
    .C(_10636_),
    .Y(_10637_));
 BUFx6f_ASAP7_75t_R _14775_ (.A(_09229_),
    .Y(_10638_));
 OA21x2_ASAP7_75t_R _14776_ (.A1(_10635_),
    .A2(_10637_),
    .B(_10638_),
    .Y(_03121_));
 NOR2x1_ASAP7_75t_R _14777_ (.A(_01793_),
    .B(_10617_),
    .Y(_10639_));
 OA21x2_ASAP7_75t_R _14778_ (.A1(_10631_),
    .A2(_10632_),
    .B(_02101_),
    .Y(_10640_));
 AOI211x1_ASAP7_75t_R _14779_ (.A1(_02143_),
    .A2(_10628_),
    .B(_10630_),
    .C(_10640_),
    .Y(_10641_));
 OA21x2_ASAP7_75t_R _14780_ (.A1(_10639_),
    .A2(_10641_),
    .B(_10638_),
    .Y(_03122_));
 NOR2x1_ASAP7_75t_R _14781_ (.A(_01792_),
    .B(_10617_),
    .Y(_10642_));
 OA21x2_ASAP7_75t_R _14782_ (.A1(_10631_),
    .A2(_10632_),
    .B(_02100_),
    .Y(_10643_));
 AOI211x1_ASAP7_75t_R _14783_ (.A1(_02142_),
    .A2(_10628_),
    .B(_10630_),
    .C(_10643_),
    .Y(_10644_));
 OA21x2_ASAP7_75t_R _14784_ (.A1(_10642_),
    .A2(_10644_),
    .B(_10638_),
    .Y(_03123_));
 NOR2x1_ASAP7_75t_R _14785_ (.A(_01791_),
    .B(_10617_),
    .Y(_10645_));
 OA21x2_ASAP7_75t_R _14786_ (.A1(_10631_),
    .A2(_10632_),
    .B(_02099_),
    .Y(_10646_));
 AOI211x1_ASAP7_75t_R _14787_ (.A1(_02141_),
    .A2(_10628_),
    .B(_10630_),
    .C(_10646_),
    .Y(_10647_));
 OA21x2_ASAP7_75t_R _14788_ (.A1(_10645_),
    .A2(_10647_),
    .B(_10638_),
    .Y(_03124_));
 NOR2x1_ASAP7_75t_R _14789_ (.A(_01790_),
    .B(_10617_),
    .Y(_10648_));
 OA21x2_ASAP7_75t_R _14790_ (.A1(_10631_),
    .A2(_10632_),
    .B(_02098_),
    .Y(_10649_));
 AOI211x1_ASAP7_75t_R _14791_ (.A1(_02140_),
    .A2(_10628_),
    .B(_10630_),
    .C(_10649_),
    .Y(_10650_));
 OA21x2_ASAP7_75t_R _14792_ (.A1(_10648_),
    .A2(_10650_),
    .B(_10638_),
    .Y(_03125_));
 OA21x2_ASAP7_75t_R _14793_ (.A1(_10631_),
    .A2(_10632_),
    .B(_02097_),
    .Y(_10651_));
 AO21x1_ASAP7_75t_R _14794_ (.A1(_02139_),
    .A2(_10628_),
    .B(_10651_),
    .Y(_10652_));
 AOI21x1_ASAP7_75t_R _14795_ (.A1(_10617_),
    .A2(_10652_),
    .B(_10530_),
    .Y(_03126_));
 NOR2x1_ASAP7_75t_R _14796_ (.A(_01788_),
    .B(_10617_),
    .Y(_10653_));
 OA21x2_ASAP7_75t_R _14797_ (.A1(_10631_),
    .A2(_10632_),
    .B(_02096_),
    .Y(_10654_));
 AOI211x1_ASAP7_75t_R _14798_ (.A1(_02138_),
    .A2(_10628_),
    .B(_10630_),
    .C(_10654_),
    .Y(_10655_));
 OA21x2_ASAP7_75t_R _14799_ (.A1(_10653_),
    .A2(_10655_),
    .B(_10638_),
    .Y(_03127_));
 NOR2x1_ASAP7_75t_R _14800_ (.A(_01787_),
    .B(_10617_),
    .Y(_10656_));
 OA21x2_ASAP7_75t_R _14801_ (.A1(_10631_),
    .A2(_10632_),
    .B(_02095_),
    .Y(_10657_));
 AOI211x1_ASAP7_75t_R _14802_ (.A1(_02137_),
    .A2(_10628_),
    .B(_10630_),
    .C(_10657_),
    .Y(_10658_));
 OA21x2_ASAP7_75t_R _14803_ (.A1(_10656_),
    .A2(_10658_),
    .B(_10638_),
    .Y(_03128_));
 NOR2x1_ASAP7_75t_R _14804_ (.A(_01786_),
    .B(_10617_),
    .Y(_10659_));
 OA21x2_ASAP7_75t_R _14805_ (.A1(_10631_),
    .A2(_10626_),
    .B(_02094_),
    .Y(_10660_));
 AOI211x1_ASAP7_75t_R _14806_ (.A1(_02136_),
    .A2(_10628_),
    .B(_10630_),
    .C(_10660_),
    .Y(_10661_));
 OA21x2_ASAP7_75t_R _14807_ (.A1(_10659_),
    .A2(_10661_),
    .B(_10638_),
    .Y(_03129_));
 AND3x1_ASAP7_75t_R _14808_ (.A(_09632_),
    .B(_10531_),
    .C(_10632_),
    .Y(_03130_));
 AOI21x1_ASAP7_75t_R _14809_ (.A1(_10536_),
    .A2(_10613_),
    .B(_10538_),
    .Y(_10662_));
 OA211x2_ASAP7_75t_R _14810_ (.A1(_10620_),
    .A2(_10662_),
    .B(_10614_),
    .C(_10627_),
    .Y(_10663_));
 NOR2x1_ASAP7_75t_R _14811_ (.A(_10013_),
    .B(_10663_),
    .Y(_03131_));
 NOR2x1_ASAP7_75t_R _14812_ (.A(_01783_),
    .B(_10616_),
    .Y(_10664_));
 OA21x2_ASAP7_75t_R _14813_ (.A1(_10571_),
    .A2(_10626_),
    .B(_02091_),
    .Y(_10665_));
 AOI211x1_ASAP7_75t_R _14814_ (.A1(_02133_),
    .A2(_10627_),
    .B(_10630_),
    .C(_10665_),
    .Y(_10666_));
 OA21x2_ASAP7_75t_R _14815_ (.A1(_10664_),
    .A2(_10666_),
    .B(_10638_),
    .Y(_03132_));
 NOR2x1_ASAP7_75t_R _14816_ (.A(_01782_),
    .B(_10616_),
    .Y(_10667_));
 OA21x2_ASAP7_75t_R _14817_ (.A1(_10571_),
    .A2(_10626_),
    .B(_02090_),
    .Y(_10668_));
 AOI211x1_ASAP7_75t_R _14818_ (.A1(_02132_),
    .A2(_10627_),
    .B(_10629_),
    .C(_10668_),
    .Y(_10669_));
 OA21x2_ASAP7_75t_R _14819_ (.A1(_10667_),
    .A2(_10669_),
    .B(_10638_),
    .Y(_03133_));
 AO21x2_ASAP7_75t_R _14820_ (.A1(_10536_),
    .A2(_10613_),
    .B(_10538_),
    .Y(_10670_));
 BUFx6f_ASAP7_75t_R _14821_ (.A(_10670_),
    .Y(_10671_));
 NOR2x1_ASAP7_75t_R _14822_ (.A(_01795_),
    .B(_10671_),
    .Y(_10672_));
 OR2x2_ASAP7_75t_R _14823_ (.A(_02134_),
    .B(_10566_),
    .Y(_10673_));
 AO21x2_ASAP7_75t_R _14824_ (.A1(_02135_),
    .A2(_10563_),
    .B(_10673_),
    .Y(_10674_));
 OA21x2_ASAP7_75t_R _14825_ (.A1(_10619_),
    .A2(_10621_),
    .B(_10536_),
    .Y(_10675_));
 OA21x2_ASAP7_75t_R _14826_ (.A1(_10566_),
    .A2(_10623_),
    .B(_10538_),
    .Y(_10676_));
 OA31x2_ASAP7_75t_R _14827_ (.A1(_10571_),
    .A2(_10675_),
    .A3(_10676_),
    .B1(_10568_),
    .Y(_10677_));
 NAND2x1_ASAP7_75t_R _14828_ (.A(_10674_),
    .B(_10677_),
    .Y(_10678_));
 BUFx6f_ASAP7_75t_R _14829_ (.A(_10678_),
    .Y(_10679_));
 BUFx6f_ASAP7_75t_R _14830_ (.A(_10674_),
    .Y(_10680_));
 BUFx6f_ASAP7_75t_R _14831_ (.A(_10677_),
    .Y(_10681_));
 AND3x1_ASAP7_75t_R _14832_ (.A(_02103_),
    .B(_10680_),
    .C(_10681_),
    .Y(_10682_));
 AOI211x1_ASAP7_75t_R _14833_ (.A1(_02145_),
    .A2(_10679_),
    .B(_10682_),
    .C(_10662_),
    .Y(_10683_));
 BUFx6f_ASAP7_75t_R _14834_ (.A(_09229_),
    .Y(_10684_));
 OA21x2_ASAP7_75t_R _14835_ (.A1(_10672_),
    .A2(_10683_),
    .B(_10684_),
    .Y(_03134_));
 NOR2x1_ASAP7_75t_R _14836_ (.A(_01794_),
    .B(_10671_),
    .Y(_10685_));
 AND3x1_ASAP7_75t_R _14837_ (.A(_02102_),
    .B(_10680_),
    .C(_10681_),
    .Y(_10686_));
 AOI211x1_ASAP7_75t_R _14838_ (.A1(_02144_),
    .A2(_10679_),
    .B(_10686_),
    .C(_10662_),
    .Y(_10687_));
 OA21x2_ASAP7_75t_R _14839_ (.A1(_10685_),
    .A2(_10687_),
    .B(_10684_),
    .Y(_03135_));
 NOR2x1_ASAP7_75t_R _14840_ (.A(_01793_),
    .B(_10671_),
    .Y(_10688_));
 AND3x1_ASAP7_75t_R _14841_ (.A(_02101_),
    .B(_10680_),
    .C(_10681_),
    .Y(_10689_));
 AOI211x1_ASAP7_75t_R _14842_ (.A1(_02143_),
    .A2(_10679_),
    .B(_10689_),
    .C(_10662_),
    .Y(_10690_));
 OA21x2_ASAP7_75t_R _14843_ (.A1(_10688_),
    .A2(_10690_),
    .B(_10684_),
    .Y(_03136_));
 NOR2x1_ASAP7_75t_R _14844_ (.A(_01792_),
    .B(_10671_),
    .Y(_10691_));
 AND3x1_ASAP7_75t_R _14845_ (.A(_02100_),
    .B(_10680_),
    .C(_10681_),
    .Y(_10692_));
 AOI211x1_ASAP7_75t_R _14846_ (.A1(_02142_),
    .A2(_10679_),
    .B(_10692_),
    .C(_10662_),
    .Y(_10693_));
 OA21x2_ASAP7_75t_R _14847_ (.A1(_10691_),
    .A2(_10693_),
    .B(_10684_),
    .Y(_03137_));
 NOR2x1_ASAP7_75t_R _14848_ (.A(_01791_),
    .B(_10671_),
    .Y(_10694_));
 AND3x1_ASAP7_75t_R _14849_ (.A(_02099_),
    .B(_10680_),
    .C(_10681_),
    .Y(_10695_));
 AOI211x1_ASAP7_75t_R _14850_ (.A1(_02141_),
    .A2(_10679_),
    .B(_10695_),
    .C(_10662_),
    .Y(_10696_));
 OA21x2_ASAP7_75t_R _14851_ (.A1(_10694_),
    .A2(_10696_),
    .B(_10684_),
    .Y(_03138_));
 NOR2x1_ASAP7_75t_R _14852_ (.A(_01790_),
    .B(_10671_),
    .Y(_10697_));
 AND3x1_ASAP7_75t_R _14853_ (.A(_02098_),
    .B(_10680_),
    .C(_10681_),
    .Y(_10698_));
 AOI211x1_ASAP7_75t_R _14854_ (.A1(_02140_),
    .A2(_10679_),
    .B(_10698_),
    .C(_10662_),
    .Y(_10699_));
 OA21x2_ASAP7_75t_R _14855_ (.A1(_10697_),
    .A2(_10699_),
    .B(_10684_),
    .Y(_03139_));
 AND2x2_ASAP7_75t_R _14856_ (.A(_10569_),
    .B(_10662_),
    .Y(_10700_));
 AO21x1_ASAP7_75t_R _14857_ (.A1(_10680_),
    .A2(_10681_),
    .B(_10564_),
    .Y(_10701_));
 OA211x2_ASAP7_75t_R _14858_ (.A1(_10544_),
    .A2(_10679_),
    .B(_10701_),
    .C(_10670_),
    .Y(_10702_));
 OA21x2_ASAP7_75t_R _14859_ (.A1(_10700_),
    .A2(_10702_),
    .B(_10684_),
    .Y(_03140_));
 NOR2x1_ASAP7_75t_R _14860_ (.A(_01788_),
    .B(_10671_),
    .Y(_10703_));
 INVx1_ASAP7_75t_R _14861_ (.A(_02096_),
    .Y(_10704_));
 AO21x1_ASAP7_75t_R _14862_ (.A1(_10674_),
    .A2(_10677_),
    .B(_10533_),
    .Y(_10705_));
 OA211x2_ASAP7_75t_R _14863_ (.A1(_10704_),
    .A2(_10679_),
    .B(_10705_),
    .C(_10670_),
    .Y(_10706_));
 OA21x2_ASAP7_75t_R _14864_ (.A1(_10703_),
    .A2(_10706_),
    .B(_10684_),
    .Y(_03141_));
 NOR2x1_ASAP7_75t_R _14865_ (.A(_01787_),
    .B(_10671_),
    .Y(_10707_));
 INVx1_ASAP7_75t_R _14866_ (.A(_02095_),
    .Y(_10708_));
 AO21x1_ASAP7_75t_R _14867_ (.A1(_10674_),
    .A2(_10677_),
    .B(_10565_),
    .Y(_10709_));
 OA211x2_ASAP7_75t_R _14868_ (.A1(_10708_),
    .A2(_10678_),
    .B(_10709_),
    .C(_10670_),
    .Y(_10710_));
 OA21x2_ASAP7_75t_R _14869_ (.A1(_10707_),
    .A2(_10710_),
    .B(_10684_),
    .Y(_03142_));
 NOR2x1_ASAP7_75t_R _14870_ (.A(_01786_),
    .B(_10671_),
    .Y(_10711_));
 INVx1_ASAP7_75t_R _14871_ (.A(_02094_),
    .Y(_10712_));
 AO21x1_ASAP7_75t_R _14872_ (.A1(_10674_),
    .A2(_10677_),
    .B(_10532_),
    .Y(_10713_));
 OA211x2_ASAP7_75t_R _14873_ (.A1(_10712_),
    .A2(_10678_),
    .B(_10713_),
    .C(_10670_),
    .Y(_10714_));
 OA21x2_ASAP7_75t_R _14874_ (.A1(_10711_),
    .A2(_10714_),
    .B(_10684_),
    .Y(_03143_));
 OR4x1_ASAP7_75t_R _14875_ (.A(_08712_),
    .B(_10538_),
    .C(_10537_),
    .D(_10613_),
    .Y(_10715_));
 INVx1_ASAP7_75t_R _14876_ (.A(_10715_),
    .Y(_03144_));
 BUFx12f_ASAP7_75t_R _14877_ (.A(_10012_),
    .Y(_10716_));
 INVx1_ASAP7_75t_R _14878_ (.A(_10681_),
    .Y(_10717_));
 AND3x1_ASAP7_75t_R _14879_ (.A(_10670_),
    .B(_10680_),
    .C(_10717_),
    .Y(_10718_));
 NOR2x1_ASAP7_75t_R _14880_ (.A(_10716_),
    .B(_10718_),
    .Y(_03145_));
 NOR2x1_ASAP7_75t_R _14881_ (.A(_01783_),
    .B(_10671_),
    .Y(_10719_));
 AND3x1_ASAP7_75t_R _14882_ (.A(_02091_),
    .B(_10680_),
    .C(_10681_),
    .Y(_10720_));
 AOI211x1_ASAP7_75t_R _14883_ (.A1(_02133_),
    .A2(_10679_),
    .B(_10720_),
    .C(_10662_),
    .Y(_10721_));
 BUFx6f_ASAP7_75t_R _14884_ (.A(_09229_),
    .Y(_10722_));
 OA21x2_ASAP7_75t_R _14885_ (.A1(_10719_),
    .A2(_10721_),
    .B(_10722_),
    .Y(_03146_));
 NOR2x1_ASAP7_75t_R _14886_ (.A(_01782_),
    .B(_10670_),
    .Y(_10723_));
 AND3x1_ASAP7_75t_R _14887_ (.A(_02090_),
    .B(_10680_),
    .C(_10681_),
    .Y(_10724_));
 AOI211x1_ASAP7_75t_R _14888_ (.A1(_02132_),
    .A2(_10679_),
    .B(_10724_),
    .C(_10662_),
    .Y(_10725_));
 OA21x2_ASAP7_75t_R _14889_ (.A1(_10723_),
    .A2(_10725_),
    .B(_10722_),
    .Y(_03147_));
 AND2x2_ASAP7_75t_R _14890_ (.A(_09957_),
    .B(_00011_),
    .Y(_03148_));
 BUFx6f_ASAP7_75t_R _14891_ (.A(_02008_),
    .Y(_10726_));
 NOR2x1_ASAP7_75t_R _14892_ (.A(_10726_),
    .B(_02009_),
    .Y(_10727_));
 NOR2x1_ASAP7_75t_R _14893_ (.A(_02053_),
    .B(_02054_),
    .Y(_10728_));
 AO21x1_ASAP7_75t_R _14894_ (.A1(_02052_),
    .A2(_10728_),
    .B(_02050_),
    .Y(_10729_));
 BUFx6f_ASAP7_75t_R _14895_ (.A(_10729_),
    .Y(_10730_));
 BUFx6f_ASAP7_75t_R _14896_ (.A(_01771_),
    .Y(_10731_));
 BUFx6f_ASAP7_75t_R _14897_ (.A(_01775_),
    .Y(_10732_));
 INVx2_ASAP7_75t_R _14898_ (.A(_10732_),
    .Y(_10733_));
 BUFx6f_ASAP7_75t_R _14899_ (.A(_01770_),
    .Y(_10734_));
 AO21x1_ASAP7_75t_R _14900_ (.A1(_10731_),
    .A2(_10733_),
    .B(_10734_),
    .Y(_10735_));
 OR2x6_ASAP7_75t_R _14901_ (.A(_02050_),
    .B(_02051_),
    .Y(_10736_));
 OA21x2_ASAP7_75t_R _14902_ (.A1(_10730_),
    .A2(_10735_),
    .B(_10736_),
    .Y(_10737_));
 INVx1_ASAP7_75t_R _14903_ (.A(_10726_),
    .Y(_10738_));
 BUFx6f_ASAP7_75t_R _14904_ (.A(_02010_),
    .Y(_10739_));
 NOR2x2_ASAP7_75t_R _14905_ (.A(_02011_),
    .B(_02012_),
    .Y(_10740_));
 AND4x1_ASAP7_75t_R _14906_ (.A(_10738_),
    .B(_10739_),
    .C(_02013_),
    .D(_10740_),
    .Y(_10741_));
 OA21x2_ASAP7_75t_R _14907_ (.A1(_10727_),
    .A2(_10737_),
    .B(_10741_),
    .Y(_10742_));
 INVx2_ASAP7_75t_R _14908_ (.A(_10734_),
    .Y(_10743_));
 AND2x2_ASAP7_75t_R _14909_ (.A(_02009_),
    .B(_10739_),
    .Y(_10744_));
 AO221x1_ASAP7_75t_R _14910_ (.A1(_10743_),
    .A2(_10732_),
    .B1(_10740_),
    .B2(_10744_),
    .C(_10726_),
    .Y(_10745_));
 AND2x2_ASAP7_75t_R _14911_ (.A(_10734_),
    .B(_10739_),
    .Y(_10746_));
 OA21x2_ASAP7_75t_R _14912_ (.A1(_00011_),
    .A2(_10726_),
    .B(_10734_),
    .Y(_10747_));
 AO21x1_ASAP7_75t_R _14913_ (.A1(_10740_),
    .A2(_10746_),
    .B(_10747_),
    .Y(_10748_));
 AO21x1_ASAP7_75t_R _14914_ (.A1(_10731_),
    .A2(_10745_),
    .B(_10748_),
    .Y(_10749_));
 OR2x6_ASAP7_75t_R _14915_ (.A(_10726_),
    .B(_02009_),
    .Y(_10750_));
 OR2x2_ASAP7_75t_R _14916_ (.A(_10734_),
    .B(_10726_),
    .Y(_10751_));
 AO221x1_ASAP7_75t_R _14917_ (.A1(_10731_),
    .A2(_10732_),
    .B1(_10739_),
    .B2(_10740_),
    .C(_10751_),
    .Y(_10752_));
 INVx1_ASAP7_75t_R _14918_ (.A(_02052_),
    .Y(_10753_));
 OR5x1_ASAP7_75t_R _14919_ (.A(_02050_),
    .B(_10753_),
    .C(_02053_),
    .D(_02054_),
    .E(_02055_),
    .Y(_10754_));
 AO21x2_ASAP7_75t_R _14920_ (.A1(_10750_),
    .A2(_10752_),
    .B(_10754_),
    .Y(_10755_));
 OA211x2_ASAP7_75t_R _14921_ (.A1(_10730_),
    .A2(_10749_),
    .B(_10755_),
    .C(_10736_),
    .Y(_10756_));
 BUFx6f_ASAP7_75t_R _14922_ (.A(_10756_),
    .Y(_10757_));
 AND2x4_ASAP7_75t_R _14923_ (.A(_10742_),
    .B(_10757_),
    .Y(_10758_));
 BUFx6f_ASAP7_75t_R _14924_ (.A(_10758_),
    .Y(_10759_));
 NAND2x1_ASAP7_75t_R _14925_ (.A(_02019_),
    .B(_10759_),
    .Y(_10760_));
 INVx2_ASAP7_75t_R _14926_ (.A(_02061_),
    .Y(_10761_));
 AO21x1_ASAP7_75t_R _14927_ (.A1(_10742_),
    .A2(_10757_),
    .B(_10761_),
    .Y(_10762_));
 BUFx12f_ASAP7_75t_R _14928_ (.A(_08571_),
    .Y(_10763_));
 AND2x4_ASAP7_75t_R _14929_ (.A(_10743_),
    .B(_10731_),
    .Y(_10764_));
 OAI21x1_ASAP7_75t_R _14930_ (.A1(_10730_),
    .A2(_10735_),
    .B(_10736_),
    .Y(_10765_));
 INVx1_ASAP7_75t_R _14931_ (.A(_10741_),
    .Y(_10766_));
 AO21x2_ASAP7_75t_R _14932_ (.A1(_10750_),
    .A2(_10765_),
    .B(_10766_),
    .Y(_10767_));
 NAND2x1_ASAP7_75t_R _14933_ (.A(_10733_),
    .B(_10750_),
    .Y(_10768_));
 NOR2x1_ASAP7_75t_R _14934_ (.A(_02050_),
    .B(_02051_),
    .Y(_10769_));
 OR3x1_ASAP7_75t_R _14935_ (.A(_10732_),
    .B(_10727_),
    .C(_10769_),
    .Y(_10770_));
 INVx1_ASAP7_75t_R _14936_ (.A(_02050_),
    .Y(_10771_));
 INVx1_ASAP7_75t_R _14937_ (.A(_02055_),
    .Y(_10772_));
 AND4x1_ASAP7_75t_R _14938_ (.A(_10771_),
    .B(_02052_),
    .C(_10772_),
    .D(_10728_),
    .Y(_10773_));
 OA22x2_ASAP7_75t_R _14939_ (.A1(_10741_),
    .A2(_10768_),
    .B1(_10770_),
    .B2(_10773_),
    .Y(_10774_));
 NAND2x1_ASAP7_75t_R _14940_ (.A(_10732_),
    .B(_10736_),
    .Y(_10775_));
 AO21x1_ASAP7_75t_R _14941_ (.A1(_10741_),
    .A2(_10730_),
    .B(_10775_),
    .Y(_10776_));
 AO21x1_ASAP7_75t_R _14942_ (.A1(_10739_),
    .A2(_10740_),
    .B(_10726_),
    .Y(_10777_));
 NAND2x1_ASAP7_75t_R _14943_ (.A(_10732_),
    .B(_10750_),
    .Y(_10778_));
 OA211x2_ASAP7_75t_R _14944_ (.A1(_10732_),
    .A2(_10777_),
    .B(_10773_),
    .C(_10778_),
    .Y(_10779_));
 AOI21x1_ASAP7_75t_R _14945_ (.A1(_10774_),
    .A2(_10776_),
    .B(_10779_),
    .Y(_10780_));
 AND5x2_ASAP7_75t_R _14946_ (.A(_10732_),
    .B(_10764_),
    .C(_10767_),
    .D(_10756_),
    .E(_10780_),
    .Y(_10781_));
 NOR2x2_ASAP7_75t_R _14947_ (.A(_10763_),
    .B(_10781_),
    .Y(_10782_));
 NOR2x1_ASAP7_75t_R _14948_ (.A(_09221_),
    .B(_01781_),
    .Y(_10783_));
 BUFx6f_ASAP7_75t_R _14949_ (.A(_10781_),
    .Y(_10784_));
 AO32x1_ASAP7_75t_R _14950_ (.A1(_10760_),
    .A2(_10762_),
    .A3(_10782_),
    .B1(_10783_),
    .B2(_10784_),
    .Y(_03149_));
 NAND2x1_ASAP7_75t_R _14951_ (.A(_02018_),
    .B(_10759_),
    .Y(_10785_));
 INVx2_ASAP7_75t_R _14952_ (.A(_02060_),
    .Y(_10786_));
 AO21x1_ASAP7_75t_R _14953_ (.A1(_10742_),
    .A2(_10757_),
    .B(_10786_),
    .Y(_10787_));
 NOR2x1_ASAP7_75t_R _14954_ (.A(_09221_),
    .B(_01780_),
    .Y(_10788_));
 AO32x1_ASAP7_75t_R _14955_ (.A1(_10782_),
    .A2(_10785_),
    .A3(_10787_),
    .B1(_10788_),
    .B2(_10784_),
    .Y(_03150_));
 NAND2x1_ASAP7_75t_R _14956_ (.A(_02017_),
    .B(_10759_),
    .Y(_10789_));
 INVx2_ASAP7_75t_R _14957_ (.A(_02059_),
    .Y(_10790_));
 AO21x1_ASAP7_75t_R _14958_ (.A1(_10742_),
    .A2(_10757_),
    .B(_10790_),
    .Y(_10791_));
 NOR2x1_ASAP7_75t_R _14959_ (.A(_09221_),
    .B(_01779_),
    .Y(_10792_));
 AO32x1_ASAP7_75t_R _14960_ (.A1(_10782_),
    .A2(_10789_),
    .A3(_10791_),
    .B1(_10792_),
    .B2(_10784_),
    .Y(_03151_));
 NAND2x1_ASAP7_75t_R _14961_ (.A(_02016_),
    .B(_10759_),
    .Y(_10793_));
 INVx2_ASAP7_75t_R _14962_ (.A(_02058_),
    .Y(_10794_));
 AO21x1_ASAP7_75t_R _14963_ (.A1(_10742_),
    .A2(_10757_),
    .B(_10794_),
    .Y(_10795_));
 NOR2x1_ASAP7_75t_R _14964_ (.A(_09221_),
    .B(_01778_),
    .Y(_10796_));
 AO32x1_ASAP7_75t_R _14965_ (.A1(_10782_),
    .A2(_10793_),
    .A3(_10795_),
    .B1(_10796_),
    .B2(_10784_),
    .Y(_03152_));
 NAND2x1_ASAP7_75t_R _14966_ (.A(_02015_),
    .B(_10759_),
    .Y(_10797_));
 INVx2_ASAP7_75t_R _14967_ (.A(_02057_),
    .Y(_10798_));
 AO21x1_ASAP7_75t_R _14968_ (.A1(_10742_),
    .A2(_10757_),
    .B(_10798_),
    .Y(_10799_));
 NOR2x1_ASAP7_75t_R _14969_ (.A(_09221_),
    .B(_01777_),
    .Y(_10800_));
 AO32x1_ASAP7_75t_R _14970_ (.A1(_10782_),
    .A2(_10797_),
    .A3(_10799_),
    .B1(_10800_),
    .B2(_10784_),
    .Y(_03153_));
 NAND2x1_ASAP7_75t_R _14971_ (.A(_02014_),
    .B(_10759_),
    .Y(_10801_));
 INVx2_ASAP7_75t_R _14972_ (.A(_02056_),
    .Y(_10802_));
 AO21x1_ASAP7_75t_R _14973_ (.A1(_10742_),
    .A2(_10757_),
    .B(_10802_),
    .Y(_10803_));
 NOR2x1_ASAP7_75t_R _14974_ (.A(_09221_),
    .B(_01776_),
    .Y(_10804_));
 AO32x1_ASAP7_75t_R _14975_ (.A1(_10782_),
    .A2(_10801_),
    .A3(_10803_),
    .B1(_10804_),
    .B2(_10784_),
    .Y(_03154_));
 OR4x1_ASAP7_75t_R _14976_ (.A(_08712_),
    .B(_02055_),
    .C(_10781_),
    .D(_10759_),
    .Y(_10805_));
 INVx1_ASAP7_75t_R _14977_ (.A(_10805_),
    .Y(_03155_));
 NAND2x1_ASAP7_75t_R _14978_ (.A(_01774_),
    .B(_10784_),
    .Y(_10806_));
 INVx1_ASAP7_75t_R _14979_ (.A(_02054_),
    .Y(_10807_));
 OR3x1_ASAP7_75t_R _14980_ (.A(_10807_),
    .B(_10781_),
    .C(_10758_),
    .Y(_10808_));
 AND3x1_ASAP7_75t_R _14981_ (.A(_09632_),
    .B(_10806_),
    .C(_10808_),
    .Y(_03156_));
 BUFx6f_ASAP7_75t_R _14982_ (.A(_08581_),
    .Y(_10809_));
 NAND2x1_ASAP7_75t_R _14983_ (.A(_01773_),
    .B(_10781_),
    .Y(_10810_));
 INVx1_ASAP7_75t_R _14984_ (.A(_02053_),
    .Y(_10811_));
 OR3x1_ASAP7_75t_R _14985_ (.A(_10811_),
    .B(_10781_),
    .C(_10758_),
    .Y(_10812_));
 AND3x1_ASAP7_75t_R _14986_ (.A(_10809_),
    .B(_10810_),
    .C(_10812_),
    .Y(_03157_));
 INVx1_ASAP7_75t_R _14987_ (.A(_01772_),
    .Y(_10813_));
 NAND2x1_ASAP7_75t_R _14988_ (.A(_10813_),
    .B(_10784_),
    .Y(_10814_));
 OR3x1_ASAP7_75t_R _14989_ (.A(_02052_),
    .B(_10781_),
    .C(_10759_),
    .Y(_10815_));
 AOI21x1_ASAP7_75t_R _14990_ (.A1(_10814_),
    .A2(_10815_),
    .B(_10530_),
    .Y(_03158_));
 OAI21x1_ASAP7_75t_R _14991_ (.A1(_10730_),
    .A2(_10749_),
    .B(_10755_),
    .Y(_10816_));
 AND3x1_ASAP7_75t_R _14992_ (.A(_10809_),
    .B(_10736_),
    .C(_10816_),
    .Y(_03159_));
 NAND2x1_ASAP7_75t_R _14993_ (.A(_10767_),
    .B(_10757_),
    .Y(_10817_));
 AND3x1_ASAP7_75t_R _14994_ (.A(_10732_),
    .B(_10764_),
    .C(_10780_),
    .Y(_10818_));
 OA21x2_ASAP7_75t_R _14995_ (.A1(_10817_),
    .A2(_10818_),
    .B(_10722_),
    .Y(_03160_));
 NAND2x1_ASAP7_75t_R _14996_ (.A(_02007_),
    .B(_10759_),
    .Y(_10819_));
 INVx2_ASAP7_75t_R _14997_ (.A(_02049_),
    .Y(_10820_));
 AO21x1_ASAP7_75t_R _14998_ (.A1(_10742_),
    .A2(_10757_),
    .B(_10820_),
    .Y(_10821_));
 NOR2x1_ASAP7_75t_R _14999_ (.A(_09221_),
    .B(_01769_),
    .Y(_10822_));
 AO32x1_ASAP7_75t_R _15000_ (.A1(_10782_),
    .A2(_10819_),
    .A3(_10821_),
    .B1(_10822_),
    .B2(_10784_),
    .Y(_03161_));
 NAND2x1_ASAP7_75t_R _15001_ (.A(_02006_),
    .B(_10759_),
    .Y(_10823_));
 INVx2_ASAP7_75t_R _15002_ (.A(_02048_),
    .Y(_10824_));
 AO21x1_ASAP7_75t_R _15003_ (.A1(_10742_),
    .A2(_10757_),
    .B(_10824_),
    .Y(_10825_));
 BUFx12f_ASAP7_75t_R _15004_ (.A(_08571_),
    .Y(_10826_));
 NOR2x1_ASAP7_75t_R _15005_ (.A(_10826_),
    .B(_01768_),
    .Y(_10827_));
 AO32x1_ASAP7_75t_R _15006_ (.A1(_10782_),
    .A2(_10823_),
    .A3(_10825_),
    .B1(_10827_),
    .B2(_10784_),
    .Y(_03162_));
 OA211x2_ASAP7_75t_R _15007_ (.A1(_10733_),
    .A2(_02050_),
    .B(_10743_),
    .C(_10731_),
    .Y(_10828_));
 AND5x1_ASAP7_75t_R _15008_ (.A(_10743_),
    .B(_10731_),
    .C(_02051_),
    .D(_02052_),
    .E(_10728_),
    .Y(_10829_));
 INVx1_ASAP7_75t_R _15009_ (.A(_00011_),
    .Y(_10830_));
 AND2x2_ASAP7_75t_R _15010_ (.A(_10734_),
    .B(_02052_),
    .Y(_10831_));
 AND2x2_ASAP7_75t_R _15011_ (.A(_10734_),
    .B(_02050_),
    .Y(_10832_));
 AO221x1_ASAP7_75t_R _15012_ (.A1(_10734_),
    .A2(_10830_),
    .B1(_10728_),
    .B2(_10831_),
    .C(_10832_),
    .Y(_10833_));
 OR4x1_ASAP7_75t_R _15013_ (.A(_10777_),
    .B(_10828_),
    .C(_10829_),
    .D(_10833_),
    .Y(_10834_));
 OA211x2_ASAP7_75t_R _15014_ (.A1(_10766_),
    .A2(_10737_),
    .B(_10834_),
    .C(_10750_),
    .Y(_10835_));
 OAI21x1_ASAP7_75t_R _15015_ (.A1(_10769_),
    .A2(_10755_),
    .B(_10773_),
    .Y(_10836_));
 AND5x2_ASAP7_75t_R _15016_ (.A(_10733_),
    .B(_10764_),
    .C(_10780_),
    .D(_10835_),
    .E(_10836_),
    .Y(_10837_));
 BUFx6f_ASAP7_75t_R _15017_ (.A(_10837_),
    .Y(_10838_));
 BUFx6f_ASAP7_75t_R _15018_ (.A(_10835_),
    .Y(_10839_));
 BUFx12f_ASAP7_75t_R _15019_ (.A(_10839_),
    .Y(_10840_));
 NAND2x1_ASAP7_75t_R _15020_ (.A(_10761_),
    .B(_10840_),
    .Y(_10841_));
 OR2x2_ASAP7_75t_R _15021_ (.A(_02019_),
    .B(_10839_),
    .Y(_10842_));
 AOI211x1_ASAP7_75t_R _15022_ (.A1(_10841_),
    .A2(_10842_),
    .B(_10021_),
    .C(_10838_),
    .Y(_10843_));
 AO21x1_ASAP7_75t_R _15023_ (.A1(_10783_),
    .A2(_10838_),
    .B(_10843_),
    .Y(_03163_));
 NAND2x1_ASAP7_75t_R _15024_ (.A(_10786_),
    .B(_10840_),
    .Y(_10844_));
 OR2x2_ASAP7_75t_R _15025_ (.A(_02018_),
    .B(_10839_),
    .Y(_10845_));
 AOI211x1_ASAP7_75t_R _15026_ (.A1(_10844_),
    .A2(_10845_),
    .B(_10021_),
    .C(_10838_),
    .Y(_10846_));
 AO21x1_ASAP7_75t_R _15027_ (.A1(_10788_),
    .A2(_10838_),
    .B(_10846_),
    .Y(_03164_));
 NAND2x1_ASAP7_75t_R _15028_ (.A(_10790_),
    .B(_10840_),
    .Y(_10847_));
 OR2x2_ASAP7_75t_R _15029_ (.A(_02017_),
    .B(_10839_),
    .Y(_10848_));
 AOI211x1_ASAP7_75t_R _15030_ (.A1(_10847_),
    .A2(_10848_),
    .B(_10021_),
    .C(_10837_),
    .Y(_10849_));
 AO21x1_ASAP7_75t_R _15031_ (.A1(_10792_),
    .A2(_10838_),
    .B(_10849_),
    .Y(_03165_));
 NAND2x1_ASAP7_75t_R _15032_ (.A(_10794_),
    .B(_10840_),
    .Y(_10850_));
 OR2x2_ASAP7_75t_R _15033_ (.A(_02016_),
    .B(_10839_),
    .Y(_10851_));
 AOI211x1_ASAP7_75t_R _15034_ (.A1(_10850_),
    .A2(_10851_),
    .B(_10021_),
    .C(_10837_),
    .Y(_10852_));
 AO21x1_ASAP7_75t_R _15035_ (.A1(_10796_),
    .A2(_10838_),
    .B(_10852_),
    .Y(_03166_));
 NAND2x1_ASAP7_75t_R _15036_ (.A(_10798_),
    .B(_10840_),
    .Y(_10853_));
 OR2x2_ASAP7_75t_R _15037_ (.A(_02015_),
    .B(_10839_),
    .Y(_10854_));
 AOI211x1_ASAP7_75t_R _15038_ (.A1(_10853_),
    .A2(_10854_),
    .B(_10021_),
    .C(_10837_),
    .Y(_10855_));
 AO21x1_ASAP7_75t_R _15039_ (.A1(_10800_),
    .A2(_10838_),
    .B(_10855_),
    .Y(_03167_));
 NAND2x1_ASAP7_75t_R _15040_ (.A(_10802_),
    .B(_10840_),
    .Y(_10856_));
 OR2x2_ASAP7_75t_R _15041_ (.A(_02014_),
    .B(_10839_),
    .Y(_10857_));
 AOI211x1_ASAP7_75t_R _15042_ (.A1(_10856_),
    .A2(_10857_),
    .B(_10021_),
    .C(_10837_),
    .Y(_10858_));
 AO21x1_ASAP7_75t_R _15043_ (.A1(_10804_),
    .A2(_10838_),
    .B(_10858_),
    .Y(_03168_));
 AND3x1_ASAP7_75t_R _15044_ (.A(_10733_),
    .B(_10764_),
    .C(_10780_),
    .Y(_10859_));
 NAND3x1_ASAP7_75t_R _15045_ (.A(_10840_),
    .B(_10836_),
    .C(_10859_),
    .Y(_10860_));
 NOR2x1_ASAP7_75t_R _15046_ (.A(_10828_),
    .B(_10829_),
    .Y(_10861_));
 NOR2x1_ASAP7_75t_R _15047_ (.A(_10777_),
    .B(_10833_),
    .Y(_10862_));
 AO221x1_ASAP7_75t_R _15048_ (.A1(_10741_),
    .A2(_10765_),
    .B1(_10861_),
    .B2(_10862_),
    .C(_10727_),
    .Y(_10863_));
 BUFx3_ASAP7_75t_R _15049_ (.A(_10863_),
    .Y(_10864_));
 AND2x2_ASAP7_75t_R _15050_ (.A(_02055_),
    .B(_10839_),
    .Y(_10865_));
 AO21x1_ASAP7_75t_R _15051_ (.A1(_02013_),
    .A2(_10864_),
    .B(_10865_),
    .Y(_10866_));
 AOI21x1_ASAP7_75t_R _15052_ (.A1(_10860_),
    .A2(_10866_),
    .B(_10530_),
    .Y(_03169_));
 NAND2x1_ASAP7_75t_R _15053_ (.A(_02012_),
    .B(_10864_),
    .Y(_10867_));
 OA211x2_ASAP7_75t_R _15054_ (.A1(_10807_),
    .A2(_10864_),
    .B(_10867_),
    .C(_09058_),
    .Y(_10868_));
 NOR2x1_ASAP7_75t_R _15055_ (.A(_08641_),
    .B(_01774_),
    .Y(_10869_));
 AND2x2_ASAP7_75t_R _15056_ (.A(_10837_),
    .B(_10869_),
    .Y(_10870_));
 AO21x1_ASAP7_75t_R _15057_ (.A1(_10860_),
    .A2(_10868_),
    .B(_10870_),
    .Y(_03170_));
 NAND2x1_ASAP7_75t_R _15058_ (.A(_02011_),
    .B(_10864_),
    .Y(_10871_));
 OA211x2_ASAP7_75t_R _15059_ (.A1(_10811_),
    .A2(_10864_),
    .B(_10871_),
    .C(_09058_),
    .Y(_10872_));
 NOR2x1_ASAP7_75t_R _15060_ (.A(_08641_),
    .B(_01773_),
    .Y(_10873_));
 AND2x2_ASAP7_75t_R _15061_ (.A(_10837_),
    .B(_10873_),
    .Y(_10874_));
 AO21x1_ASAP7_75t_R _15062_ (.A1(_10860_),
    .A2(_10872_),
    .B(_10874_),
    .Y(_03171_));
 NAND2x1_ASAP7_75t_R _15063_ (.A(_10739_),
    .B(_10864_),
    .Y(_10875_));
 OA211x2_ASAP7_75t_R _15064_ (.A1(_10753_),
    .A2(_10864_),
    .B(_10875_),
    .C(_08584_),
    .Y(_10876_));
 NOR2x1_ASAP7_75t_R _15065_ (.A(_08641_),
    .B(_01772_),
    .Y(_10877_));
 AND2x2_ASAP7_75t_R _15066_ (.A(_10837_),
    .B(_10877_),
    .Y(_10878_));
 AO21x1_ASAP7_75t_R _15067_ (.A1(_10860_),
    .A2(_10876_),
    .B(_10878_),
    .Y(_03172_));
 OA21x2_ASAP7_75t_R _15068_ (.A1(_10766_),
    .A2(_10737_),
    .B(_10834_),
    .Y(_10879_));
 OR3x1_ASAP7_75t_R _15069_ (.A(_08642_),
    .B(_10727_),
    .C(_10879_),
    .Y(_10880_));
 INVx1_ASAP7_75t_R _15070_ (.A(_10880_),
    .Y(_03173_));
 NAND2x1_ASAP7_75t_R _15071_ (.A(_10840_),
    .B(_10836_),
    .Y(_10881_));
 OA21x2_ASAP7_75t_R _15072_ (.A1(_10881_),
    .A2(_10859_),
    .B(_10722_),
    .Y(_03174_));
 NAND2x1_ASAP7_75t_R _15073_ (.A(_10820_),
    .B(_10840_),
    .Y(_10882_));
 OR2x2_ASAP7_75t_R _15074_ (.A(_02007_),
    .B(_10839_),
    .Y(_10883_));
 AOI211x1_ASAP7_75t_R _15075_ (.A1(_10882_),
    .A2(_10883_),
    .B(_10021_),
    .C(_10837_),
    .Y(_10884_));
 AO21x1_ASAP7_75t_R _15076_ (.A1(_10822_),
    .A2(_10838_),
    .B(_10884_),
    .Y(_03175_));
 NAND2x1_ASAP7_75t_R _15077_ (.A(_10824_),
    .B(_10840_),
    .Y(_10885_));
 OR2x2_ASAP7_75t_R _15078_ (.A(_02006_),
    .B(_10839_),
    .Y(_10886_));
 AOI211x1_ASAP7_75t_R _15079_ (.A1(_10885_),
    .A2(_10886_),
    .B(_10021_),
    .C(_10837_),
    .Y(_10887_));
 AO21x1_ASAP7_75t_R _15080_ (.A1(_10827_),
    .A2(_10838_),
    .B(_10887_),
    .Y(_03176_));
 INVx1_ASAP7_75t_R _15081_ (.A(_02009_),
    .Y(_10888_));
 AOI211x1_ASAP7_75t_R _15082_ (.A1(_10731_),
    .A2(_10745_),
    .B(_10748_),
    .C(_10769_),
    .Y(_10889_));
 AOI21x1_ASAP7_75t_R _15083_ (.A1(_10739_),
    .A2(_10740_),
    .B(_10726_),
    .Y(_10890_));
 OA221x2_ASAP7_75t_R _15084_ (.A1(_10888_),
    .A2(_10834_),
    .B1(_10889_),
    .B2(_10730_),
    .C(_10890_),
    .Y(_10891_));
 BUFx6f_ASAP7_75t_R _15085_ (.A(_10891_),
    .Y(_10892_));
 NAND2x1_ASAP7_75t_R _15086_ (.A(_02019_),
    .B(_10892_),
    .Y(_10893_));
 BUFx6f_ASAP7_75t_R _15087_ (.A(_10891_),
    .Y(_10894_));
 OR2x2_ASAP7_75t_R _15088_ (.A(_10761_),
    .B(_10894_),
    .Y(_10895_));
 AOI21x1_ASAP7_75t_R _15089_ (.A1(_10731_),
    .A2(_10780_),
    .B(_10734_),
    .Y(_10896_));
 NOR2x1_ASAP7_75t_R _15090_ (.A(_08683_),
    .B(_10896_),
    .Y(_10897_));
 BUFx6f_ASAP7_75t_R _15091_ (.A(_10896_),
    .Y(_10898_));
 AO32x1_ASAP7_75t_R _15092_ (.A1(_10893_),
    .A2(_10895_),
    .A3(_10897_),
    .B1(_10898_),
    .B2(_10783_),
    .Y(_03177_));
 BUFx6f_ASAP7_75t_R _15093_ (.A(_10897_),
    .Y(_10899_));
 NAND2x1_ASAP7_75t_R _15094_ (.A(_02018_),
    .B(_10892_),
    .Y(_10900_));
 OR2x2_ASAP7_75t_R _15095_ (.A(_10786_),
    .B(_10894_),
    .Y(_10901_));
 AO32x1_ASAP7_75t_R _15096_ (.A1(_10899_),
    .A2(_10900_),
    .A3(_10901_),
    .B1(_10898_),
    .B2(_10788_),
    .Y(_03178_));
 NAND2x1_ASAP7_75t_R _15097_ (.A(_02017_),
    .B(_10892_),
    .Y(_10902_));
 OR2x2_ASAP7_75t_R _15098_ (.A(_10790_),
    .B(_10894_),
    .Y(_10903_));
 AO32x1_ASAP7_75t_R _15099_ (.A1(_10899_),
    .A2(_10902_),
    .A3(_10903_),
    .B1(_10898_),
    .B2(_10792_),
    .Y(_03179_));
 NAND2x1_ASAP7_75t_R _15100_ (.A(_02016_),
    .B(_10892_),
    .Y(_10904_));
 OR2x2_ASAP7_75t_R _15101_ (.A(_10794_),
    .B(_10894_),
    .Y(_10905_));
 AO32x1_ASAP7_75t_R _15102_ (.A1(_10899_),
    .A2(_10904_),
    .A3(_10905_),
    .B1(_10898_),
    .B2(_10796_),
    .Y(_03180_));
 NAND2x1_ASAP7_75t_R _15103_ (.A(_02015_),
    .B(_10892_),
    .Y(_10906_));
 OR2x2_ASAP7_75t_R _15104_ (.A(_10798_),
    .B(_10894_),
    .Y(_10907_));
 AO32x1_ASAP7_75t_R _15105_ (.A1(_10899_),
    .A2(_10906_),
    .A3(_10907_),
    .B1(_10898_),
    .B2(_10800_),
    .Y(_03181_));
 NAND2x1_ASAP7_75t_R _15106_ (.A(_02014_),
    .B(_10892_),
    .Y(_10908_));
 OR2x2_ASAP7_75t_R _15107_ (.A(_10802_),
    .B(_10894_),
    .Y(_10909_));
 AO32x1_ASAP7_75t_R _15108_ (.A1(_10899_),
    .A2(_10908_),
    .A3(_10909_),
    .B1(_10898_),
    .B2(_10804_),
    .Y(_03182_));
 NAND2x1_ASAP7_75t_R _15109_ (.A(_02013_),
    .B(_10894_),
    .Y(_10910_));
 OA21x2_ASAP7_75t_R _15110_ (.A1(_10772_),
    .A2(_10894_),
    .B(_10910_),
    .Y(_10911_));
 AND3x1_ASAP7_75t_R _15111_ (.A(_08599_),
    .B(_10733_),
    .C(_10896_),
    .Y(_10912_));
 AO21x1_ASAP7_75t_R _15112_ (.A1(_10899_),
    .A2(_10911_),
    .B(_10912_),
    .Y(_03183_));
 NAND2x1_ASAP7_75t_R _15113_ (.A(_02012_),
    .B(_10892_),
    .Y(_10913_));
 OR2x2_ASAP7_75t_R _15114_ (.A(_10807_),
    .B(_10894_),
    .Y(_10914_));
 AO32x1_ASAP7_75t_R _15115_ (.A1(_10899_),
    .A2(_10913_),
    .A3(_10914_),
    .B1(_10898_),
    .B2(_10869_),
    .Y(_03184_));
 NAND2x1_ASAP7_75t_R _15116_ (.A(_02011_),
    .B(_10892_),
    .Y(_10915_));
 OR2x2_ASAP7_75t_R _15117_ (.A(_10811_),
    .B(_10891_),
    .Y(_10916_));
 AO32x1_ASAP7_75t_R _15118_ (.A1(_10899_),
    .A2(_10915_),
    .A3(_10916_),
    .B1(_10898_),
    .B2(_10873_),
    .Y(_03185_));
 NAND2x1_ASAP7_75t_R _15119_ (.A(_10739_),
    .B(_10892_),
    .Y(_10917_));
 OR2x2_ASAP7_75t_R _15120_ (.A(_10753_),
    .B(_10891_),
    .Y(_10918_));
 AO32x1_ASAP7_75t_R _15121_ (.A1(_10899_),
    .A2(_10917_),
    .A3(_10918_),
    .B1(_10898_),
    .B2(_10877_),
    .Y(_03186_));
 INVx1_ASAP7_75t_R _15122_ (.A(_10731_),
    .Y(_10919_));
 OR4x1_ASAP7_75t_R _15123_ (.A(_08712_),
    .B(_10734_),
    .C(_10919_),
    .D(_10780_),
    .Y(_10920_));
 INVx1_ASAP7_75t_R _15124_ (.A(_10920_),
    .Y(_03187_));
 OAI21x1_ASAP7_75t_R _15125_ (.A1(_10888_),
    .A2(_10834_),
    .B(_10890_),
    .Y(_10921_));
 OAI21x1_ASAP7_75t_R _15126_ (.A1(_10730_),
    .A2(_10889_),
    .B(_10921_),
    .Y(_10922_));
 OA21x2_ASAP7_75t_R _15127_ (.A1(_10898_),
    .A2(_10922_),
    .B(_10722_),
    .Y(_03188_));
 NAND2x1_ASAP7_75t_R _15128_ (.A(_02007_),
    .B(_10892_),
    .Y(_10923_));
 OR2x2_ASAP7_75t_R _15129_ (.A(_10820_),
    .B(_10891_),
    .Y(_10924_));
 AO32x1_ASAP7_75t_R _15130_ (.A1(_10899_),
    .A2(_10923_),
    .A3(_10924_),
    .B1(_10896_),
    .B2(_10822_),
    .Y(_03189_));
 NAND2x1_ASAP7_75t_R _15131_ (.A(_02006_),
    .B(_10894_),
    .Y(_10925_));
 OR2x2_ASAP7_75t_R _15132_ (.A(_10824_),
    .B(_10891_),
    .Y(_10926_));
 AO32x1_ASAP7_75t_R _15133_ (.A1(_10897_),
    .A2(_10925_),
    .A3(_10926_),
    .B1(_10896_),
    .B2(_10827_),
    .Y(_03190_));
 BUFx6f_ASAP7_75t_R _15134_ (.A(_08722_),
    .Y(_10927_));
 AND2x2_ASAP7_75t_R _15135_ (.A(_10927_),
    .B(_00012_),
    .Y(_03191_));
 BUFx6f_ASAP7_75t_R _15136_ (.A(_01924_),
    .Y(_10928_));
 INVx1_ASAP7_75t_R _15137_ (.A(_01928_),
    .Y(_10929_));
 BUFx6f_ASAP7_75t_R _15138_ (.A(_01926_),
    .Y(_10930_));
 BUFx6f_ASAP7_75t_R _15139_ (.A(_01927_),
    .Y(_10931_));
 NAND2x1_ASAP7_75t_R _15140_ (.A(_10930_),
    .B(_10931_),
    .Y(_10932_));
 OR3x1_ASAP7_75t_R _15141_ (.A(_10928_),
    .B(_10929_),
    .C(_10932_),
    .Y(_10933_));
 BUFx6f_ASAP7_75t_R _15142_ (.A(_01966_),
    .Y(_10934_));
 NOR2x2_ASAP7_75t_R _15143_ (.A(_10934_),
    .B(_01967_),
    .Y(_10935_));
 BUFx6f_ASAP7_75t_R _15144_ (.A(_01743_),
    .Y(_10936_));
 INVx1_ASAP7_75t_R _15145_ (.A(_10936_),
    .Y(_10937_));
 BUFx6f_ASAP7_75t_R _15146_ (.A(_01746_),
    .Y(_10938_));
 AOI21x1_ASAP7_75t_R _15147_ (.A1(_01968_),
    .A2(_01969_),
    .B(_10934_),
    .Y(_10939_));
 INVx1_ASAP7_75t_R _15148_ (.A(_01742_),
    .Y(_10940_));
 OA211x2_ASAP7_75t_R _15149_ (.A1(_10937_),
    .A2(_10938_),
    .B(_10939_),
    .C(_10940_),
    .Y(_10941_));
 INVx1_ASAP7_75t_R _15150_ (.A(_10928_),
    .Y(_10942_));
 AND4x1_ASAP7_75t_R _15151_ (.A(_10942_),
    .B(_10930_),
    .C(_10931_),
    .D(_01928_),
    .Y(_10943_));
 NOR2x2_ASAP7_75t_R _15152_ (.A(_10928_),
    .B(_01925_),
    .Y(_10944_));
 INVx1_ASAP7_75t_R _15153_ (.A(_10944_),
    .Y(_10945_));
 OA211x2_ASAP7_75t_R _15154_ (.A1(_10935_),
    .A2(_10941_),
    .B(_10943_),
    .C(_10945_),
    .Y(_10946_));
 OA21x2_ASAP7_75t_R _15155_ (.A1(_10937_),
    .A2(_10938_),
    .B(_10940_),
    .Y(_10947_));
 AND3x1_ASAP7_75t_R _15156_ (.A(_01742_),
    .B(_00012_),
    .C(_10939_),
    .Y(_10948_));
 AO21x2_ASAP7_75t_R _15157_ (.A1(_10930_),
    .A2(_10931_),
    .B(_10928_),
    .Y(_10949_));
 NOR2x1_ASAP7_75t_R _15158_ (.A(_10949_),
    .B(_10944_),
    .Y(_10950_));
 AND3x1_ASAP7_75t_R _15159_ (.A(_01967_),
    .B(_01968_),
    .C(_01969_),
    .Y(_10951_));
 OAI21x1_ASAP7_75t_R _15160_ (.A1(_10934_),
    .A2(_10951_),
    .B(_10936_),
    .Y(_10952_));
 OA211x2_ASAP7_75t_R _15161_ (.A1(_10947_),
    .A2(_10948_),
    .B(_10950_),
    .C(_10952_),
    .Y(_10953_));
 NOR3x1_ASAP7_75t_R _15162_ (.A(_10933_),
    .B(_10946_),
    .C(_10953_),
    .Y(_10954_));
 INVx1_ASAP7_75t_R _15163_ (.A(_10934_),
    .Y(_10955_));
 INVx2_ASAP7_75t_R _15164_ (.A(_01970_),
    .Y(_10956_));
 AND4x1_ASAP7_75t_R _15165_ (.A(_10955_),
    .B(_01968_),
    .C(_01969_),
    .D(_10956_),
    .Y(_10957_));
 AO21x2_ASAP7_75t_R _15166_ (.A1(_01968_),
    .A2(_01969_),
    .B(_10934_),
    .Y(_10958_));
 INVx1_ASAP7_75t_R _15167_ (.A(_10938_),
    .Y(_10959_));
 AO221x1_ASAP7_75t_R _15168_ (.A1(_10957_),
    .A2(_10944_),
    .B1(_10943_),
    .B2(_10958_),
    .C(_10959_),
    .Y(_10960_));
 OAI21x1_ASAP7_75t_R _15169_ (.A1(_10934_),
    .A2(_01967_),
    .B(_10938_),
    .Y(_10961_));
 OA21x2_ASAP7_75t_R _15170_ (.A1(_10938_),
    .A2(_10944_),
    .B(_10961_),
    .Y(_10962_));
 NAND2x1_ASAP7_75t_R _15171_ (.A(_10940_),
    .B(_10936_),
    .Y(_10963_));
 AO211x2_ASAP7_75t_R _15172_ (.A1(_10957_),
    .A2(_10943_),
    .B(_10962_),
    .C(_10963_),
    .Y(_10964_));
 OR2x6_ASAP7_75t_R _15173_ (.A(_10960_),
    .B(_10964_),
    .Y(_10965_));
 INVx1_ASAP7_75t_R _15174_ (.A(_10965_),
    .Y(_10966_));
 AO31x2_ASAP7_75t_R _15175_ (.A1(_01925_),
    .A2(_10930_),
    .A3(_10931_),
    .B(_10928_),
    .Y(_10967_));
 NAND2x1_ASAP7_75t_R _15176_ (.A(_10936_),
    .B(_10967_),
    .Y(_10968_));
 INVx1_ASAP7_75t_R _15177_ (.A(_00012_),
    .Y(_10969_));
 AOI21x1_ASAP7_75t_R _15178_ (.A1(_10930_),
    .A2(_10931_),
    .B(_10928_),
    .Y(_10970_));
 AOI21x1_ASAP7_75t_R _15179_ (.A1(_10936_),
    .A2(_10938_),
    .B(_01742_),
    .Y(_10971_));
 AO31x2_ASAP7_75t_R _15180_ (.A1(_01742_),
    .A2(_10969_),
    .A3(_10970_),
    .B(_10971_),
    .Y(_10972_));
 AO21x1_ASAP7_75t_R _15181_ (.A1(_10971_),
    .A2(_10970_),
    .B(_10944_),
    .Y(_10973_));
 AO32x2_ASAP7_75t_R _15182_ (.A1(_10968_),
    .A2(_10972_),
    .A3(_10939_),
    .B1(_10957_),
    .B2(_10973_),
    .Y(_10974_));
 NOR2x1_ASAP7_75t_R _15183_ (.A(_10935_),
    .B(_10974_),
    .Y(_10975_));
 OAI21x1_ASAP7_75t_R _15184_ (.A1(_10954_),
    .A2(_10966_),
    .B(_10975_),
    .Y(_10976_));
 BUFx6f_ASAP7_75t_R _15185_ (.A(_10954_),
    .Y(_10977_));
 NAND2x1_ASAP7_75t_R _15186_ (.A(_01935_),
    .B(_10977_),
    .Y(_10978_));
 INVx1_ASAP7_75t_R _15187_ (.A(_01753_),
    .Y(_10979_));
 BUFx6f_ASAP7_75t_R _15188_ (.A(_10954_),
    .Y(_10980_));
 BUFx6f_ASAP7_75t_R _15189_ (.A(_10965_),
    .Y(_10981_));
 OR3x1_ASAP7_75t_R _15190_ (.A(_10979_),
    .B(_10980_),
    .C(_10981_),
    .Y(_10982_));
 OR2x6_ASAP7_75t_R _15191_ (.A(_10935_),
    .B(_10974_),
    .Y(_10983_));
 BUFx12f_ASAP7_75t_R _15192_ (.A(_10983_),
    .Y(_10984_));
 AOI21x1_ASAP7_75t_R _15193_ (.A1(_10978_),
    .A2(_10982_),
    .B(_10984_),
    .Y(_10985_));
 BUFx12f_ASAP7_75t_R _15194_ (.A(_09818_),
    .Y(_10986_));
 AOI211x1_ASAP7_75t_R _15195_ (.A1(_01977_),
    .A2(_10976_),
    .B(_10985_),
    .C(_10986_),
    .Y(_03192_));
 NAND2x1_ASAP7_75t_R _15196_ (.A(_01934_),
    .B(_10977_),
    .Y(_10987_));
 INVx1_ASAP7_75t_R _15197_ (.A(_01752_),
    .Y(_10988_));
 OR3x1_ASAP7_75t_R _15198_ (.A(_10988_),
    .B(_10980_),
    .C(_10981_),
    .Y(_10989_));
 AOI21x1_ASAP7_75t_R _15199_ (.A1(_10987_),
    .A2(_10989_),
    .B(_10984_),
    .Y(_10990_));
 AOI211x1_ASAP7_75t_R _15200_ (.A1(_01976_),
    .A2(_10976_),
    .B(_10990_),
    .C(_10986_),
    .Y(_03193_));
 NAND2x1_ASAP7_75t_R _15201_ (.A(_01933_),
    .B(_10977_),
    .Y(_10991_));
 INVx1_ASAP7_75t_R _15202_ (.A(_01751_),
    .Y(_10992_));
 OR3x1_ASAP7_75t_R _15203_ (.A(_10992_),
    .B(_10980_),
    .C(_10981_),
    .Y(_10993_));
 AOI21x1_ASAP7_75t_R _15204_ (.A1(_10991_),
    .A2(_10993_),
    .B(_10984_),
    .Y(_10994_));
 BUFx12f_ASAP7_75t_R _15205_ (.A(_09818_),
    .Y(_10995_));
 AOI211x1_ASAP7_75t_R _15206_ (.A1(_01975_),
    .A2(_10976_),
    .B(_10994_),
    .C(_10995_),
    .Y(_03194_));
 NAND2x1_ASAP7_75t_R _15207_ (.A(_01932_),
    .B(_10977_),
    .Y(_10996_));
 INVx1_ASAP7_75t_R _15208_ (.A(_01750_),
    .Y(_10997_));
 OR3x1_ASAP7_75t_R _15209_ (.A(_10997_),
    .B(_10980_),
    .C(_10981_),
    .Y(_10998_));
 AOI21x1_ASAP7_75t_R _15210_ (.A1(_10996_),
    .A2(_10998_),
    .B(_10984_),
    .Y(_10999_));
 AOI211x1_ASAP7_75t_R _15211_ (.A1(_01974_),
    .A2(_10976_),
    .B(_10999_),
    .C(_10995_),
    .Y(_03195_));
 NAND2x1_ASAP7_75t_R _15212_ (.A(_01931_),
    .B(_10977_),
    .Y(_11000_));
 INVx1_ASAP7_75t_R _15213_ (.A(_01749_),
    .Y(_11001_));
 OR3x1_ASAP7_75t_R _15214_ (.A(_11001_),
    .B(_10980_),
    .C(_10981_),
    .Y(_11002_));
 AOI21x1_ASAP7_75t_R _15215_ (.A1(_11000_),
    .A2(_11002_),
    .B(_10984_),
    .Y(_11003_));
 AOI211x1_ASAP7_75t_R _15216_ (.A1(_01973_),
    .A2(_10976_),
    .B(_11003_),
    .C(_10995_),
    .Y(_03196_));
 NAND2x1_ASAP7_75t_R _15217_ (.A(_01930_),
    .B(_10977_),
    .Y(_11004_));
 INVx1_ASAP7_75t_R _15218_ (.A(_01748_),
    .Y(_11005_));
 OR3x1_ASAP7_75t_R _15219_ (.A(_11005_),
    .B(_10980_),
    .C(_10981_),
    .Y(_11006_));
 AOI21x1_ASAP7_75t_R _15220_ (.A1(_11004_),
    .A2(_11006_),
    .B(_10984_),
    .Y(_11007_));
 AOI211x1_ASAP7_75t_R _15221_ (.A1(_01972_),
    .A2(_10976_),
    .B(_11007_),
    .C(_10995_),
    .Y(_03197_));
 NAND2x1_ASAP7_75t_R _15222_ (.A(_01929_),
    .B(_10977_),
    .Y(_11008_));
 INVx1_ASAP7_75t_R _15223_ (.A(_01747_),
    .Y(_11009_));
 OR3x1_ASAP7_75t_R _15224_ (.A(_11009_),
    .B(_10980_),
    .C(_10981_),
    .Y(_11010_));
 AOI21x1_ASAP7_75t_R _15225_ (.A1(_11008_),
    .A2(_11010_),
    .B(_10984_),
    .Y(_11011_));
 AOI211x1_ASAP7_75t_R _15226_ (.A1(_01971_),
    .A2(_10976_),
    .B(_11011_),
    .C(_10995_),
    .Y(_03198_));
 AND3x1_ASAP7_75t_R _15227_ (.A(_10809_),
    .B(_10956_),
    .C(_10976_),
    .Y(_03199_));
 OR3x1_ASAP7_75t_R _15228_ (.A(_01745_),
    .B(_10960_),
    .C(_10964_),
    .Y(_11012_));
 INVx2_ASAP7_75t_R _15229_ (.A(_01969_),
    .Y(_11013_));
 NAND2x1_ASAP7_75t_R _15230_ (.A(_11013_),
    .B(_10981_),
    .Y(_11014_));
 AO21x1_ASAP7_75t_R _15231_ (.A1(_11012_),
    .A2(_11014_),
    .B(_10977_),
    .Y(_11015_));
 NAND2x1_ASAP7_75t_R _15232_ (.A(_11013_),
    .B(_10984_),
    .Y(_11016_));
 AOI21x1_ASAP7_75t_R _15233_ (.A1(_11015_),
    .A2(_11016_),
    .B(_10530_),
    .Y(_03200_));
 OR3x1_ASAP7_75t_R _15234_ (.A(_01744_),
    .B(_10960_),
    .C(_10964_),
    .Y(_11017_));
 INVx2_ASAP7_75t_R _15235_ (.A(_01968_),
    .Y(_11018_));
 NAND2x1_ASAP7_75t_R _15236_ (.A(_11018_),
    .B(_10981_),
    .Y(_11019_));
 AO21x1_ASAP7_75t_R _15237_ (.A1(_11017_),
    .A2(_11019_),
    .B(_10977_),
    .Y(_11020_));
 NAND2x1_ASAP7_75t_R _15238_ (.A(_11018_),
    .B(_10984_),
    .Y(_11021_));
 AOI21x1_ASAP7_75t_R _15239_ (.A1(_11020_),
    .A2(_11021_),
    .B(_10530_),
    .Y(_03201_));
 OAI21x1_ASAP7_75t_R _15240_ (.A1(_10934_),
    .A2(_01967_),
    .B(_10974_),
    .Y(_11022_));
 NOR2x1_ASAP7_75t_R _15241_ (.A(_10716_),
    .B(_11022_),
    .Y(_03202_));
 OR3x1_ASAP7_75t_R _15242_ (.A(_10983_),
    .B(_10980_),
    .C(_10966_),
    .Y(_11023_));
 AND2x2_ASAP7_75t_R _15243_ (.A(_10927_),
    .B(_11023_),
    .Y(_03203_));
 NAND2x1_ASAP7_75t_R _15244_ (.A(_01923_),
    .B(_10977_),
    .Y(_11024_));
 INVx1_ASAP7_75t_R _15245_ (.A(_01741_),
    .Y(_11025_));
 OR3x1_ASAP7_75t_R _15246_ (.A(_11025_),
    .B(_10980_),
    .C(_10981_),
    .Y(_11026_));
 AOI21x1_ASAP7_75t_R _15247_ (.A1(_11024_),
    .A2(_11026_),
    .B(_10984_),
    .Y(_11027_));
 AOI211x1_ASAP7_75t_R _15248_ (.A1(_01965_),
    .A2(_10976_),
    .B(_11027_),
    .C(_10995_),
    .Y(_03204_));
 NAND2x1_ASAP7_75t_R _15249_ (.A(_01922_),
    .B(_10980_),
    .Y(_11028_));
 INVx1_ASAP7_75t_R _15250_ (.A(_01740_),
    .Y(_11029_));
 OR3x1_ASAP7_75t_R _15251_ (.A(_11029_),
    .B(_10954_),
    .C(_10965_),
    .Y(_11030_));
 AOI21x1_ASAP7_75t_R _15252_ (.A1(_11028_),
    .A2(_11030_),
    .B(_10983_),
    .Y(_11031_));
 AOI211x1_ASAP7_75t_R _15253_ (.A1(_01964_),
    .A2(_10976_),
    .B(_11031_),
    .C(_10995_),
    .Y(_03205_));
 AO221x1_ASAP7_75t_R _15254_ (.A1(_10949_),
    .A2(_10957_),
    .B1(_10943_),
    .B2(_10935_),
    .C(_10938_),
    .Y(_11032_));
 OR2x6_ASAP7_75t_R _15255_ (.A(_10964_),
    .B(_11032_),
    .Y(_11033_));
 OA211x2_ASAP7_75t_R _15256_ (.A1(_10947_),
    .A2(_10948_),
    .B(_10970_),
    .C(_10952_),
    .Y(_11034_));
 OA21x2_ASAP7_75t_R _15257_ (.A1(_10935_),
    .A2(_10941_),
    .B(_10943_),
    .Y(_11035_));
 OR3x1_ASAP7_75t_R _15258_ (.A(_10944_),
    .B(_11034_),
    .C(_11035_),
    .Y(_11036_));
 BUFx6f_ASAP7_75t_R _15259_ (.A(_11036_),
    .Y(_11037_));
 AO211x2_ASAP7_75t_R _15260_ (.A1(_10957_),
    .A2(_11022_),
    .B(_11033_),
    .C(_11037_),
    .Y(_11038_));
 BUFx12f_ASAP7_75t_R _15261_ (.A(_11038_),
    .Y(_11039_));
 NOR2x1_ASAP7_75t_R _15262_ (.A(_01753_),
    .B(_11039_),
    .Y(_11040_));
 INVx1_ASAP7_75t_R _15263_ (.A(_01977_),
    .Y(_11041_));
 BUFx6f_ASAP7_75t_R _15264_ (.A(_11037_),
    .Y(_11042_));
 BUFx6f_ASAP7_75t_R _15265_ (.A(_11038_),
    .Y(_11043_));
 BUFx6f_ASAP7_75t_R _15266_ (.A(_11037_),
    .Y(_11044_));
 NAND2x1_ASAP7_75t_R _15267_ (.A(_01935_),
    .B(_11044_),
    .Y(_11045_));
 OA211x2_ASAP7_75t_R _15268_ (.A1(_11041_),
    .A2(_11042_),
    .B(_11043_),
    .C(_11045_),
    .Y(_11046_));
 OA21x2_ASAP7_75t_R _15269_ (.A1(_11040_),
    .A2(_11046_),
    .B(_10722_),
    .Y(_03206_));
 NOR2x1_ASAP7_75t_R _15270_ (.A(_01752_),
    .B(_11039_),
    .Y(_11047_));
 INVx1_ASAP7_75t_R _15271_ (.A(_01976_),
    .Y(_11048_));
 NAND2x1_ASAP7_75t_R _15272_ (.A(_01934_),
    .B(_11044_),
    .Y(_11049_));
 OA211x2_ASAP7_75t_R _15273_ (.A1(_11048_),
    .A2(_11042_),
    .B(_11043_),
    .C(_11049_),
    .Y(_11050_));
 OA21x2_ASAP7_75t_R _15274_ (.A1(_11047_),
    .A2(_11050_),
    .B(_10722_),
    .Y(_03207_));
 NOR2x1_ASAP7_75t_R _15275_ (.A(_01751_),
    .B(_11039_),
    .Y(_11051_));
 INVx1_ASAP7_75t_R _15276_ (.A(_01975_),
    .Y(_11052_));
 NAND2x1_ASAP7_75t_R _15277_ (.A(_01933_),
    .B(_11044_),
    .Y(_11053_));
 OA211x2_ASAP7_75t_R _15278_ (.A1(_11052_),
    .A2(_11042_),
    .B(_11043_),
    .C(_11053_),
    .Y(_11054_));
 OA21x2_ASAP7_75t_R _15279_ (.A1(_11051_),
    .A2(_11054_),
    .B(_10722_),
    .Y(_03208_));
 NOR2x1_ASAP7_75t_R _15280_ (.A(_01750_),
    .B(_11039_),
    .Y(_11055_));
 INVx1_ASAP7_75t_R _15281_ (.A(_01974_),
    .Y(_11056_));
 NAND2x1_ASAP7_75t_R _15282_ (.A(_01932_),
    .B(_11044_),
    .Y(_11057_));
 OA211x2_ASAP7_75t_R _15283_ (.A1(_11056_),
    .A2(_11042_),
    .B(_11043_),
    .C(_11057_),
    .Y(_11058_));
 OA21x2_ASAP7_75t_R _15284_ (.A1(_11055_),
    .A2(_11058_),
    .B(_10722_),
    .Y(_03209_));
 NOR2x1_ASAP7_75t_R _15285_ (.A(_01749_),
    .B(_11039_),
    .Y(_11059_));
 INVx1_ASAP7_75t_R _15286_ (.A(_01973_),
    .Y(_11060_));
 NAND2x1_ASAP7_75t_R _15287_ (.A(_01931_),
    .B(_11044_),
    .Y(_11061_));
 OA211x2_ASAP7_75t_R _15288_ (.A1(_11060_),
    .A2(_11042_),
    .B(_11043_),
    .C(_11061_),
    .Y(_11062_));
 OA21x2_ASAP7_75t_R _15289_ (.A1(_11059_),
    .A2(_11062_),
    .B(_10722_),
    .Y(_03210_));
 NOR2x1_ASAP7_75t_R _15290_ (.A(_01748_),
    .B(_11039_),
    .Y(_11063_));
 INVx1_ASAP7_75t_R _15291_ (.A(_01972_),
    .Y(_11064_));
 NAND2x1_ASAP7_75t_R _15292_ (.A(_01930_),
    .B(_11044_),
    .Y(_11065_));
 OA211x2_ASAP7_75t_R _15293_ (.A1(_11064_),
    .A2(_11042_),
    .B(_11043_),
    .C(_11065_),
    .Y(_11066_));
 BUFx6f_ASAP7_75t_R _15294_ (.A(_09229_),
    .Y(_11067_));
 OA21x2_ASAP7_75t_R _15295_ (.A1(_11063_),
    .A2(_11066_),
    .B(_11067_),
    .Y(_03211_));
 NOR2x1_ASAP7_75t_R _15296_ (.A(_01747_),
    .B(_11039_),
    .Y(_11068_));
 INVx1_ASAP7_75t_R _15297_ (.A(_01971_),
    .Y(_11069_));
 NAND2x1_ASAP7_75t_R _15298_ (.A(_01929_),
    .B(_11037_),
    .Y(_11070_));
 OA211x2_ASAP7_75t_R _15299_ (.A1(_11069_),
    .A2(_11042_),
    .B(_11043_),
    .C(_11070_),
    .Y(_11071_));
 OA21x2_ASAP7_75t_R _15300_ (.A1(_11068_),
    .A2(_11071_),
    .B(_11067_),
    .Y(_03212_));
 NOR2x1_ASAP7_75t_R _15301_ (.A(_10956_),
    .B(_11042_),
    .Y(_11072_));
 AO21x1_ASAP7_75t_R _15302_ (.A1(_01928_),
    .A2(_11042_),
    .B(_11072_),
    .Y(_11073_));
 AOI21x1_ASAP7_75t_R _15303_ (.A1(_11039_),
    .A2(_11073_),
    .B(_10530_),
    .Y(_03213_));
 NOR2x1_ASAP7_75t_R _15304_ (.A(_01745_),
    .B(_11039_),
    .Y(_11074_));
 NAND2x1_ASAP7_75t_R _15305_ (.A(_10931_),
    .B(_11037_),
    .Y(_11075_));
 OA211x2_ASAP7_75t_R _15306_ (.A1(_11013_),
    .A2(_11044_),
    .B(_11043_),
    .C(_11075_),
    .Y(_11076_));
 OA21x2_ASAP7_75t_R _15307_ (.A1(_11074_),
    .A2(_11076_),
    .B(_11067_),
    .Y(_03214_));
 NOR2x1_ASAP7_75t_R _15308_ (.A(_01744_),
    .B(_11039_),
    .Y(_11077_));
 NAND2x1_ASAP7_75t_R _15309_ (.A(_10930_),
    .B(_11037_),
    .Y(_11078_));
 OA211x2_ASAP7_75t_R _15310_ (.A1(_11018_),
    .A2(_11044_),
    .B(_11038_),
    .C(_11078_),
    .Y(_11079_));
 OA21x2_ASAP7_75t_R _15311_ (.A1(_11077_),
    .A2(_11079_),
    .B(_11067_),
    .Y(_03215_));
 OA21x2_ASAP7_75t_R _15312_ (.A1(_10946_),
    .A2(_10953_),
    .B(_11067_),
    .Y(_03216_));
 AO21x1_ASAP7_75t_R _15313_ (.A1(_10957_),
    .A2(_11022_),
    .B(_11042_),
    .Y(_11080_));
 INVx1_ASAP7_75t_R _15314_ (.A(_11080_),
    .Y(_11081_));
 AOI21x1_ASAP7_75t_R _15315_ (.A1(_11033_),
    .A2(_11081_),
    .B(_09081_),
    .Y(_03217_));
 NOR2x1_ASAP7_75t_R _15316_ (.A(_01741_),
    .B(_11043_),
    .Y(_11082_));
 INVx1_ASAP7_75t_R _15317_ (.A(_01965_),
    .Y(_11083_));
 NAND2x1_ASAP7_75t_R _15318_ (.A(_01923_),
    .B(_11037_),
    .Y(_11084_));
 OA211x2_ASAP7_75t_R _15319_ (.A1(_11083_),
    .A2(_11044_),
    .B(_11038_),
    .C(_11084_),
    .Y(_11085_));
 OA21x2_ASAP7_75t_R _15320_ (.A1(_11082_),
    .A2(_11085_),
    .B(_11067_),
    .Y(_03218_));
 NOR2x1_ASAP7_75t_R _15321_ (.A(_01740_),
    .B(_11043_),
    .Y(_11086_));
 INVx1_ASAP7_75t_R _15322_ (.A(_01964_),
    .Y(_11087_));
 NAND2x1_ASAP7_75t_R _15323_ (.A(_01922_),
    .B(_11037_),
    .Y(_11088_));
 OA211x2_ASAP7_75t_R _15324_ (.A1(_11087_),
    .A2(_11044_),
    .B(_11038_),
    .C(_11088_),
    .Y(_11089_));
 OA21x2_ASAP7_75t_R _15325_ (.A1(_11086_),
    .A2(_11089_),
    .B(_11067_),
    .Y(_03219_));
 AOI221x1_ASAP7_75t_R _15326_ (.A1(_10957_),
    .A2(_10943_),
    .B1(_10960_),
    .B2(_11032_),
    .C(_10962_),
    .Y(_11090_));
 AO21x2_ASAP7_75t_R _15327_ (.A1(_10936_),
    .A2(_11090_),
    .B(_01742_),
    .Y(_11091_));
 OR2x6_ASAP7_75t_R _15328_ (.A(_09220_),
    .B(_11091_),
    .Y(_11092_));
 BUFx12f_ASAP7_75t_R _15329_ (.A(_11092_),
    .Y(_11093_));
 NAND2x2_ASAP7_75t_R _15330_ (.A(_08876_),
    .B(_11091_),
    .Y(_11094_));
 BUFx12f_ASAP7_75t_R _15331_ (.A(_11094_),
    .Y(_11095_));
 AND5x1_ASAP7_75t_R _15332_ (.A(_10955_),
    .B(_01967_),
    .C(_01968_),
    .D(_01969_),
    .E(_10956_),
    .Y(_11096_));
 AOI211x1_ASAP7_75t_R _15333_ (.A1(_10936_),
    .A2(_10967_),
    .B(_10958_),
    .C(_10935_),
    .Y(_11097_));
 AOI221x1_ASAP7_75t_R _15334_ (.A1(_10973_),
    .A2(_11096_),
    .B1(_11097_),
    .B2(_10972_),
    .C(_10958_),
    .Y(_11098_));
 OR3x1_ASAP7_75t_R _15335_ (.A(_10949_),
    .B(_10946_),
    .C(_10953_),
    .Y(_11099_));
 NOR2x1_ASAP7_75t_R _15336_ (.A(_11098_),
    .B(_11099_),
    .Y(_11100_));
 BUFx6f_ASAP7_75t_R _15337_ (.A(_11100_),
    .Y(_11101_));
 OR4x1_ASAP7_75t_R _15338_ (.A(_10949_),
    .B(_10946_),
    .C(_10953_),
    .D(_11098_),
    .Y(_11102_));
 BUFx6f_ASAP7_75t_R _15339_ (.A(_11102_),
    .Y(_11103_));
 AND2x2_ASAP7_75t_R _15340_ (.A(_01977_),
    .B(_11103_),
    .Y(_11104_));
 AO21x1_ASAP7_75t_R _15341_ (.A1(_01935_),
    .A2(_11101_),
    .B(_11104_),
    .Y(_11105_));
 OAI22x1_ASAP7_75t_R _15342_ (.A1(_01753_),
    .A2(_11093_),
    .B1(_11095_),
    .B2(_11105_),
    .Y(_03220_));
 AND2x2_ASAP7_75t_R _15343_ (.A(_01976_),
    .B(_11103_),
    .Y(_11106_));
 AO21x1_ASAP7_75t_R _15344_ (.A1(_01934_),
    .A2(_11101_),
    .B(_11106_),
    .Y(_11107_));
 OAI22x1_ASAP7_75t_R _15345_ (.A1(_01752_),
    .A2(_11093_),
    .B1(_11095_),
    .B2(_11107_),
    .Y(_03221_));
 AND2x2_ASAP7_75t_R _15346_ (.A(_01975_),
    .B(_11103_),
    .Y(_11108_));
 AO21x1_ASAP7_75t_R _15347_ (.A1(_01933_),
    .A2(_11101_),
    .B(_11108_),
    .Y(_11109_));
 OAI22x1_ASAP7_75t_R _15348_ (.A1(_01751_),
    .A2(_11093_),
    .B1(_11095_),
    .B2(_11109_),
    .Y(_03222_));
 AND2x2_ASAP7_75t_R _15349_ (.A(_01974_),
    .B(_11103_),
    .Y(_11110_));
 AO21x1_ASAP7_75t_R _15350_ (.A1(_01932_),
    .A2(_11101_),
    .B(_11110_),
    .Y(_11111_));
 OAI22x1_ASAP7_75t_R _15351_ (.A1(_01750_),
    .A2(_11093_),
    .B1(_11095_),
    .B2(_11111_),
    .Y(_03223_));
 AND2x2_ASAP7_75t_R _15352_ (.A(_01973_),
    .B(_11103_),
    .Y(_11112_));
 AO21x1_ASAP7_75t_R _15353_ (.A1(_01931_),
    .A2(_11101_),
    .B(_11112_),
    .Y(_11113_));
 OAI22x1_ASAP7_75t_R _15354_ (.A1(_01749_),
    .A2(_11093_),
    .B1(_11095_),
    .B2(_11113_),
    .Y(_03224_));
 AND2x2_ASAP7_75t_R _15355_ (.A(_01972_),
    .B(_11103_),
    .Y(_11114_));
 AO21x1_ASAP7_75t_R _15356_ (.A1(_01930_),
    .A2(_11101_),
    .B(_11114_),
    .Y(_11115_));
 OAI22x1_ASAP7_75t_R _15357_ (.A1(_01748_),
    .A2(_11093_),
    .B1(_11095_),
    .B2(_11115_),
    .Y(_03225_));
 AND2x2_ASAP7_75t_R _15358_ (.A(_01971_),
    .B(_11103_),
    .Y(_11116_));
 AO21x1_ASAP7_75t_R _15359_ (.A1(_01929_),
    .A2(_11101_),
    .B(_11116_),
    .Y(_11117_));
 OAI22x1_ASAP7_75t_R _15360_ (.A1(_01747_),
    .A2(_11093_),
    .B1(_11095_),
    .B2(_11117_),
    .Y(_03226_));
 AND2x2_ASAP7_75t_R _15361_ (.A(_01970_),
    .B(_11103_),
    .Y(_11118_));
 AO21x1_ASAP7_75t_R _15362_ (.A1(_01928_),
    .A2(_11101_),
    .B(_11118_),
    .Y(_11119_));
 OR3x1_ASAP7_75t_R _15363_ (.A(_09118_),
    .B(_10938_),
    .C(_11091_),
    .Y(_11120_));
 OAI21x1_ASAP7_75t_R _15364_ (.A1(_11095_),
    .A2(_11119_),
    .B(_11120_),
    .Y(_03227_));
 AND2x2_ASAP7_75t_R _15365_ (.A(_01969_),
    .B(_11103_),
    .Y(_11121_));
 AO21x1_ASAP7_75t_R _15366_ (.A1(_10931_),
    .A2(_11101_),
    .B(_11121_),
    .Y(_11122_));
 OR3x1_ASAP7_75t_R _15367_ (.A(_09118_),
    .B(_01745_),
    .C(_11091_),
    .Y(_11123_));
 OAI21x1_ASAP7_75t_R _15368_ (.A1(_11095_),
    .A2(_11122_),
    .B(_11123_),
    .Y(_03228_));
 AND2x2_ASAP7_75t_R _15369_ (.A(_01968_),
    .B(_11103_),
    .Y(_11124_));
 AO21x1_ASAP7_75t_R _15370_ (.A1(_10930_),
    .A2(_11101_),
    .B(_11124_),
    .Y(_11125_));
 BUFx6f_ASAP7_75t_R _15371_ (.A(_08656_),
    .Y(_11126_));
 OR3x1_ASAP7_75t_R _15372_ (.A(_11126_),
    .B(_01744_),
    .C(_11091_),
    .Y(_11127_));
 OAI21x1_ASAP7_75t_R _15373_ (.A1(_11095_),
    .A2(_11125_),
    .B(_11127_),
    .Y(_03229_));
 OR3x1_ASAP7_75t_R _15374_ (.A(_08642_),
    .B(_10963_),
    .C(_11090_),
    .Y(_11128_));
 INVx1_ASAP7_75t_R _15375_ (.A(_11128_),
    .Y(_03230_));
 NAND2x1_ASAP7_75t_R _15376_ (.A(_11091_),
    .B(_11099_),
    .Y(_11129_));
 OA21x2_ASAP7_75t_R _15377_ (.A1(_11098_),
    .A2(_11129_),
    .B(_11067_),
    .Y(_03231_));
 AND2x2_ASAP7_75t_R _15378_ (.A(_01965_),
    .B(_11102_),
    .Y(_11130_));
 AO21x1_ASAP7_75t_R _15379_ (.A1(_01923_),
    .A2(_11100_),
    .B(_11130_),
    .Y(_11131_));
 OAI22x1_ASAP7_75t_R _15380_ (.A1(_01741_),
    .A2(_11093_),
    .B1(_11094_),
    .B2(_11131_),
    .Y(_03232_));
 AND2x2_ASAP7_75t_R _15381_ (.A(_01964_),
    .B(_11102_),
    .Y(_11132_));
 AO21x1_ASAP7_75t_R _15382_ (.A1(_01922_),
    .A2(_11100_),
    .B(_11132_),
    .Y(_11133_));
 OAI22x1_ASAP7_75t_R _15383_ (.A1(_01740_),
    .A2(_11093_),
    .B1(_11094_),
    .B2(_11133_),
    .Y(_03233_));
 AND2x2_ASAP7_75t_R _15384_ (.A(_10927_),
    .B(_00013_),
    .Y(_03234_));
 INVx2_ASAP7_75t_R _15385_ (.A(_01884_),
    .Y(_11134_));
 OR4x1_ASAP7_75t_R _15386_ (.A(_01882_),
    .B(_11134_),
    .C(_01885_),
    .D(_01886_),
    .Y(_11135_));
 INVx1_ASAP7_75t_R _15387_ (.A(_01843_),
    .Y(_11136_));
 AO21x2_ASAP7_75t_R _15388_ (.A1(_01842_),
    .A2(_11136_),
    .B(_01840_),
    .Y(_11137_));
 BUFx6f_ASAP7_75t_R _15389_ (.A(_01732_),
    .Y(_11138_));
 AO21x1_ASAP7_75t_R _15390_ (.A1(_01729_),
    .A2(_11138_),
    .B(_01728_),
    .Y(_11139_));
 OR2x2_ASAP7_75t_R _15391_ (.A(_01840_),
    .B(_01841_),
    .Y(_11140_));
 BUFx3_ASAP7_75t_R _15392_ (.A(_11140_),
    .Y(_11141_));
 OA21x2_ASAP7_75t_R _15393_ (.A1(_11137_),
    .A2(_11139_),
    .B(_11141_),
    .Y(_11142_));
 AND3x1_ASAP7_75t_R _15394_ (.A(_01841_),
    .B(_01842_),
    .C(_11136_),
    .Y(_11143_));
 INVx3_ASAP7_75t_R _15395_ (.A(_01728_),
    .Y(_11144_));
 AO21x1_ASAP7_75t_R _15396_ (.A1(_11144_),
    .A2(_11138_),
    .B(_01840_),
    .Y(_11145_));
 OA21x2_ASAP7_75t_R _15397_ (.A1(_11143_),
    .A2(_11145_),
    .B(_01729_),
    .Y(_11146_));
 INVx1_ASAP7_75t_R _15398_ (.A(_01842_),
    .Y(_11147_));
 INVx1_ASAP7_75t_R _15399_ (.A(_00013_),
    .Y(_11148_));
 INVx1_ASAP7_75t_R _15400_ (.A(_01840_),
    .Y(_11149_));
 OA211x2_ASAP7_75t_R _15401_ (.A1(_11147_),
    .A2(_01843_),
    .B(_11148_),
    .C(_11149_),
    .Y(_11150_));
 INVx2_ASAP7_75t_R _15402_ (.A(_01882_),
    .Y(_11151_));
 OA21x2_ASAP7_75t_R _15403_ (.A1(_11134_),
    .A2(_01885_),
    .B(_11151_),
    .Y(_11152_));
 BUFx6f_ASAP7_75t_R _15404_ (.A(_11152_),
    .Y(_11153_));
 OAI21x1_ASAP7_75t_R _15405_ (.A1(_11144_),
    .A2(_11150_),
    .B(_11153_),
    .Y(_11154_));
 OA222x2_ASAP7_75t_R _15406_ (.A1(_01882_),
    .A2(_01883_),
    .B1(_11135_),
    .B2(_11142_),
    .C1(_11146_),
    .C2(_11154_),
    .Y(_11155_));
 INVx1_ASAP7_75t_R _15407_ (.A(_01729_),
    .Y(_11156_));
 OA21x2_ASAP7_75t_R _15408_ (.A1(_11156_),
    .A2(_11138_),
    .B(_11144_),
    .Y(_11157_));
 NOR2x1_ASAP7_75t_R _15409_ (.A(_01882_),
    .B(_01883_),
    .Y(_11158_));
 AO21x2_ASAP7_75t_R _15410_ (.A1(_11153_),
    .A2(_11157_),
    .B(_11158_),
    .Y(_11159_));
 INVx1_ASAP7_75t_R _15411_ (.A(_01883_),
    .Y(_11160_));
 OR3x1_ASAP7_75t_R _15412_ (.A(_11160_),
    .B(_11134_),
    .C(_01885_),
    .Y(_11161_));
 OA21x2_ASAP7_75t_R _15413_ (.A1(_01728_),
    .A2(_11138_),
    .B(_11151_),
    .Y(_11162_));
 AO21x2_ASAP7_75t_R _15414_ (.A1(_11161_),
    .A2(_11162_),
    .B(_11156_),
    .Y(_11163_));
 OA211x2_ASAP7_75t_R _15415_ (.A1(_11134_),
    .A2(_01885_),
    .B(_00013_),
    .C(_11151_),
    .Y(_11164_));
 OA21x2_ASAP7_75t_R _15416_ (.A1(_11147_),
    .A2(_01843_),
    .B(_11149_),
    .Y(_11165_));
 OA211x2_ASAP7_75t_R _15417_ (.A1(_11144_),
    .A2(_11164_),
    .B(_11165_),
    .C(_11141_),
    .Y(_11166_));
 INVx1_ASAP7_75t_R _15418_ (.A(_01844_),
    .Y(_11167_));
 OR4x1_ASAP7_75t_R _15419_ (.A(_01840_),
    .B(_11147_),
    .C(_01843_),
    .D(_11167_),
    .Y(_11168_));
 AOI221x1_ASAP7_75t_R _15420_ (.A1(_11141_),
    .A2(_11159_),
    .B1(_11163_),
    .B2(_11166_),
    .C(_11168_),
    .Y(_11169_));
 AND2x4_ASAP7_75t_R _15421_ (.A(_11155_),
    .B(_11169_),
    .Y(_11170_));
 BUFx6f_ASAP7_75t_R _15422_ (.A(_11170_),
    .Y(_11171_));
 NAND2x1_ASAP7_75t_R _15423_ (.A(_01851_),
    .B(_11171_),
    .Y(_11172_));
 BUFx6f_ASAP7_75t_R _15424_ (.A(_11155_),
    .Y(_11173_));
 BUFx6f_ASAP7_75t_R _15425_ (.A(_11169_),
    .Y(_11174_));
 INVx1_ASAP7_75t_R _15426_ (.A(_01893_),
    .Y(_11175_));
 AO21x1_ASAP7_75t_R _15427_ (.A1(_11173_),
    .A2(_11174_),
    .B(_11175_),
    .Y(_11176_));
 BUFx12f_ASAP7_75t_R _15428_ (.A(_08571_),
    .Y(_11177_));
 OA221x2_ASAP7_75t_R _15429_ (.A1(_11153_),
    .A2(_11168_),
    .B1(_11135_),
    .B2(_11141_),
    .C(_11138_),
    .Y(_11178_));
 AND4x1_ASAP7_75t_R _15430_ (.A(_11149_),
    .B(_01842_),
    .C(_11136_),
    .D(_01844_),
    .Y(_11179_));
 INVx2_ASAP7_75t_R _15431_ (.A(_01885_),
    .Y(_11180_));
 INVx2_ASAP7_75t_R _15432_ (.A(_01886_),
    .Y(_11181_));
 AND4x1_ASAP7_75t_R _15433_ (.A(_11151_),
    .B(_01884_),
    .C(_11180_),
    .D(_11181_),
    .Y(_11182_));
 NOR2x1_ASAP7_75t_R _15434_ (.A(_11138_),
    .B(_11141_),
    .Y(_11183_));
 AOI221x1_ASAP7_75t_R _15435_ (.A1(_11179_),
    .A2(_11182_),
    .B1(_11158_),
    .B2(_11138_),
    .C(_11183_),
    .Y(_11184_));
 AND2x4_ASAP7_75t_R _15436_ (.A(_11144_),
    .B(_01729_),
    .Y(_11185_));
 NAND3x1_ASAP7_75t_R _15437_ (.A(_11178_),
    .B(_11184_),
    .C(_11185_),
    .Y(_11186_));
 NOR2x2_ASAP7_75t_R _15438_ (.A(_11186_),
    .B(_11169_),
    .Y(_11187_));
 NOR2x2_ASAP7_75t_R _15439_ (.A(_11177_),
    .B(_11187_),
    .Y(_11188_));
 NOR2x1_ASAP7_75t_R _15440_ (.A(_08587_),
    .B(_01739_),
    .Y(_11189_));
 BUFx3_ASAP7_75t_R _15441_ (.A(_11187_),
    .Y(_11190_));
 AO32x1_ASAP7_75t_R _15442_ (.A1(_11172_),
    .A2(_11176_),
    .A3(_11188_),
    .B1(_11189_),
    .B2(_11190_),
    .Y(_03235_));
 NAND2x1_ASAP7_75t_R _15443_ (.A(_01850_),
    .B(_11171_),
    .Y(_11191_));
 INVx1_ASAP7_75t_R _15444_ (.A(_01892_),
    .Y(_11192_));
 AO21x1_ASAP7_75t_R _15445_ (.A1(_11173_),
    .A2(_11174_),
    .B(_11192_),
    .Y(_11193_));
 NOR2x1_ASAP7_75t_R _15446_ (.A(_08587_),
    .B(_01738_),
    .Y(_11194_));
 AO32x1_ASAP7_75t_R _15447_ (.A1(_11188_),
    .A2(_11191_),
    .A3(_11193_),
    .B1(_11194_),
    .B2(_11190_),
    .Y(_03236_));
 NAND2x1_ASAP7_75t_R _15448_ (.A(_01849_),
    .B(_11171_),
    .Y(_11195_));
 INVx1_ASAP7_75t_R _15449_ (.A(_01891_),
    .Y(_11196_));
 AO21x1_ASAP7_75t_R _15450_ (.A1(_11173_),
    .A2(_11174_),
    .B(_11196_),
    .Y(_11197_));
 NOR2x1_ASAP7_75t_R _15451_ (.A(_08587_),
    .B(_01737_),
    .Y(_11198_));
 AO32x1_ASAP7_75t_R _15452_ (.A1(_11188_),
    .A2(_11195_),
    .A3(_11197_),
    .B1(_11198_),
    .B2(_11190_),
    .Y(_03237_));
 NAND2x1_ASAP7_75t_R _15453_ (.A(_01848_),
    .B(_11171_),
    .Y(_11199_));
 INVx1_ASAP7_75t_R _15454_ (.A(_01890_),
    .Y(_11200_));
 AO21x1_ASAP7_75t_R _15455_ (.A1(_11173_),
    .A2(_11174_),
    .B(_11200_),
    .Y(_11201_));
 NOR2x1_ASAP7_75t_R _15456_ (.A(_09223_),
    .B(_01736_),
    .Y(_11202_));
 AO32x1_ASAP7_75t_R _15457_ (.A1(_11188_),
    .A2(_11199_),
    .A3(_11201_),
    .B1(_11202_),
    .B2(_11190_),
    .Y(_03238_));
 NAND2x1_ASAP7_75t_R _15458_ (.A(_01847_),
    .B(_11171_),
    .Y(_11203_));
 INVx1_ASAP7_75t_R _15459_ (.A(_01889_),
    .Y(_11204_));
 AO21x1_ASAP7_75t_R _15460_ (.A1(_11173_),
    .A2(_11174_),
    .B(_11204_),
    .Y(_11205_));
 NOR2x1_ASAP7_75t_R _15461_ (.A(_09223_),
    .B(_01735_),
    .Y(_11206_));
 AO32x1_ASAP7_75t_R _15462_ (.A1(_11188_),
    .A2(_11203_),
    .A3(_11205_),
    .B1(_11206_),
    .B2(_11190_),
    .Y(_03239_));
 NAND2x1_ASAP7_75t_R _15463_ (.A(_01846_),
    .B(_11171_),
    .Y(_11207_));
 INVx1_ASAP7_75t_R _15464_ (.A(_01888_),
    .Y(_11208_));
 AO21x1_ASAP7_75t_R _15465_ (.A1(_11173_),
    .A2(_11174_),
    .B(_11208_),
    .Y(_11209_));
 NOR2x1_ASAP7_75t_R _15466_ (.A(_09223_),
    .B(_01734_),
    .Y(_11210_));
 AO32x1_ASAP7_75t_R _15467_ (.A1(_11188_),
    .A2(_11207_),
    .A3(_11209_),
    .B1(_11210_),
    .B2(_11190_),
    .Y(_03240_));
 NAND2x1_ASAP7_75t_R _15468_ (.A(_01845_),
    .B(_11171_),
    .Y(_11211_));
 INVx1_ASAP7_75t_R _15469_ (.A(_01887_),
    .Y(_11212_));
 AO21x1_ASAP7_75t_R _15470_ (.A1(_11173_),
    .A2(_11174_),
    .B(_11212_),
    .Y(_11213_));
 NOR2x1_ASAP7_75t_R _15471_ (.A(_09223_),
    .B(_01733_),
    .Y(_11214_));
 AO32x1_ASAP7_75t_R _15472_ (.A1(_11188_),
    .A2(_11211_),
    .A3(_11213_),
    .B1(_11214_),
    .B2(_11190_),
    .Y(_03241_));
 OR4x1_ASAP7_75t_R _15473_ (.A(_08684_),
    .B(_01886_),
    .C(_11187_),
    .D(_11170_),
    .Y(_11215_));
 INVx1_ASAP7_75t_R _15474_ (.A(_11215_),
    .Y(_03242_));
 OR3x1_ASAP7_75t_R _15475_ (.A(_11180_),
    .B(_11187_),
    .C(_11170_),
    .Y(_11216_));
 NAND2x1_ASAP7_75t_R _15476_ (.A(_01731_),
    .B(_11190_),
    .Y(_11217_));
 AND3x1_ASAP7_75t_R _15477_ (.A(_10809_),
    .B(_11216_),
    .C(_11217_),
    .Y(_03243_));
 OR3x1_ASAP7_75t_R _15478_ (.A(_01730_),
    .B(_11186_),
    .C(_11174_),
    .Y(_11218_));
 OR3x1_ASAP7_75t_R _15479_ (.A(_01884_),
    .B(_11187_),
    .C(_11171_),
    .Y(_11219_));
 AOI21x1_ASAP7_75t_R _15480_ (.A1(_11218_),
    .A2(_11219_),
    .B(_09081_),
    .Y(_03244_));
 NOR2x1_ASAP7_75t_R _15481_ (.A(_11144_),
    .B(_11150_),
    .Y(_11220_));
 OAI21x1_ASAP7_75t_R _15482_ (.A1(_01882_),
    .A2(_01883_),
    .B(_11153_),
    .Y(_11221_));
 OA33x2_ASAP7_75t_R _15483_ (.A1(_11135_),
    .A2(_11158_),
    .A3(_11142_),
    .B1(_11146_),
    .B2(_11220_),
    .B3(_11221_),
    .Y(_11222_));
 NOR2x1_ASAP7_75t_R _15484_ (.A(_10716_),
    .B(_11222_),
    .Y(_03245_));
 INVx1_ASAP7_75t_R _15485_ (.A(_11173_),
    .Y(_11223_));
 NOR2x1_ASAP7_75t_R _15486_ (.A(_11223_),
    .B(_11174_),
    .Y(_11224_));
 AOI21x1_ASAP7_75t_R _15487_ (.A1(_11186_),
    .A2(_11224_),
    .B(_09081_),
    .Y(_03246_));
 NAND2x1_ASAP7_75t_R _15488_ (.A(_01839_),
    .B(_11171_),
    .Y(_11225_));
 INVx1_ASAP7_75t_R _15489_ (.A(_01881_),
    .Y(_11226_));
 AO21x1_ASAP7_75t_R _15490_ (.A1(_11173_),
    .A2(_11174_),
    .B(_11226_),
    .Y(_11227_));
 NOR2x1_ASAP7_75t_R _15491_ (.A(_09223_),
    .B(_01727_),
    .Y(_11228_));
 AO32x1_ASAP7_75t_R _15492_ (.A1(_11188_),
    .A2(_11225_),
    .A3(_11227_),
    .B1(_11228_),
    .B2(_11190_),
    .Y(_03247_));
 NAND2x1_ASAP7_75t_R _15493_ (.A(_01838_),
    .B(_11171_),
    .Y(_11229_));
 INVx1_ASAP7_75t_R _15494_ (.A(_01880_),
    .Y(_11230_));
 AO21x1_ASAP7_75t_R _15495_ (.A1(_11173_),
    .A2(_11169_),
    .B(_11230_),
    .Y(_11231_));
 NOR2x1_ASAP7_75t_R _15496_ (.A(_09223_),
    .B(_02356_),
    .Y(_11232_));
 AO32x1_ASAP7_75t_R _15497_ (.A1(_11188_),
    .A2(_11229_),
    .A3(_11231_),
    .B1(_11232_),
    .B2(_11190_),
    .Y(_03248_));
 OA21x2_ASAP7_75t_R _15498_ (.A1(_11144_),
    .A2(_11164_),
    .B(_11165_),
    .Y(_11233_));
 INVx1_ASAP7_75t_R _15499_ (.A(_11141_),
    .Y(_11234_));
 AO221x1_ASAP7_75t_R _15500_ (.A1(_11179_),
    .A2(_11159_),
    .B1(_11163_),
    .B2(_11233_),
    .C(_11234_),
    .Y(_11235_));
 BUFx6f_ASAP7_75t_R _15501_ (.A(_11235_),
    .Y(_11236_));
 AOI221x1_ASAP7_75t_R _15502_ (.A1(_11179_),
    .A2(_11158_),
    .B1(_11137_),
    .B2(_11182_),
    .C(_11138_),
    .Y(_11237_));
 NAND3x1_ASAP7_75t_R _15503_ (.A(_11184_),
    .B(_11185_),
    .C(_11237_),
    .Y(_11238_));
 AO211x2_ASAP7_75t_R _15504_ (.A1(_11182_),
    .A2(_11222_),
    .B(_11236_),
    .C(_11238_),
    .Y(_11239_));
 BUFx12f_ASAP7_75t_R _15505_ (.A(_11239_),
    .Y(_11240_));
 NOR2x1_ASAP7_75t_R _15506_ (.A(_01739_),
    .B(_11240_),
    .Y(_11241_));
 BUFx6f_ASAP7_75t_R _15507_ (.A(_11236_),
    .Y(_11242_));
 BUFx6f_ASAP7_75t_R _15508_ (.A(_11239_),
    .Y(_11243_));
 BUFx6f_ASAP7_75t_R _15509_ (.A(_11236_),
    .Y(_11244_));
 NAND2x1_ASAP7_75t_R _15510_ (.A(_01851_),
    .B(_11244_),
    .Y(_11245_));
 OA211x2_ASAP7_75t_R _15511_ (.A1(_11175_),
    .A2(_11242_),
    .B(_11243_),
    .C(_11245_),
    .Y(_11246_));
 OA21x2_ASAP7_75t_R _15512_ (.A1(_11241_),
    .A2(_11246_),
    .B(_11067_),
    .Y(_03249_));
 NOR2x1_ASAP7_75t_R _15513_ (.A(_01738_),
    .B(_11240_),
    .Y(_11247_));
 NAND2x1_ASAP7_75t_R _15514_ (.A(_01850_),
    .B(_11244_),
    .Y(_11248_));
 OA211x2_ASAP7_75t_R _15515_ (.A1(_11192_),
    .A2(_11242_),
    .B(_11243_),
    .C(_11248_),
    .Y(_11249_));
 OA21x2_ASAP7_75t_R _15516_ (.A1(_11247_),
    .A2(_11249_),
    .B(_11067_),
    .Y(_03250_));
 NOR2x1_ASAP7_75t_R _15517_ (.A(_01737_),
    .B(_11240_),
    .Y(_11250_));
 NAND2x1_ASAP7_75t_R _15518_ (.A(_01849_),
    .B(_11244_),
    .Y(_11251_));
 OA211x2_ASAP7_75t_R _15519_ (.A1(_11196_),
    .A2(_11242_),
    .B(_11243_),
    .C(_11251_),
    .Y(_11252_));
 BUFx6f_ASAP7_75t_R _15520_ (.A(_09229_),
    .Y(_11253_));
 OA21x2_ASAP7_75t_R _15521_ (.A1(_11250_),
    .A2(_11252_),
    .B(_11253_),
    .Y(_03251_));
 NOR2x1_ASAP7_75t_R _15522_ (.A(_01736_),
    .B(_11240_),
    .Y(_11254_));
 NAND2x1_ASAP7_75t_R _15523_ (.A(_01848_),
    .B(_11244_),
    .Y(_11255_));
 OA211x2_ASAP7_75t_R _15524_ (.A1(_11200_),
    .A2(_11242_),
    .B(_11243_),
    .C(_11255_),
    .Y(_11256_));
 OA21x2_ASAP7_75t_R _15525_ (.A1(_11254_),
    .A2(_11256_),
    .B(_11253_),
    .Y(_03252_));
 NOR2x1_ASAP7_75t_R _15526_ (.A(_01735_),
    .B(_11240_),
    .Y(_11257_));
 NAND2x1_ASAP7_75t_R _15527_ (.A(_01847_),
    .B(_11244_),
    .Y(_11258_));
 OA211x2_ASAP7_75t_R _15528_ (.A1(_11204_),
    .A2(_11242_),
    .B(_11243_),
    .C(_11258_),
    .Y(_11259_));
 OA21x2_ASAP7_75t_R _15529_ (.A1(_11257_),
    .A2(_11259_),
    .B(_11253_),
    .Y(_03253_));
 NOR2x1_ASAP7_75t_R _15530_ (.A(_01734_),
    .B(_11240_),
    .Y(_11260_));
 NAND2x1_ASAP7_75t_R _15531_ (.A(_01846_),
    .B(_11244_),
    .Y(_11261_));
 OA211x2_ASAP7_75t_R _15532_ (.A1(_11208_),
    .A2(_11242_),
    .B(_11243_),
    .C(_11261_),
    .Y(_11262_));
 OA21x2_ASAP7_75t_R _15533_ (.A1(_11260_),
    .A2(_11262_),
    .B(_11253_),
    .Y(_03254_));
 NOR2x1_ASAP7_75t_R _15534_ (.A(_01733_),
    .B(_11240_),
    .Y(_11263_));
 NAND2x1_ASAP7_75t_R _15535_ (.A(_01845_),
    .B(_11236_),
    .Y(_11264_));
 OA211x2_ASAP7_75t_R _15536_ (.A1(_11212_),
    .A2(_11242_),
    .B(_11243_),
    .C(_11264_),
    .Y(_11265_));
 OA21x2_ASAP7_75t_R _15537_ (.A1(_11263_),
    .A2(_11265_),
    .B(_11253_),
    .Y(_03255_));
 NOR2x1_ASAP7_75t_R _15538_ (.A(_11181_),
    .B(_11242_),
    .Y(_11266_));
 AO21x1_ASAP7_75t_R _15539_ (.A1(_01844_),
    .A2(_11242_),
    .B(_11266_),
    .Y(_11267_));
 AOI21x1_ASAP7_75t_R _15540_ (.A1(_11240_),
    .A2(_11267_),
    .B(_09081_),
    .Y(_03256_));
 NOR2x1_ASAP7_75t_R _15541_ (.A(_01731_),
    .B(_11240_),
    .Y(_11268_));
 NAND2x1_ASAP7_75t_R _15542_ (.A(_01843_),
    .B(_11236_),
    .Y(_11269_));
 OA211x2_ASAP7_75t_R _15543_ (.A1(_11180_),
    .A2(_11244_),
    .B(_11243_),
    .C(_11269_),
    .Y(_11270_));
 OA21x2_ASAP7_75t_R _15544_ (.A1(_11268_),
    .A2(_11270_),
    .B(_11253_),
    .Y(_03257_));
 NOR2x1_ASAP7_75t_R _15545_ (.A(_01730_),
    .B(_11240_),
    .Y(_11271_));
 NAND2x1_ASAP7_75t_R _15546_ (.A(_01842_),
    .B(_11236_),
    .Y(_11272_));
 OA211x2_ASAP7_75t_R _15547_ (.A1(_11134_),
    .A2(_11244_),
    .B(_11239_),
    .C(_11272_),
    .Y(_11273_));
 OA21x2_ASAP7_75t_R _15548_ (.A1(_11271_),
    .A2(_11273_),
    .B(_11253_),
    .Y(_03258_));
 AND2x2_ASAP7_75t_R _15549_ (.A(_11179_),
    .B(_11141_),
    .Y(_11274_));
 AOI22x1_ASAP7_75t_R _15550_ (.A1(_11163_),
    .A2(_11166_),
    .B1(_11274_),
    .B2(_11159_),
    .Y(_11275_));
 NOR2x1_ASAP7_75t_R _15551_ (.A(_10716_),
    .B(_11275_),
    .Y(_03259_));
 AOI21x1_ASAP7_75t_R _15552_ (.A1(_11182_),
    .A2(_11222_),
    .B(_11242_),
    .Y(_11276_));
 AOI21x1_ASAP7_75t_R _15553_ (.A1(_11276_),
    .A2(_11238_),
    .B(_09081_),
    .Y(_03260_));
 NOR2x1_ASAP7_75t_R _15554_ (.A(_01727_),
    .B(_11243_),
    .Y(_11277_));
 NAND2x1_ASAP7_75t_R _15555_ (.A(_01839_),
    .B(_11236_),
    .Y(_11278_));
 OA211x2_ASAP7_75t_R _15556_ (.A1(_11226_),
    .A2(_11244_),
    .B(_11239_),
    .C(_11278_),
    .Y(_11279_));
 OA21x2_ASAP7_75t_R _15557_ (.A1(_11277_),
    .A2(_11279_),
    .B(_11253_),
    .Y(_03261_));
 NOR2x1_ASAP7_75t_R _15558_ (.A(_02356_),
    .B(_11243_),
    .Y(_11280_));
 NAND2x1_ASAP7_75t_R _15559_ (.A(_01838_),
    .B(_11236_),
    .Y(_11281_));
 OA211x2_ASAP7_75t_R _15560_ (.A1(_11230_),
    .A2(_11244_),
    .B(_11239_),
    .C(_11281_),
    .Y(_11282_));
 OA21x2_ASAP7_75t_R _15561_ (.A1(_11280_),
    .A2(_11282_),
    .B(_11253_),
    .Y(_03262_));
 AO221x1_ASAP7_75t_R _15562_ (.A1(_11163_),
    .A2(_11166_),
    .B1(_11274_),
    .B2(_11159_),
    .C(_11137_),
    .Y(_11283_));
 AOI21x1_ASAP7_75t_R _15563_ (.A1(_11153_),
    .A2(_11222_),
    .B(_11283_),
    .Y(_11284_));
 BUFx6f_ASAP7_75t_R _15564_ (.A(_11284_),
    .Y(_11285_));
 NAND2x1_ASAP7_75t_R _15565_ (.A(_01851_),
    .B(_11285_),
    .Y(_11286_));
 BUFx6f_ASAP7_75t_R _15566_ (.A(_11284_),
    .Y(_11287_));
 OR2x2_ASAP7_75t_R _15567_ (.A(_11175_),
    .B(_11287_),
    .Y(_11288_));
 OA21x2_ASAP7_75t_R _15568_ (.A1(_11178_),
    .A2(_11237_),
    .B(_11184_),
    .Y(_11289_));
 AOI21x1_ASAP7_75t_R _15569_ (.A1(_01729_),
    .A2(_11289_),
    .B(_01728_),
    .Y(_11290_));
 NOR2x1_ASAP7_75t_R _15570_ (.A(_08572_),
    .B(_11290_),
    .Y(_11291_));
 BUFx3_ASAP7_75t_R _15571_ (.A(_11290_),
    .Y(_11292_));
 AO32x1_ASAP7_75t_R _15572_ (.A1(_11286_),
    .A2(_11288_),
    .A3(_11291_),
    .B1(_11292_),
    .B2(_11189_),
    .Y(_03263_));
 BUFx6f_ASAP7_75t_R _15573_ (.A(_11291_),
    .Y(_11293_));
 NAND2x1_ASAP7_75t_R _15574_ (.A(_01850_),
    .B(_11285_),
    .Y(_11294_));
 OR2x2_ASAP7_75t_R _15575_ (.A(_11192_),
    .B(_11287_),
    .Y(_11295_));
 AO32x1_ASAP7_75t_R _15576_ (.A1(_11293_),
    .A2(_11294_),
    .A3(_11295_),
    .B1(_11292_),
    .B2(_11194_),
    .Y(_03264_));
 NAND2x1_ASAP7_75t_R _15577_ (.A(_01849_),
    .B(_11285_),
    .Y(_11296_));
 OR2x2_ASAP7_75t_R _15578_ (.A(_11196_),
    .B(_11287_),
    .Y(_11297_));
 AO32x1_ASAP7_75t_R _15579_ (.A1(_11293_),
    .A2(_11296_),
    .A3(_11297_),
    .B1(_11292_),
    .B2(_11198_),
    .Y(_03265_));
 NAND2x1_ASAP7_75t_R _15580_ (.A(_01848_),
    .B(_11285_),
    .Y(_11298_));
 OR2x2_ASAP7_75t_R _15581_ (.A(_11200_),
    .B(_11287_),
    .Y(_11299_));
 AO32x1_ASAP7_75t_R _15582_ (.A1(_11293_),
    .A2(_11298_),
    .A3(_11299_),
    .B1(_11292_),
    .B2(_11202_),
    .Y(_03266_));
 NAND2x1_ASAP7_75t_R _15583_ (.A(_01847_),
    .B(_11285_),
    .Y(_11300_));
 OR2x2_ASAP7_75t_R _15584_ (.A(_11204_),
    .B(_11287_),
    .Y(_11301_));
 AO32x1_ASAP7_75t_R _15585_ (.A1(_11293_),
    .A2(_11300_),
    .A3(_11301_),
    .B1(_11292_),
    .B2(_11206_),
    .Y(_03267_));
 NAND2x1_ASAP7_75t_R _15586_ (.A(_01846_),
    .B(_11285_),
    .Y(_11302_));
 OR2x2_ASAP7_75t_R _15587_ (.A(_11208_),
    .B(_11287_),
    .Y(_11303_));
 AO32x1_ASAP7_75t_R _15588_ (.A1(_11293_),
    .A2(_11302_),
    .A3(_11303_),
    .B1(_11292_),
    .B2(_11210_),
    .Y(_03268_));
 NAND2x1_ASAP7_75t_R _15589_ (.A(_01845_),
    .B(_11285_),
    .Y(_11304_));
 OR2x2_ASAP7_75t_R _15590_ (.A(_11212_),
    .B(_11287_),
    .Y(_11305_));
 AO32x1_ASAP7_75t_R _15591_ (.A1(_11293_),
    .A2(_11304_),
    .A3(_11305_),
    .B1(_11290_),
    .B2(_11214_),
    .Y(_03269_));
 NAND2x1_ASAP7_75t_R _15592_ (.A(_01844_),
    .B(_11285_),
    .Y(_11306_));
 OR2x2_ASAP7_75t_R _15593_ (.A(_11181_),
    .B(_11287_),
    .Y(_11307_));
 NOR2x1_ASAP7_75t_R _15594_ (.A(_09934_),
    .B(_11138_),
    .Y(_11308_));
 AO32x1_ASAP7_75t_R _15595_ (.A1(_11293_),
    .A2(_11306_),
    .A3(_11307_),
    .B1(_11308_),
    .B2(_11292_),
    .Y(_03270_));
 NAND2x1_ASAP7_75t_R _15596_ (.A(_01843_),
    .B(_11285_),
    .Y(_11309_));
 OR2x2_ASAP7_75t_R _15597_ (.A(_11180_),
    .B(_11284_),
    .Y(_11310_));
 NOR2x1_ASAP7_75t_R _15598_ (.A(_09934_),
    .B(_01731_),
    .Y(_11311_));
 AO32x1_ASAP7_75t_R _15599_ (.A1(_11293_),
    .A2(_11309_),
    .A3(_11310_),
    .B1(_11311_),
    .B2(_11292_),
    .Y(_03271_));
 NAND2x1_ASAP7_75t_R _15600_ (.A(_01842_),
    .B(_11285_),
    .Y(_11312_));
 OR2x2_ASAP7_75t_R _15601_ (.A(_11134_),
    .B(_11284_),
    .Y(_11313_));
 NOR2x1_ASAP7_75t_R _15602_ (.A(_09934_),
    .B(_01730_),
    .Y(_11314_));
 AO32x1_ASAP7_75t_R _15603_ (.A1(_11293_),
    .A2(_11312_),
    .A3(_11313_),
    .B1(_11314_),
    .B2(_11292_),
    .Y(_03272_));
 OR4x1_ASAP7_75t_R _15604_ (.A(_08684_),
    .B(_01728_),
    .C(_11156_),
    .D(_11289_),
    .Y(_11315_));
 INVx1_ASAP7_75t_R _15605_ (.A(_11315_),
    .Y(_03273_));
 AO22x1_ASAP7_75t_R _15606_ (.A1(_11165_),
    .A2(_11275_),
    .B1(_11222_),
    .B2(_11153_),
    .Y(_11316_));
 OA21x2_ASAP7_75t_R _15607_ (.A1(_11292_),
    .A2(_11316_),
    .B(_11253_),
    .Y(_03274_));
 NAND2x1_ASAP7_75t_R _15608_ (.A(_01839_),
    .B(_11287_),
    .Y(_11317_));
 OR2x2_ASAP7_75t_R _15609_ (.A(_11226_),
    .B(_11284_),
    .Y(_11318_));
 AO32x1_ASAP7_75t_R _15610_ (.A1(_11293_),
    .A2(_11317_),
    .A3(_11318_),
    .B1(_11290_),
    .B2(_11228_),
    .Y(_03275_));
 NAND2x1_ASAP7_75t_R _15611_ (.A(_01838_),
    .B(_11287_),
    .Y(_11319_));
 OR2x2_ASAP7_75t_R _15612_ (.A(_11230_),
    .B(_11284_),
    .Y(_11320_));
 AO32x1_ASAP7_75t_R _15613_ (.A1(_11291_),
    .A2(_11319_),
    .A3(_11320_),
    .B1(_11290_),
    .B2(_11232_),
    .Y(_03276_));
 AND2x2_ASAP7_75t_R _15614_ (.A(_10927_),
    .B(_00014_),
    .Y(_03277_));
 BUFx6f_ASAP7_75t_R _15615_ (.A(_02351_),
    .Y(_11321_));
 INVx2_ASAP7_75t_R _15616_ (.A(_02354_),
    .Y(_11322_));
 BUFx6f_ASAP7_75t_R _15617_ (.A(_01756_),
    .Y(_11323_));
 AO221x1_ASAP7_75t_R _15618_ (.A1(_01757_),
    .A2(_01758_),
    .B1(_11321_),
    .B2(_11322_),
    .C(_11323_),
    .Y(_11324_));
 INVx1_ASAP7_75t_R _15619_ (.A(_00014_),
    .Y(_11325_));
 NOR2x1_ASAP7_75t_R _15620_ (.A(_11323_),
    .B(_01758_),
    .Y(_11326_));
 AOI21x1_ASAP7_75t_R _15621_ (.A1(_11325_),
    .A2(_11326_),
    .B(_11322_),
    .Y(_11327_));
 AO21x2_ASAP7_75t_R _15622_ (.A1(_02353_),
    .A2(_11324_),
    .B(_11327_),
    .Y(_11328_));
 BUFx6f_ASAP7_75t_R _15623_ (.A(_01798_),
    .Y(_11329_));
 BUFx6f_ASAP7_75t_R _15624_ (.A(_01800_),
    .Y(_11330_));
 OR2x6_ASAP7_75t_R _15625_ (.A(_11329_),
    .B(_11330_),
    .Y(_11331_));
 BUFx6f_ASAP7_75t_R _15626_ (.A(_01799_),
    .Y(_11332_));
 AO211x2_ASAP7_75t_R _15627_ (.A1(_11321_),
    .A2(_02353_),
    .B(_02354_),
    .C(_01758_),
    .Y(_11333_));
 AO21x2_ASAP7_75t_R _15628_ (.A1(_01757_),
    .A2(_11333_),
    .B(_11323_),
    .Y(_11334_));
 INVx1_ASAP7_75t_R _15629_ (.A(_11330_),
    .Y(_11335_));
 OR3x2_ASAP7_75t_R _15630_ (.A(_11329_),
    .B(_11335_),
    .C(_01801_),
    .Y(_11336_));
 OA22x2_ASAP7_75t_R _15631_ (.A1(_11329_),
    .A2(_11332_),
    .B1(_11334_),
    .B2(_11336_),
    .Y(_11337_));
 INVx2_ASAP7_75t_R _15632_ (.A(_11323_),
    .Y(_11338_));
 AND2x4_ASAP7_75t_R _15633_ (.A(_01758_),
    .B(_01759_),
    .Y(_11339_));
 NAND2x1_ASAP7_75t_R _15634_ (.A(_11338_),
    .B(_11339_),
    .Y(_11340_));
 INVx1_ASAP7_75t_R _15635_ (.A(_11321_),
    .Y(_11341_));
 OR2x2_ASAP7_75t_R _15636_ (.A(_02354_),
    .B(_11330_),
    .Y(_11342_));
 AO21x1_ASAP7_75t_R _15637_ (.A1(_11341_),
    .A2(_02353_),
    .B(_11342_),
    .Y(_11343_));
 NOR2x1_ASAP7_75t_R _15638_ (.A(_11323_),
    .B(_01757_),
    .Y(_11344_));
 AOI211x1_ASAP7_75t_R _15639_ (.A1(_11332_),
    .A2(_11343_),
    .B(_11344_),
    .C(_11329_),
    .Y(_11345_));
 NOR2x1_ASAP7_75t_R _15640_ (.A(_11340_),
    .B(_11345_),
    .Y(_11346_));
 OA211x2_ASAP7_75t_R _15641_ (.A1(_11328_),
    .A2(_11331_),
    .B(_11337_),
    .C(_11346_),
    .Y(_11347_));
 BUFx6f_ASAP7_75t_R _15642_ (.A(_11347_),
    .Y(_11348_));
 NOR2x1_ASAP7_75t_R _15643_ (.A(_11329_),
    .B(_11332_),
    .Y(_11349_));
 AOI211x1_ASAP7_75t_R _15644_ (.A1(_02353_),
    .A2(_11324_),
    .B(_11327_),
    .C(_11331_),
    .Y(_11350_));
 NOR2x1_ASAP7_75t_R _15645_ (.A(_11334_),
    .B(_11336_),
    .Y(_11351_));
 OR5x2_ASAP7_75t_R _15646_ (.A(_11349_),
    .B(_11340_),
    .C(_11345_),
    .D(_11350_),
    .E(_11351_),
    .Y(_11352_));
 AND2x2_ASAP7_75t_R _15647_ (.A(_01809_),
    .B(_11352_),
    .Y(_11353_));
 AO21x1_ASAP7_75t_R _15648_ (.A1(_01767_),
    .A2(_11348_),
    .B(_11353_),
    .Y(_11354_));
 INVx1_ASAP7_75t_R _15649_ (.A(_11329_),
    .Y(_11355_));
 INVx1_ASAP7_75t_R _15650_ (.A(_01801_),
    .Y(_11356_));
 AO32x1_ASAP7_75t_R _15651_ (.A1(_11338_),
    .A2(_11321_),
    .A3(_11339_),
    .B1(_11355_),
    .B2(_11356_),
    .Y(_11357_));
 INVx1_ASAP7_75t_R _15652_ (.A(_01757_),
    .Y(_11358_));
 OA211x2_ASAP7_75t_R _15653_ (.A1(_11358_),
    .A2(_11339_),
    .B(_11330_),
    .C(_11338_),
    .Y(_11359_));
 INVx1_ASAP7_75t_R _15654_ (.A(_02353_),
    .Y(_11360_));
 AO211x2_ASAP7_75t_R _15655_ (.A1(_11321_),
    .A2(_11349_),
    .B(_11360_),
    .C(_02354_),
    .Y(_11361_));
 AND2x2_ASAP7_75t_R _15656_ (.A(_11329_),
    .B(_11321_),
    .Y(_11362_));
 OA211x2_ASAP7_75t_R _15657_ (.A1(_11349_),
    .A2(_11362_),
    .B(_11339_),
    .C(_11338_),
    .Y(_11363_));
 AOI211x1_ASAP7_75t_R _15658_ (.A1(_11357_),
    .A2(_11359_),
    .B(_11361_),
    .C(_11363_),
    .Y(_11364_));
 AND2x4_ASAP7_75t_R _15659_ (.A(_11321_),
    .B(_11364_),
    .Y(_11365_));
 OA221x2_ASAP7_75t_R _15660_ (.A1(_11340_),
    .A2(_11345_),
    .B1(_11328_),
    .B2(_11331_),
    .C(_11337_),
    .Y(_11366_));
 AO21x2_ASAP7_75t_R _15661_ (.A1(_11365_),
    .A2(_11366_),
    .B(_08641_),
    .Y(_11367_));
 BUFx12f_ASAP7_75t_R _15662_ (.A(_11367_),
    .Y(_11368_));
 NAND2x1_ASAP7_75t_R _15663_ (.A(_11365_),
    .B(_11366_),
    .Y(_11369_));
 BUFx6f_ASAP7_75t_R _15664_ (.A(_11369_),
    .Y(_11370_));
 OR3x1_ASAP7_75t_R _15665_ (.A(_11126_),
    .B(_02343_),
    .C(_11370_),
    .Y(_11371_));
 OAI21x1_ASAP7_75t_R _15666_ (.A1(_11354_),
    .A2(_11368_),
    .B(_11371_),
    .Y(_03278_));
 BUFx6f_ASAP7_75t_R _15667_ (.A(_11352_),
    .Y(_11372_));
 AND2x2_ASAP7_75t_R _15668_ (.A(_01808_),
    .B(_11372_),
    .Y(_11373_));
 AO21x1_ASAP7_75t_R _15669_ (.A1(_01766_),
    .A2(_11348_),
    .B(_11373_),
    .Y(_11374_));
 OR3x1_ASAP7_75t_R _15670_ (.A(_11126_),
    .B(_02344_),
    .C(_11370_),
    .Y(_11375_));
 OAI21x1_ASAP7_75t_R _15671_ (.A1(_11368_),
    .A2(_11374_),
    .B(_11375_),
    .Y(_03279_));
 AND2x2_ASAP7_75t_R _15672_ (.A(_01807_),
    .B(_11372_),
    .Y(_11376_));
 AO21x1_ASAP7_75t_R _15673_ (.A1(_01765_),
    .A2(_11348_),
    .B(_11376_),
    .Y(_11377_));
 OR3x1_ASAP7_75t_R _15674_ (.A(_11126_),
    .B(_02345_),
    .C(_11370_),
    .Y(_11378_));
 OAI21x1_ASAP7_75t_R _15675_ (.A1(_11368_),
    .A2(_11377_),
    .B(_11378_),
    .Y(_03280_));
 AND2x2_ASAP7_75t_R _15676_ (.A(_01806_),
    .B(_11372_),
    .Y(_11379_));
 AO21x1_ASAP7_75t_R _15677_ (.A1(_01764_),
    .A2(_11348_),
    .B(_11379_),
    .Y(_11380_));
 OR3x1_ASAP7_75t_R _15678_ (.A(_11126_),
    .B(_02346_),
    .C(_11370_),
    .Y(_11381_));
 OAI21x1_ASAP7_75t_R _15679_ (.A1(_11368_),
    .A2(_11380_),
    .B(_11381_),
    .Y(_03281_));
 AND2x2_ASAP7_75t_R _15680_ (.A(_01805_),
    .B(_11372_),
    .Y(_11382_));
 AO21x1_ASAP7_75t_R _15681_ (.A1(_01763_),
    .A2(_11348_),
    .B(_11382_),
    .Y(_11383_));
 OR3x1_ASAP7_75t_R _15682_ (.A(_11126_),
    .B(_02347_),
    .C(_11370_),
    .Y(_11384_));
 OAI21x1_ASAP7_75t_R _15683_ (.A1(_11368_),
    .A2(_11383_),
    .B(_11384_),
    .Y(_03282_));
 AND2x2_ASAP7_75t_R _15684_ (.A(_01804_),
    .B(_11372_),
    .Y(_11385_));
 AO21x1_ASAP7_75t_R _15685_ (.A1(_01762_),
    .A2(_11348_),
    .B(_11385_),
    .Y(_11386_));
 OR3x1_ASAP7_75t_R _15686_ (.A(_11126_),
    .B(_02348_),
    .C(_11370_),
    .Y(_11387_));
 OAI21x1_ASAP7_75t_R _15687_ (.A1(_11368_),
    .A2(_11386_),
    .B(_11387_),
    .Y(_03283_));
 AND2x2_ASAP7_75t_R _15688_ (.A(_01803_),
    .B(_11372_),
    .Y(_11388_));
 AO21x1_ASAP7_75t_R _15689_ (.A1(_01761_),
    .A2(_11348_),
    .B(_11388_),
    .Y(_11389_));
 OR3x1_ASAP7_75t_R _15690_ (.A(_11126_),
    .B(_02349_),
    .C(_11370_),
    .Y(_11390_));
 OAI21x1_ASAP7_75t_R _15691_ (.A1(_11368_),
    .A2(_11389_),
    .B(_11390_),
    .Y(_03284_));
 AND2x2_ASAP7_75t_R _15692_ (.A(_01802_),
    .B(_11372_),
    .Y(_11391_));
 AO21x1_ASAP7_75t_R _15693_ (.A1(_01760_),
    .A2(_11348_),
    .B(_11391_),
    .Y(_11392_));
 OR3x1_ASAP7_75t_R _15694_ (.A(_11126_),
    .B(_02350_),
    .C(_11370_),
    .Y(_11393_));
 OAI21x1_ASAP7_75t_R _15695_ (.A1(_11368_),
    .A2(_11392_),
    .B(_11393_),
    .Y(_03285_));
 AND4x1_ASAP7_75t_R _15696_ (.A(_08999_),
    .B(_11356_),
    .C(_11370_),
    .D(_11372_),
    .Y(_03286_));
 INVx1_ASAP7_75t_R _15697_ (.A(_02352_),
    .Y(_11394_));
 AND3x1_ASAP7_75t_R _15698_ (.A(_11394_),
    .B(_11365_),
    .C(_11366_),
    .Y(_11395_));
 AND3x1_ASAP7_75t_R _15699_ (.A(_11335_),
    .B(_11369_),
    .C(_11372_),
    .Y(_11396_));
 BUFx12f_ASAP7_75t_R _15700_ (.A(_09229_),
    .Y(_11397_));
 OA21x2_ASAP7_75t_R _15701_ (.A1(_11395_),
    .A2(_11396_),
    .B(_11397_),
    .Y(_03287_));
 NAND2x1_ASAP7_75t_R _15702_ (.A(_11330_),
    .B(_11356_),
    .Y(_11398_));
 OAI22x1_ASAP7_75t_R _15703_ (.A1(_11330_),
    .A2(_11328_),
    .B1(_11334_),
    .B2(_11398_),
    .Y(_11399_));
 AND4x1_ASAP7_75t_R _15704_ (.A(_08999_),
    .B(_11355_),
    .C(_11332_),
    .D(_11399_),
    .Y(_03288_));
 INVx1_ASAP7_75t_R _15705_ (.A(_11365_),
    .Y(_11400_));
 AOI21x1_ASAP7_75t_R _15706_ (.A1(_11400_),
    .A2(_11366_),
    .B(_09081_),
    .Y(_03289_));
 AND2x2_ASAP7_75t_R _15707_ (.A(_01797_),
    .B(_11372_),
    .Y(_11401_));
 AO21x1_ASAP7_75t_R _15708_ (.A1(_01755_),
    .A2(_11348_),
    .B(_11401_),
    .Y(_11402_));
 OR3x1_ASAP7_75t_R _15709_ (.A(_11126_),
    .B(_02355_),
    .C(_11370_),
    .Y(_11403_));
 OAI21x1_ASAP7_75t_R _15710_ (.A1(_11368_),
    .A2(_11402_),
    .B(_11403_),
    .Y(_03290_));
 AND2x2_ASAP7_75t_R _15711_ (.A(_01796_),
    .B(_11352_),
    .Y(_11404_));
 AO21x1_ASAP7_75t_R _15712_ (.A1(_01754_),
    .A2(_11348_),
    .B(_11404_),
    .Y(_11405_));
 BUFx6f_ASAP7_75t_R _15713_ (.A(_08656_),
    .Y(_11406_));
 OR3x1_ASAP7_75t_R _15714_ (.A(_11406_),
    .B(_02342_),
    .C(_11369_),
    .Y(_11407_));
 OAI21x1_ASAP7_75t_R _15715_ (.A1(_11368_),
    .A2(_11405_),
    .B(_11407_),
    .Y(_03291_));
 OR2x2_ASAP7_75t_R _15716_ (.A(_11323_),
    .B(_01757_),
    .Y(_11408_));
 OA211x2_ASAP7_75t_R _15717_ (.A1(_11326_),
    .A2(_11336_),
    .B(_11341_),
    .C(_11408_),
    .Y(_11409_));
 NAND2x1_ASAP7_75t_R _15718_ (.A(_11332_),
    .B(_11330_),
    .Y(_11410_));
 AND2x2_ASAP7_75t_R _15719_ (.A(_02354_),
    .B(_00014_),
    .Y(_11411_));
 AO32x1_ASAP7_75t_R _15720_ (.A1(_11322_),
    .A2(_11321_),
    .A3(_11410_),
    .B1(_11411_),
    .B2(_11335_),
    .Y(_11412_));
 AO22x2_ASAP7_75t_R _15721_ (.A1(_11322_),
    .A2(_11360_),
    .B1(_11412_),
    .B2(_11355_),
    .Y(_11413_));
 AOI211x1_ASAP7_75t_R _15722_ (.A1(_11332_),
    .A2(_11343_),
    .B(_11340_),
    .C(_11329_),
    .Y(_11414_));
 AO221x1_ASAP7_75t_R _15723_ (.A1(_11338_),
    .A2(_11358_),
    .B1(_11326_),
    .B2(_11413_),
    .C(_11414_),
    .Y(_11415_));
 AOI21x1_ASAP7_75t_R _15724_ (.A1(_01757_),
    .A2(_11333_),
    .B(_11323_),
    .Y(_11416_));
 AOI21x1_ASAP7_75t_R _15725_ (.A1(_11332_),
    .A2(_11416_),
    .B(_11336_),
    .Y(_11417_));
 NOR2x1_ASAP7_75t_R _15726_ (.A(_11415_),
    .B(_11417_),
    .Y(_11418_));
 AND3x4_ASAP7_75t_R _15727_ (.A(_11364_),
    .B(_11409_),
    .C(_11418_),
    .Y(_11419_));
 BUFx12f_ASAP7_75t_R _15728_ (.A(_11419_),
    .Y(_11420_));
 BUFx6f_ASAP7_75t_R _15729_ (.A(_11415_),
    .Y(_11421_));
 AOI211x1_ASAP7_75t_R _15730_ (.A1(_11326_),
    .A2(_11413_),
    .B(_11414_),
    .C(_11344_),
    .Y(_11422_));
 BUFx6f_ASAP7_75t_R _15731_ (.A(_11422_),
    .Y(_11423_));
 AO21x1_ASAP7_75t_R _15732_ (.A1(_01809_),
    .A2(_11423_),
    .B(_10826_),
    .Y(_11424_));
 AO21x1_ASAP7_75t_R _15733_ (.A1(_01767_),
    .A2(_11421_),
    .B(_11424_),
    .Y(_11425_));
 NAND2x1_ASAP7_75t_R _15734_ (.A(_11364_),
    .B(_11409_),
    .Y(_11426_));
 OR3x2_ASAP7_75t_R _15735_ (.A(_11426_),
    .B(_11415_),
    .C(_11417_),
    .Y(_11427_));
 BUFx6f_ASAP7_75t_R _15736_ (.A(_11427_),
    .Y(_11428_));
 OR3x1_ASAP7_75t_R _15737_ (.A(_11406_),
    .B(_02343_),
    .C(_11428_),
    .Y(_11429_));
 OAI21x1_ASAP7_75t_R _15738_ (.A1(_11420_),
    .A2(_11425_),
    .B(_11429_),
    .Y(_03292_));
 AO21x1_ASAP7_75t_R _15739_ (.A1(_01808_),
    .A2(_11423_),
    .B(_10826_),
    .Y(_11430_));
 AO21x1_ASAP7_75t_R _15740_ (.A1(_01766_),
    .A2(_11421_),
    .B(_11430_),
    .Y(_11431_));
 OR3x1_ASAP7_75t_R _15741_ (.A(_11406_),
    .B(_02344_),
    .C(_11428_),
    .Y(_11432_));
 OAI21x1_ASAP7_75t_R _15742_ (.A1(_11420_),
    .A2(_11431_),
    .B(_11432_),
    .Y(_03293_));
 AO21x1_ASAP7_75t_R _15743_ (.A1(_01807_),
    .A2(_11423_),
    .B(_10826_),
    .Y(_11433_));
 AO21x1_ASAP7_75t_R _15744_ (.A1(_01765_),
    .A2(_11421_),
    .B(_11433_),
    .Y(_11434_));
 OR3x1_ASAP7_75t_R _15745_ (.A(_11406_),
    .B(_02345_),
    .C(_11428_),
    .Y(_11435_));
 OAI21x1_ASAP7_75t_R _15746_ (.A1(_11420_),
    .A2(_11434_),
    .B(_11435_),
    .Y(_03294_));
 AO21x1_ASAP7_75t_R _15747_ (.A1(_01806_),
    .A2(_11423_),
    .B(_08765_),
    .Y(_11436_));
 AO21x1_ASAP7_75t_R _15748_ (.A1(_01764_),
    .A2(_11421_),
    .B(_11436_),
    .Y(_11437_));
 OR3x1_ASAP7_75t_R _15749_ (.A(_11406_),
    .B(_02346_),
    .C(_11428_),
    .Y(_11438_));
 OAI21x1_ASAP7_75t_R _15750_ (.A1(_11420_),
    .A2(_11437_),
    .B(_11438_),
    .Y(_03295_));
 AO21x1_ASAP7_75t_R _15751_ (.A1(_01805_),
    .A2(_11423_),
    .B(_08765_),
    .Y(_11439_));
 AO21x1_ASAP7_75t_R _15752_ (.A1(_01763_),
    .A2(_11421_),
    .B(_11439_),
    .Y(_11440_));
 OR3x1_ASAP7_75t_R _15753_ (.A(_11406_),
    .B(_02347_),
    .C(_11428_),
    .Y(_11441_));
 OAI21x1_ASAP7_75t_R _15754_ (.A1(_11420_),
    .A2(_11440_),
    .B(_11441_),
    .Y(_03296_));
 AO21x1_ASAP7_75t_R _15755_ (.A1(_01804_),
    .A2(_11423_),
    .B(_08765_),
    .Y(_11442_));
 AO21x1_ASAP7_75t_R _15756_ (.A1(_01762_),
    .A2(_11421_),
    .B(_11442_),
    .Y(_11443_));
 OR3x1_ASAP7_75t_R _15757_ (.A(_11406_),
    .B(_02348_),
    .C(_11428_),
    .Y(_11444_));
 OAI21x1_ASAP7_75t_R _15758_ (.A1(_11420_),
    .A2(_11443_),
    .B(_11444_),
    .Y(_03297_));
 AO21x1_ASAP7_75t_R _15759_ (.A1(_01803_),
    .A2(_11423_),
    .B(_08765_),
    .Y(_11445_));
 AO21x1_ASAP7_75t_R _15760_ (.A1(_01761_),
    .A2(_11421_),
    .B(_11445_),
    .Y(_11446_));
 OR3x1_ASAP7_75t_R _15761_ (.A(_11406_),
    .B(_02349_),
    .C(_11428_),
    .Y(_11447_));
 OAI21x1_ASAP7_75t_R _15762_ (.A1(_11420_),
    .A2(_11446_),
    .B(_11447_),
    .Y(_03298_));
 AO21x1_ASAP7_75t_R _15763_ (.A1(_01802_),
    .A2(_11423_),
    .B(_08765_),
    .Y(_11448_));
 AO21x1_ASAP7_75t_R _15764_ (.A1(_01760_),
    .A2(_11421_),
    .B(_11448_),
    .Y(_11449_));
 OR3x1_ASAP7_75t_R _15765_ (.A(_11406_),
    .B(_02350_),
    .C(_11428_),
    .Y(_11450_));
 OAI21x1_ASAP7_75t_R _15766_ (.A1(_11420_),
    .A2(_11449_),
    .B(_11450_),
    .Y(_03299_));
 AND2x2_ASAP7_75t_R _15767_ (.A(_01801_),
    .B(_11422_),
    .Y(_11451_));
 AO21x1_ASAP7_75t_R _15768_ (.A1(_01759_),
    .A2(_11421_),
    .B(_11451_),
    .Y(_11452_));
 AOI21x1_ASAP7_75t_R _15769_ (.A1(_11428_),
    .A2(_11452_),
    .B(_09081_),
    .Y(_03300_));
 OA21x2_ASAP7_75t_R _15770_ (.A1(_11344_),
    .A2(_11414_),
    .B(_01758_),
    .Y(_11453_));
 AO21x1_ASAP7_75t_R _15771_ (.A1(_11330_),
    .A2(_11422_),
    .B(_11453_),
    .Y(_11454_));
 NAND2x1_ASAP7_75t_R _15772_ (.A(_11427_),
    .B(_11454_),
    .Y(_11455_));
 OA211x2_ASAP7_75t_R _15773_ (.A1(_11394_),
    .A2(_11428_),
    .B(_11455_),
    .C(_09830_),
    .Y(_03301_));
 AO21x1_ASAP7_75t_R _15774_ (.A1(_11326_),
    .A2(_11413_),
    .B(_11414_),
    .Y(_11456_));
 AND3x1_ASAP7_75t_R _15775_ (.A(_10809_),
    .B(_11408_),
    .C(_11456_),
    .Y(_03302_));
 AOI21x1_ASAP7_75t_R _15776_ (.A1(_11426_),
    .A2(_11418_),
    .B(_09081_),
    .Y(_03303_));
 AO21x1_ASAP7_75t_R _15777_ (.A1(_01797_),
    .A2(_11423_),
    .B(_08765_),
    .Y(_11457_));
 AO21x1_ASAP7_75t_R _15778_ (.A1(_01755_),
    .A2(_11421_),
    .B(_11457_),
    .Y(_11458_));
 OR3x1_ASAP7_75t_R _15779_ (.A(_11406_),
    .B(_02355_),
    .C(_11427_),
    .Y(_11459_));
 OAI21x1_ASAP7_75t_R _15780_ (.A1(_11420_),
    .A2(_11458_),
    .B(_11459_),
    .Y(_03304_));
 AO21x1_ASAP7_75t_R _15781_ (.A1(_01796_),
    .A2(_11423_),
    .B(_08765_),
    .Y(_11460_));
 AO21x1_ASAP7_75t_R _15782_ (.A1(_01754_),
    .A2(_11415_),
    .B(_11460_),
    .Y(_11461_));
 OR3x1_ASAP7_75t_R _15783_ (.A(_08941_),
    .B(_02342_),
    .C(_11427_),
    .Y(_11462_));
 OAI21x1_ASAP7_75t_R _15784_ (.A1(_11420_),
    .A2(_11461_),
    .B(_11462_),
    .Y(_03305_));
 OR4x1_ASAP7_75t_R _15785_ (.A(net4),
    .B(net3),
    .C(net6),
    .D(net5),
    .Y(_11463_));
 OR3x1_ASAP7_75t_R _15786_ (.A(net2),
    .B(net1),
    .C(_11463_),
    .Y(_11464_));
 AND2x6_ASAP7_75t_R _15787_ (.A(_08526_),
    .B(_11464_),
    .Y(_11465_));
 BUFx12f_ASAP7_75t_R _15788_ (.A(_11465_),
    .Y(_11466_));
 BUFx6f_ASAP7_75t_R _15789_ (.A(_01717_),
    .Y(_11467_));
 AND4x1_ASAP7_75t_R _15790_ (.A(_01688_),
    .B(_01716_),
    .C(_11467_),
    .D(_01718_),
    .Y(_11468_));
 AND5x1_ASAP7_75t_R _15791_ (.A(_01707_),
    .B(_01712_),
    .C(_01713_),
    .D(_01715_),
    .E(_11468_),
    .Y(_11469_));
 AND5x2_ASAP7_75t_R _15792_ (.A(_01709_),
    .B(_01710_),
    .C(_01711_),
    .D(_11466_),
    .E(_11469_),
    .Y(_11470_));
 BUFx6f_ASAP7_75t_R _15793_ (.A(_01700_),
    .Y(_11471_));
 AND4x1_ASAP7_75t_R _15794_ (.A(_01702_),
    .B(_01703_),
    .C(_01704_),
    .D(_01705_),
    .Y(_11472_));
 AND4x1_ASAP7_75t_R _15795_ (.A(_01696_),
    .B(_01698_),
    .C(_01699_),
    .D(_01706_),
    .Y(_11473_));
 AND5x1_ASAP7_75t_R _15796_ (.A(_01689_),
    .B(_01690_),
    .C(_01695_),
    .D(_01714_),
    .E(_11473_),
    .Y(_11474_));
 BUFx6f_ASAP7_75t_R _15797_ (.A(_01692_),
    .Y(_11475_));
 AND3x1_ASAP7_75t_R _15798_ (.A(_01693_),
    .B(_01694_),
    .C(_01697_),
    .Y(_11476_));
 OR3x1_ASAP7_75t_R _15799_ (.A(_01691_),
    .B(_11475_),
    .C(_11476_),
    .Y(_11477_));
 AND5x2_ASAP7_75t_R _15800_ (.A(_11471_),
    .B(_01701_),
    .C(_11472_),
    .D(_11474_),
    .E(_11477_),
    .Y(_11478_));
 NAND2x2_ASAP7_75t_R _15801_ (.A(_11470_),
    .B(_11478_),
    .Y(_11479_));
 NOR2x1_ASAP7_75t_R _15802_ (.A(_01645_),
    .B(_11479_),
    .Y(_03306_));
 NOR2x1_ASAP7_75t_R _15803_ (.A(_01648_),
    .B(_11479_),
    .Y(_03307_));
 NOR2x1_ASAP7_75t_R _15804_ (.A(_01647_),
    .B(_11479_),
    .Y(_03308_));
 NOR2x1_ASAP7_75t_R _15805_ (.A(_01646_),
    .B(_11479_),
    .Y(_03309_));
 NOR2x1_ASAP7_75t_R _15806_ (.A(_01644_),
    .B(_11479_),
    .Y(_03310_));
 NOR2x1_ASAP7_75t_R _15807_ (.A(_01643_),
    .B(_11479_),
    .Y(_03311_));
 INVx1_ASAP7_75t_R _15808_ (.A(_11479_),
    .Y(_03312_));
 AND2x2_ASAP7_75t_R _15809_ (.A(_10927_),
    .B(_00031_),
    .Y(_03313_));
 OR4x1_ASAP7_75t_R _15810_ (.A(_01693_),
    .B(_01694_),
    .C(_01697_),
    .D(_02631_),
    .Y(_11480_));
 OR4x1_ASAP7_75t_R _15811_ (.A(_01689_),
    .B(_01690_),
    .C(_01691_),
    .D(_11475_),
    .Y(_11481_));
 OR4x1_ASAP7_75t_R _15812_ (.A(_01688_),
    .B(_01718_),
    .C(_11480_),
    .D(_11481_),
    .Y(_11482_));
 BUFx6f_ASAP7_75t_R _15813_ (.A(_11482_),
    .Y(_11483_));
 OR3x1_ASAP7_75t_R _15814_ (.A(_01688_),
    .B(_11480_),
    .C(_11481_),
    .Y(_11484_));
 NAND2x1_ASAP7_75t_R _15815_ (.A(_01718_),
    .B(_11484_),
    .Y(_11485_));
 AND3x1_ASAP7_75t_R _15816_ (.A(_10809_),
    .B(_11483_),
    .C(_11485_),
    .Y(_03314_));
 OR4x1_ASAP7_75t_R _15817_ (.A(_01688_),
    .B(_01689_),
    .C(_01691_),
    .D(_11475_),
    .Y(_11486_));
 OR3x1_ASAP7_75t_R _15818_ (.A(_01697_),
    .B(_01708_),
    .C(_00031_),
    .Y(_11487_));
 OR3x2_ASAP7_75t_R _15819_ (.A(_01693_),
    .B(_01694_),
    .C(_11487_),
    .Y(_11488_));
 OR4x1_ASAP7_75t_R _15820_ (.A(_01690_),
    .B(_01718_),
    .C(_11486_),
    .D(_11488_),
    .Y(_11489_));
 XOR2x2_ASAP7_75t_R _15821_ (.A(_11467_),
    .B(_11489_),
    .Y(_11490_));
 AND2x2_ASAP7_75t_R _15822_ (.A(_10927_),
    .B(_11490_),
    .Y(_03315_));
 OR3x1_ASAP7_75t_R _15823_ (.A(_01716_),
    .B(_11467_),
    .C(_11483_),
    .Y(_11491_));
 OAI21x1_ASAP7_75t_R _15824_ (.A1(_11467_),
    .A2(_11483_),
    .B(_01716_),
    .Y(_11492_));
 AND3x1_ASAP7_75t_R _15825_ (.A(_10809_),
    .B(_11491_),
    .C(_11492_),
    .Y(_03316_));
 OR3x1_ASAP7_75t_R _15826_ (.A(_01716_),
    .B(_11467_),
    .C(_11489_),
    .Y(_11493_));
 XOR2x2_ASAP7_75t_R _15827_ (.A(_01715_),
    .B(_11493_),
    .Y(_11494_));
 AND2x2_ASAP7_75t_R _15828_ (.A(_10927_),
    .B(_11494_),
    .Y(_03317_));
 OR4x1_ASAP7_75t_R _15829_ (.A(_01715_),
    .B(_01716_),
    .C(_11467_),
    .D(_11483_),
    .Y(_11495_));
 XOR2x2_ASAP7_75t_R _15830_ (.A(_01714_),
    .B(_11495_),
    .Y(_11496_));
 AND2x2_ASAP7_75t_R _15831_ (.A(_10927_),
    .B(_11496_),
    .Y(_03318_));
 OR5x1_ASAP7_75t_R _15832_ (.A(_01714_),
    .B(_01715_),
    .C(_01716_),
    .D(_11467_),
    .E(_11489_),
    .Y(_11497_));
 XOR2x2_ASAP7_75t_R _15833_ (.A(_01713_),
    .B(_11497_),
    .Y(_11498_));
 AND2x2_ASAP7_75t_R _15834_ (.A(_10927_),
    .B(_11498_),
    .Y(_03319_));
 OR5x2_ASAP7_75t_R _15835_ (.A(_01713_),
    .B(_01714_),
    .C(_01715_),
    .D(_01716_),
    .E(_11467_),
    .Y(_11499_));
 OR3x1_ASAP7_75t_R _15836_ (.A(_01712_),
    .B(_11483_),
    .C(_11499_),
    .Y(_11500_));
 OAI21x1_ASAP7_75t_R _15837_ (.A1(_11483_),
    .A2(_11499_),
    .B(_01712_),
    .Y(_11501_));
 AND3x1_ASAP7_75t_R _15838_ (.A(_10809_),
    .B(_11500_),
    .C(_11501_),
    .Y(_03320_));
 OR3x1_ASAP7_75t_R _15839_ (.A(_01712_),
    .B(_11489_),
    .C(_11499_),
    .Y(_11502_));
 XOR2x2_ASAP7_75t_R _15840_ (.A(_01711_),
    .B(_11502_),
    .Y(_11503_));
 AND2x2_ASAP7_75t_R _15841_ (.A(_10927_),
    .B(_11503_),
    .Y(_03321_));
 OR4x1_ASAP7_75t_R _15842_ (.A(_01710_),
    .B(_01711_),
    .C(_01712_),
    .D(_11499_),
    .Y(_11504_));
 OR4x1_ASAP7_75t_R _15843_ (.A(_01711_),
    .B(_01712_),
    .C(_11483_),
    .D(_11499_),
    .Y(_11505_));
 NAND2x1_ASAP7_75t_R _15844_ (.A(_01710_),
    .B(_11505_),
    .Y(_11506_));
 OA211x2_ASAP7_75t_R _15845_ (.A1(_11483_),
    .A2(_11504_),
    .B(_11506_),
    .C(_09830_),
    .Y(_03322_));
 BUFx12f_ASAP7_75t_R _15846_ (.A(_08598_),
    .Y(_11507_));
 BUFx6f_ASAP7_75t_R _15847_ (.A(_11507_),
    .Y(_11508_));
 OR2x6_ASAP7_75t_R _15848_ (.A(_11489_),
    .B(_11504_),
    .Y(_11509_));
 XOR2x2_ASAP7_75t_R _15849_ (.A(_01709_),
    .B(_11509_),
    .Y(_11510_));
 AND2x2_ASAP7_75t_R _15850_ (.A(_11508_),
    .B(_11510_),
    .Y(_03323_));
 NOR2x1_ASAP7_75t_R _15851_ (.A(_10716_),
    .B(_02632_),
    .Y(_03324_));
 OR3x1_ASAP7_75t_R _15852_ (.A(_01709_),
    .B(_11483_),
    .C(_11504_),
    .Y(_11511_));
 XOR2x2_ASAP7_75t_R _15853_ (.A(_01707_),
    .B(_11511_),
    .Y(_11512_));
 AND2x2_ASAP7_75t_R _15854_ (.A(_11508_),
    .B(_11512_),
    .Y(_03325_));
 OR3x1_ASAP7_75t_R _15855_ (.A(_01707_),
    .B(_01709_),
    .C(_11509_),
    .Y(_11513_));
 XOR2x2_ASAP7_75t_R _15856_ (.A(_01706_),
    .B(_11513_),
    .Y(_11514_));
 AND2x2_ASAP7_75t_R _15857_ (.A(_11508_),
    .B(_11514_),
    .Y(_03326_));
 OR5x1_ASAP7_75t_R _15858_ (.A(_01706_),
    .B(_01707_),
    .C(_01709_),
    .D(_11483_),
    .E(_11504_),
    .Y(_11515_));
 XOR2x2_ASAP7_75t_R _15859_ (.A(_01705_),
    .B(_11515_),
    .Y(_11516_));
 AND2x2_ASAP7_75t_R _15860_ (.A(_11508_),
    .B(_11516_),
    .Y(_03327_));
 OR5x1_ASAP7_75t_R _15861_ (.A(_01704_),
    .B(_01705_),
    .C(_01706_),
    .D(_01707_),
    .E(_01709_),
    .Y(_11517_));
 OR3x2_ASAP7_75t_R _15862_ (.A(_11489_),
    .B(_11504_),
    .C(_11517_),
    .Y(_11518_));
 OR5x1_ASAP7_75t_R _15863_ (.A(_01705_),
    .B(_01706_),
    .C(_01707_),
    .D(_01709_),
    .E(_11509_),
    .Y(_11519_));
 NAND2x1_ASAP7_75t_R _15864_ (.A(_01704_),
    .B(_11519_),
    .Y(_11520_));
 AND3x1_ASAP7_75t_R _15865_ (.A(_10809_),
    .B(_11518_),
    .C(_11520_),
    .Y(_03328_));
 OR3x2_ASAP7_75t_R _15866_ (.A(_11482_),
    .B(_11504_),
    .C(_11517_),
    .Y(_11521_));
 XOR2x2_ASAP7_75t_R _15867_ (.A(_01703_),
    .B(_11521_),
    .Y(_11522_));
 AND2x2_ASAP7_75t_R _15868_ (.A(_11508_),
    .B(_11522_),
    .Y(_03329_));
 OR3x1_ASAP7_75t_R _15869_ (.A(_01702_),
    .B(_01703_),
    .C(_11518_),
    .Y(_11523_));
 OAI21x1_ASAP7_75t_R _15870_ (.A1(_01703_),
    .A2(_11518_),
    .B(_01702_),
    .Y(_11524_));
 AND3x1_ASAP7_75t_R _15871_ (.A(_10809_),
    .B(_11523_),
    .C(_11524_),
    .Y(_03330_));
 BUFx6f_ASAP7_75t_R _15872_ (.A(_08581_),
    .Y(_11525_));
 OR3x2_ASAP7_75t_R _15873_ (.A(_01701_),
    .B(_01702_),
    .C(_01703_),
    .Y(_11526_));
 OR2x6_ASAP7_75t_R _15874_ (.A(_11521_),
    .B(_11526_),
    .Y(_11527_));
 OR3x1_ASAP7_75t_R _15875_ (.A(_01702_),
    .B(_01703_),
    .C(_11521_),
    .Y(_11528_));
 NAND2x1_ASAP7_75t_R _15876_ (.A(_01701_),
    .B(_11528_),
    .Y(_11529_));
 AND3x1_ASAP7_75t_R _15877_ (.A(_11525_),
    .B(_11527_),
    .C(_11529_),
    .Y(_03331_));
 OR2x6_ASAP7_75t_R _15878_ (.A(_11518_),
    .B(_11526_),
    .Y(_11530_));
 XNOR2x2_ASAP7_75t_R _15879_ (.A(_11471_),
    .B(_11530_),
    .Y(_11531_));
 NOR2x1_ASAP7_75t_R _15880_ (.A(_10716_),
    .B(_11531_),
    .Y(_03332_));
 OR3x1_ASAP7_75t_R _15881_ (.A(_01699_),
    .B(_11471_),
    .C(_11527_),
    .Y(_11532_));
 OAI21x1_ASAP7_75t_R _15882_ (.A1(_11471_),
    .A2(_11527_),
    .B(_01699_),
    .Y(_11533_));
 AND3x1_ASAP7_75t_R _15883_ (.A(_11525_),
    .B(_11532_),
    .C(_11533_),
    .Y(_03333_));
 OR4x1_ASAP7_75t_R _15884_ (.A(_01699_),
    .B(_11471_),
    .C(_11518_),
    .D(_11526_),
    .Y(_11534_));
 XOR2x2_ASAP7_75t_R _15885_ (.A(_01698_),
    .B(_11534_),
    .Y(_11535_));
 AND2x2_ASAP7_75t_R _15886_ (.A(_11508_),
    .B(_11535_),
    .Y(_03334_));
 XOR2x2_ASAP7_75t_R _15887_ (.A(_01697_),
    .B(_02631_),
    .Y(_11536_));
 AND2x2_ASAP7_75t_R _15888_ (.A(_11508_),
    .B(_11536_),
    .Y(_03335_));
 OR4x1_ASAP7_75t_R _15889_ (.A(_01698_),
    .B(_01699_),
    .C(_11471_),
    .D(_11527_),
    .Y(_11537_));
 XOR2x2_ASAP7_75t_R _15890_ (.A(_01696_),
    .B(_11537_),
    .Y(_11538_));
 AND2x2_ASAP7_75t_R _15891_ (.A(_11508_),
    .B(_11538_),
    .Y(_03336_));
 OR4x1_ASAP7_75t_R _15892_ (.A(_01696_),
    .B(_01698_),
    .C(_01699_),
    .D(_11471_),
    .Y(_11539_));
 OR3x1_ASAP7_75t_R _15893_ (.A(_01695_),
    .B(_11530_),
    .C(_11539_),
    .Y(_11540_));
 OAI21x1_ASAP7_75t_R _15894_ (.A1(_11530_),
    .A2(_11539_),
    .B(_01695_),
    .Y(_11541_));
 AND3x1_ASAP7_75t_R _15895_ (.A(_11525_),
    .B(_11540_),
    .C(_11541_),
    .Y(_03337_));
 XOR2x2_ASAP7_75t_R _15896_ (.A(_01694_),
    .B(_11487_),
    .Y(_11542_));
 AND2x2_ASAP7_75t_R _15897_ (.A(_11508_),
    .B(_11542_),
    .Y(_03338_));
 OR3x1_ASAP7_75t_R _15898_ (.A(_01694_),
    .B(_01697_),
    .C(_02631_),
    .Y(_11543_));
 NAND2x1_ASAP7_75t_R _15899_ (.A(_01693_),
    .B(_11543_),
    .Y(_11544_));
 AND3x1_ASAP7_75t_R _15900_ (.A(_11525_),
    .B(_11480_),
    .C(_11544_),
    .Y(_03339_));
 XOR2x2_ASAP7_75t_R _15901_ (.A(_11475_),
    .B(_11488_),
    .Y(_11545_));
 AND2x2_ASAP7_75t_R _15902_ (.A(_11508_),
    .B(_11545_),
    .Y(_03340_));
 OR3x1_ASAP7_75t_R _15903_ (.A(_01691_),
    .B(_11475_),
    .C(_11480_),
    .Y(_11546_));
 OAI21x1_ASAP7_75t_R _15904_ (.A1(_11475_),
    .A2(_11480_),
    .B(_01691_),
    .Y(_11547_));
 AND3x1_ASAP7_75t_R _15905_ (.A(_11525_),
    .B(_11546_),
    .C(_11547_),
    .Y(_03341_));
 BUFx6f_ASAP7_75t_R _15906_ (.A(_11507_),
    .Y(_11548_));
 OR3x1_ASAP7_75t_R _15907_ (.A(_01691_),
    .B(_11475_),
    .C(_11488_),
    .Y(_11549_));
 XOR2x2_ASAP7_75t_R _15908_ (.A(_01690_),
    .B(_11549_),
    .Y(_11550_));
 AND2x2_ASAP7_75t_R _15909_ (.A(_11548_),
    .B(_11550_),
    .Y(_03342_));
 OR4x1_ASAP7_75t_R _15910_ (.A(_01690_),
    .B(_01691_),
    .C(_11475_),
    .D(_11480_),
    .Y(_11551_));
 NAND2x1_ASAP7_75t_R _15911_ (.A(_01689_),
    .B(_11551_),
    .Y(_11552_));
 OA211x2_ASAP7_75t_R _15912_ (.A1(_11480_),
    .A2(_11481_),
    .B(_11552_),
    .C(_09830_),
    .Y(_03343_));
 OR3x1_ASAP7_75t_R _15913_ (.A(_01688_),
    .B(_11481_),
    .C(_11488_),
    .Y(_11553_));
 OAI21x1_ASAP7_75t_R _15914_ (.A1(_11481_),
    .A2(_11488_),
    .B(_01688_),
    .Y(_11554_));
 AND3x1_ASAP7_75t_R _15915_ (.A(_11525_),
    .B(_11553_),
    .C(_11554_),
    .Y(_03344_));
 BUFx3_ASAP7_75t_R _15916_ (.A(_01649_),
    .Y(_11555_));
 AND4x1_ASAP7_75t_R _15917_ (.A(_11555_),
    .B(_01677_),
    .C(_01678_),
    .D(_01679_),
    .Y(_11556_));
 AND5x1_ASAP7_75t_R _15918_ (.A(_01668_),
    .B(_01673_),
    .C(_01674_),
    .D(_01676_),
    .E(_11556_),
    .Y(_11557_));
 AND5x1_ASAP7_75t_R _15919_ (.A(_01670_),
    .B(_01671_),
    .C(_01672_),
    .D(_11466_),
    .E(_11557_),
    .Y(_11558_));
 BUFx3_ASAP7_75t_R _15920_ (.A(_01665_),
    .Y(_11559_));
 AND4x1_ASAP7_75t_R _15921_ (.A(_01663_),
    .B(_01664_),
    .C(_11559_),
    .D(_01666_),
    .Y(_11560_));
 AND4x1_ASAP7_75t_R _15922_ (.A(_01657_),
    .B(_01659_),
    .C(_01660_),
    .D(_01667_),
    .Y(_11561_));
 AND5x1_ASAP7_75t_R _15923_ (.A(_01650_),
    .B(_01651_),
    .C(_01656_),
    .D(_01675_),
    .E(_11561_),
    .Y(_11562_));
 AND3x1_ASAP7_75t_R _15924_ (.A(_01654_),
    .B(_01655_),
    .C(_01658_),
    .Y(_11563_));
 OR3x1_ASAP7_75t_R _15925_ (.A(_01652_),
    .B(_01653_),
    .C(_11563_),
    .Y(_11564_));
 AND5x2_ASAP7_75t_R _15926_ (.A(_01661_),
    .B(_01662_),
    .C(_11560_),
    .D(_11562_),
    .E(_11564_),
    .Y(_11565_));
 NAND2x2_ASAP7_75t_R _15927_ (.A(_11558_),
    .B(_11565_),
    .Y(_11566_));
 NOR2x1_ASAP7_75t_R _15928_ (.A(_01639_),
    .B(_11566_),
    .Y(_03345_));
 INVx1_ASAP7_75t_R _15929_ (.A(_11566_),
    .Y(_03346_));
 NOR2x1_ASAP7_75t_R _15930_ (.A(_01642_),
    .B(_11566_),
    .Y(_03347_));
 NOR2x1_ASAP7_75t_R _15931_ (.A(_01641_),
    .B(_11566_),
    .Y(_03348_));
 NOR2x1_ASAP7_75t_R _15932_ (.A(_01640_),
    .B(_11566_),
    .Y(_03349_));
 NOR2x1_ASAP7_75t_R _15933_ (.A(_01638_),
    .B(_11566_),
    .Y(_03350_));
 NOR2x1_ASAP7_75t_R _15934_ (.A(_01637_),
    .B(_11566_),
    .Y(_03351_));
 INVx1_ASAP7_75t_R _15935_ (.A(_11566_),
    .Y(_03352_));
 AND2x2_ASAP7_75t_R _15936_ (.A(_11548_),
    .B(_00032_),
    .Y(_03353_));
 OR4x1_ASAP7_75t_R _15937_ (.A(_01654_),
    .B(_01655_),
    .C(_01658_),
    .D(_02623_),
    .Y(_11567_));
 OR4x1_ASAP7_75t_R _15938_ (.A(_01650_),
    .B(_01651_),
    .C(_01652_),
    .D(_01653_),
    .Y(_11568_));
 OR2x6_ASAP7_75t_R _15939_ (.A(_11567_),
    .B(_11568_),
    .Y(_11569_));
 OR3x1_ASAP7_75t_R _15940_ (.A(_11555_),
    .B(_01679_),
    .C(_11569_),
    .Y(_11570_));
 OAI21x1_ASAP7_75t_R _15941_ (.A1(_11555_),
    .A2(_11569_),
    .B(_01679_),
    .Y(_11571_));
 AND3x1_ASAP7_75t_R _15942_ (.A(_11525_),
    .B(_11570_),
    .C(_11571_),
    .Y(_03354_));
 OR5x2_ASAP7_75t_R _15943_ (.A(_01654_),
    .B(_01655_),
    .C(_01658_),
    .D(_01669_),
    .E(_00032_),
    .Y(_11572_));
 OR2x2_ASAP7_75t_R _15944_ (.A(_11568_),
    .B(_11572_),
    .Y(_11573_));
 OR3x1_ASAP7_75t_R _15945_ (.A(_11555_),
    .B(_01679_),
    .C(_11573_),
    .Y(_11574_));
 XOR2x2_ASAP7_75t_R _15946_ (.A(_01678_),
    .B(_11574_),
    .Y(_11575_));
 AND2x2_ASAP7_75t_R _15947_ (.A(_11548_),
    .B(_11575_),
    .Y(_03355_));
 OR4x1_ASAP7_75t_R _15948_ (.A(_11555_),
    .B(_01677_),
    .C(_01678_),
    .D(_01679_),
    .Y(_11576_));
 OR3x2_ASAP7_75t_R _15949_ (.A(_11567_),
    .B(_11568_),
    .C(_11576_),
    .Y(_11577_));
 OR4x1_ASAP7_75t_R _15950_ (.A(_11555_),
    .B(_01678_),
    .C(_01679_),
    .D(_11569_),
    .Y(_11578_));
 NAND2x1_ASAP7_75t_R _15951_ (.A(_01677_),
    .B(_11578_),
    .Y(_11579_));
 AND3x1_ASAP7_75t_R _15952_ (.A(_11525_),
    .B(_11577_),
    .C(_11579_),
    .Y(_03356_));
 OR3x2_ASAP7_75t_R _15953_ (.A(_11568_),
    .B(_11572_),
    .C(_11576_),
    .Y(_11580_));
 XOR2x2_ASAP7_75t_R _15954_ (.A(_01676_),
    .B(_11580_),
    .Y(_11581_));
 AND2x2_ASAP7_75t_R _15955_ (.A(_11548_),
    .B(_11581_),
    .Y(_03357_));
 OR3x1_ASAP7_75t_R _15956_ (.A(_01675_),
    .B(_01676_),
    .C(_11577_),
    .Y(_11582_));
 OAI21x1_ASAP7_75t_R _15957_ (.A1(_01676_),
    .A2(_11577_),
    .B(_01675_),
    .Y(_11583_));
 AND3x1_ASAP7_75t_R _15958_ (.A(_11525_),
    .B(_11582_),
    .C(_11583_),
    .Y(_03358_));
 OR3x1_ASAP7_75t_R _15959_ (.A(_01675_),
    .B(_01676_),
    .C(_11580_),
    .Y(_11584_));
 XOR2x2_ASAP7_75t_R _15960_ (.A(_01674_),
    .B(_11584_),
    .Y(_11585_));
 AND2x2_ASAP7_75t_R _15961_ (.A(_11548_),
    .B(_11585_),
    .Y(_03359_));
 OR4x1_ASAP7_75t_R _15962_ (.A(_01673_),
    .B(_01674_),
    .C(_01675_),
    .D(_01676_),
    .Y(_11586_));
 OR4x1_ASAP7_75t_R _15963_ (.A(_01674_),
    .B(_01675_),
    .C(_01676_),
    .D(_11577_),
    .Y(_11587_));
 NAND2x1_ASAP7_75t_R _15964_ (.A(_01673_),
    .B(_11587_),
    .Y(_11588_));
 BUFx12f_ASAP7_75t_R _15965_ (.A(_08876_),
    .Y(_11589_));
 OA211x2_ASAP7_75t_R _15966_ (.A1(_11577_),
    .A2(_11586_),
    .B(_11588_),
    .C(_11589_),
    .Y(_03360_));
 OR3x1_ASAP7_75t_R _15967_ (.A(_01672_),
    .B(_11580_),
    .C(_11586_),
    .Y(_11590_));
 OAI21x1_ASAP7_75t_R _15968_ (.A1(_11580_),
    .A2(_11586_),
    .B(_01672_),
    .Y(_11591_));
 AND3x1_ASAP7_75t_R _15969_ (.A(_11525_),
    .B(_11590_),
    .C(_11591_),
    .Y(_03361_));
 OR3x1_ASAP7_75t_R _15970_ (.A(_01672_),
    .B(_11577_),
    .C(_11586_),
    .Y(_11592_));
 XOR2x2_ASAP7_75t_R _15971_ (.A(_01671_),
    .B(_11592_),
    .Y(_11593_));
 AND2x2_ASAP7_75t_R _15972_ (.A(_11548_),
    .B(_11593_),
    .Y(_03362_));
 BUFx6f_ASAP7_75t_R _15973_ (.A(_08581_),
    .Y(_11594_));
 OR5x2_ASAP7_75t_R _15974_ (.A(_01670_),
    .B(_01671_),
    .C(_01672_),
    .D(_11580_),
    .E(_11586_),
    .Y(_11595_));
 OR4x1_ASAP7_75t_R _15975_ (.A(_01671_),
    .B(_01672_),
    .C(_11580_),
    .D(_11586_),
    .Y(_11596_));
 NAND2x1_ASAP7_75t_R _15976_ (.A(_01670_),
    .B(_11596_),
    .Y(_11597_));
 AND3x1_ASAP7_75t_R _15977_ (.A(_11594_),
    .B(_11595_),
    .C(_11597_),
    .Y(_03363_));
 NOR2x1_ASAP7_75t_R _15978_ (.A(_10716_),
    .B(_02624_),
    .Y(_03364_));
 OR5x2_ASAP7_75t_R _15979_ (.A(_01670_),
    .B(_01671_),
    .C(_01672_),
    .D(_11577_),
    .E(_11586_),
    .Y(_11598_));
 XOR2x2_ASAP7_75t_R _15980_ (.A(_01668_),
    .B(_11598_),
    .Y(_11599_));
 AND2x2_ASAP7_75t_R _15981_ (.A(_11548_),
    .B(_11599_),
    .Y(_03365_));
 OR3x1_ASAP7_75t_R _15982_ (.A(_01667_),
    .B(_01668_),
    .C(_11595_),
    .Y(_11600_));
 OAI21x1_ASAP7_75t_R _15983_ (.A1(_01668_),
    .A2(_11595_),
    .B(_01667_),
    .Y(_11601_));
 AND3x1_ASAP7_75t_R _15984_ (.A(_11594_),
    .B(_11600_),
    .C(_11601_),
    .Y(_03366_));
 OR4x1_ASAP7_75t_R _15985_ (.A(_01666_),
    .B(_01667_),
    .C(_01668_),
    .D(_11598_),
    .Y(_11602_));
 OR3x1_ASAP7_75t_R _15986_ (.A(_01667_),
    .B(_01668_),
    .C(_11598_),
    .Y(_11603_));
 NAND2x1_ASAP7_75t_R _15987_ (.A(_01666_),
    .B(_11603_),
    .Y(_11604_));
 AND3x1_ASAP7_75t_R _15988_ (.A(_11594_),
    .B(_11602_),
    .C(_11604_),
    .Y(_03367_));
 OR4x1_ASAP7_75t_R _15989_ (.A(_01666_),
    .B(_01667_),
    .C(_01668_),
    .D(_11595_),
    .Y(_11605_));
 XOR2x2_ASAP7_75t_R _15990_ (.A(_11559_),
    .B(_11605_),
    .Y(_11606_));
 AND2x2_ASAP7_75t_R _15991_ (.A(_11548_),
    .B(_11606_),
    .Y(_03368_));
 OR3x1_ASAP7_75t_R _15992_ (.A(_01664_),
    .B(_11559_),
    .C(_11602_),
    .Y(_11607_));
 OAI21x1_ASAP7_75t_R _15993_ (.A1(_11559_),
    .A2(_11602_),
    .B(_01664_),
    .Y(_11608_));
 AND3x1_ASAP7_75t_R _15994_ (.A(_11594_),
    .B(_11607_),
    .C(_11608_),
    .Y(_03369_));
 OR3x1_ASAP7_75t_R _15995_ (.A(_01664_),
    .B(_11559_),
    .C(_11605_),
    .Y(_11609_));
 XOR2x2_ASAP7_75t_R _15996_ (.A(_01663_),
    .B(_11609_),
    .Y(_11610_));
 AND2x2_ASAP7_75t_R _15997_ (.A(_11548_),
    .B(_11610_),
    .Y(_03370_));
 OR4x1_ASAP7_75t_R _15998_ (.A(_01663_),
    .B(_01664_),
    .C(_11559_),
    .D(_11602_),
    .Y(_11611_));
 XOR2x2_ASAP7_75t_R _15999_ (.A(_01662_),
    .B(_11611_),
    .Y(_11612_));
 AND2x2_ASAP7_75t_R _16000_ (.A(_11548_),
    .B(_11612_),
    .Y(_03371_));
 BUFx6f_ASAP7_75t_R _16001_ (.A(_11507_),
    .Y(_11613_));
 OR5x1_ASAP7_75t_R _16002_ (.A(_01662_),
    .B(_01663_),
    .C(_01664_),
    .D(_11559_),
    .E(_11605_),
    .Y(_11614_));
 XOR2x2_ASAP7_75t_R _16003_ (.A(_01661_),
    .B(_11614_),
    .Y(_11615_));
 AND2x2_ASAP7_75t_R _16004_ (.A(_11613_),
    .B(_11615_),
    .Y(_03372_));
 OR5x2_ASAP7_75t_R _16005_ (.A(_01661_),
    .B(_01662_),
    .C(_01663_),
    .D(_01664_),
    .E(_11559_),
    .Y(_11616_));
 OR3x1_ASAP7_75t_R _16006_ (.A(_01660_),
    .B(_11602_),
    .C(_11616_),
    .Y(_11617_));
 OAI21x1_ASAP7_75t_R _16007_ (.A1(_11602_),
    .A2(_11616_),
    .B(_01660_),
    .Y(_11618_));
 AND3x1_ASAP7_75t_R _16008_ (.A(_11594_),
    .B(_11617_),
    .C(_11618_),
    .Y(_03373_));
 OR3x1_ASAP7_75t_R _16009_ (.A(_01660_),
    .B(_11605_),
    .C(_11616_),
    .Y(_11619_));
 XOR2x2_ASAP7_75t_R _16010_ (.A(_01659_),
    .B(_11619_),
    .Y(_11620_));
 AND2x2_ASAP7_75t_R _16011_ (.A(_11613_),
    .B(_11620_),
    .Y(_03374_));
 XOR2x2_ASAP7_75t_R _16012_ (.A(_01658_),
    .B(_02623_),
    .Y(_11621_));
 AND2x2_ASAP7_75t_R _16013_ (.A(_11613_),
    .B(_11621_),
    .Y(_03375_));
 OR4x1_ASAP7_75t_R _16014_ (.A(_01659_),
    .B(_01660_),
    .C(_11602_),
    .D(_11616_),
    .Y(_11622_));
 XOR2x2_ASAP7_75t_R _16015_ (.A(_01657_),
    .B(_11622_),
    .Y(_11623_));
 AND2x2_ASAP7_75t_R _16016_ (.A(_11613_),
    .B(_11623_),
    .Y(_03376_));
 OR5x1_ASAP7_75t_R _16017_ (.A(_01657_),
    .B(_01659_),
    .C(_01660_),
    .D(_11605_),
    .E(_11616_),
    .Y(_11624_));
 XOR2x2_ASAP7_75t_R _16018_ (.A(_01656_),
    .B(_11624_),
    .Y(_11625_));
 AND2x2_ASAP7_75t_R _16019_ (.A(_11613_),
    .B(_11625_),
    .Y(_03377_));
 OR3x1_ASAP7_75t_R _16020_ (.A(_01658_),
    .B(_01669_),
    .C(_00032_),
    .Y(_11626_));
 XOR2x2_ASAP7_75t_R _16021_ (.A(_01655_),
    .B(_11626_),
    .Y(_11627_));
 AND2x2_ASAP7_75t_R _16022_ (.A(_11613_),
    .B(_11627_),
    .Y(_03378_));
 OR3x1_ASAP7_75t_R _16023_ (.A(_01655_),
    .B(_01658_),
    .C(_02623_),
    .Y(_11628_));
 NAND2x1_ASAP7_75t_R _16024_ (.A(_01654_),
    .B(_11628_),
    .Y(_11629_));
 AND3x1_ASAP7_75t_R _16025_ (.A(_11594_),
    .B(_11567_),
    .C(_11629_),
    .Y(_03379_));
 XOR2x2_ASAP7_75t_R _16026_ (.A(_01653_),
    .B(_11572_),
    .Y(_11630_));
 AND2x2_ASAP7_75t_R _16027_ (.A(_11613_),
    .B(_11630_),
    .Y(_03380_));
 OR3x1_ASAP7_75t_R _16028_ (.A(_01652_),
    .B(_01653_),
    .C(_11567_),
    .Y(_11631_));
 OAI21x1_ASAP7_75t_R _16029_ (.A1(_01653_),
    .A2(_11567_),
    .B(_01652_),
    .Y(_11632_));
 AND3x1_ASAP7_75t_R _16030_ (.A(_11594_),
    .B(_11631_),
    .C(_11632_),
    .Y(_03381_));
 OR3x1_ASAP7_75t_R _16031_ (.A(_01652_),
    .B(_01653_),
    .C(_11572_),
    .Y(_11633_));
 XOR2x2_ASAP7_75t_R _16032_ (.A(_01651_),
    .B(_11633_),
    .Y(_11634_));
 AND2x2_ASAP7_75t_R _16033_ (.A(_11613_),
    .B(_11634_),
    .Y(_03382_));
 OR4x1_ASAP7_75t_R _16034_ (.A(_01651_),
    .B(_01652_),
    .C(_01653_),
    .D(_11567_),
    .Y(_11635_));
 NAND2x1_ASAP7_75t_R _16035_ (.A(_01650_),
    .B(_11635_),
    .Y(_11636_));
 AND3x1_ASAP7_75t_R _16036_ (.A(_11594_),
    .B(_11569_),
    .C(_11636_),
    .Y(_03383_));
 XOR2x2_ASAP7_75t_R _16037_ (.A(_11555_),
    .B(_11573_),
    .Y(_11637_));
 AND2x2_ASAP7_75t_R _16038_ (.A(_11613_),
    .B(_11637_),
    .Y(_03384_));
 AND2x2_ASAP7_75t_R _16039_ (.A(_11613_),
    .B(_00015_),
    .Y(_03385_));
 BUFx6f_ASAP7_75t_R _16040_ (.A(_02330_),
    .Y(_11638_));
 INVx1_ASAP7_75t_R _16041_ (.A(_02331_),
    .Y(_11639_));
 INVx2_ASAP7_75t_R _16042_ (.A(_02337_),
    .Y(_11640_));
 AND4x1_ASAP7_75t_R _16043_ (.A(_01681_),
    .B(_01682_),
    .C(_01683_),
    .D(_01684_),
    .Y(_05017_));
 AND3x4_ASAP7_75t_R _16044_ (.A(\xs[0].cli1.i[39] ),
    .B(_01685_),
    .C(_05017_),
    .Y(_05018_));
 OA21x2_ASAP7_75t_R _16045_ (.A1(_01680_),
    .A2(_05017_),
    .B(_11640_),
    .Y(_05019_));
 AND4x1_ASAP7_75t_R _16046_ (.A(_01720_),
    .B(_01721_),
    .C(_01722_),
    .D(_01723_),
    .Y(_05020_));
 AND3x1_ASAP7_75t_R _16047_ (.A(\peo[0][39] ),
    .B(\peo[0][32] ),
    .C(_05020_),
    .Y(_05021_));
 OA21x2_ASAP7_75t_R _16048_ (.A1(_05018_),
    .A2(_05019_),
    .B(_05021_),
    .Y(_05022_));
 OR2x2_ASAP7_75t_R _16049_ (.A(_01719_),
    .B(_05020_),
    .Y(_05023_));
 BUFx3_ASAP7_75t_R _16050_ (.A(_05023_),
    .Y(_05024_));
 AND3x1_ASAP7_75t_R _16051_ (.A(_02337_),
    .B(_05018_),
    .C(_05024_),
    .Y(_05025_));
 INVx1_ASAP7_75t_R _16052_ (.A(_11638_),
    .Y(_05026_));
 OA21x2_ASAP7_75t_R _16053_ (.A1(_05022_),
    .A2(_05025_),
    .B(_05026_),
    .Y(_05027_));
 OR4x1_ASAP7_75t_R _16054_ (.A(_11638_),
    .B(_11639_),
    .C(_11640_),
    .D(_05027_),
    .Y(_05028_));
 NOR2x1_ASAP7_75t_R _16055_ (.A(_02341_),
    .B(_05028_),
    .Y(_05029_));
 OR2x6_ASAP7_75t_R _16056_ (.A(_01680_),
    .B(_05017_),
    .Y(_05030_));
 NAND2x1_ASAP7_75t_R _16057_ (.A(_11638_),
    .B(_00015_),
    .Y(_05031_));
 AO21x1_ASAP7_75t_R _16058_ (.A1(_02331_),
    .A2(_11640_),
    .B(_11638_),
    .Y(_05032_));
 OA21x2_ASAP7_75t_R _16059_ (.A1(_05030_),
    .A2(_05031_),
    .B(_05032_),
    .Y(_05033_));
 OA21x2_ASAP7_75t_R _16060_ (.A1(_05024_),
    .A2(_05033_),
    .B(_05018_),
    .Y(_05034_));
 NAND2x1_ASAP7_75t_R _16061_ (.A(_01687_),
    .B(_05034_),
    .Y(_05035_));
 OA211x2_ASAP7_75t_R _16062_ (.A1(\peo[0][0] ),
    .A2(_05034_),
    .B(_05035_),
    .C(_05028_),
    .Y(_05036_));
 OA21x2_ASAP7_75t_R _16063_ (.A1(_05029_),
    .A2(_05036_),
    .B(_11397_),
    .Y(_03386_));
 OR2x2_ASAP7_75t_R _16064_ (.A(_08683_),
    .B(_05028_),
    .Y(_05037_));
 BUFx3_ASAP7_75t_R _16065_ (.A(_05037_),
    .Y(_05038_));
 NOR2x1_ASAP7_75t_R _16066_ (.A(_02340_),
    .B(_05038_),
    .Y(_03387_));
 NOR2x1_ASAP7_75t_R _16067_ (.A(_02339_),
    .B(_05038_),
    .Y(_03388_));
 NOR2x1_ASAP7_75t_R _16068_ (.A(_02338_),
    .B(_05038_),
    .Y(_03389_));
 NOR2x1_ASAP7_75t_R _16069_ (.A(_02329_),
    .B(_05038_),
    .Y(_03390_));
 NOR2x1_ASAP7_75t_R _16070_ (.A(_02328_),
    .B(_05038_),
    .Y(_03391_));
 OA21x2_ASAP7_75t_R _16071_ (.A1(_11640_),
    .A2(_05024_),
    .B(_02331_),
    .Y(_05039_));
 OAI22x1_ASAP7_75t_R _16072_ (.A1(_05024_),
    .A2(_05031_),
    .B1(_05039_),
    .B2(_11638_),
    .Y(_05040_));
 NOR2x1_ASAP7_75t_R _16073_ (.A(_05024_),
    .B(_05032_),
    .Y(_05041_));
 NOR2x2_ASAP7_75t_R _16074_ (.A(_01680_),
    .B(_05017_),
    .Y(_05042_));
 AO21x1_ASAP7_75t_R _16075_ (.A1(_05018_),
    .A2(_05041_),
    .B(_05042_),
    .Y(_05043_));
 AND3x1_ASAP7_75t_R _16076_ (.A(_01687_),
    .B(_05040_),
    .C(_05043_),
    .Y(_05044_));
 INVx1_ASAP7_75t_R _16077_ (.A(_05044_),
    .Y(_05045_));
 AO21x1_ASAP7_75t_R _16078_ (.A1(_05040_),
    .A2(_05043_),
    .B(\peo[0][0] ),
    .Y(_05046_));
 OR3x1_ASAP7_75t_R _16079_ (.A(_11638_),
    .B(_11639_),
    .C(_02337_),
    .Y(_05047_));
 AOI21x1_ASAP7_75t_R _16080_ (.A1(_05021_),
    .A2(_05030_),
    .B(_05047_),
    .Y(_05048_));
 NOR2x1_ASAP7_75t_R _16081_ (.A(_09314_),
    .B(_05048_),
    .Y(_05049_));
 NOR2x1_ASAP7_75t_R _16082_ (.A(_09934_),
    .B(_02341_),
    .Y(_05050_));
 AO32x1_ASAP7_75t_R _16083_ (.A1(_05045_),
    .A2(_05046_),
    .A3(_05049_),
    .B1(_05050_),
    .B2(_05048_),
    .Y(_03392_));
 OR3x2_ASAP7_75t_R _16084_ (.A(_10763_),
    .B(_05027_),
    .C(_05047_),
    .Y(_05051_));
 NOR2x1_ASAP7_75t_R _16085_ (.A(_02340_),
    .B(_05051_),
    .Y(_03393_));
 NOR2x1_ASAP7_75t_R _16086_ (.A(_02339_),
    .B(_05051_),
    .Y(_03394_));
 NOR2x1_ASAP7_75t_R _16087_ (.A(_02338_),
    .B(_05051_),
    .Y(_03395_));
 NOR2x1_ASAP7_75t_R _16088_ (.A(_02329_),
    .B(_05051_),
    .Y(_03396_));
 NOR2x1_ASAP7_75t_R _16089_ (.A(_02328_),
    .B(_05051_),
    .Y(_03397_));
 OA22x2_ASAP7_75t_R _16090_ (.A1(_05024_),
    .A2(_05031_),
    .B1(_05039_),
    .B2(_11638_),
    .Y(_05052_));
 NAND2x1_ASAP7_75t_R _16091_ (.A(_05042_),
    .B(_05052_),
    .Y(_05053_));
 AND3x1_ASAP7_75t_R _16092_ (.A(_01687_),
    .B(_05042_),
    .C(_05052_),
    .Y(_05054_));
 AO21x1_ASAP7_75t_R _16093_ (.A1(_01725_),
    .A2(_05053_),
    .B(_05054_),
    .Y(_05055_));
 AOI21x1_ASAP7_75t_R _16094_ (.A1(_05026_),
    .A2(_11639_),
    .B(_05027_),
    .Y(_05056_));
 NAND2x2_ASAP7_75t_R _16095_ (.A(_08528_),
    .B(_05056_),
    .Y(_05057_));
 OR3x1_ASAP7_75t_R _16096_ (.A(_08941_),
    .B(_02341_),
    .C(_05056_),
    .Y(_05058_));
 OAI21x1_ASAP7_75t_R _16097_ (.A1(_05055_),
    .A2(_05057_),
    .B(_05058_),
    .Y(_03398_));
 OR2x2_ASAP7_75t_R _16098_ (.A(_09220_),
    .B(_05056_),
    .Y(_05059_));
 BUFx6f_ASAP7_75t_R _16099_ (.A(_05059_),
    .Y(_05060_));
 NOR2x1_ASAP7_75t_R _16100_ (.A(_02340_),
    .B(_05060_),
    .Y(_03399_));
 NOR2x1_ASAP7_75t_R _16101_ (.A(_02339_),
    .B(_05060_),
    .Y(_03400_));
 NOR2x1_ASAP7_75t_R _16102_ (.A(_02338_),
    .B(_05060_),
    .Y(_03401_));
 AND3x1_ASAP7_75t_R _16103_ (.A(_01685_),
    .B(_05042_),
    .C(_05052_),
    .Y(_05061_));
 AO21x1_ASAP7_75t_R _16104_ (.A1(_01724_),
    .A2(_05053_),
    .B(_05061_),
    .Y(_05062_));
 OR3x1_ASAP7_75t_R _16105_ (.A(_08941_),
    .B(_02337_),
    .C(_05056_),
    .Y(_05063_));
 OAI21x1_ASAP7_75t_R _16106_ (.A1(_05057_),
    .A2(_05062_),
    .B(_05063_),
    .Y(_03402_));
 AND3x1_ASAP7_75t_R _16107_ (.A(_01684_),
    .B(_05042_),
    .C(_05052_),
    .Y(_05064_));
 AO21x1_ASAP7_75t_R _16108_ (.A1(_01723_),
    .A2(_05053_),
    .B(_05064_),
    .Y(_05065_));
 OR3x1_ASAP7_75t_R _16109_ (.A(_08941_),
    .B(_02336_),
    .C(_05056_),
    .Y(_05066_));
 OAI21x1_ASAP7_75t_R _16110_ (.A1(_05057_),
    .A2(_05065_),
    .B(_05066_),
    .Y(_03403_));
 AND3x1_ASAP7_75t_R _16111_ (.A(_01683_),
    .B(_05042_),
    .C(_05052_),
    .Y(_05067_));
 AO21x1_ASAP7_75t_R _16112_ (.A1(_01722_),
    .A2(_05053_),
    .B(_05067_),
    .Y(_05068_));
 OR3x1_ASAP7_75t_R _16113_ (.A(_08941_),
    .B(_02335_),
    .C(_05056_),
    .Y(_05069_));
 OAI21x1_ASAP7_75t_R _16114_ (.A1(_05057_),
    .A2(_05068_),
    .B(_05069_),
    .Y(_03404_));
 AND3x1_ASAP7_75t_R _16115_ (.A(_01682_),
    .B(_05042_),
    .C(_05052_),
    .Y(_05070_));
 AO21x1_ASAP7_75t_R _16116_ (.A1(_01721_),
    .A2(_05053_),
    .B(_05070_),
    .Y(_05071_));
 OR3x1_ASAP7_75t_R _16117_ (.A(_08941_),
    .B(_02334_),
    .C(_05056_),
    .Y(_05072_));
 OAI21x1_ASAP7_75t_R _16118_ (.A1(_05057_),
    .A2(_05071_),
    .B(_05072_),
    .Y(_03405_));
 AND3x1_ASAP7_75t_R _16119_ (.A(_01681_),
    .B(_05042_),
    .C(_05052_),
    .Y(_05073_));
 AO21x1_ASAP7_75t_R _16120_ (.A1(_01720_),
    .A2(_05053_),
    .B(_05073_),
    .Y(_05074_));
 OR3x1_ASAP7_75t_R _16121_ (.A(_08941_),
    .B(_02333_),
    .C(_05056_),
    .Y(_05075_));
 OAI21x1_ASAP7_75t_R _16122_ (.A1(_05057_),
    .A2(_05074_),
    .B(_05075_),
    .Y(_03406_));
 NOR2x1_ASAP7_75t_R _16123_ (.A(_02332_),
    .B(_05060_),
    .Y(_03407_));
 OA211x2_ASAP7_75t_R _16124_ (.A1(_11638_),
    .A2(_02331_),
    .B(_05027_),
    .C(_11589_),
    .Y(_03408_));
 AND3x1_ASAP7_75t_R _16125_ (.A(_05030_),
    .B(_05024_),
    .C(_05056_),
    .Y(_05076_));
 NOR2x1_ASAP7_75t_R _16126_ (.A(_10716_),
    .B(_05076_),
    .Y(_03409_));
 NOR2x1_ASAP7_75t_R _16127_ (.A(_02329_),
    .B(_05060_),
    .Y(_03410_));
 NOR2x1_ASAP7_75t_R _16128_ (.A(_02328_),
    .B(_05060_),
    .Y(_03411_));
 BUFx6f_ASAP7_75t_R _16129_ (.A(_01612_),
    .Y(_05077_));
 AND4x1_ASAP7_75t_R _16130_ (.A(_01584_),
    .B(_05077_),
    .C(_01613_),
    .D(_01614_),
    .Y(_05078_));
 AND5x1_ASAP7_75t_R _16131_ (.A(_01603_),
    .B(_01608_),
    .C(_01609_),
    .D(_01611_),
    .E(_05078_),
    .Y(_05079_));
 AND5x2_ASAP7_75t_R _16132_ (.A(_01605_),
    .B(_01606_),
    .C(_01607_),
    .D(_11466_),
    .E(_05079_),
    .Y(_05080_));
 AND4x1_ASAP7_75t_R _16133_ (.A(_01598_),
    .B(_01599_),
    .C(_01600_),
    .D(_01601_),
    .Y(_05081_));
 AND4x1_ASAP7_75t_R _16134_ (.A(_01592_),
    .B(_01594_),
    .C(_01595_),
    .D(_01602_),
    .Y(_05082_));
 AND5x1_ASAP7_75t_R _16135_ (.A(_01585_),
    .B(_01586_),
    .C(_01591_),
    .D(_01610_),
    .E(_05082_),
    .Y(_05083_));
 BUFx3_ASAP7_75t_R _16136_ (.A(_01588_),
    .Y(_05084_));
 AND3x1_ASAP7_75t_R _16137_ (.A(_01589_),
    .B(_01590_),
    .C(_01593_),
    .Y(_05085_));
 OR3x1_ASAP7_75t_R _16138_ (.A(_01587_),
    .B(_05084_),
    .C(_05085_),
    .Y(_05086_));
 AND5x2_ASAP7_75t_R _16139_ (.A(_01596_),
    .B(_01597_),
    .C(_05081_),
    .D(_05083_),
    .E(_05086_),
    .Y(_05087_));
 NAND2x2_ASAP7_75t_R _16140_ (.A(_05080_),
    .B(_05087_),
    .Y(_05088_));
 NOR2x1_ASAP7_75t_R _16141_ (.A(_01541_),
    .B(_05088_),
    .Y(_03412_));
 INVx1_ASAP7_75t_R _16142_ (.A(_05088_),
    .Y(_03413_));
 NOR2x1_ASAP7_75t_R _16143_ (.A(_01544_),
    .B(_05088_),
    .Y(_03414_));
 NOR2x1_ASAP7_75t_R _16144_ (.A(_01543_),
    .B(_05088_),
    .Y(_03415_));
 NOR2x1_ASAP7_75t_R _16145_ (.A(_01542_),
    .B(_05088_),
    .Y(_03416_));
 NOR2x1_ASAP7_75t_R _16146_ (.A(_01540_),
    .B(_05088_),
    .Y(_03417_));
 NOR2x1_ASAP7_75t_R _16147_ (.A(_01539_),
    .B(_05088_),
    .Y(_03418_));
 INVx1_ASAP7_75t_R _16148_ (.A(_05088_),
    .Y(_03419_));
 BUFx6f_ASAP7_75t_R _16149_ (.A(_11507_),
    .Y(_05089_));
 AND2x2_ASAP7_75t_R _16150_ (.A(_05089_),
    .B(_00033_),
    .Y(_03420_));
 OR4x1_ASAP7_75t_R _16151_ (.A(_01589_),
    .B(_01590_),
    .C(_01593_),
    .D(_02627_),
    .Y(_05090_));
 OR5x2_ASAP7_75t_R _16152_ (.A(_01584_),
    .B(_01585_),
    .C(_01586_),
    .D(_01587_),
    .E(_05084_),
    .Y(_05091_));
 OR3x1_ASAP7_75t_R _16153_ (.A(_01614_),
    .B(_05090_),
    .C(_05091_),
    .Y(_05092_));
 OAI21x1_ASAP7_75t_R _16154_ (.A1(_05090_),
    .A2(_05091_),
    .B(_01614_),
    .Y(_05093_));
 AND3x1_ASAP7_75t_R _16155_ (.A(_11594_),
    .B(_05092_),
    .C(_05093_),
    .Y(_03421_));
 OR5x2_ASAP7_75t_R _16156_ (.A(_01589_),
    .B(_01590_),
    .C(_01593_),
    .D(_01604_),
    .E(_00033_),
    .Y(_05094_));
 OR4x1_ASAP7_75t_R _16157_ (.A(_01613_),
    .B(_01614_),
    .C(_05091_),
    .D(_05094_),
    .Y(_05095_));
 OR3x1_ASAP7_75t_R _16158_ (.A(_01614_),
    .B(_05091_),
    .C(_05094_),
    .Y(_05096_));
 NAND2x1_ASAP7_75t_R _16159_ (.A(_01613_),
    .B(_05096_),
    .Y(_05097_));
 AND3x1_ASAP7_75t_R _16160_ (.A(_11594_),
    .B(_05095_),
    .C(_05097_),
    .Y(_03422_));
 OR4x1_ASAP7_75t_R _16161_ (.A(_01613_),
    .B(_01614_),
    .C(_05090_),
    .D(_05091_),
    .Y(_05098_));
 XOR2x2_ASAP7_75t_R _16162_ (.A(_05077_),
    .B(_05098_),
    .Y(_05099_));
 AND2x2_ASAP7_75t_R _16163_ (.A(_05089_),
    .B(_05099_),
    .Y(_03423_));
 BUFx6f_ASAP7_75t_R _16164_ (.A(_08581_),
    .Y(_05100_));
 OR3x1_ASAP7_75t_R _16165_ (.A(_01611_),
    .B(_05077_),
    .C(_05095_),
    .Y(_05101_));
 OAI21x1_ASAP7_75t_R _16166_ (.A1(_05077_),
    .A2(_05095_),
    .B(_01611_),
    .Y(_05102_));
 AND3x1_ASAP7_75t_R _16167_ (.A(_05100_),
    .B(_05101_),
    .C(_05102_),
    .Y(_03424_));
 OR3x1_ASAP7_75t_R _16168_ (.A(_01611_),
    .B(_05077_),
    .C(_05098_),
    .Y(_05103_));
 XOR2x2_ASAP7_75t_R _16169_ (.A(_01610_),
    .B(_05103_),
    .Y(_05104_));
 AND2x2_ASAP7_75t_R _16170_ (.A(_05089_),
    .B(_05104_),
    .Y(_03425_));
 OR4x1_ASAP7_75t_R _16171_ (.A(_01610_),
    .B(_01611_),
    .C(_05077_),
    .D(_05095_),
    .Y(_05105_));
 XOR2x2_ASAP7_75t_R _16172_ (.A(_01609_),
    .B(_05105_),
    .Y(_05106_));
 AND2x2_ASAP7_75t_R _16173_ (.A(_05089_),
    .B(_05106_),
    .Y(_03426_));
 OR5x1_ASAP7_75t_R _16174_ (.A(_01609_),
    .B(_01610_),
    .C(_01611_),
    .D(_05077_),
    .E(_05098_),
    .Y(_05107_));
 XOR2x2_ASAP7_75t_R _16175_ (.A(_01608_),
    .B(_05107_),
    .Y(_05108_));
 AND2x2_ASAP7_75t_R _16176_ (.A(_05089_),
    .B(_05108_),
    .Y(_03427_));
 OR5x2_ASAP7_75t_R _16177_ (.A(_01608_),
    .B(_01609_),
    .C(_01610_),
    .D(_01611_),
    .E(_05077_),
    .Y(_05109_));
 OR3x1_ASAP7_75t_R _16178_ (.A(_01607_),
    .B(_05095_),
    .C(_05109_),
    .Y(_05110_));
 OAI21x1_ASAP7_75t_R _16179_ (.A1(_05095_),
    .A2(_05109_),
    .B(_01607_),
    .Y(_05111_));
 AND3x1_ASAP7_75t_R _16180_ (.A(_05100_),
    .B(_05110_),
    .C(_05111_),
    .Y(_03428_));
 OR3x2_ASAP7_75t_R _16181_ (.A(_01607_),
    .B(_05098_),
    .C(_05109_),
    .Y(_05112_));
 XOR2x2_ASAP7_75t_R _16182_ (.A(_01606_),
    .B(_05112_),
    .Y(_05113_));
 AND2x2_ASAP7_75t_R _16183_ (.A(_05089_),
    .B(_05113_),
    .Y(_03429_));
 OR4x1_ASAP7_75t_R _16184_ (.A(_01606_),
    .B(_01607_),
    .C(_05095_),
    .D(_05109_),
    .Y(_05114_));
 XOR2x2_ASAP7_75t_R _16185_ (.A(_01605_),
    .B(_05114_),
    .Y(_05115_));
 AND2x2_ASAP7_75t_R _16186_ (.A(_05089_),
    .B(_05115_),
    .Y(_03430_));
 NOR2x1_ASAP7_75t_R _16187_ (.A(_10716_),
    .B(_02628_),
    .Y(_03431_));
 OR3x1_ASAP7_75t_R _16188_ (.A(_01605_),
    .B(_01606_),
    .C(_05112_),
    .Y(_05116_));
 XOR2x2_ASAP7_75t_R _16189_ (.A(_01603_),
    .B(_05116_),
    .Y(_05117_));
 AND2x2_ASAP7_75t_R _16190_ (.A(_05089_),
    .B(_05117_),
    .Y(_03432_));
 OR3x1_ASAP7_75t_R _16191_ (.A(_01603_),
    .B(_01605_),
    .C(_05114_),
    .Y(_05118_));
 XOR2x2_ASAP7_75t_R _16192_ (.A(_01602_),
    .B(_05118_),
    .Y(_05119_));
 AND2x2_ASAP7_75t_R _16193_ (.A(_05089_),
    .B(_05119_),
    .Y(_03433_));
 OR2x2_ASAP7_75t_R _16194_ (.A(_01606_),
    .B(_05112_),
    .Y(_05120_));
 OR4x1_ASAP7_75t_R _16195_ (.A(_01602_),
    .B(_01603_),
    .C(_01605_),
    .D(_05120_),
    .Y(_05121_));
 XOR2x2_ASAP7_75t_R _16196_ (.A(_01601_),
    .B(_05121_),
    .Y(_05122_));
 AND2x2_ASAP7_75t_R _16197_ (.A(_05089_),
    .B(_05122_),
    .Y(_03434_));
 OR5x2_ASAP7_75t_R _16198_ (.A(_01600_),
    .B(_01601_),
    .C(_01602_),
    .D(_01603_),
    .E(_01605_),
    .Y(_05123_));
 OR5x1_ASAP7_75t_R _16199_ (.A(_01601_),
    .B(_01602_),
    .C(_01603_),
    .D(_01605_),
    .E(_05114_),
    .Y(_05124_));
 NAND2x1_ASAP7_75t_R _16200_ (.A(_01600_),
    .B(_05124_),
    .Y(_05125_));
 OA211x2_ASAP7_75t_R _16201_ (.A1(_05114_),
    .A2(_05123_),
    .B(_05125_),
    .C(_11589_),
    .Y(_03435_));
 BUFx6f_ASAP7_75t_R _16202_ (.A(_11507_),
    .Y(_05126_));
 OR5x2_ASAP7_75t_R _16203_ (.A(_01606_),
    .B(_01607_),
    .C(_05098_),
    .D(_05109_),
    .E(_05123_),
    .Y(_05127_));
 XOR2x2_ASAP7_75t_R _16204_ (.A(_01599_),
    .B(_05127_),
    .Y(_05128_));
 AND2x2_ASAP7_75t_R _16205_ (.A(_05126_),
    .B(_05128_),
    .Y(_03436_));
 OR3x1_ASAP7_75t_R _16206_ (.A(_01599_),
    .B(_05114_),
    .C(_05123_),
    .Y(_05129_));
 XOR2x2_ASAP7_75t_R _16207_ (.A(_01598_),
    .B(_05129_),
    .Y(_05130_));
 AND2x2_ASAP7_75t_R _16208_ (.A(_05126_),
    .B(_05130_),
    .Y(_03437_));
 OR4x1_ASAP7_75t_R _16209_ (.A(_01597_),
    .B(_01598_),
    .C(_01599_),
    .D(_05127_),
    .Y(_05131_));
 OR3x1_ASAP7_75t_R _16210_ (.A(_01598_),
    .B(_01599_),
    .C(_05127_),
    .Y(_05132_));
 NAND2x1_ASAP7_75t_R _16211_ (.A(_01597_),
    .B(_05132_),
    .Y(_05133_));
 AND3x1_ASAP7_75t_R _16212_ (.A(_05100_),
    .B(_05131_),
    .C(_05133_),
    .Y(_03438_));
 OR5x2_ASAP7_75t_R _16213_ (.A(_01597_),
    .B(_01598_),
    .C(_01599_),
    .D(_05114_),
    .E(_05123_),
    .Y(_05134_));
 XOR2x2_ASAP7_75t_R _16214_ (.A(_01596_),
    .B(_05134_),
    .Y(_05135_));
 AND2x2_ASAP7_75t_R _16215_ (.A(_05126_),
    .B(_05135_),
    .Y(_03439_));
 OR3x1_ASAP7_75t_R _16216_ (.A(_01595_),
    .B(_01596_),
    .C(_05131_),
    .Y(_05136_));
 OAI21x1_ASAP7_75t_R _16217_ (.A1(_01596_),
    .A2(_05131_),
    .B(_01595_),
    .Y(_05137_));
 AND3x1_ASAP7_75t_R _16218_ (.A(_05100_),
    .B(_05136_),
    .C(_05137_),
    .Y(_03440_));
 OR3x1_ASAP7_75t_R _16219_ (.A(_01595_),
    .B(_01596_),
    .C(_05134_),
    .Y(_05138_));
 XOR2x2_ASAP7_75t_R _16220_ (.A(_01594_),
    .B(_05138_),
    .Y(_05139_));
 AND2x2_ASAP7_75t_R _16221_ (.A(_05126_),
    .B(_05139_),
    .Y(_03441_));
 XOR2x2_ASAP7_75t_R _16222_ (.A(_01593_),
    .B(_02627_),
    .Y(_05140_));
 AND2x2_ASAP7_75t_R _16223_ (.A(_05126_),
    .B(_05140_),
    .Y(_03442_));
 OR4x1_ASAP7_75t_R _16224_ (.A(_01594_),
    .B(_01595_),
    .C(_01596_),
    .D(_05131_),
    .Y(_05141_));
 XOR2x2_ASAP7_75t_R _16225_ (.A(_01592_),
    .B(_05141_),
    .Y(_05142_));
 AND2x2_ASAP7_75t_R _16226_ (.A(_05126_),
    .B(_05142_),
    .Y(_03443_));
 OR5x1_ASAP7_75t_R _16227_ (.A(_01592_),
    .B(_01594_),
    .C(_01595_),
    .D(_01596_),
    .E(_05134_),
    .Y(_05143_));
 XOR2x2_ASAP7_75t_R _16228_ (.A(_01591_),
    .B(_05143_),
    .Y(_05144_));
 AND2x2_ASAP7_75t_R _16229_ (.A(_05126_),
    .B(_05144_),
    .Y(_03444_));
 OR3x1_ASAP7_75t_R _16230_ (.A(_01593_),
    .B(_01604_),
    .C(_00033_),
    .Y(_05145_));
 XOR2x2_ASAP7_75t_R _16231_ (.A(_01590_),
    .B(_05145_),
    .Y(_05146_));
 AND2x2_ASAP7_75t_R _16232_ (.A(_05126_),
    .B(_05146_),
    .Y(_03445_));
 OR3x1_ASAP7_75t_R _16233_ (.A(_01590_),
    .B(_01593_),
    .C(_02627_),
    .Y(_05147_));
 NAND2x1_ASAP7_75t_R _16234_ (.A(_01589_),
    .B(_05147_),
    .Y(_05148_));
 AND3x1_ASAP7_75t_R _16235_ (.A(_05100_),
    .B(_05090_),
    .C(_05148_),
    .Y(_03446_));
 XOR2x2_ASAP7_75t_R _16236_ (.A(_05084_),
    .B(_05094_),
    .Y(_05149_));
 AND2x2_ASAP7_75t_R _16237_ (.A(_05126_),
    .B(_05149_),
    .Y(_03447_));
 OR3x1_ASAP7_75t_R _16238_ (.A(_01587_),
    .B(_05084_),
    .C(_05090_),
    .Y(_05150_));
 OAI21x1_ASAP7_75t_R _16239_ (.A1(_05084_),
    .A2(_05090_),
    .B(_01587_),
    .Y(_05151_));
 AND3x1_ASAP7_75t_R _16240_ (.A(_05100_),
    .B(_05150_),
    .C(_05151_),
    .Y(_03448_));
 OR3x1_ASAP7_75t_R _16241_ (.A(_01587_),
    .B(_05084_),
    .C(_05094_),
    .Y(_05152_));
 XOR2x2_ASAP7_75t_R _16242_ (.A(_01586_),
    .B(_05152_),
    .Y(_05153_));
 AND2x2_ASAP7_75t_R _16243_ (.A(_05126_),
    .B(_05153_),
    .Y(_03449_));
 BUFx6f_ASAP7_75t_R _16244_ (.A(_11507_),
    .Y(_05154_));
 OR4x1_ASAP7_75t_R _16245_ (.A(_01586_),
    .B(_01587_),
    .C(_05084_),
    .D(_05090_),
    .Y(_05155_));
 XOR2x2_ASAP7_75t_R _16246_ (.A(_01585_),
    .B(_05155_),
    .Y(_05156_));
 AND2x2_ASAP7_75t_R _16247_ (.A(_05154_),
    .B(_05156_),
    .Y(_03450_));
 OR5x1_ASAP7_75t_R _16248_ (.A(_01585_),
    .B(_01586_),
    .C(_01587_),
    .D(_05084_),
    .E(_05094_),
    .Y(_05157_));
 XOR2x2_ASAP7_75t_R _16249_ (.A(_01584_),
    .B(_05157_),
    .Y(_05158_));
 AND2x2_ASAP7_75t_R _16250_ (.A(_05154_),
    .B(_05158_),
    .Y(_03451_));
 BUFx6f_ASAP7_75t_R _16251_ (.A(_01568_),
    .Y(_05159_));
 BUFx3_ASAP7_75t_R _16252_ (.A(_01545_),
    .Y(_05160_));
 AND4x1_ASAP7_75t_R _16253_ (.A(_05160_),
    .B(_01573_),
    .C(_01574_),
    .D(_01575_),
    .Y(_05161_));
 AND5x1_ASAP7_75t_R _16254_ (.A(_01564_),
    .B(_01569_),
    .C(_01570_),
    .D(_01572_),
    .E(_05161_),
    .Y(_05162_));
 AND5x2_ASAP7_75t_R _16255_ (.A(_01566_),
    .B(_01567_),
    .C(_05159_),
    .D(_11466_),
    .E(_05162_),
    .Y(_05163_));
 BUFx6f_ASAP7_75t_R _16256_ (.A(_01560_),
    .Y(_05164_));
 AND4x1_ASAP7_75t_R _16257_ (.A(_01559_),
    .B(_05164_),
    .C(_01561_),
    .D(_01562_),
    .Y(_05165_));
 AND4x1_ASAP7_75t_R _16258_ (.A(_01553_),
    .B(_01555_),
    .C(_01556_),
    .D(_01563_),
    .Y(_05166_));
 AND5x1_ASAP7_75t_R _16259_ (.A(_01546_),
    .B(_01547_),
    .C(_01552_),
    .D(_01571_),
    .E(_05166_),
    .Y(_05167_));
 BUFx3_ASAP7_75t_R _16260_ (.A(_01549_),
    .Y(_05168_));
 AND3x1_ASAP7_75t_R _16261_ (.A(_01550_),
    .B(_01551_),
    .C(_01554_),
    .Y(_05169_));
 OR3x1_ASAP7_75t_R _16262_ (.A(_01548_),
    .B(_05168_),
    .C(_05169_),
    .Y(_05170_));
 AND5x2_ASAP7_75t_R _16263_ (.A(_01557_),
    .B(_01558_),
    .C(_05165_),
    .D(_05167_),
    .E(_05170_),
    .Y(_05171_));
 NAND2x2_ASAP7_75t_R _16264_ (.A(_05163_),
    .B(_05171_),
    .Y(_05172_));
 NOR2x1_ASAP7_75t_R _16265_ (.A(_01535_),
    .B(_05172_),
    .Y(_03452_));
 INVx1_ASAP7_75t_R _16266_ (.A(_05172_),
    .Y(_03453_));
 NOR2x1_ASAP7_75t_R _16267_ (.A(_01538_),
    .B(_05172_),
    .Y(_03454_));
 NOR2x1_ASAP7_75t_R _16268_ (.A(_01537_),
    .B(_05172_),
    .Y(_03455_));
 NOR2x1_ASAP7_75t_R _16269_ (.A(_01536_),
    .B(_05172_),
    .Y(_03456_));
 NOR2x1_ASAP7_75t_R _16270_ (.A(_01534_),
    .B(_05172_),
    .Y(_03457_));
 NOR2x1_ASAP7_75t_R _16271_ (.A(_01533_),
    .B(_05172_),
    .Y(_03458_));
 INVx1_ASAP7_75t_R _16272_ (.A(_05172_),
    .Y(_03459_));
 AND2x2_ASAP7_75t_R _16273_ (.A(_05154_),
    .B(_00034_),
    .Y(_03460_));
 OR4x1_ASAP7_75t_R _16274_ (.A(_01550_),
    .B(_01551_),
    .C(_01554_),
    .D(_02635_),
    .Y(_05173_));
 OR5x1_ASAP7_75t_R _16275_ (.A(_01546_),
    .B(_01547_),
    .C(_01548_),
    .D(_05168_),
    .E(_05173_),
    .Y(_05174_));
 BUFx3_ASAP7_75t_R _16276_ (.A(_05174_),
    .Y(_05175_));
 OR3x1_ASAP7_75t_R _16277_ (.A(_05160_),
    .B(_01575_),
    .C(_05175_),
    .Y(_05176_));
 OAI21x1_ASAP7_75t_R _16278_ (.A1(_05160_),
    .A2(_05175_),
    .B(_01575_),
    .Y(_05177_));
 AND3x1_ASAP7_75t_R _16279_ (.A(_05100_),
    .B(_05176_),
    .C(_05177_),
    .Y(_03461_));
 OR5x2_ASAP7_75t_R _16280_ (.A(_01550_),
    .B(_01551_),
    .C(_01554_),
    .D(_01565_),
    .E(_00034_),
    .Y(_05178_));
 OR5x2_ASAP7_75t_R _16281_ (.A(_01546_),
    .B(_01547_),
    .C(_01548_),
    .D(_05168_),
    .E(_05178_),
    .Y(_05179_));
 OR3x1_ASAP7_75t_R _16282_ (.A(_05160_),
    .B(_01575_),
    .C(_05179_),
    .Y(_05180_));
 XOR2x2_ASAP7_75t_R _16283_ (.A(_01574_),
    .B(_05180_),
    .Y(_05181_));
 AND2x2_ASAP7_75t_R _16284_ (.A(_05154_),
    .B(_05181_),
    .Y(_03462_));
 OR4x1_ASAP7_75t_R _16285_ (.A(_05160_),
    .B(_01574_),
    .C(_01575_),
    .D(_05175_),
    .Y(_05182_));
 XOR2x2_ASAP7_75t_R _16286_ (.A(_01573_),
    .B(_05182_),
    .Y(_05183_));
 AND2x2_ASAP7_75t_R _16287_ (.A(_05154_),
    .B(_05183_),
    .Y(_03463_));
 OR4x1_ASAP7_75t_R _16288_ (.A(_05160_),
    .B(_01573_),
    .C(_01574_),
    .D(_01575_),
    .Y(_05184_));
 OR3x1_ASAP7_75t_R _16289_ (.A(_01572_),
    .B(_05179_),
    .C(_05184_),
    .Y(_05185_));
 OAI21x1_ASAP7_75t_R _16290_ (.A1(_05179_),
    .A2(_05184_),
    .B(_01572_),
    .Y(_05186_));
 AND3x1_ASAP7_75t_R _16291_ (.A(_05100_),
    .B(_05185_),
    .C(_05186_),
    .Y(_03464_));
 OR3x1_ASAP7_75t_R _16292_ (.A(_01572_),
    .B(_05175_),
    .C(_05184_),
    .Y(_05187_));
 XOR2x2_ASAP7_75t_R _16293_ (.A(_01571_),
    .B(_05187_),
    .Y(_05188_));
 AND2x2_ASAP7_75t_R _16294_ (.A(_05154_),
    .B(_05188_),
    .Y(_03465_));
 OR4x1_ASAP7_75t_R _16295_ (.A(_01571_),
    .B(_01572_),
    .C(_05179_),
    .D(_05184_),
    .Y(_05189_));
 XOR2x2_ASAP7_75t_R _16296_ (.A(_01570_),
    .B(_05189_),
    .Y(_05190_));
 AND2x2_ASAP7_75t_R _16297_ (.A(_05154_),
    .B(_05190_),
    .Y(_03466_));
 OR4x1_ASAP7_75t_R _16298_ (.A(_01570_),
    .B(_01571_),
    .C(_01572_),
    .D(_05184_),
    .Y(_05191_));
 OR3x2_ASAP7_75t_R _16299_ (.A(_01569_),
    .B(_05175_),
    .C(_05191_),
    .Y(_05192_));
 OAI21x1_ASAP7_75t_R _16300_ (.A1(_05175_),
    .A2(_05191_),
    .B(_01569_),
    .Y(_05193_));
 AND3x1_ASAP7_75t_R _16301_ (.A(_05100_),
    .B(_05192_),
    .C(_05193_),
    .Y(_03467_));
 OR3x2_ASAP7_75t_R _16302_ (.A(_01569_),
    .B(_05179_),
    .C(_05191_),
    .Y(_05194_));
 XOR2x2_ASAP7_75t_R _16303_ (.A(_05159_),
    .B(_05194_),
    .Y(_05195_));
 AND2x2_ASAP7_75t_R _16304_ (.A(_05154_),
    .B(_05195_),
    .Y(_03468_));
 OR3x1_ASAP7_75t_R _16305_ (.A(_01567_),
    .B(_05159_),
    .C(_05192_),
    .Y(_05196_));
 OAI21x1_ASAP7_75t_R _16306_ (.A1(_05159_),
    .A2(_05192_),
    .B(_01567_),
    .Y(_05197_));
 AND3x1_ASAP7_75t_R _16307_ (.A(_05100_),
    .B(_05196_),
    .C(_05197_),
    .Y(_03469_));
 OR3x1_ASAP7_75t_R _16308_ (.A(_01567_),
    .B(_05159_),
    .C(_05194_),
    .Y(_05198_));
 XOR2x2_ASAP7_75t_R _16309_ (.A(_01566_),
    .B(_05198_),
    .Y(_05199_));
 AND2x2_ASAP7_75t_R _16310_ (.A(_05154_),
    .B(_05199_),
    .Y(_03470_));
 NOR2x1_ASAP7_75t_R _16311_ (.A(_10716_),
    .B(_02636_),
    .Y(_03471_));
 OR4x1_ASAP7_75t_R _16312_ (.A(_01566_),
    .B(_01567_),
    .C(_05159_),
    .D(_05192_),
    .Y(_05200_));
 XOR2x2_ASAP7_75t_R _16313_ (.A(_01564_),
    .B(_05200_),
    .Y(_05201_));
 AND2x2_ASAP7_75t_R _16314_ (.A(_05154_),
    .B(_05201_),
    .Y(_03472_));
 BUFx6f_ASAP7_75t_R _16315_ (.A(_11507_),
    .Y(_05202_));
 OR5x1_ASAP7_75t_R _16316_ (.A(_01564_),
    .B(_01566_),
    .C(_01567_),
    .D(_05159_),
    .E(_05194_),
    .Y(_05203_));
 XOR2x2_ASAP7_75t_R _16317_ (.A(_01563_),
    .B(_05203_),
    .Y(_05204_));
 AND2x2_ASAP7_75t_R _16318_ (.A(_05202_),
    .B(_05204_),
    .Y(_03473_));
 BUFx6f_ASAP7_75t_R _16319_ (.A(_08581_),
    .Y(_05205_));
 OR5x2_ASAP7_75t_R _16320_ (.A(_01563_),
    .B(_01564_),
    .C(_01566_),
    .D(_01567_),
    .E(_05159_),
    .Y(_05206_));
 OR3x1_ASAP7_75t_R _16321_ (.A(_01562_),
    .B(_05192_),
    .C(_05206_),
    .Y(_05207_));
 OAI21x1_ASAP7_75t_R _16322_ (.A1(_05192_),
    .A2(_05206_),
    .B(_01562_),
    .Y(_05208_));
 AND3x1_ASAP7_75t_R _16323_ (.A(_05205_),
    .B(_05207_),
    .C(_05208_),
    .Y(_03474_));
 OR4x1_ASAP7_75t_R _16324_ (.A(_01561_),
    .B(_01562_),
    .C(_05194_),
    .D(_05206_),
    .Y(_05209_));
 OR3x1_ASAP7_75t_R _16325_ (.A(_01562_),
    .B(_05194_),
    .C(_05206_),
    .Y(_05210_));
 NAND2x1_ASAP7_75t_R _16326_ (.A(_01561_),
    .B(_05210_),
    .Y(_05211_));
 AND3x1_ASAP7_75t_R _16327_ (.A(_05205_),
    .B(_05209_),
    .C(_05211_),
    .Y(_03475_));
 OR4x1_ASAP7_75t_R _16328_ (.A(_01561_),
    .B(_01562_),
    .C(_05192_),
    .D(_05206_),
    .Y(_05212_));
 XOR2x2_ASAP7_75t_R _16329_ (.A(_05164_),
    .B(_05212_),
    .Y(_05213_));
 AND2x2_ASAP7_75t_R _16330_ (.A(_05202_),
    .B(_05213_),
    .Y(_03476_));
 OR3x1_ASAP7_75t_R _16331_ (.A(_01559_),
    .B(_05164_),
    .C(_05209_),
    .Y(_05214_));
 OAI21x1_ASAP7_75t_R _16332_ (.A1(_05164_),
    .A2(_05209_),
    .B(_01559_),
    .Y(_05215_));
 AND3x1_ASAP7_75t_R _16333_ (.A(_05205_),
    .B(_05214_),
    .C(_05215_),
    .Y(_03477_));
 OR3x1_ASAP7_75t_R _16334_ (.A(_01559_),
    .B(_05164_),
    .C(_05212_),
    .Y(_05216_));
 XOR2x2_ASAP7_75t_R _16335_ (.A(_01558_),
    .B(_05216_),
    .Y(_05217_));
 AND2x2_ASAP7_75t_R _16336_ (.A(_05202_),
    .B(_05217_),
    .Y(_03478_));
 OR4x1_ASAP7_75t_R _16337_ (.A(_01558_),
    .B(_01559_),
    .C(_05164_),
    .D(_05209_),
    .Y(_05218_));
 XOR2x2_ASAP7_75t_R _16338_ (.A(_01557_),
    .B(_05218_),
    .Y(_05219_));
 AND2x2_ASAP7_75t_R _16339_ (.A(_05202_),
    .B(_05219_),
    .Y(_03479_));
 OR5x1_ASAP7_75t_R _16340_ (.A(_01557_),
    .B(_01558_),
    .C(_01559_),
    .D(_05164_),
    .E(_05212_),
    .Y(_05220_));
 XOR2x2_ASAP7_75t_R _16341_ (.A(_01556_),
    .B(_05220_),
    .Y(_05221_));
 AND2x2_ASAP7_75t_R _16342_ (.A(_05202_),
    .B(_05221_),
    .Y(_03480_));
 OR5x2_ASAP7_75t_R _16343_ (.A(_01556_),
    .B(_01557_),
    .C(_01558_),
    .D(_01559_),
    .E(_05164_),
    .Y(_05222_));
 OR3x1_ASAP7_75t_R _16344_ (.A(_01555_),
    .B(_05209_),
    .C(_05222_),
    .Y(_05223_));
 OAI21x1_ASAP7_75t_R _16345_ (.A1(_05209_),
    .A2(_05222_),
    .B(_01555_),
    .Y(_05224_));
 AND3x1_ASAP7_75t_R _16346_ (.A(_05205_),
    .B(_05223_),
    .C(_05224_),
    .Y(_03481_));
 XOR2x2_ASAP7_75t_R _16347_ (.A(_01554_),
    .B(_02635_),
    .Y(_05225_));
 AND2x2_ASAP7_75t_R _16348_ (.A(_05202_),
    .B(_05225_),
    .Y(_03482_));
 OR3x1_ASAP7_75t_R _16349_ (.A(_01555_),
    .B(_05212_),
    .C(_05222_),
    .Y(_05226_));
 XOR2x2_ASAP7_75t_R _16350_ (.A(_01553_),
    .B(_05226_),
    .Y(_05227_));
 AND2x2_ASAP7_75t_R _16351_ (.A(_05202_),
    .B(_05227_),
    .Y(_03483_));
 OR4x1_ASAP7_75t_R _16352_ (.A(_01553_),
    .B(_01555_),
    .C(_05209_),
    .D(_05222_),
    .Y(_05228_));
 XOR2x2_ASAP7_75t_R _16353_ (.A(_01552_),
    .B(_05228_),
    .Y(_05229_));
 AND2x2_ASAP7_75t_R _16354_ (.A(_05202_),
    .B(_05229_),
    .Y(_03484_));
 OR3x1_ASAP7_75t_R _16355_ (.A(_01554_),
    .B(_01565_),
    .C(_00034_),
    .Y(_05230_));
 XOR2x2_ASAP7_75t_R _16356_ (.A(_01551_),
    .B(_05230_),
    .Y(_05231_));
 AND2x2_ASAP7_75t_R _16357_ (.A(_05202_),
    .B(_05231_),
    .Y(_03485_));
 OR3x1_ASAP7_75t_R _16358_ (.A(_01551_),
    .B(_01554_),
    .C(_02635_),
    .Y(_05232_));
 NAND2x1_ASAP7_75t_R _16359_ (.A(_01550_),
    .B(_05232_),
    .Y(_05233_));
 AND3x1_ASAP7_75t_R _16360_ (.A(_05205_),
    .B(_05173_),
    .C(_05233_),
    .Y(_03486_));
 XOR2x2_ASAP7_75t_R _16361_ (.A(_05168_),
    .B(_05178_),
    .Y(_05234_));
 AND2x2_ASAP7_75t_R _16362_ (.A(_05202_),
    .B(_05234_),
    .Y(_03487_));
 OR3x1_ASAP7_75t_R _16363_ (.A(_01548_),
    .B(_05168_),
    .C(_05173_),
    .Y(_05235_));
 OAI21x1_ASAP7_75t_R _16364_ (.A1(_05168_),
    .A2(_05173_),
    .B(_01548_),
    .Y(_05236_));
 AND3x1_ASAP7_75t_R _16365_ (.A(_05205_),
    .B(_05235_),
    .C(_05236_),
    .Y(_03488_));
 BUFx6f_ASAP7_75t_R _16366_ (.A(_11507_),
    .Y(_05237_));
 OR3x1_ASAP7_75t_R _16367_ (.A(_01548_),
    .B(_05168_),
    .C(_05178_),
    .Y(_05238_));
 XOR2x2_ASAP7_75t_R _16368_ (.A(_01547_),
    .B(_05238_),
    .Y(_05239_));
 AND2x2_ASAP7_75t_R _16369_ (.A(_05237_),
    .B(_05239_),
    .Y(_03489_));
 OR4x1_ASAP7_75t_R _16370_ (.A(_01547_),
    .B(_01548_),
    .C(_05168_),
    .D(_05173_),
    .Y(_05240_));
 NAND2x1_ASAP7_75t_R _16371_ (.A(_01546_),
    .B(_05240_),
    .Y(_05241_));
 AND3x1_ASAP7_75t_R _16372_ (.A(_05205_),
    .B(_05175_),
    .C(_05241_),
    .Y(_03490_));
 XOR2x2_ASAP7_75t_R _16373_ (.A(_05160_),
    .B(_05179_),
    .Y(_05242_));
 AND2x2_ASAP7_75t_R _16374_ (.A(_05237_),
    .B(_05242_),
    .Y(_03491_));
 AND2x2_ASAP7_75t_R _16375_ (.A(_05237_),
    .B(_00016_),
    .Y(_03492_));
 INVx1_ASAP7_75t_R _16376_ (.A(_02131_),
    .Y(_05243_));
 BUFx6f_ASAP7_75t_R _16377_ (.A(_02127_),
    .Y(_05244_));
 INVx1_ASAP7_75t_R _16378_ (.A(_05244_),
    .Y(_05245_));
 OR2x2_ASAP7_75t_R _16379_ (.A(_01615_),
    .B(_01620_),
    .Y(_05246_));
 OR4x1_ASAP7_75t_R _16380_ (.A(_01577_),
    .B(\xs[10].cli1.i[35] ),
    .C(_01579_),
    .D(\xs[10].cli1.i[33] ),
    .Y(_05247_));
 OR3x2_ASAP7_75t_R _16381_ (.A(_01576_),
    .B(\peo[21][32] ),
    .C(_05247_),
    .Y(_05248_));
 AO21x1_ASAP7_75t_R _16382_ (.A1(\xs[10].cli1.i[39] ),
    .A2(_05247_),
    .B(_05244_),
    .Y(_05249_));
 AND4x1_ASAP7_75t_R _16383_ (.A(\peo[20][36] ),
    .B(_01617_),
    .C(\peo[20][34] ),
    .D(_01619_),
    .Y(_05250_));
 NOR2x1_ASAP7_75t_R _16384_ (.A(_01615_),
    .B(_05250_),
    .Y(_05251_));
 AO221x1_ASAP7_75t_R _16385_ (.A1(_05245_),
    .A2(_05246_),
    .B1(_05248_),
    .B2(_05249_),
    .C(_05251_),
    .Y(_05252_));
 INVx2_ASAP7_75t_R _16386_ (.A(_02120_),
    .Y(_05253_));
 AND2x4_ASAP7_75t_R _16387_ (.A(_05253_),
    .B(_02121_),
    .Y(_05254_));
 AND3x4_ASAP7_75t_R _16388_ (.A(_05244_),
    .B(_05252_),
    .C(_05254_),
    .Y(_05255_));
 AND2x2_ASAP7_75t_R _16389_ (.A(_05243_),
    .B(_05255_),
    .Y(_05256_));
 NOR2x1_ASAP7_75t_R _16390_ (.A(\peo[21][0] ),
    .B(_05248_),
    .Y(_05257_));
 OA211x2_ASAP7_75t_R _16391_ (.A1(_01581_),
    .A2(_05247_),
    .B(_05244_),
    .C(\xs[10].cli1.i[39] ),
    .Y(_05258_));
 AND4x1_ASAP7_75t_R _16392_ (.A(_02120_),
    .B(_00016_),
    .C(\xs[10].cli1.i[39] ),
    .D(_05247_),
    .Y(_05259_));
 AOI21x1_ASAP7_75t_R _16393_ (.A1(_05253_),
    .A2(_05258_),
    .B(_05259_),
    .Y(_05260_));
 OR2x6_ASAP7_75t_R _16394_ (.A(_01615_),
    .B(_05250_),
    .Y(_05261_));
 NAND2x1_ASAP7_75t_R _16395_ (.A(\xs[10].cli1.i[39] ),
    .B(_05247_),
    .Y(_05262_));
 OA21x2_ASAP7_75t_R _16396_ (.A1(_05261_),
    .A2(_05248_),
    .B(_05262_),
    .Y(_05263_));
 OA33x2_ASAP7_75t_R _16397_ (.A1(_01615_),
    .A2(_05250_),
    .A3(_05260_),
    .B1(_05263_),
    .B2(_02121_),
    .B3(_02120_),
    .Y(_05264_));
 INVx1_ASAP7_75t_R _16398_ (.A(_02121_),
    .Y(_05265_));
 OA21x2_ASAP7_75t_R _16399_ (.A1(_05265_),
    .A2(_05244_),
    .B(_05253_),
    .Y(_05266_));
 OA21x2_ASAP7_75t_R _16400_ (.A1(_05259_),
    .A2(_05266_),
    .B(_05251_),
    .Y(_05267_));
 OA21x2_ASAP7_75t_R _16401_ (.A1(_05248_),
    .A2(_05267_),
    .B(_01622_),
    .Y(_05268_));
 AOI211x1_ASAP7_75t_R _16402_ (.A1(_05257_),
    .A2(_05264_),
    .B(_05268_),
    .C(_05255_),
    .Y(_05269_));
 OA21x2_ASAP7_75t_R _16403_ (.A1(_05256_),
    .A2(_05269_),
    .B(_11397_),
    .Y(_03493_));
 NAND2x2_ASAP7_75t_R _16404_ (.A(_09229_),
    .B(_05255_),
    .Y(_05270_));
 NOR2x1_ASAP7_75t_R _16405_ (.A(_02130_),
    .B(_05270_),
    .Y(_03494_));
 NOR2x1_ASAP7_75t_R _16406_ (.A(_02129_),
    .B(_05270_),
    .Y(_03495_));
 NOR2x1_ASAP7_75t_R _16407_ (.A(_02128_),
    .B(_05270_),
    .Y(_03496_));
 NOR2x1_ASAP7_75t_R _16408_ (.A(_02119_),
    .B(_05270_),
    .Y(_03497_));
 NOR2x1_ASAP7_75t_R _16409_ (.A(_02118_),
    .B(_05270_),
    .Y(_03498_));
 NAND2x1_ASAP7_75t_R _16410_ (.A(_05252_),
    .B(_05254_),
    .Y(_05271_));
 OAI21x1_ASAP7_75t_R _16411_ (.A1(_05244_),
    .A2(_05271_),
    .B(_01622_),
    .Y(_05272_));
 OR3x1_ASAP7_75t_R _16412_ (.A(_05244_),
    .B(_05243_),
    .C(_05271_),
    .Y(_05273_));
 AND2x2_ASAP7_75t_R _16413_ (.A(_08584_),
    .B(_05264_),
    .Y(_05274_));
 NOR2x1_ASAP7_75t_R _16414_ (.A(_09934_),
    .B(_01583_),
    .Y(_05275_));
 INVx1_ASAP7_75t_R _16415_ (.A(_05264_),
    .Y(_05276_));
 AO32x1_ASAP7_75t_R _16416_ (.A1(_05272_),
    .A2(_05273_),
    .A3(_05274_),
    .B1(_05275_),
    .B2(_05276_),
    .Y(_03499_));
 OR3x2_ASAP7_75t_R _16417_ (.A(_10763_),
    .B(_05244_),
    .C(_05271_),
    .Y(_05277_));
 NOR2x1_ASAP7_75t_R _16418_ (.A(_02130_),
    .B(_05277_),
    .Y(_03500_));
 NOR2x1_ASAP7_75t_R _16419_ (.A(_02129_),
    .B(_05277_),
    .Y(_03501_));
 NOR2x1_ASAP7_75t_R _16420_ (.A(_02128_),
    .B(_05277_),
    .Y(_03502_));
 NOR2x1_ASAP7_75t_R _16421_ (.A(_02119_),
    .B(_05277_),
    .Y(_03503_));
 NOR2x1_ASAP7_75t_R _16422_ (.A(_02118_),
    .B(_05277_),
    .Y(_03504_));
 OA211x2_ASAP7_75t_R _16423_ (.A1(_02120_),
    .A2(_02121_),
    .B(_05247_),
    .C(\xs[10].cli1.i[39] ),
    .Y(_05278_));
 OAI21x1_ASAP7_75t_R _16424_ (.A1(_05261_),
    .A2(_05260_),
    .B(_05278_),
    .Y(_05279_));
 NAND2x1_ASAP7_75t_R _16425_ (.A(_01622_),
    .B(_05279_),
    .Y(_05280_));
 OA21x2_ASAP7_75t_R _16426_ (.A1(_05261_),
    .A2(_05260_),
    .B(_05278_),
    .Y(_05281_));
 NAND2x1_ASAP7_75t_R _16427_ (.A(_01583_),
    .B(_05281_),
    .Y(_05282_));
 AOI21x1_ASAP7_75t_R _16428_ (.A1(_02121_),
    .A2(_05252_),
    .B(_02120_),
    .Y(_05283_));
 NOR2x1_ASAP7_75t_R _16429_ (.A(_10826_),
    .B(_05283_),
    .Y(_05284_));
 NOR2x1_ASAP7_75t_R _16430_ (.A(_09934_),
    .B(_02131_),
    .Y(_05285_));
 AO32x1_ASAP7_75t_R _16431_ (.A1(_05280_),
    .A2(_05282_),
    .A3(_05284_),
    .B1(_05285_),
    .B2(_05283_),
    .Y(_03505_));
 NAND2x2_ASAP7_75t_R _16432_ (.A(_08876_),
    .B(_05283_),
    .Y(_05286_));
 NOR2x1_ASAP7_75t_R _16433_ (.A(_02130_),
    .B(_05286_),
    .Y(_03506_));
 NOR2x1_ASAP7_75t_R _16434_ (.A(_02129_),
    .B(_05286_),
    .Y(_03507_));
 NOR2x1_ASAP7_75t_R _16435_ (.A(_02128_),
    .B(_05286_),
    .Y(_03508_));
 NAND2x1_ASAP7_75t_R _16436_ (.A(_01620_),
    .B(_05279_),
    .Y(_05287_));
 NAND2x1_ASAP7_75t_R _16437_ (.A(_01581_),
    .B(_05281_),
    .Y(_05288_));
 NOR2x1_ASAP7_75t_R _16438_ (.A(_09934_),
    .B(_05244_),
    .Y(_05289_));
 AO32x1_ASAP7_75t_R _16439_ (.A1(_05284_),
    .A2(_05287_),
    .A3(_05288_),
    .B1(_05289_),
    .B2(_05283_),
    .Y(_03509_));
 NAND2x1_ASAP7_75t_R _16440_ (.A(_01619_),
    .B(_05279_),
    .Y(_05290_));
 NAND2x1_ASAP7_75t_R _16441_ (.A(_01580_),
    .B(_05281_),
    .Y(_05291_));
 NOR2x1_ASAP7_75t_R _16442_ (.A(_09934_),
    .B(_02126_),
    .Y(_05292_));
 AO32x1_ASAP7_75t_R _16443_ (.A1(_05284_),
    .A2(_05290_),
    .A3(_05291_),
    .B1(_05292_),
    .B2(_05283_),
    .Y(_03510_));
 AO32x1_ASAP7_75t_R _16444_ (.A1(\xs[10].cli1.i[39] ),
    .A2(_01579_),
    .A3(_05264_),
    .B1(_05279_),
    .B2(_01618_),
    .Y(_05293_));
 OR2x6_ASAP7_75t_R _16445_ (.A(_10826_),
    .B(_05283_),
    .Y(_05294_));
 OAI22x1_ASAP7_75t_R _16446_ (.A1(_02125_),
    .A2(_05286_),
    .B1(_05293_),
    .B2(_05294_),
    .Y(_03511_));
 NAND2x1_ASAP7_75t_R _16447_ (.A(_01617_),
    .B(_05279_),
    .Y(_05295_));
 NAND2x1_ASAP7_75t_R _16448_ (.A(_01578_),
    .B(_05281_),
    .Y(_05296_));
 NOR2x1_ASAP7_75t_R _16449_ (.A(_09934_),
    .B(_02124_),
    .Y(_05297_));
 AO32x1_ASAP7_75t_R _16450_ (.A1(_05284_),
    .A2(_05295_),
    .A3(_05296_),
    .B1(_05297_),
    .B2(_05283_),
    .Y(_03512_));
 AO32x1_ASAP7_75t_R _16451_ (.A1(\xs[10].cli1.i[39] ),
    .A2(_01577_),
    .A3(_05264_),
    .B1(_05279_),
    .B2(_01616_),
    .Y(_05298_));
 OAI22x1_ASAP7_75t_R _16452_ (.A1(_02123_),
    .A2(_05286_),
    .B1(_05298_),
    .B2(_05294_),
    .Y(_03513_));
 NOR2x1_ASAP7_75t_R _16453_ (.A(_02122_),
    .B(_05286_),
    .Y(_03514_));
 OR4x1_ASAP7_75t_R _16454_ (.A(_08684_),
    .B(_02120_),
    .C(_05265_),
    .D(_05252_),
    .Y(_05299_));
 INVx1_ASAP7_75t_R _16455_ (.A(_05299_),
    .Y(_03515_));
 BUFx12f_ASAP7_75t_R _16456_ (.A(_10012_),
    .Y(_05300_));
 AOI211x1_ASAP7_75t_R _16457_ (.A1(\xs[10].cli1.i[39] ),
    .A2(_05247_),
    .B(_05283_),
    .C(_05251_),
    .Y(_05301_));
 NOR2x1_ASAP7_75t_R _16458_ (.A(_05300_),
    .B(_05301_),
    .Y(_03516_));
 NOR2x1_ASAP7_75t_R _16459_ (.A(_02119_),
    .B(_05286_),
    .Y(_03517_));
 NOR2x1_ASAP7_75t_R _16460_ (.A(_02118_),
    .B(_05286_),
    .Y(_03518_));
 BUFx3_ASAP7_75t_R _16461_ (.A(_01507_),
    .Y(_05302_));
 BUFx3_ASAP7_75t_R _16462_ (.A(_01480_),
    .Y(_05303_));
 AND4x1_ASAP7_75t_R _16463_ (.A(_05303_),
    .B(_01508_),
    .C(_01509_),
    .D(_01510_),
    .Y(_05304_));
 AND5x1_ASAP7_75t_R _16464_ (.A(_01499_),
    .B(_01504_),
    .C(_01505_),
    .D(_05302_),
    .E(_05304_),
    .Y(_05305_));
 AND5x2_ASAP7_75t_R _16465_ (.A(_01501_),
    .B(_01502_),
    .C(_01503_),
    .D(_11466_),
    .E(_05305_),
    .Y(_05306_));
 AND4x1_ASAP7_75t_R _16466_ (.A(_01494_),
    .B(_01495_),
    .C(_01496_),
    .D(_01497_),
    .Y(_05307_));
 AND4x1_ASAP7_75t_R _16467_ (.A(_01488_),
    .B(_01490_),
    .C(_01491_),
    .D(_01498_),
    .Y(_05308_));
 AND5x1_ASAP7_75t_R _16468_ (.A(_01481_),
    .B(_01482_),
    .C(_01487_),
    .D(_01506_),
    .E(_05308_),
    .Y(_05309_));
 AND3x1_ASAP7_75t_R _16469_ (.A(_01485_),
    .B(_01486_),
    .C(_01489_),
    .Y(_05310_));
 OR3x1_ASAP7_75t_R _16470_ (.A(_01483_),
    .B(_01484_),
    .C(_05310_),
    .Y(_05311_));
 AND5x2_ASAP7_75t_R _16471_ (.A(_01492_),
    .B(_01493_),
    .C(_05307_),
    .D(_05309_),
    .E(_05311_),
    .Y(_05312_));
 NAND2x2_ASAP7_75t_R _16472_ (.A(_05306_),
    .B(_05312_),
    .Y(_05313_));
 NOR2x1_ASAP7_75t_R _16473_ (.A(_01437_),
    .B(_05313_),
    .Y(_03519_));
 INVx1_ASAP7_75t_R _16474_ (.A(_05313_),
    .Y(_03520_));
 NOR2x1_ASAP7_75t_R _16475_ (.A(_01440_),
    .B(_05313_),
    .Y(_03521_));
 NOR2x1_ASAP7_75t_R _16476_ (.A(_01439_),
    .B(_05313_),
    .Y(_03522_));
 NOR2x1_ASAP7_75t_R _16477_ (.A(_01438_),
    .B(_05313_),
    .Y(_03523_));
 NOR2x1_ASAP7_75t_R _16478_ (.A(_01436_),
    .B(_05313_),
    .Y(_03524_));
 NOR2x1_ASAP7_75t_R _16479_ (.A(_01435_),
    .B(_05313_),
    .Y(_03525_));
 INVx1_ASAP7_75t_R _16480_ (.A(_05313_),
    .Y(_03526_));
 AND2x2_ASAP7_75t_R _16481_ (.A(_05237_),
    .B(_00035_),
    .Y(_03527_));
 OR4x1_ASAP7_75t_R _16482_ (.A(_01485_),
    .B(_01486_),
    .C(_01489_),
    .D(_02637_),
    .Y(_05314_));
 OR4x1_ASAP7_75t_R _16483_ (.A(_01481_),
    .B(_01482_),
    .C(_01483_),
    .D(_01484_),
    .Y(_05315_));
 OR2x6_ASAP7_75t_R _16484_ (.A(_05314_),
    .B(_05315_),
    .Y(_05316_));
 OR3x1_ASAP7_75t_R _16485_ (.A(_05303_),
    .B(_01510_),
    .C(_05316_),
    .Y(_05317_));
 OAI21x1_ASAP7_75t_R _16486_ (.A1(_05303_),
    .A2(_05316_),
    .B(_01510_),
    .Y(_05318_));
 AND3x1_ASAP7_75t_R _16487_ (.A(_05205_),
    .B(_05317_),
    .C(_05318_),
    .Y(_03528_));
 OR5x2_ASAP7_75t_R _16488_ (.A(_01485_),
    .B(_01486_),
    .C(_01489_),
    .D(_01500_),
    .E(_00035_),
    .Y(_05319_));
 OR2x2_ASAP7_75t_R _16489_ (.A(_05315_),
    .B(_05319_),
    .Y(_05320_));
 OR3x1_ASAP7_75t_R _16490_ (.A(_05303_),
    .B(_01510_),
    .C(_05320_),
    .Y(_05321_));
 XOR2x2_ASAP7_75t_R _16491_ (.A(_01509_),
    .B(_05321_),
    .Y(_05322_));
 AND2x2_ASAP7_75t_R _16492_ (.A(_05237_),
    .B(_05322_),
    .Y(_03529_));
 OR4x1_ASAP7_75t_R _16493_ (.A(_05303_),
    .B(_01508_),
    .C(_01509_),
    .D(_01510_),
    .Y(_05323_));
 OR3x2_ASAP7_75t_R _16494_ (.A(_05314_),
    .B(_05315_),
    .C(_05323_),
    .Y(_05324_));
 OR4x1_ASAP7_75t_R _16495_ (.A(_05303_),
    .B(_01509_),
    .C(_01510_),
    .D(_05316_),
    .Y(_05325_));
 NAND2x1_ASAP7_75t_R _16496_ (.A(_01508_),
    .B(_05325_),
    .Y(_05326_));
 AND3x1_ASAP7_75t_R _16497_ (.A(_05205_),
    .B(_05324_),
    .C(_05326_),
    .Y(_03530_));
 OR3x2_ASAP7_75t_R _16498_ (.A(_05315_),
    .B(_05319_),
    .C(_05323_),
    .Y(_05327_));
 XOR2x2_ASAP7_75t_R _16499_ (.A(_05302_),
    .B(_05327_),
    .Y(_05328_));
 AND2x2_ASAP7_75t_R _16500_ (.A(_05237_),
    .B(_05328_),
    .Y(_03531_));
 OR3x1_ASAP7_75t_R _16501_ (.A(_01506_),
    .B(_05302_),
    .C(_05324_),
    .Y(_05329_));
 OAI21x1_ASAP7_75t_R _16502_ (.A1(_05302_),
    .A2(_05324_),
    .B(_01506_),
    .Y(_05330_));
 AND3x1_ASAP7_75t_R _16503_ (.A(_05205_),
    .B(_05329_),
    .C(_05330_),
    .Y(_03532_));
 OR3x1_ASAP7_75t_R _16504_ (.A(_01506_),
    .B(_05302_),
    .C(_05327_),
    .Y(_05331_));
 XOR2x2_ASAP7_75t_R _16505_ (.A(_01505_),
    .B(_05331_),
    .Y(_05332_));
 AND2x2_ASAP7_75t_R _16506_ (.A(_05237_),
    .B(_05332_),
    .Y(_03533_));
 OR4x1_ASAP7_75t_R _16507_ (.A(_01505_),
    .B(_01506_),
    .C(_05302_),
    .D(_05324_),
    .Y(_05333_));
 XOR2x2_ASAP7_75t_R _16508_ (.A(_01504_),
    .B(_05333_),
    .Y(_05334_));
 AND2x2_ASAP7_75t_R _16509_ (.A(_05237_),
    .B(_05334_),
    .Y(_03534_));
 OR5x1_ASAP7_75t_R _16510_ (.A(_01504_),
    .B(_01505_),
    .C(_01506_),
    .D(_05302_),
    .E(_05327_),
    .Y(_05335_));
 XOR2x2_ASAP7_75t_R _16511_ (.A(_01503_),
    .B(_05335_),
    .Y(_05336_));
 AND2x2_ASAP7_75t_R _16512_ (.A(_05237_),
    .B(_05336_),
    .Y(_03535_));
 BUFx12f_ASAP7_75t_R _16513_ (.A(_08527_),
    .Y(_05337_));
 BUFx6f_ASAP7_75t_R _16514_ (.A(_05337_),
    .Y(_05338_));
 OR5x2_ASAP7_75t_R _16515_ (.A(_01503_),
    .B(_01504_),
    .C(_01505_),
    .D(_01506_),
    .E(_05302_),
    .Y(_05339_));
 OR3x2_ASAP7_75t_R _16516_ (.A(_01502_),
    .B(_05324_),
    .C(_05339_),
    .Y(_05340_));
 OAI21x1_ASAP7_75t_R _16517_ (.A1(_05324_),
    .A2(_05339_),
    .B(_01502_),
    .Y(_05341_));
 AND3x1_ASAP7_75t_R _16518_ (.A(_05338_),
    .B(_05340_),
    .C(_05341_),
    .Y(_03536_));
 OR3x2_ASAP7_75t_R _16519_ (.A(_01502_),
    .B(_05327_),
    .C(_05339_),
    .Y(_05342_));
 XOR2x2_ASAP7_75t_R _16520_ (.A(_01501_),
    .B(_05342_),
    .Y(_05343_));
 AND2x2_ASAP7_75t_R _16521_ (.A(_05237_),
    .B(_05343_),
    .Y(_03537_));
 NOR2x1_ASAP7_75t_R _16522_ (.A(_05300_),
    .B(_02638_),
    .Y(_03538_));
 OR3x1_ASAP7_75t_R _16523_ (.A(_01499_),
    .B(_01501_),
    .C(_05340_),
    .Y(_05344_));
 OAI21x1_ASAP7_75t_R _16524_ (.A1(_01501_),
    .A2(_05340_),
    .B(_01499_),
    .Y(_05345_));
 AND3x1_ASAP7_75t_R _16525_ (.A(_05338_),
    .B(_05344_),
    .C(_05345_),
    .Y(_03539_));
 BUFx6f_ASAP7_75t_R _16526_ (.A(_11507_),
    .Y(_05346_));
 OR3x1_ASAP7_75t_R _16527_ (.A(_01499_),
    .B(_01501_),
    .C(_05342_),
    .Y(_05347_));
 XOR2x2_ASAP7_75t_R _16528_ (.A(_01498_),
    .B(_05347_),
    .Y(_05348_));
 AND2x2_ASAP7_75t_R _16529_ (.A(_05346_),
    .B(_05348_),
    .Y(_03540_));
 OR4x1_ASAP7_75t_R _16530_ (.A(_01498_),
    .B(_01499_),
    .C(_01501_),
    .D(_05340_),
    .Y(_05349_));
 XOR2x2_ASAP7_75t_R _16531_ (.A(_01497_),
    .B(_05349_),
    .Y(_05350_));
 AND2x2_ASAP7_75t_R _16532_ (.A(_05346_),
    .B(_05350_),
    .Y(_03541_));
 OR4x1_ASAP7_75t_R _16533_ (.A(_01497_),
    .B(_01498_),
    .C(_01499_),
    .D(_01501_),
    .Y(_05351_));
 OR3x2_ASAP7_75t_R _16534_ (.A(_01496_),
    .B(_05342_),
    .C(_05351_),
    .Y(_05352_));
 OAI21x1_ASAP7_75t_R _16535_ (.A1(_05342_),
    .A2(_05351_),
    .B(_01496_),
    .Y(_05353_));
 AND3x1_ASAP7_75t_R _16536_ (.A(_05338_),
    .B(_05352_),
    .C(_05353_),
    .Y(_03542_));
 OR3x2_ASAP7_75t_R _16537_ (.A(_01496_),
    .B(_05340_),
    .C(_05351_),
    .Y(_05354_));
 XOR2x2_ASAP7_75t_R _16538_ (.A(_01495_),
    .B(_05354_),
    .Y(_05355_));
 AND2x2_ASAP7_75t_R _16539_ (.A(_05346_),
    .B(_05355_),
    .Y(_03543_));
 OR3x1_ASAP7_75t_R _16540_ (.A(_01494_),
    .B(_01495_),
    .C(_05352_),
    .Y(_05356_));
 OAI21x1_ASAP7_75t_R _16541_ (.A1(_01495_),
    .A2(_05352_),
    .B(_01494_),
    .Y(_05357_));
 AND3x1_ASAP7_75t_R _16542_ (.A(_05338_),
    .B(_05356_),
    .C(_05357_),
    .Y(_03544_));
 OR3x1_ASAP7_75t_R _16543_ (.A(_01494_),
    .B(_01495_),
    .C(_05354_),
    .Y(_05358_));
 XOR2x2_ASAP7_75t_R _16544_ (.A(_01493_),
    .B(_05358_),
    .Y(_05359_));
 AND2x2_ASAP7_75t_R _16545_ (.A(_05346_),
    .B(_05359_),
    .Y(_03545_));
 OR4x1_ASAP7_75t_R _16546_ (.A(_01493_),
    .B(_01494_),
    .C(_01495_),
    .D(_05352_),
    .Y(_05360_));
 XOR2x2_ASAP7_75t_R _16547_ (.A(_01492_),
    .B(_05360_),
    .Y(_05361_));
 AND2x2_ASAP7_75t_R _16548_ (.A(_05346_),
    .B(_05361_),
    .Y(_03546_));
 OR4x1_ASAP7_75t_R _16549_ (.A(_01492_),
    .B(_01493_),
    .C(_01494_),
    .D(_01495_),
    .Y(_05362_));
 OR3x1_ASAP7_75t_R _16550_ (.A(_01491_),
    .B(_05354_),
    .C(_05362_),
    .Y(_05363_));
 OAI21x1_ASAP7_75t_R _16551_ (.A1(_05354_),
    .A2(_05362_),
    .B(_01491_),
    .Y(_05364_));
 AND3x1_ASAP7_75t_R _16552_ (.A(_05338_),
    .B(_05363_),
    .C(_05364_),
    .Y(_03547_));
 OR3x1_ASAP7_75t_R _16553_ (.A(_01491_),
    .B(_05352_),
    .C(_05362_),
    .Y(_05365_));
 XOR2x2_ASAP7_75t_R _16554_ (.A(_01490_),
    .B(_05365_),
    .Y(_05366_));
 AND2x2_ASAP7_75t_R _16555_ (.A(_05346_),
    .B(_05366_),
    .Y(_03548_));
 XOR2x2_ASAP7_75t_R _16556_ (.A(_01489_),
    .B(_02637_),
    .Y(_05367_));
 AND2x2_ASAP7_75t_R _16557_ (.A(_05346_),
    .B(_05367_),
    .Y(_03549_));
 OR4x1_ASAP7_75t_R _16558_ (.A(_01490_),
    .B(_01491_),
    .C(_05354_),
    .D(_05362_),
    .Y(_05368_));
 XOR2x2_ASAP7_75t_R _16559_ (.A(_01488_),
    .B(_05368_),
    .Y(_05369_));
 AND2x2_ASAP7_75t_R _16560_ (.A(_05346_),
    .B(_05369_),
    .Y(_03550_));
 OR5x1_ASAP7_75t_R _16561_ (.A(_01488_),
    .B(_01490_),
    .C(_01491_),
    .D(_05352_),
    .E(_05362_),
    .Y(_05370_));
 XOR2x2_ASAP7_75t_R _16562_ (.A(_01487_),
    .B(_05370_),
    .Y(_05371_));
 AND2x2_ASAP7_75t_R _16563_ (.A(_05346_),
    .B(_05371_),
    .Y(_03551_));
 OR3x1_ASAP7_75t_R _16564_ (.A(_01489_),
    .B(_01500_),
    .C(_00035_),
    .Y(_05372_));
 XOR2x2_ASAP7_75t_R _16565_ (.A(_01486_),
    .B(_05372_),
    .Y(_05373_));
 AND2x2_ASAP7_75t_R _16566_ (.A(_05346_),
    .B(_05373_),
    .Y(_03552_));
 OR3x1_ASAP7_75t_R _16567_ (.A(_01486_),
    .B(_01489_),
    .C(_02637_),
    .Y(_05374_));
 NAND2x1_ASAP7_75t_R _16568_ (.A(_01485_),
    .B(_05374_),
    .Y(_05375_));
 AND3x1_ASAP7_75t_R _16569_ (.A(_05338_),
    .B(_05314_),
    .C(_05375_),
    .Y(_03553_));
 BUFx6f_ASAP7_75t_R _16570_ (.A(_11507_),
    .Y(_05376_));
 XOR2x2_ASAP7_75t_R _16571_ (.A(_01484_),
    .B(_05319_),
    .Y(_05377_));
 AND2x2_ASAP7_75t_R _16572_ (.A(_05376_),
    .B(_05377_),
    .Y(_03554_));
 OR3x1_ASAP7_75t_R _16573_ (.A(_01483_),
    .B(_01484_),
    .C(_05314_),
    .Y(_05378_));
 OAI21x1_ASAP7_75t_R _16574_ (.A1(_01484_),
    .A2(_05314_),
    .B(_01483_),
    .Y(_05379_));
 AND3x1_ASAP7_75t_R _16575_ (.A(_05338_),
    .B(_05378_),
    .C(_05379_),
    .Y(_03555_));
 OR3x1_ASAP7_75t_R _16576_ (.A(_01483_),
    .B(_01484_),
    .C(_05319_),
    .Y(_05380_));
 XOR2x2_ASAP7_75t_R _16577_ (.A(_01482_),
    .B(_05380_),
    .Y(_05381_));
 AND2x2_ASAP7_75t_R _16578_ (.A(_05376_),
    .B(_05381_),
    .Y(_03556_));
 OR4x1_ASAP7_75t_R _16579_ (.A(_01482_),
    .B(_01483_),
    .C(_01484_),
    .D(_05314_),
    .Y(_05382_));
 NAND2x1_ASAP7_75t_R _16580_ (.A(_01481_),
    .B(_05382_),
    .Y(_05383_));
 AND3x1_ASAP7_75t_R _16581_ (.A(_05338_),
    .B(_05316_),
    .C(_05383_),
    .Y(_03557_));
 XOR2x2_ASAP7_75t_R _16582_ (.A(_05303_),
    .B(_05320_),
    .Y(_05384_));
 AND2x2_ASAP7_75t_R _16583_ (.A(_05376_),
    .B(_05384_),
    .Y(_03558_));
 BUFx6f_ASAP7_75t_R _16584_ (.A(_01464_),
    .Y(_05385_));
 BUFx6f_ASAP7_75t_R _16585_ (.A(_01441_),
    .Y(_05386_));
 AND4x1_ASAP7_75t_R _16586_ (.A(_05386_),
    .B(_01469_),
    .C(_01470_),
    .D(_01471_),
    .Y(_05387_));
 AND5x1_ASAP7_75t_R _16587_ (.A(_01460_),
    .B(_01465_),
    .C(_01466_),
    .D(_01468_),
    .E(_05387_),
    .Y(_05388_));
 AND5x2_ASAP7_75t_R _16588_ (.A(_01462_),
    .B(_01463_),
    .C(_05385_),
    .D(_11466_),
    .E(_05388_),
    .Y(_05389_));
 BUFx6f_ASAP7_75t_R _16589_ (.A(_01456_),
    .Y(_05390_));
 AND4x1_ASAP7_75t_R _16590_ (.A(_01455_),
    .B(_05390_),
    .C(_01457_),
    .D(_01458_),
    .Y(_05391_));
 AND4x1_ASAP7_75t_R _16591_ (.A(_01449_),
    .B(_01451_),
    .C(_01452_),
    .D(_01459_),
    .Y(_05392_));
 AND5x1_ASAP7_75t_R _16592_ (.A(_01442_),
    .B(_01443_),
    .C(_01448_),
    .D(_01467_),
    .E(_05392_),
    .Y(_05393_));
 AND3x1_ASAP7_75t_R _16593_ (.A(_01446_),
    .B(_01447_),
    .C(_01450_),
    .Y(_05394_));
 OR3x1_ASAP7_75t_R _16594_ (.A(_01444_),
    .B(_01445_),
    .C(_05394_),
    .Y(_05395_));
 AND5x2_ASAP7_75t_R _16595_ (.A(_01453_),
    .B(_01454_),
    .C(_05391_),
    .D(_05393_),
    .E(_05395_),
    .Y(_05396_));
 NAND2x2_ASAP7_75t_R _16596_ (.A(_05389_),
    .B(_05396_),
    .Y(_05397_));
 NOR2x1_ASAP7_75t_R _16597_ (.A(_01431_),
    .B(_05397_),
    .Y(_03559_));
 INVx1_ASAP7_75t_R _16598_ (.A(_05397_),
    .Y(_03560_));
 NOR2x1_ASAP7_75t_R _16599_ (.A(_01434_),
    .B(_05397_),
    .Y(_03561_));
 NOR2x1_ASAP7_75t_R _16600_ (.A(_01433_),
    .B(_05397_),
    .Y(_03562_));
 NOR2x1_ASAP7_75t_R _16601_ (.A(_01432_),
    .B(_05397_),
    .Y(_03563_));
 NOR2x1_ASAP7_75t_R _16602_ (.A(_01430_),
    .B(_05397_),
    .Y(_03564_));
 NOR2x1_ASAP7_75t_R _16603_ (.A(_01429_),
    .B(_05397_),
    .Y(_03565_));
 INVx1_ASAP7_75t_R _16604_ (.A(_05397_),
    .Y(_03566_));
 AND2x2_ASAP7_75t_R _16605_ (.A(_05376_),
    .B(_00036_),
    .Y(_03567_));
 OR4x1_ASAP7_75t_R _16606_ (.A(_01446_),
    .B(_01447_),
    .C(_01450_),
    .D(_02643_),
    .Y(_05398_));
 OR4x1_ASAP7_75t_R _16607_ (.A(_01442_),
    .B(_01443_),
    .C(_01444_),
    .D(_01445_),
    .Y(_05399_));
 OR2x6_ASAP7_75t_R _16608_ (.A(_05398_),
    .B(_05399_),
    .Y(_05400_));
 OR3x1_ASAP7_75t_R _16609_ (.A(_05386_),
    .B(_01471_),
    .C(_05400_),
    .Y(_05401_));
 OAI21x1_ASAP7_75t_R _16610_ (.A1(_05386_),
    .A2(_05400_),
    .B(_01471_),
    .Y(_05402_));
 AND3x1_ASAP7_75t_R _16611_ (.A(_05338_),
    .B(_05401_),
    .C(_05402_),
    .Y(_03568_));
 OR5x2_ASAP7_75t_R _16612_ (.A(_01446_),
    .B(_01447_),
    .C(_01450_),
    .D(_01461_),
    .E(_00036_),
    .Y(_05403_));
 OR2x6_ASAP7_75t_R _16613_ (.A(_05399_),
    .B(_05403_),
    .Y(_05404_));
 OR3x1_ASAP7_75t_R _16614_ (.A(_05386_),
    .B(_01471_),
    .C(_05404_),
    .Y(_05405_));
 XOR2x2_ASAP7_75t_R _16615_ (.A(_01470_),
    .B(_05405_),
    .Y(_05406_));
 AND2x2_ASAP7_75t_R _16616_ (.A(_05376_),
    .B(_05406_),
    .Y(_03569_));
 OR4x1_ASAP7_75t_R _16617_ (.A(_05386_),
    .B(_01470_),
    .C(_01471_),
    .D(_05400_),
    .Y(_05407_));
 XOR2x2_ASAP7_75t_R _16618_ (.A(_01469_),
    .B(_05407_),
    .Y(_05408_));
 AND2x2_ASAP7_75t_R _16619_ (.A(_05376_),
    .B(_05408_),
    .Y(_03570_));
 OR5x2_ASAP7_75t_R _16620_ (.A(_05386_),
    .B(_01468_),
    .C(_01469_),
    .D(_01470_),
    .E(_01471_),
    .Y(_05409_));
 OR5x1_ASAP7_75t_R _16621_ (.A(_05386_),
    .B(_01469_),
    .C(_01470_),
    .D(_01471_),
    .E(_05404_),
    .Y(_05410_));
 NAND2x1_ASAP7_75t_R _16622_ (.A(_01468_),
    .B(_05410_),
    .Y(_05411_));
 OA211x2_ASAP7_75t_R _16623_ (.A1(_05404_),
    .A2(_05409_),
    .B(_05411_),
    .C(_11589_),
    .Y(_03571_));
 OR3x2_ASAP7_75t_R _16624_ (.A(_05398_),
    .B(_05399_),
    .C(_05409_),
    .Y(_05412_));
 XOR2x2_ASAP7_75t_R _16625_ (.A(_01467_),
    .B(_05412_),
    .Y(_05413_));
 AND2x2_ASAP7_75t_R _16626_ (.A(_05376_),
    .B(_05413_),
    .Y(_03572_));
 OR3x1_ASAP7_75t_R _16627_ (.A(_01467_),
    .B(_05404_),
    .C(_05409_),
    .Y(_05414_));
 XOR2x2_ASAP7_75t_R _16628_ (.A(_01466_),
    .B(_05414_),
    .Y(_05415_));
 AND2x2_ASAP7_75t_R _16629_ (.A(_05376_),
    .B(_05415_),
    .Y(_03573_));
 OR4x1_ASAP7_75t_R _16630_ (.A(_01465_),
    .B(_01466_),
    .C(_01467_),
    .D(_05412_),
    .Y(_05416_));
 OR3x1_ASAP7_75t_R _16631_ (.A(_01466_),
    .B(_01467_),
    .C(_05412_),
    .Y(_05417_));
 NAND2x1_ASAP7_75t_R _16632_ (.A(_01465_),
    .B(_05417_),
    .Y(_05418_));
 AND3x1_ASAP7_75t_R _16633_ (.A(_05338_),
    .B(_05416_),
    .C(_05418_),
    .Y(_03574_));
 OR5x2_ASAP7_75t_R _16634_ (.A(_01465_),
    .B(_01466_),
    .C(_01467_),
    .D(_05404_),
    .E(_05409_),
    .Y(_05419_));
 XOR2x2_ASAP7_75t_R _16635_ (.A(_05385_),
    .B(_05419_),
    .Y(_05420_));
 AND2x2_ASAP7_75t_R _16636_ (.A(_05376_),
    .B(_05420_),
    .Y(_03575_));
 BUFx6f_ASAP7_75t_R _16637_ (.A(_05337_),
    .Y(_05421_));
 OR3x1_ASAP7_75t_R _16638_ (.A(_01463_),
    .B(_05385_),
    .C(_05416_),
    .Y(_05422_));
 OAI21x1_ASAP7_75t_R _16639_ (.A1(_05385_),
    .A2(_05416_),
    .B(_01463_),
    .Y(_05423_));
 AND3x1_ASAP7_75t_R _16640_ (.A(_05421_),
    .B(_05422_),
    .C(_05423_),
    .Y(_03576_));
 OR3x1_ASAP7_75t_R _16641_ (.A(_01463_),
    .B(_05385_),
    .C(_05419_),
    .Y(_05424_));
 XOR2x2_ASAP7_75t_R _16642_ (.A(_01462_),
    .B(_05424_),
    .Y(_05425_));
 AND2x2_ASAP7_75t_R _16643_ (.A(_05376_),
    .B(_05425_),
    .Y(_03577_));
 NOR2x1_ASAP7_75t_R _16644_ (.A(_05300_),
    .B(_02644_),
    .Y(_03578_));
 BUFx12f_ASAP7_75t_R _16645_ (.A(_08598_),
    .Y(_05426_));
 BUFx6f_ASAP7_75t_R _16646_ (.A(_05426_),
    .Y(_05427_));
 OR4x1_ASAP7_75t_R _16647_ (.A(_01462_),
    .B(_01463_),
    .C(_05385_),
    .D(_05416_),
    .Y(_05428_));
 XOR2x2_ASAP7_75t_R _16648_ (.A(_01460_),
    .B(_05428_),
    .Y(_05429_));
 AND2x2_ASAP7_75t_R _16649_ (.A(_05427_),
    .B(_05429_),
    .Y(_03579_));
 OR5x1_ASAP7_75t_R _16650_ (.A(_01460_),
    .B(_01462_),
    .C(_01463_),
    .D(_05385_),
    .E(_05419_),
    .Y(_05430_));
 XOR2x2_ASAP7_75t_R _16651_ (.A(_01459_),
    .B(_05430_),
    .Y(_05431_));
 AND2x2_ASAP7_75t_R _16652_ (.A(_05427_),
    .B(_05431_),
    .Y(_03580_));
 OR5x2_ASAP7_75t_R _16653_ (.A(_01459_),
    .B(_01460_),
    .C(_01462_),
    .D(_01463_),
    .E(_05385_),
    .Y(_05432_));
 OR3x1_ASAP7_75t_R _16654_ (.A(_01458_),
    .B(_05416_),
    .C(_05432_),
    .Y(_05433_));
 OAI21x1_ASAP7_75t_R _16655_ (.A1(_05416_),
    .A2(_05432_),
    .B(_01458_),
    .Y(_05434_));
 AND3x1_ASAP7_75t_R _16656_ (.A(_05421_),
    .B(_05433_),
    .C(_05434_),
    .Y(_03581_));
 OR4x1_ASAP7_75t_R _16657_ (.A(_01457_),
    .B(_01458_),
    .C(_05419_),
    .D(_05432_),
    .Y(_05435_));
 OR3x1_ASAP7_75t_R _16658_ (.A(_01458_),
    .B(_05419_),
    .C(_05432_),
    .Y(_05436_));
 NAND2x1_ASAP7_75t_R _16659_ (.A(_01457_),
    .B(_05436_),
    .Y(_05437_));
 AND3x1_ASAP7_75t_R _16660_ (.A(_05421_),
    .B(_05435_),
    .C(_05437_),
    .Y(_03582_));
 OR4x1_ASAP7_75t_R _16661_ (.A(_01457_),
    .B(_01458_),
    .C(_05416_),
    .D(_05432_),
    .Y(_05438_));
 XOR2x2_ASAP7_75t_R _16662_ (.A(_05390_),
    .B(_05438_),
    .Y(_05439_));
 AND2x2_ASAP7_75t_R _16663_ (.A(_05427_),
    .B(_05439_),
    .Y(_03583_));
 OR3x1_ASAP7_75t_R _16664_ (.A(_01455_),
    .B(_05390_),
    .C(_05435_),
    .Y(_05440_));
 OAI21x1_ASAP7_75t_R _16665_ (.A1(_05390_),
    .A2(_05435_),
    .B(_01455_),
    .Y(_05441_));
 AND3x1_ASAP7_75t_R _16666_ (.A(_05421_),
    .B(_05440_),
    .C(_05441_),
    .Y(_03584_));
 OR3x1_ASAP7_75t_R _16667_ (.A(_01455_),
    .B(_05390_),
    .C(_05438_),
    .Y(_05442_));
 XOR2x2_ASAP7_75t_R _16668_ (.A(_01454_),
    .B(_05442_),
    .Y(_05443_));
 AND2x2_ASAP7_75t_R _16669_ (.A(_05427_),
    .B(_05443_),
    .Y(_03585_));
 OR4x1_ASAP7_75t_R _16670_ (.A(_01454_),
    .B(_01455_),
    .C(_05390_),
    .D(_05435_),
    .Y(_05444_));
 XOR2x2_ASAP7_75t_R _16671_ (.A(_01453_),
    .B(_05444_),
    .Y(_05445_));
 AND2x2_ASAP7_75t_R _16672_ (.A(_05427_),
    .B(_05445_),
    .Y(_03586_));
 OR5x1_ASAP7_75t_R _16673_ (.A(_01453_),
    .B(_01454_),
    .C(_01455_),
    .D(_05390_),
    .E(_05438_),
    .Y(_05446_));
 XOR2x2_ASAP7_75t_R _16674_ (.A(_01452_),
    .B(_05446_),
    .Y(_05447_));
 AND2x2_ASAP7_75t_R _16675_ (.A(_05427_),
    .B(_05447_),
    .Y(_03587_));
 OR5x2_ASAP7_75t_R _16676_ (.A(_01452_),
    .B(_01453_),
    .C(_01454_),
    .D(_01455_),
    .E(_05390_),
    .Y(_05448_));
 OR3x1_ASAP7_75t_R _16677_ (.A(_01451_),
    .B(_05435_),
    .C(_05448_),
    .Y(_05449_));
 OAI21x1_ASAP7_75t_R _16678_ (.A1(_05435_),
    .A2(_05448_),
    .B(_01451_),
    .Y(_05450_));
 AND3x1_ASAP7_75t_R _16679_ (.A(_05421_),
    .B(_05449_),
    .C(_05450_),
    .Y(_03588_));
 XOR2x2_ASAP7_75t_R _16680_ (.A(_01450_),
    .B(_02643_),
    .Y(_05451_));
 AND2x2_ASAP7_75t_R _16681_ (.A(_05427_),
    .B(_05451_),
    .Y(_03589_));
 OR3x1_ASAP7_75t_R _16682_ (.A(_01451_),
    .B(_05438_),
    .C(_05448_),
    .Y(_05452_));
 XOR2x2_ASAP7_75t_R _16683_ (.A(_01449_),
    .B(_05452_),
    .Y(_05453_));
 AND2x2_ASAP7_75t_R _16684_ (.A(_05427_),
    .B(_05453_),
    .Y(_03590_));
 OR4x1_ASAP7_75t_R _16685_ (.A(_01449_),
    .B(_01451_),
    .C(_05435_),
    .D(_05448_),
    .Y(_05454_));
 XOR2x2_ASAP7_75t_R _16686_ (.A(_01448_),
    .B(_05454_),
    .Y(_05455_));
 AND2x2_ASAP7_75t_R _16687_ (.A(_05427_),
    .B(_05455_),
    .Y(_03591_));
 OR3x1_ASAP7_75t_R _16688_ (.A(_01450_),
    .B(_01461_),
    .C(_00036_),
    .Y(_05456_));
 XOR2x2_ASAP7_75t_R _16689_ (.A(_01447_),
    .B(_05456_),
    .Y(_05457_));
 AND2x2_ASAP7_75t_R _16690_ (.A(_05427_),
    .B(_05457_),
    .Y(_03592_));
 OR3x1_ASAP7_75t_R _16691_ (.A(_01447_),
    .B(_01450_),
    .C(_02643_),
    .Y(_05458_));
 NAND2x1_ASAP7_75t_R _16692_ (.A(_01446_),
    .B(_05458_),
    .Y(_05459_));
 AND3x1_ASAP7_75t_R _16693_ (.A(_05421_),
    .B(_05398_),
    .C(_05459_),
    .Y(_03593_));
 BUFx6f_ASAP7_75t_R _16694_ (.A(_05426_),
    .Y(_05460_));
 XOR2x2_ASAP7_75t_R _16695_ (.A(_01445_),
    .B(_05403_),
    .Y(_05461_));
 AND2x2_ASAP7_75t_R _16696_ (.A(_05460_),
    .B(_05461_),
    .Y(_03594_));
 OR3x1_ASAP7_75t_R _16697_ (.A(_01444_),
    .B(_01445_),
    .C(_05398_),
    .Y(_05462_));
 OAI21x1_ASAP7_75t_R _16698_ (.A1(_01445_),
    .A2(_05398_),
    .B(_01444_),
    .Y(_05463_));
 AND3x1_ASAP7_75t_R _16699_ (.A(_05421_),
    .B(_05462_),
    .C(_05463_),
    .Y(_03595_));
 OR3x1_ASAP7_75t_R _16700_ (.A(_01444_),
    .B(_01445_),
    .C(_05403_),
    .Y(_05464_));
 XOR2x2_ASAP7_75t_R _16701_ (.A(_01443_),
    .B(_05464_),
    .Y(_05465_));
 AND2x2_ASAP7_75t_R _16702_ (.A(_05460_),
    .B(_05465_),
    .Y(_03596_));
 OR4x1_ASAP7_75t_R _16703_ (.A(_01443_),
    .B(_01444_),
    .C(_01445_),
    .D(_05398_),
    .Y(_05466_));
 NAND2x1_ASAP7_75t_R _16704_ (.A(_01442_),
    .B(_05466_),
    .Y(_05467_));
 AND3x1_ASAP7_75t_R _16705_ (.A(_05421_),
    .B(_05400_),
    .C(_05467_),
    .Y(_03597_));
 XOR2x2_ASAP7_75t_R _16706_ (.A(_05386_),
    .B(_05404_),
    .Y(_05468_));
 AND2x2_ASAP7_75t_R _16707_ (.A(_05460_),
    .B(_05468_),
    .Y(_03598_));
 AND2x2_ASAP7_75t_R _16708_ (.A(_05460_),
    .B(_00017_),
    .Y(_03599_));
 BUFx6f_ASAP7_75t_R _16709_ (.A(_02106_),
    .Y(_05469_));
 INVx1_ASAP7_75t_R _16710_ (.A(_02113_),
    .Y(_05470_));
 OR2x2_ASAP7_75t_R _16711_ (.A(_01511_),
    .B(_01516_),
    .Y(_05471_));
 OR2x2_ASAP7_75t_R _16712_ (.A(_01514_),
    .B(_01515_),
    .Y(_05472_));
 OA31x2_ASAP7_75t_R _16713_ (.A1(_01512_),
    .A2(\peo[22][35] ),
    .A3(_05472_),
    .B1(\peo[22][39] ),
    .Y(_05473_));
 AO21x1_ASAP7_75t_R _16714_ (.A1(_05470_),
    .A2(_05471_),
    .B(_05473_),
    .Y(_05474_));
 OR2x2_ASAP7_75t_R _16715_ (.A(_01475_),
    .B(_01476_),
    .Y(_05475_));
 OA31x2_ASAP7_75t_R _16716_ (.A1(_01473_),
    .A2(\xs[11].cli1.i[35] ),
    .A3(_05475_),
    .B1(\xs[11].cli1.i[39] ),
    .Y(_05476_));
 OR5x2_ASAP7_75t_R _16717_ (.A(_01472_),
    .B(_01473_),
    .C(\xs[11].cli1.i[35] ),
    .D(\peo[23][32] ),
    .E(_05475_),
    .Y(_05477_));
 OA21x2_ASAP7_75t_R _16718_ (.A1(_02113_),
    .A2(_05476_),
    .B(_05477_),
    .Y(_05478_));
 OA21x2_ASAP7_75t_R _16719_ (.A1(_05474_),
    .A2(_05478_),
    .B(_02107_),
    .Y(_05479_));
 INVx2_ASAP7_75t_R _16720_ (.A(_05479_),
    .Y(_05480_));
 OR4x1_ASAP7_75t_R _16721_ (.A(_09220_),
    .B(_05469_),
    .C(_05470_),
    .D(_05480_),
    .Y(_05481_));
 BUFx6f_ASAP7_75t_R _16722_ (.A(_05481_),
    .Y(_05482_));
 INVx3_ASAP7_75t_R _16723_ (.A(_05469_),
    .Y(_05483_));
 AND3x1_ASAP7_75t_R _16724_ (.A(_05483_),
    .B(_02113_),
    .C(_05479_),
    .Y(_05484_));
 AO21x1_ASAP7_75t_R _16725_ (.A1(_00017_),
    .A2(_05476_),
    .B(_05483_),
    .Y(_05485_));
 INVx1_ASAP7_75t_R _16726_ (.A(_02107_),
    .Y(_05486_));
 OR3x1_ASAP7_75t_R _16727_ (.A(_05469_),
    .B(_05486_),
    .C(_02113_),
    .Y(_05487_));
 AND3x1_ASAP7_75t_R _16728_ (.A(_05473_),
    .B(_05485_),
    .C(_05487_),
    .Y(_05488_));
 OA21x2_ASAP7_75t_R _16729_ (.A1(_05477_),
    .A2(_05488_),
    .B(_01518_),
    .Y(_05489_));
 OR3x1_ASAP7_75t_R _16730_ (.A(_08941_),
    .B(_05484_),
    .C(_05489_),
    .Y(_05490_));
 NOR2x1_ASAP7_75t_R _16731_ (.A(_01475_),
    .B(_01476_),
    .Y(_05491_));
 AND5x1_ASAP7_75t_R _16732_ (.A(\xs[11].cli1.i[39] ),
    .B(\xs[11].cli1.i[36] ),
    .C(_01474_),
    .D(_01477_),
    .E(_05491_),
    .Y(_05492_));
 AO21x1_ASAP7_75t_R _16733_ (.A1(_05473_),
    .A2(_05492_),
    .B(_05476_),
    .Y(_05493_));
 OA21x2_ASAP7_75t_R _16734_ (.A1(_05492_),
    .A2(_05476_),
    .B(_02113_),
    .Y(_05494_));
 AND3x1_ASAP7_75t_R _16735_ (.A(_05469_),
    .B(_00017_),
    .C(_05476_),
    .Y(_05495_));
 AO21x1_ASAP7_75t_R _16736_ (.A1(_05483_),
    .A2(_05494_),
    .B(_05495_),
    .Y(_05496_));
 AO32x1_ASAP7_75t_R _16737_ (.A1(_05483_),
    .A2(_05486_),
    .A3(_05493_),
    .B1(_05496_),
    .B2(_05473_),
    .Y(_05497_));
 BUFx3_ASAP7_75t_R _16738_ (.A(_05497_),
    .Y(_05498_));
 NOR3x1_ASAP7_75t_R _16739_ (.A(\peo[23][0] ),
    .B(_05477_),
    .C(_05498_),
    .Y(_05499_));
 OAI22x1_ASAP7_75t_R _16740_ (.A1(_02117_),
    .A2(_05482_),
    .B1(_05490_),
    .B2(_05499_),
    .Y(_03600_));
 NOR2x1_ASAP7_75t_R _16741_ (.A(_02116_),
    .B(_05482_),
    .Y(_03601_));
 NOR2x1_ASAP7_75t_R _16742_ (.A(_02115_),
    .B(_05482_),
    .Y(_03602_));
 NOR2x1_ASAP7_75t_R _16743_ (.A(_02114_),
    .B(_05482_),
    .Y(_03603_));
 NOR2x1_ASAP7_75t_R _16744_ (.A(_02105_),
    .B(_05482_),
    .Y(_03604_));
 NOR2x1_ASAP7_75t_R _16745_ (.A(_02104_),
    .B(_05482_),
    .Y(_03605_));
 NOR2x1_ASAP7_75t_R _16746_ (.A(_05474_),
    .B(_05478_),
    .Y(_05500_));
 OAI21x1_ASAP7_75t_R _16747_ (.A1(_05500_),
    .A2(_05487_),
    .B(_01518_),
    .Y(_05501_));
 INVx1_ASAP7_75t_R _16748_ (.A(_02117_),
    .Y(_05502_));
 OR3x1_ASAP7_75t_R _16749_ (.A(_05502_),
    .B(_05500_),
    .C(_05487_),
    .Y(_05503_));
 AO21x1_ASAP7_75t_R _16750_ (.A1(_05501_),
    .A2(_05503_),
    .B(_05498_),
    .Y(_05504_));
 NAND2x1_ASAP7_75t_R _16751_ (.A(_01479_),
    .B(_05498_),
    .Y(_05505_));
 AND3x1_ASAP7_75t_R _16752_ (.A(_05421_),
    .B(_05504_),
    .C(_05505_),
    .Y(_03606_));
 OR4x1_ASAP7_75t_R _16753_ (.A(_11177_),
    .B(_05469_),
    .C(_02113_),
    .D(_05480_),
    .Y(_05506_));
 NOR2x1_ASAP7_75t_R _16754_ (.A(_02116_),
    .B(_05506_),
    .Y(_03607_));
 NOR2x1_ASAP7_75t_R _16755_ (.A(_02115_),
    .B(_05506_),
    .Y(_03608_));
 NOR2x1_ASAP7_75t_R _16756_ (.A(_02114_),
    .B(_05506_),
    .Y(_03609_));
 NOR2x1_ASAP7_75t_R _16757_ (.A(_02105_),
    .B(_05506_),
    .Y(_03610_));
 NOR2x1_ASAP7_75t_R _16758_ (.A(_02104_),
    .B(_05506_),
    .Y(_03611_));
 OA21x2_ASAP7_75t_R _16759_ (.A1(_05469_),
    .A2(_05479_),
    .B(_08584_),
    .Y(_05507_));
 OAI21x1_ASAP7_75t_R _16760_ (.A1(_05469_),
    .A2(_02107_),
    .B(_05476_),
    .Y(_05508_));
 AO21x1_ASAP7_75t_R _16761_ (.A1(_05473_),
    .A2(_05496_),
    .B(_05508_),
    .Y(_05509_));
 BUFx6f_ASAP7_75t_R _16762_ (.A(_05509_),
    .Y(_05510_));
 OR2x2_ASAP7_75t_R _16763_ (.A(\peo[23][0] ),
    .B(_05510_),
    .Y(_05511_));
 NAND2x1_ASAP7_75t_R _16764_ (.A(_01518_),
    .B(_05510_),
    .Y(_05512_));
 AND3x4_ASAP7_75t_R _16765_ (.A(_08876_),
    .B(_05483_),
    .C(_05480_),
    .Y(_05513_));
 AO32x1_ASAP7_75t_R _16766_ (.A1(_05507_),
    .A2(_05511_),
    .A3(_05512_),
    .B1(_05513_),
    .B2(_05502_),
    .Y(_03612_));
 OR3x1_ASAP7_75t_R _16767_ (.A(_08578_),
    .B(_05469_),
    .C(_05479_),
    .Y(_05514_));
 BUFx6f_ASAP7_75t_R _16768_ (.A(_05514_),
    .Y(_05515_));
 NOR2x1_ASAP7_75t_R _16769_ (.A(_02116_),
    .B(_05515_),
    .Y(_03613_));
 NOR2x1_ASAP7_75t_R _16770_ (.A(_02115_),
    .B(_05515_),
    .Y(_03614_));
 NOR2x1_ASAP7_75t_R _16771_ (.A(_02114_),
    .B(_05515_),
    .Y(_03615_));
 OR2x2_ASAP7_75t_R _16772_ (.A(\peo[23][32] ),
    .B(_05510_),
    .Y(_05516_));
 NAND2x1_ASAP7_75t_R _16773_ (.A(_01516_),
    .B(_05510_),
    .Y(_05517_));
 AO32x1_ASAP7_75t_R _16774_ (.A1(_05507_),
    .A2(_05516_),
    .A3(_05517_),
    .B1(_05513_),
    .B2(_05470_),
    .Y(_03616_));
 NAND2x1_ASAP7_75t_R _16775_ (.A(_01515_),
    .B(_05510_),
    .Y(_05518_));
 OR3x1_ASAP7_75t_R _16776_ (.A(_01472_),
    .B(\xs[11].cli1.i[33] ),
    .C(_05498_),
    .Y(_05519_));
 INVx1_ASAP7_75t_R _16777_ (.A(_02112_),
    .Y(_05520_));
 AO32x1_ASAP7_75t_R _16778_ (.A1(_05507_),
    .A2(_05518_),
    .A3(_05519_),
    .B1(_05513_),
    .B2(_05520_),
    .Y(_03617_));
 NAND2x1_ASAP7_75t_R _16779_ (.A(_01514_),
    .B(_05510_),
    .Y(_05521_));
 OR3x1_ASAP7_75t_R _16780_ (.A(_01472_),
    .B(\xs[11].cli1.i[34] ),
    .C(_05498_),
    .Y(_05522_));
 INVx1_ASAP7_75t_R _16781_ (.A(_02111_),
    .Y(_05523_));
 AO32x1_ASAP7_75t_R _16782_ (.A1(_05507_),
    .A2(_05521_),
    .A3(_05522_),
    .B1(_05513_),
    .B2(_05523_),
    .Y(_03618_));
 OR2x2_ASAP7_75t_R _16783_ (.A(\xs[11].cli1.i[35] ),
    .B(_05510_),
    .Y(_05524_));
 NAND2x1_ASAP7_75t_R _16784_ (.A(_01513_),
    .B(_05510_),
    .Y(_05525_));
 INVx1_ASAP7_75t_R _16785_ (.A(_02110_),
    .Y(_05526_));
 AO32x1_ASAP7_75t_R _16786_ (.A1(_05507_),
    .A2(_05524_),
    .A3(_05525_),
    .B1(_05513_),
    .B2(_05526_),
    .Y(_03619_));
 NAND2x1_ASAP7_75t_R _16787_ (.A(_01512_),
    .B(_05510_),
    .Y(_05527_));
 OR3x1_ASAP7_75t_R _16788_ (.A(_01472_),
    .B(\xs[11].cli1.i[36] ),
    .C(_05498_),
    .Y(_05528_));
 INVx1_ASAP7_75t_R _16789_ (.A(_02109_),
    .Y(_05529_));
 AO32x1_ASAP7_75t_R _16790_ (.A1(_05507_),
    .A2(_05527_),
    .A3(_05528_),
    .B1(_05513_),
    .B2(_05529_),
    .Y(_03620_));
 NOR2x1_ASAP7_75t_R _16791_ (.A(_02108_),
    .B(_05515_),
    .Y(_03621_));
 AND4x1_ASAP7_75t_R _16792_ (.A(_08999_),
    .B(_05483_),
    .C(_02107_),
    .D(_05500_),
    .Y(_03622_));
 AOI211x1_ASAP7_75t_R _16793_ (.A1(_05483_),
    .A2(_05480_),
    .B(_05476_),
    .C(_05473_),
    .Y(_05530_));
 NOR2x1_ASAP7_75t_R _16794_ (.A(_05300_),
    .B(_05530_),
    .Y(_03623_));
 NOR2x1_ASAP7_75t_R _16795_ (.A(_02105_),
    .B(_05515_),
    .Y(_03624_));
 NOR2x1_ASAP7_75t_R _16796_ (.A(_02104_),
    .B(_05515_),
    .Y(_03625_));
 BUFx3_ASAP7_75t_R _16797_ (.A(_01403_),
    .Y(_05531_));
 BUFx3_ASAP7_75t_R _16798_ (.A(_01376_),
    .Y(_05532_));
 AND4x1_ASAP7_75t_R _16799_ (.A(_05532_),
    .B(_01404_),
    .C(_01405_),
    .D(_01406_),
    .Y(_05533_));
 AND5x1_ASAP7_75t_R _16800_ (.A(_01395_),
    .B(_01400_),
    .C(_01401_),
    .D(_05531_),
    .E(_05533_),
    .Y(_05534_));
 AND5x2_ASAP7_75t_R _16801_ (.A(_01397_),
    .B(_01398_),
    .C(_01399_),
    .D(_11466_),
    .E(_05534_),
    .Y(_05535_));
 AND4x1_ASAP7_75t_R _16802_ (.A(_01390_),
    .B(_01391_),
    .C(_01392_),
    .D(_01393_),
    .Y(_05536_));
 AND4x1_ASAP7_75t_R _16803_ (.A(_01384_),
    .B(_01386_),
    .C(_01387_),
    .D(_01394_),
    .Y(_05537_));
 AND5x1_ASAP7_75t_R _16804_ (.A(_01377_),
    .B(_01378_),
    .C(_01383_),
    .D(_01402_),
    .E(_05537_),
    .Y(_05538_));
 AND3x1_ASAP7_75t_R _16805_ (.A(_01381_),
    .B(_01382_),
    .C(_01385_),
    .Y(_05539_));
 OR3x1_ASAP7_75t_R _16806_ (.A(_01379_),
    .B(_01380_),
    .C(_05539_),
    .Y(_05540_));
 AND5x2_ASAP7_75t_R _16807_ (.A(_01388_),
    .B(_01389_),
    .C(_05536_),
    .D(_05538_),
    .E(_05540_),
    .Y(_05541_));
 NAND2x2_ASAP7_75t_R _16808_ (.A(_05535_),
    .B(_05541_),
    .Y(_05542_));
 NOR2x1_ASAP7_75t_R _16809_ (.A(_01333_),
    .B(_05542_),
    .Y(_03626_));
 INVx1_ASAP7_75t_R _16810_ (.A(_05542_),
    .Y(_03627_));
 NOR2x1_ASAP7_75t_R _16811_ (.A(_01336_),
    .B(_05542_),
    .Y(_03628_));
 NOR2x1_ASAP7_75t_R _16812_ (.A(_01335_),
    .B(_05542_),
    .Y(_03629_));
 NOR2x1_ASAP7_75t_R _16813_ (.A(_01334_),
    .B(_05542_),
    .Y(_03630_));
 NOR2x1_ASAP7_75t_R _16814_ (.A(_01332_),
    .B(_05542_),
    .Y(_03631_));
 NOR2x1_ASAP7_75t_R _16815_ (.A(_01331_),
    .B(_05542_),
    .Y(_03632_));
 INVx1_ASAP7_75t_R _16816_ (.A(_05542_),
    .Y(_03633_));
 AND2x2_ASAP7_75t_R _16817_ (.A(_05460_),
    .B(_00037_),
    .Y(_03634_));
 OR4x1_ASAP7_75t_R _16818_ (.A(_01381_),
    .B(_01382_),
    .C(_01385_),
    .D(_02655_),
    .Y(_05543_));
 OR4x1_ASAP7_75t_R _16819_ (.A(_01377_),
    .B(_01378_),
    .C(_01379_),
    .D(_01380_),
    .Y(_05544_));
 OR2x6_ASAP7_75t_R _16820_ (.A(_05543_),
    .B(_05544_),
    .Y(_05545_));
 OR3x1_ASAP7_75t_R _16821_ (.A(_05532_),
    .B(_01406_),
    .C(_05545_),
    .Y(_05546_));
 OAI21x1_ASAP7_75t_R _16822_ (.A1(_05532_),
    .A2(_05545_),
    .B(_01406_),
    .Y(_05547_));
 AND3x1_ASAP7_75t_R _16823_ (.A(_05421_),
    .B(_05546_),
    .C(_05547_),
    .Y(_03635_));
 OR5x2_ASAP7_75t_R _16824_ (.A(_01381_),
    .B(_01382_),
    .C(_01385_),
    .D(_01396_),
    .E(_00037_),
    .Y(_05548_));
 OR2x2_ASAP7_75t_R _16825_ (.A(_05544_),
    .B(_05548_),
    .Y(_05549_));
 OR3x1_ASAP7_75t_R _16826_ (.A(_05532_),
    .B(_01406_),
    .C(_05549_),
    .Y(_05550_));
 XOR2x2_ASAP7_75t_R _16827_ (.A(_01405_),
    .B(_05550_),
    .Y(_05551_));
 AND2x2_ASAP7_75t_R _16828_ (.A(_05460_),
    .B(_05551_),
    .Y(_03636_));
 BUFx6f_ASAP7_75t_R _16829_ (.A(_05337_),
    .Y(_05552_));
 OR4x1_ASAP7_75t_R _16830_ (.A(_05532_),
    .B(_01404_),
    .C(_01405_),
    .D(_01406_),
    .Y(_05553_));
 OR3x2_ASAP7_75t_R _16831_ (.A(_05543_),
    .B(_05544_),
    .C(_05553_),
    .Y(_05554_));
 OR4x1_ASAP7_75t_R _16832_ (.A(_05532_),
    .B(_01405_),
    .C(_01406_),
    .D(_05545_),
    .Y(_05555_));
 NAND2x1_ASAP7_75t_R _16833_ (.A(_01404_),
    .B(_05555_),
    .Y(_05556_));
 AND3x1_ASAP7_75t_R _16834_ (.A(_05552_),
    .B(_05554_),
    .C(_05556_),
    .Y(_03637_));
 OR3x2_ASAP7_75t_R _16835_ (.A(_05544_),
    .B(_05548_),
    .C(_05553_),
    .Y(_05557_));
 XOR2x2_ASAP7_75t_R _16836_ (.A(_05531_),
    .B(_05557_),
    .Y(_05558_));
 AND2x2_ASAP7_75t_R _16837_ (.A(_05460_),
    .B(_05558_),
    .Y(_03638_));
 OR3x1_ASAP7_75t_R _16838_ (.A(_01402_),
    .B(_05531_),
    .C(_05554_),
    .Y(_05559_));
 OAI21x1_ASAP7_75t_R _16839_ (.A1(_05531_),
    .A2(_05554_),
    .B(_01402_),
    .Y(_05560_));
 AND3x1_ASAP7_75t_R _16840_ (.A(_05552_),
    .B(_05559_),
    .C(_05560_),
    .Y(_03639_));
 OR3x1_ASAP7_75t_R _16841_ (.A(_01402_),
    .B(_05531_),
    .C(_05557_),
    .Y(_05561_));
 XOR2x2_ASAP7_75t_R _16842_ (.A(_01401_),
    .B(_05561_),
    .Y(_05562_));
 AND2x2_ASAP7_75t_R _16843_ (.A(_05460_),
    .B(_05562_),
    .Y(_03640_));
 OR4x1_ASAP7_75t_R _16844_ (.A(_01401_),
    .B(_01402_),
    .C(_05531_),
    .D(_05554_),
    .Y(_05563_));
 XOR2x2_ASAP7_75t_R _16845_ (.A(_01400_),
    .B(_05563_),
    .Y(_05564_));
 AND2x2_ASAP7_75t_R _16846_ (.A(_05460_),
    .B(_05564_),
    .Y(_03641_));
 OR5x1_ASAP7_75t_R _16847_ (.A(_01400_),
    .B(_01401_),
    .C(_01402_),
    .D(_05531_),
    .E(_05557_),
    .Y(_05565_));
 XOR2x2_ASAP7_75t_R _16848_ (.A(_01399_),
    .B(_05565_),
    .Y(_05566_));
 AND2x2_ASAP7_75t_R _16849_ (.A(_05460_),
    .B(_05566_),
    .Y(_03642_));
 OR5x2_ASAP7_75t_R _16850_ (.A(_01399_),
    .B(_01400_),
    .C(_01401_),
    .D(_01402_),
    .E(_05531_),
    .Y(_05567_));
 OR3x2_ASAP7_75t_R _16851_ (.A(_01398_),
    .B(_05554_),
    .C(_05567_),
    .Y(_05568_));
 OAI21x1_ASAP7_75t_R _16852_ (.A1(_05554_),
    .A2(_05567_),
    .B(_01398_),
    .Y(_05569_));
 AND3x1_ASAP7_75t_R _16853_ (.A(_05552_),
    .B(_05568_),
    .C(_05569_),
    .Y(_03643_));
 BUFx6f_ASAP7_75t_R _16854_ (.A(_05426_),
    .Y(_05570_));
 OR3x2_ASAP7_75t_R _16855_ (.A(_01398_),
    .B(_05557_),
    .C(_05567_),
    .Y(_05571_));
 XOR2x2_ASAP7_75t_R _16856_ (.A(_01397_),
    .B(_05571_),
    .Y(_05572_));
 AND2x2_ASAP7_75t_R _16857_ (.A(_05570_),
    .B(_05572_),
    .Y(_03644_));
 NOR2x1_ASAP7_75t_R _16858_ (.A(_05300_),
    .B(_02656_),
    .Y(_03645_));
 OR3x1_ASAP7_75t_R _16859_ (.A(_01395_),
    .B(_01397_),
    .C(_05568_),
    .Y(_05573_));
 OAI21x1_ASAP7_75t_R _16860_ (.A1(_01397_),
    .A2(_05568_),
    .B(_01395_),
    .Y(_05574_));
 AND3x1_ASAP7_75t_R _16861_ (.A(_05552_),
    .B(_05573_),
    .C(_05574_),
    .Y(_03646_));
 OR3x1_ASAP7_75t_R _16862_ (.A(_01395_),
    .B(_01397_),
    .C(_05571_),
    .Y(_05575_));
 XOR2x2_ASAP7_75t_R _16863_ (.A(_01394_),
    .B(_05575_),
    .Y(_05576_));
 AND2x2_ASAP7_75t_R _16864_ (.A(_05570_),
    .B(_05576_),
    .Y(_03647_));
 OR4x1_ASAP7_75t_R _16865_ (.A(_01394_),
    .B(_01395_),
    .C(_01397_),
    .D(_05568_),
    .Y(_05577_));
 XOR2x2_ASAP7_75t_R _16866_ (.A(_01393_),
    .B(_05577_),
    .Y(_05578_));
 AND2x2_ASAP7_75t_R _16867_ (.A(_05570_),
    .B(_05578_),
    .Y(_03648_));
 OR4x1_ASAP7_75t_R _16868_ (.A(_01393_),
    .B(_01394_),
    .C(_01395_),
    .D(_01397_),
    .Y(_05579_));
 OR3x2_ASAP7_75t_R _16869_ (.A(_01392_),
    .B(_05571_),
    .C(_05579_),
    .Y(_05580_));
 OAI21x1_ASAP7_75t_R _16870_ (.A1(_05571_),
    .A2(_05579_),
    .B(_01392_),
    .Y(_05581_));
 AND3x1_ASAP7_75t_R _16871_ (.A(_05552_),
    .B(_05580_),
    .C(_05581_),
    .Y(_03649_));
 OR3x2_ASAP7_75t_R _16872_ (.A(_01392_),
    .B(_05568_),
    .C(_05579_),
    .Y(_05582_));
 XOR2x2_ASAP7_75t_R _16873_ (.A(_01391_),
    .B(_05582_),
    .Y(_05583_));
 AND2x2_ASAP7_75t_R _16874_ (.A(_05570_),
    .B(_05583_),
    .Y(_03650_));
 OR3x1_ASAP7_75t_R _16875_ (.A(_01390_),
    .B(_01391_),
    .C(_05580_),
    .Y(_05584_));
 OAI21x1_ASAP7_75t_R _16876_ (.A1(_01391_),
    .A2(_05580_),
    .B(_01390_),
    .Y(_05585_));
 AND3x1_ASAP7_75t_R _16877_ (.A(_05552_),
    .B(_05584_),
    .C(_05585_),
    .Y(_03651_));
 OR3x1_ASAP7_75t_R _16878_ (.A(_01390_),
    .B(_01391_),
    .C(_05582_),
    .Y(_05586_));
 XOR2x2_ASAP7_75t_R _16879_ (.A(_01389_),
    .B(_05586_),
    .Y(_05587_));
 AND2x2_ASAP7_75t_R _16880_ (.A(_05570_),
    .B(_05587_),
    .Y(_03652_));
 OR4x1_ASAP7_75t_R _16881_ (.A(_01389_),
    .B(_01390_),
    .C(_01391_),
    .D(_05580_),
    .Y(_05588_));
 XOR2x2_ASAP7_75t_R _16882_ (.A(_01388_),
    .B(_05588_),
    .Y(_05589_));
 AND2x2_ASAP7_75t_R _16883_ (.A(_05570_),
    .B(_05589_),
    .Y(_03653_));
 OR4x1_ASAP7_75t_R _16884_ (.A(_01388_),
    .B(_01389_),
    .C(_01390_),
    .D(_01391_),
    .Y(_05590_));
 OR3x1_ASAP7_75t_R _16885_ (.A(_01387_),
    .B(_05582_),
    .C(_05590_),
    .Y(_05591_));
 OAI21x1_ASAP7_75t_R _16886_ (.A1(_05582_),
    .A2(_05590_),
    .B(_01387_),
    .Y(_05592_));
 AND3x1_ASAP7_75t_R _16887_ (.A(_05552_),
    .B(_05591_),
    .C(_05592_),
    .Y(_03654_));
 OR3x1_ASAP7_75t_R _16888_ (.A(_01387_),
    .B(_05580_),
    .C(_05590_),
    .Y(_05593_));
 XOR2x2_ASAP7_75t_R _16889_ (.A(_01386_),
    .B(_05593_),
    .Y(_05594_));
 AND2x2_ASAP7_75t_R _16890_ (.A(_05570_),
    .B(_05594_),
    .Y(_03655_));
 XOR2x2_ASAP7_75t_R _16891_ (.A(_01385_),
    .B(_02655_),
    .Y(_05595_));
 AND2x2_ASAP7_75t_R _16892_ (.A(_05570_),
    .B(_05595_),
    .Y(_03656_));
 OR4x1_ASAP7_75t_R _16893_ (.A(_01386_),
    .B(_01387_),
    .C(_05582_),
    .D(_05590_),
    .Y(_05596_));
 XOR2x2_ASAP7_75t_R _16894_ (.A(_01384_),
    .B(_05596_),
    .Y(_05597_));
 AND2x2_ASAP7_75t_R _16895_ (.A(_05570_),
    .B(_05597_),
    .Y(_03657_));
 OR5x1_ASAP7_75t_R _16896_ (.A(_01384_),
    .B(_01386_),
    .C(_01387_),
    .D(_05580_),
    .E(_05590_),
    .Y(_05598_));
 XOR2x2_ASAP7_75t_R _16897_ (.A(_01383_),
    .B(_05598_),
    .Y(_05599_));
 AND2x2_ASAP7_75t_R _16898_ (.A(_05570_),
    .B(_05599_),
    .Y(_03658_));
 BUFx6f_ASAP7_75t_R _16899_ (.A(_05426_),
    .Y(_05600_));
 OR3x1_ASAP7_75t_R _16900_ (.A(_01385_),
    .B(_01396_),
    .C(_00037_),
    .Y(_05601_));
 XOR2x2_ASAP7_75t_R _16901_ (.A(_01382_),
    .B(_05601_),
    .Y(_05602_));
 AND2x2_ASAP7_75t_R _16902_ (.A(_05600_),
    .B(_05602_),
    .Y(_03659_));
 OR3x1_ASAP7_75t_R _16903_ (.A(_01382_),
    .B(_01385_),
    .C(_02655_),
    .Y(_05603_));
 NAND2x1_ASAP7_75t_R _16904_ (.A(_01381_),
    .B(_05603_),
    .Y(_05604_));
 AND3x1_ASAP7_75t_R _16905_ (.A(_05552_),
    .B(_05543_),
    .C(_05604_),
    .Y(_03660_));
 XOR2x2_ASAP7_75t_R _16906_ (.A(_01380_),
    .B(_05548_),
    .Y(_05605_));
 AND2x2_ASAP7_75t_R _16907_ (.A(_05600_),
    .B(_05605_),
    .Y(_03661_));
 OR3x1_ASAP7_75t_R _16908_ (.A(_01379_),
    .B(_01380_),
    .C(_05543_),
    .Y(_05606_));
 OAI21x1_ASAP7_75t_R _16909_ (.A1(_01380_),
    .A2(_05543_),
    .B(_01379_),
    .Y(_05607_));
 AND3x1_ASAP7_75t_R _16910_ (.A(_05552_),
    .B(_05606_),
    .C(_05607_),
    .Y(_03662_));
 OR3x1_ASAP7_75t_R _16911_ (.A(_01379_),
    .B(_01380_),
    .C(_05548_),
    .Y(_05608_));
 XOR2x2_ASAP7_75t_R _16912_ (.A(_01378_),
    .B(_05608_),
    .Y(_05609_));
 AND2x2_ASAP7_75t_R _16913_ (.A(_05600_),
    .B(_05609_),
    .Y(_03663_));
 OR4x1_ASAP7_75t_R _16914_ (.A(_01378_),
    .B(_01379_),
    .C(_01380_),
    .D(_05543_),
    .Y(_05610_));
 NAND2x1_ASAP7_75t_R _16915_ (.A(_01377_),
    .B(_05610_),
    .Y(_05611_));
 AND3x1_ASAP7_75t_R _16916_ (.A(_05552_),
    .B(_05545_),
    .C(_05611_),
    .Y(_03664_));
 XOR2x2_ASAP7_75t_R _16917_ (.A(_05532_),
    .B(_05549_),
    .Y(_05612_));
 AND2x2_ASAP7_75t_R _16918_ (.A(_05600_),
    .B(_05612_),
    .Y(_03665_));
 BUFx6f_ASAP7_75t_R _16919_ (.A(_01360_),
    .Y(_05613_));
 BUFx6f_ASAP7_75t_R _16920_ (.A(_01337_),
    .Y(_05614_));
 AND4x1_ASAP7_75t_R _16921_ (.A(_05614_),
    .B(_01365_),
    .C(_01366_),
    .D(_01367_),
    .Y(_05615_));
 AND5x1_ASAP7_75t_R _16922_ (.A(_01356_),
    .B(_01361_),
    .C(_01362_),
    .D(_01364_),
    .E(_05615_),
    .Y(_05616_));
 AND5x2_ASAP7_75t_R _16923_ (.A(_01358_),
    .B(_01359_),
    .C(_05613_),
    .D(_11466_),
    .E(_05616_),
    .Y(_05617_));
 BUFx3_ASAP7_75t_R _16924_ (.A(_01352_),
    .Y(_05618_));
 AND4x1_ASAP7_75t_R _16925_ (.A(_01351_),
    .B(_05618_),
    .C(_01353_),
    .D(_01354_),
    .Y(_05619_));
 AND4x1_ASAP7_75t_R _16926_ (.A(_01345_),
    .B(_01347_),
    .C(_01348_),
    .D(_01355_),
    .Y(_05620_));
 AND5x1_ASAP7_75t_R _16927_ (.A(_01338_),
    .B(_01339_),
    .C(_01344_),
    .D(_01363_),
    .E(_05620_),
    .Y(_05621_));
 AND3x1_ASAP7_75t_R _16928_ (.A(_01342_),
    .B(_01343_),
    .C(_01346_),
    .Y(_05622_));
 OR3x1_ASAP7_75t_R _16929_ (.A(_01340_),
    .B(_01341_),
    .C(_05622_),
    .Y(_05623_));
 AND5x2_ASAP7_75t_R _16930_ (.A(_01349_),
    .B(_01350_),
    .C(_05619_),
    .D(_05621_),
    .E(_05623_),
    .Y(_05624_));
 NAND2x2_ASAP7_75t_R _16931_ (.A(_05617_),
    .B(_05624_),
    .Y(_05625_));
 NOR2x1_ASAP7_75t_R _16932_ (.A(_01327_),
    .B(_05625_),
    .Y(_03666_));
 INVx1_ASAP7_75t_R _16933_ (.A(_05625_),
    .Y(_03667_));
 NOR2x1_ASAP7_75t_R _16934_ (.A(_01330_),
    .B(_05625_),
    .Y(_03668_));
 NOR2x1_ASAP7_75t_R _16935_ (.A(_01329_),
    .B(_05625_),
    .Y(_03669_));
 NOR2x1_ASAP7_75t_R _16936_ (.A(_01328_),
    .B(_05625_),
    .Y(_03670_));
 NOR2x1_ASAP7_75t_R _16937_ (.A(_01326_),
    .B(_05625_),
    .Y(_03671_));
 NOR2x1_ASAP7_75t_R _16938_ (.A(_01325_),
    .B(_05625_),
    .Y(_03672_));
 INVx1_ASAP7_75t_R _16939_ (.A(_05625_),
    .Y(_03673_));
 AND2x2_ASAP7_75t_R _16940_ (.A(_05600_),
    .B(_00038_),
    .Y(_03674_));
 BUFx6f_ASAP7_75t_R _16941_ (.A(_05337_),
    .Y(_05626_));
 OR4x1_ASAP7_75t_R _16942_ (.A(_01342_),
    .B(_01343_),
    .C(_01346_),
    .D(_02625_),
    .Y(_05627_));
 OR4x1_ASAP7_75t_R _16943_ (.A(_01338_),
    .B(_01339_),
    .C(_01340_),
    .D(_01341_),
    .Y(_05628_));
 OR2x6_ASAP7_75t_R _16944_ (.A(_05627_),
    .B(_05628_),
    .Y(_05629_));
 OR3x1_ASAP7_75t_R _16945_ (.A(_05614_),
    .B(_01367_),
    .C(_05629_),
    .Y(_05630_));
 OAI21x1_ASAP7_75t_R _16946_ (.A1(_05614_),
    .A2(_05629_),
    .B(_01367_),
    .Y(_05631_));
 AND3x1_ASAP7_75t_R _16947_ (.A(_05626_),
    .B(_05630_),
    .C(_05631_),
    .Y(_03675_));
 OR5x2_ASAP7_75t_R _16948_ (.A(_01342_),
    .B(_01343_),
    .C(_01346_),
    .D(_01357_),
    .E(_00038_),
    .Y(_05632_));
 OR2x6_ASAP7_75t_R _16949_ (.A(_05628_),
    .B(_05632_),
    .Y(_05633_));
 OR3x1_ASAP7_75t_R _16950_ (.A(_05614_),
    .B(_01367_),
    .C(_05633_),
    .Y(_05634_));
 XOR2x2_ASAP7_75t_R _16951_ (.A(_01366_),
    .B(_05634_),
    .Y(_05635_));
 AND2x2_ASAP7_75t_R _16952_ (.A(_05600_),
    .B(_05635_),
    .Y(_03676_));
 OR4x1_ASAP7_75t_R _16953_ (.A(_05614_),
    .B(_01366_),
    .C(_01367_),
    .D(_05629_),
    .Y(_05636_));
 XOR2x2_ASAP7_75t_R _16954_ (.A(_01365_),
    .B(_05636_),
    .Y(_05637_));
 AND2x2_ASAP7_75t_R _16955_ (.A(_05600_),
    .B(_05637_),
    .Y(_03677_));
 OR5x2_ASAP7_75t_R _16956_ (.A(_05614_),
    .B(_01364_),
    .C(_01365_),
    .D(_01366_),
    .E(_01367_),
    .Y(_05638_));
 OR5x1_ASAP7_75t_R _16957_ (.A(_05614_),
    .B(_01365_),
    .C(_01366_),
    .D(_01367_),
    .E(_05633_),
    .Y(_05639_));
 NAND2x1_ASAP7_75t_R _16958_ (.A(_01364_),
    .B(_05639_),
    .Y(_05640_));
 OA211x2_ASAP7_75t_R _16959_ (.A1(_05633_),
    .A2(_05638_),
    .B(_05640_),
    .C(_11589_),
    .Y(_03678_));
 OR3x2_ASAP7_75t_R _16960_ (.A(_05627_),
    .B(_05628_),
    .C(_05638_),
    .Y(_05641_));
 XOR2x2_ASAP7_75t_R _16961_ (.A(_01363_),
    .B(_05641_),
    .Y(_05642_));
 AND2x2_ASAP7_75t_R _16962_ (.A(_05600_),
    .B(_05642_),
    .Y(_03679_));
 OR3x1_ASAP7_75t_R _16963_ (.A(_01363_),
    .B(_05633_),
    .C(_05638_),
    .Y(_05643_));
 XOR2x2_ASAP7_75t_R _16964_ (.A(_01362_),
    .B(_05643_),
    .Y(_05644_));
 AND2x2_ASAP7_75t_R _16965_ (.A(_05600_),
    .B(_05644_),
    .Y(_03680_));
 OR4x1_ASAP7_75t_R _16966_ (.A(_01361_),
    .B(_01362_),
    .C(_01363_),
    .D(_05641_),
    .Y(_05645_));
 OR3x1_ASAP7_75t_R _16967_ (.A(_01362_),
    .B(_01363_),
    .C(_05641_),
    .Y(_05646_));
 NAND2x1_ASAP7_75t_R _16968_ (.A(_01361_),
    .B(_05646_),
    .Y(_05647_));
 AND3x1_ASAP7_75t_R _16969_ (.A(_05626_),
    .B(_05645_),
    .C(_05647_),
    .Y(_03681_));
 OR5x2_ASAP7_75t_R _16970_ (.A(_01361_),
    .B(_01362_),
    .C(_01363_),
    .D(_05633_),
    .E(_05638_),
    .Y(_05648_));
 XOR2x2_ASAP7_75t_R _16971_ (.A(_05613_),
    .B(_05648_),
    .Y(_05649_));
 AND2x2_ASAP7_75t_R _16972_ (.A(_05600_),
    .B(_05649_),
    .Y(_03682_));
 OR3x1_ASAP7_75t_R _16973_ (.A(_01359_),
    .B(_05613_),
    .C(_05645_),
    .Y(_05650_));
 OAI21x1_ASAP7_75t_R _16974_ (.A1(_05613_),
    .A2(_05645_),
    .B(_01359_),
    .Y(_05651_));
 AND3x1_ASAP7_75t_R _16975_ (.A(_05626_),
    .B(_05650_),
    .C(_05651_),
    .Y(_03683_));
 BUFx6f_ASAP7_75t_R _16976_ (.A(_05426_),
    .Y(_05652_));
 OR3x1_ASAP7_75t_R _16977_ (.A(_01359_),
    .B(_05613_),
    .C(_05648_),
    .Y(_05653_));
 XOR2x2_ASAP7_75t_R _16978_ (.A(_01358_),
    .B(_05653_),
    .Y(_05654_));
 AND2x2_ASAP7_75t_R _16979_ (.A(_05652_),
    .B(_05654_),
    .Y(_03684_));
 NOR2x1_ASAP7_75t_R _16980_ (.A(_05300_),
    .B(_02626_),
    .Y(_03685_));
 OR4x1_ASAP7_75t_R _16981_ (.A(_01358_),
    .B(_01359_),
    .C(_05613_),
    .D(_05645_),
    .Y(_05655_));
 XOR2x2_ASAP7_75t_R _16982_ (.A(_01356_),
    .B(_05655_),
    .Y(_05656_));
 AND2x2_ASAP7_75t_R _16983_ (.A(_05652_),
    .B(_05656_),
    .Y(_03686_));
 OR5x1_ASAP7_75t_R _16984_ (.A(_01356_),
    .B(_01358_),
    .C(_01359_),
    .D(_05613_),
    .E(_05648_),
    .Y(_05657_));
 XOR2x2_ASAP7_75t_R _16985_ (.A(_01355_),
    .B(_05657_),
    .Y(_05658_));
 AND2x2_ASAP7_75t_R _16986_ (.A(_05652_),
    .B(_05658_),
    .Y(_03687_));
 OR5x2_ASAP7_75t_R _16987_ (.A(_01355_),
    .B(_01356_),
    .C(_01358_),
    .D(_01359_),
    .E(_05613_),
    .Y(_05659_));
 OR3x1_ASAP7_75t_R _16988_ (.A(_01354_),
    .B(_05645_),
    .C(_05659_),
    .Y(_05660_));
 OAI21x1_ASAP7_75t_R _16989_ (.A1(_05645_),
    .A2(_05659_),
    .B(_01354_),
    .Y(_05661_));
 AND3x1_ASAP7_75t_R _16990_ (.A(_05626_),
    .B(_05660_),
    .C(_05661_),
    .Y(_03688_));
 OR4x1_ASAP7_75t_R _16991_ (.A(_01353_),
    .B(_01354_),
    .C(_05648_),
    .D(_05659_),
    .Y(_05662_));
 OR3x1_ASAP7_75t_R _16992_ (.A(_01354_),
    .B(_05648_),
    .C(_05659_),
    .Y(_05663_));
 NAND2x1_ASAP7_75t_R _16993_ (.A(_01353_),
    .B(_05663_),
    .Y(_05664_));
 AND3x1_ASAP7_75t_R _16994_ (.A(_05626_),
    .B(_05662_),
    .C(_05664_),
    .Y(_03689_));
 OR4x1_ASAP7_75t_R _16995_ (.A(_01353_),
    .B(_01354_),
    .C(_05645_),
    .D(_05659_),
    .Y(_05665_));
 XOR2x2_ASAP7_75t_R _16996_ (.A(_05618_),
    .B(_05665_),
    .Y(_05666_));
 AND2x2_ASAP7_75t_R _16997_ (.A(_05652_),
    .B(_05666_),
    .Y(_03690_));
 OR3x1_ASAP7_75t_R _16998_ (.A(_01351_),
    .B(_05618_),
    .C(_05662_),
    .Y(_05667_));
 OAI21x1_ASAP7_75t_R _16999_ (.A1(_05618_),
    .A2(_05662_),
    .B(_01351_),
    .Y(_05668_));
 AND3x1_ASAP7_75t_R _17000_ (.A(_05626_),
    .B(_05667_),
    .C(_05668_),
    .Y(_03691_));
 OR3x1_ASAP7_75t_R _17001_ (.A(_01351_),
    .B(_05618_),
    .C(_05665_),
    .Y(_05669_));
 XOR2x2_ASAP7_75t_R _17002_ (.A(_01350_),
    .B(_05669_),
    .Y(_05670_));
 AND2x2_ASAP7_75t_R _17003_ (.A(_05652_),
    .B(_05670_),
    .Y(_03692_));
 OR4x1_ASAP7_75t_R _17004_ (.A(_01350_),
    .B(_01351_),
    .C(_05618_),
    .D(_05662_),
    .Y(_05671_));
 XOR2x2_ASAP7_75t_R _17005_ (.A(_01349_),
    .B(_05671_),
    .Y(_05672_));
 AND2x2_ASAP7_75t_R _17006_ (.A(_05652_),
    .B(_05672_),
    .Y(_03693_));
 OR5x1_ASAP7_75t_R _17007_ (.A(_01349_),
    .B(_01350_),
    .C(_01351_),
    .D(_05618_),
    .E(_05665_),
    .Y(_05673_));
 XOR2x2_ASAP7_75t_R _17008_ (.A(_01348_),
    .B(_05673_),
    .Y(_05674_));
 AND2x2_ASAP7_75t_R _17009_ (.A(_05652_),
    .B(_05674_),
    .Y(_03694_));
 OR5x2_ASAP7_75t_R _17010_ (.A(_01348_),
    .B(_01349_),
    .C(_01350_),
    .D(_01351_),
    .E(_05618_),
    .Y(_05675_));
 OR3x1_ASAP7_75t_R _17011_ (.A(_01347_),
    .B(_05662_),
    .C(_05675_),
    .Y(_05676_));
 OAI21x1_ASAP7_75t_R _17012_ (.A1(_05662_),
    .A2(_05675_),
    .B(_01347_),
    .Y(_05677_));
 AND3x1_ASAP7_75t_R _17013_ (.A(_05626_),
    .B(_05676_),
    .C(_05677_),
    .Y(_03695_));
 XOR2x2_ASAP7_75t_R _17014_ (.A(_01346_),
    .B(_02625_),
    .Y(_05678_));
 AND2x2_ASAP7_75t_R _17015_ (.A(_05652_),
    .B(_05678_),
    .Y(_03696_));
 OR3x1_ASAP7_75t_R _17016_ (.A(_01347_),
    .B(_05665_),
    .C(_05675_),
    .Y(_05679_));
 XOR2x2_ASAP7_75t_R _17017_ (.A(_01345_),
    .B(_05679_),
    .Y(_05680_));
 AND2x2_ASAP7_75t_R _17018_ (.A(_05652_),
    .B(_05680_),
    .Y(_03697_));
 OR4x1_ASAP7_75t_R _17019_ (.A(_01345_),
    .B(_01347_),
    .C(_05662_),
    .D(_05675_),
    .Y(_05681_));
 XOR2x2_ASAP7_75t_R _17020_ (.A(_01344_),
    .B(_05681_),
    .Y(_05682_));
 AND2x2_ASAP7_75t_R _17021_ (.A(_05652_),
    .B(_05682_),
    .Y(_03698_));
 BUFx6f_ASAP7_75t_R _17022_ (.A(_05426_),
    .Y(_05683_));
 OR3x1_ASAP7_75t_R _17023_ (.A(_01346_),
    .B(_01357_),
    .C(_00038_),
    .Y(_05684_));
 XOR2x2_ASAP7_75t_R _17024_ (.A(_01343_),
    .B(_05684_),
    .Y(_05685_));
 AND2x2_ASAP7_75t_R _17025_ (.A(_05683_),
    .B(_05685_),
    .Y(_03699_));
 OR3x1_ASAP7_75t_R _17026_ (.A(_01343_),
    .B(_01346_),
    .C(_02625_),
    .Y(_05686_));
 NAND2x1_ASAP7_75t_R _17027_ (.A(_01342_),
    .B(_05686_),
    .Y(_05687_));
 AND3x1_ASAP7_75t_R _17028_ (.A(_05626_),
    .B(_05627_),
    .C(_05687_),
    .Y(_03700_));
 XOR2x2_ASAP7_75t_R _17029_ (.A(_01341_),
    .B(_05632_),
    .Y(_05688_));
 AND2x2_ASAP7_75t_R _17030_ (.A(_05683_),
    .B(_05688_),
    .Y(_03701_));
 OR3x1_ASAP7_75t_R _17031_ (.A(_01340_),
    .B(_01341_),
    .C(_05627_),
    .Y(_05689_));
 OAI21x1_ASAP7_75t_R _17032_ (.A1(_01341_),
    .A2(_05627_),
    .B(_01340_),
    .Y(_05690_));
 AND3x1_ASAP7_75t_R _17033_ (.A(_05626_),
    .B(_05689_),
    .C(_05690_),
    .Y(_03702_));
 OR3x1_ASAP7_75t_R _17034_ (.A(_01340_),
    .B(_01341_),
    .C(_05632_),
    .Y(_05691_));
 XOR2x2_ASAP7_75t_R _17035_ (.A(_01339_),
    .B(_05691_),
    .Y(_05692_));
 AND2x2_ASAP7_75t_R _17036_ (.A(_05683_),
    .B(_05692_),
    .Y(_03703_));
 OR4x1_ASAP7_75t_R _17037_ (.A(_01339_),
    .B(_01340_),
    .C(_01341_),
    .D(_05627_),
    .Y(_05693_));
 NAND2x1_ASAP7_75t_R _17038_ (.A(_01338_),
    .B(_05693_),
    .Y(_05694_));
 AND3x1_ASAP7_75t_R _17039_ (.A(_05626_),
    .B(_05629_),
    .C(_05694_),
    .Y(_03704_));
 XOR2x2_ASAP7_75t_R _17040_ (.A(_05614_),
    .B(_05633_),
    .Y(_05695_));
 AND2x2_ASAP7_75t_R _17041_ (.A(_05683_),
    .B(_05695_),
    .Y(_03705_));
 AND2x2_ASAP7_75t_R _17042_ (.A(_05683_),
    .B(_00018_),
    .Y(_03706_));
 BUFx6f_ASAP7_75t_R _17043_ (.A(_02078_),
    .Y(_05696_));
 NAND2x1_ASAP7_75t_R _17044_ (.A(_01371_),
    .B(_01372_),
    .Y(_05697_));
 OR2x6_ASAP7_75t_R _17045_ (.A(_01369_),
    .B(_01370_),
    .Y(_05698_));
 OAI21x1_ASAP7_75t_R _17046_ (.A1(_05697_),
    .A2(_05698_),
    .B(\xs[12].cli1.i[39] ),
    .Y(_05699_));
 BUFx6f_ASAP7_75t_R _17047_ (.A(_02085_),
    .Y(_05700_));
 INVx1_ASAP7_75t_R _17048_ (.A(_05700_),
    .Y(_05701_));
 AND2x4_ASAP7_75t_R _17049_ (.A(_01410_),
    .B(_01411_),
    .Y(_05702_));
 NOR2x1_ASAP7_75t_R _17050_ (.A(_01408_),
    .B(_01409_),
    .Y(_05703_));
 AO21x2_ASAP7_75t_R _17051_ (.A1(_05702_),
    .A2(_05703_),
    .B(_01407_),
    .Y(_05704_));
 AO21x1_ASAP7_75t_R _17052_ (.A1(_02079_),
    .A2(_05701_),
    .B(_05704_),
    .Y(_05705_));
 OA21x2_ASAP7_75t_R _17053_ (.A1(_02079_),
    .A2(_05699_),
    .B(_05705_),
    .Y(_05706_));
 OR4x1_ASAP7_75t_R _17054_ (.A(_01368_),
    .B(\peo[25][32] ),
    .C(_05697_),
    .D(_05698_),
    .Y(_05707_));
 INVx1_ASAP7_75t_R _17055_ (.A(_05707_),
    .Y(_05708_));
 OA21x2_ASAP7_75t_R _17056_ (.A1(_05696_),
    .A2(_05706_),
    .B(_05708_),
    .Y(_05709_));
 INVx2_ASAP7_75t_R _17057_ (.A(_05696_),
    .Y(_05710_));
 AND2x4_ASAP7_75t_R _17058_ (.A(_05710_),
    .B(_02079_),
    .Y(_05711_));
 AOI21x1_ASAP7_75t_R _17059_ (.A1(_05702_),
    .A2(_05703_),
    .B(_01407_),
    .Y(_05712_));
 NAND2x1_ASAP7_75t_R _17060_ (.A(_05710_),
    .B(_05700_),
    .Y(_05713_));
 OR3x1_ASAP7_75t_R _17061_ (.A(_05696_),
    .B(_01407_),
    .C(_01412_),
    .Y(_05714_));
 NAND2x1_ASAP7_75t_R _17062_ (.A(_05702_),
    .B(_05703_),
    .Y(_05715_));
 OA22x2_ASAP7_75t_R _17063_ (.A1(_05712_),
    .A2(_05713_),
    .B1(_05714_),
    .B2(_05715_),
    .Y(_05716_));
 OA21x2_ASAP7_75t_R _17064_ (.A1(_05697_),
    .A2(_05698_),
    .B(\xs[12].cli1.i[39] ),
    .Y(_05717_));
 OR4x1_ASAP7_75t_R _17065_ (.A(_05700_),
    .B(_05715_),
    .C(_05717_),
    .D(_05714_),
    .Y(_05718_));
 OA21x2_ASAP7_75t_R _17066_ (.A1(_05707_),
    .A2(_05716_),
    .B(_05718_),
    .Y(_05719_));
 NAND3x1_ASAP7_75t_R _17067_ (.A(_05700_),
    .B(_05711_),
    .C(_05719_),
    .Y(_05720_));
 AND4x1_ASAP7_75t_R _17068_ (.A(_05700_),
    .B(_02089_),
    .C(_05711_),
    .D(_05719_),
    .Y(_05721_));
 AOI21x1_ASAP7_75t_R _17069_ (.A1(_01414_),
    .A2(_05720_),
    .B(_05721_),
    .Y(_05722_));
 NAND2x1_ASAP7_75t_R _17070_ (.A(_01375_),
    .B(_05709_),
    .Y(_05723_));
 OA211x2_ASAP7_75t_R _17071_ (.A1(_05709_),
    .A2(_05722_),
    .B(_05723_),
    .C(_11589_),
    .Y(_03707_));
 NAND2x1_ASAP7_75t_R _17072_ (.A(_05711_),
    .B(_05719_),
    .Y(_05724_));
 OR3x2_ASAP7_75t_R _17073_ (.A(_10763_),
    .B(_05701_),
    .C(_05724_),
    .Y(_05725_));
 NOR2x1_ASAP7_75t_R _17074_ (.A(_02088_),
    .B(_05725_),
    .Y(_03708_));
 NOR2x1_ASAP7_75t_R _17075_ (.A(_02087_),
    .B(_05725_),
    .Y(_03709_));
 NOR2x1_ASAP7_75t_R _17076_ (.A(_02086_),
    .B(_05725_),
    .Y(_03710_));
 NOR2x1_ASAP7_75t_R _17077_ (.A(_02077_),
    .B(_05725_),
    .Y(_03711_));
 NOR2x1_ASAP7_75t_R _17078_ (.A(_02076_),
    .B(_05725_),
    .Y(_03712_));
 OAI21x1_ASAP7_75t_R _17079_ (.A1(_05700_),
    .A2(_05724_),
    .B(_01414_),
    .Y(_05726_));
 INVx1_ASAP7_75t_R _17080_ (.A(_02089_),
    .Y(_05727_));
 OR3x1_ASAP7_75t_R _17081_ (.A(_05700_),
    .B(_05727_),
    .C(_05724_),
    .Y(_05728_));
 AND2x2_ASAP7_75t_R _17082_ (.A(_05696_),
    .B(_05717_),
    .Y(_05729_));
 OA21x2_ASAP7_75t_R _17083_ (.A1(_05701_),
    .A2(_05704_),
    .B(_02079_),
    .Y(_05730_));
 OA21x2_ASAP7_75t_R _17084_ (.A1(_05707_),
    .A2(_05704_),
    .B(_05699_),
    .Y(_05731_));
 NOR2x1_ASAP7_75t_R _17085_ (.A(_05730_),
    .B(_05731_),
    .Y(_05732_));
 AO32x1_ASAP7_75t_R _17086_ (.A1(_00018_),
    .A2(_05712_),
    .A3(_05729_),
    .B1(_05732_),
    .B2(_05710_),
    .Y(_05733_));
 NOR2x1_ASAP7_75t_R _17087_ (.A(_09314_),
    .B(_05733_),
    .Y(_05734_));
 NOR2x1_ASAP7_75t_R _17088_ (.A(_09924_),
    .B(_01375_),
    .Y(_05735_));
 AO32x1_ASAP7_75t_R _17089_ (.A1(_05726_),
    .A2(_05728_),
    .A3(_05734_),
    .B1(_05733_),
    .B2(_05735_),
    .Y(_03713_));
 OR3x2_ASAP7_75t_R _17090_ (.A(_10763_),
    .B(_05700_),
    .C(_05724_),
    .Y(_05736_));
 NOR2x1_ASAP7_75t_R _17091_ (.A(_02088_),
    .B(_05736_),
    .Y(_03714_));
 NOR2x1_ASAP7_75t_R _17092_ (.A(_02087_),
    .B(_05736_),
    .Y(_03715_));
 NOR2x1_ASAP7_75t_R _17093_ (.A(_02086_),
    .B(_05736_),
    .Y(_03716_));
 NOR2x1_ASAP7_75t_R _17094_ (.A(_02077_),
    .B(_05736_),
    .Y(_03717_));
 NOR2x1_ASAP7_75t_R _17095_ (.A(_02076_),
    .B(_05736_),
    .Y(_03718_));
 OAI21x1_ASAP7_75t_R _17096_ (.A1(_05696_),
    .A2(_02079_),
    .B(_05719_),
    .Y(_05737_));
 NAND2x1_ASAP7_75t_R _17097_ (.A(_00018_),
    .B(_05712_),
    .Y(_05738_));
 OA211x2_ASAP7_75t_R _17098_ (.A1(_05701_),
    .A2(_05704_),
    .B(_05717_),
    .C(_05711_),
    .Y(_05739_));
 AOI21x1_ASAP7_75t_R _17099_ (.A1(_05738_),
    .A2(_05729_),
    .B(_05739_),
    .Y(_05740_));
 BUFx6f_ASAP7_75t_R _17100_ (.A(_05740_),
    .Y(_05741_));
 NAND2x1_ASAP7_75t_R _17101_ (.A(\peo[24][0] ),
    .B(_05741_),
    .Y(_05742_));
 OA21x2_ASAP7_75t_R _17102_ (.A1(_05696_),
    .A2(_02079_),
    .B(_05719_),
    .Y(_05743_));
 OA211x2_ASAP7_75t_R _17103_ (.A1(_01375_),
    .A2(_05741_),
    .B(_05742_),
    .C(_05743_),
    .Y(_05744_));
 AOI211x1_ASAP7_75t_R _17104_ (.A1(_02089_),
    .A2(_05737_),
    .B(_05744_),
    .C(_10995_),
    .Y(_03719_));
 NAND2x2_ASAP7_75t_R _17105_ (.A(_09029_),
    .B(_05737_),
    .Y(_05745_));
 NOR2x1_ASAP7_75t_R _17106_ (.A(_02088_),
    .B(_05745_),
    .Y(_03720_));
 NOR2x1_ASAP7_75t_R _17107_ (.A(_02087_),
    .B(_05745_),
    .Y(_03721_));
 NOR2x1_ASAP7_75t_R _17108_ (.A(_02086_),
    .B(_05745_),
    .Y(_03722_));
 NAND2x1_ASAP7_75t_R _17109_ (.A(\peo[24][32] ),
    .B(_05741_),
    .Y(_05746_));
 OA211x2_ASAP7_75t_R _17110_ (.A1(_01373_),
    .A2(_05741_),
    .B(_05746_),
    .C(_05743_),
    .Y(_05747_));
 AOI211x1_ASAP7_75t_R _17111_ (.A1(_05700_),
    .A2(_05737_),
    .B(_05747_),
    .C(_10995_),
    .Y(_03723_));
 NAND2x1_ASAP7_75t_R _17112_ (.A(\peo[24][33] ),
    .B(_05741_),
    .Y(_05748_));
 OA211x2_ASAP7_75t_R _17113_ (.A1(_01372_),
    .A2(_05741_),
    .B(_05748_),
    .C(_05743_),
    .Y(_05749_));
 AOI211x1_ASAP7_75t_R _17114_ (.A1(_02084_),
    .A2(_05737_),
    .B(_05749_),
    .C(_10995_),
    .Y(_03724_));
 NAND2x1_ASAP7_75t_R _17115_ (.A(\peo[24][34] ),
    .B(_05741_),
    .Y(_05750_));
 OA211x2_ASAP7_75t_R _17116_ (.A1(_01371_),
    .A2(_05741_),
    .B(_05750_),
    .C(_05743_),
    .Y(_05751_));
 AOI211x1_ASAP7_75t_R _17117_ (.A1(_02083_),
    .A2(_05737_),
    .B(_05751_),
    .C(_09145_),
    .Y(_03725_));
 NAND2x1_ASAP7_75t_R _17118_ (.A(\peo[24][35] ),
    .B(_05740_),
    .Y(_05752_));
 OA211x2_ASAP7_75t_R _17119_ (.A1(_01370_),
    .A2(_05741_),
    .B(_05752_),
    .C(_05743_),
    .Y(_05753_));
 AOI211x1_ASAP7_75t_R _17120_ (.A1(_02082_),
    .A2(_05737_),
    .B(_05753_),
    .C(_09145_),
    .Y(_03726_));
 NAND2x1_ASAP7_75t_R _17121_ (.A(\peo[24][36] ),
    .B(_05740_),
    .Y(_05754_));
 OA211x2_ASAP7_75t_R _17122_ (.A1(_01369_),
    .A2(_05741_),
    .B(_05754_),
    .C(_05743_),
    .Y(_05755_));
 AOI211x1_ASAP7_75t_R _17123_ (.A1(_02081_),
    .A2(_05737_),
    .B(_05755_),
    .C(_09145_),
    .Y(_03727_));
 NOR2x1_ASAP7_75t_R _17124_ (.A(_02080_),
    .B(_05745_),
    .Y(_03728_));
 OR2x2_ASAP7_75t_R _17125_ (.A(_05707_),
    .B(_05713_),
    .Y(_05756_));
 OA21x2_ASAP7_75t_R _17126_ (.A1(_05700_),
    .A2(_05717_),
    .B(_05707_),
    .Y(_05757_));
 OR3x1_ASAP7_75t_R _17127_ (.A(_05696_),
    .B(_01412_),
    .C(_05757_),
    .Y(_05758_));
 AO21x1_ASAP7_75t_R _17128_ (.A1(_01407_),
    .A2(_05756_),
    .B(_05712_),
    .Y(_05759_));
 AOI21x1_ASAP7_75t_R _17129_ (.A1(_05756_),
    .A2(_05758_),
    .B(_05759_),
    .Y(_05760_));
 OA211x2_ASAP7_75t_R _17130_ (.A1(_05696_),
    .A2(_02079_),
    .B(_05760_),
    .C(_11589_),
    .Y(_03729_));
 OR3x1_ASAP7_75t_R _17131_ (.A(_05712_),
    .B(_05717_),
    .C(_05737_),
    .Y(_05761_));
 AND2x2_ASAP7_75t_R _17132_ (.A(_05683_),
    .B(_05761_),
    .Y(_03730_));
 NOR2x1_ASAP7_75t_R _17133_ (.A(_02077_),
    .B(_05745_),
    .Y(_03731_));
 NOR2x1_ASAP7_75t_R _17134_ (.A(_02076_),
    .B(_05745_),
    .Y(_03732_));
 BUFx3_ASAP7_75t_R _17135_ (.A(_01299_),
    .Y(_05762_));
 BUFx3_ASAP7_75t_R _17136_ (.A(_01272_),
    .Y(_05763_));
 AND4x1_ASAP7_75t_R _17137_ (.A(_05763_),
    .B(_01300_),
    .C(_01301_),
    .D(_01302_),
    .Y(_05764_));
 AND5x1_ASAP7_75t_R _17138_ (.A(_01291_),
    .B(_01296_),
    .C(_01297_),
    .D(_05762_),
    .E(_05764_),
    .Y(_05765_));
 AND5x2_ASAP7_75t_R _17139_ (.A(_01293_),
    .B(_01294_),
    .C(_01295_),
    .D(_11466_),
    .E(_05765_),
    .Y(_05766_));
 AND4x1_ASAP7_75t_R _17140_ (.A(_01286_),
    .B(_01287_),
    .C(_01288_),
    .D(_01289_),
    .Y(_05767_));
 AND4x1_ASAP7_75t_R _17141_ (.A(_01280_),
    .B(_01282_),
    .C(_01283_),
    .D(_01290_),
    .Y(_05768_));
 AND5x1_ASAP7_75t_R _17142_ (.A(_01273_),
    .B(_01274_),
    .C(_01279_),
    .D(_01298_),
    .E(_05768_),
    .Y(_05769_));
 AND3x1_ASAP7_75t_R _17143_ (.A(_01277_),
    .B(_01278_),
    .C(_01281_),
    .Y(_05770_));
 OR3x1_ASAP7_75t_R _17144_ (.A(_01275_),
    .B(_01276_),
    .C(_05770_),
    .Y(_05771_));
 AND5x2_ASAP7_75t_R _17145_ (.A(_01284_),
    .B(_01285_),
    .C(_05767_),
    .D(_05769_),
    .E(_05771_),
    .Y(_05772_));
 NAND2x2_ASAP7_75t_R _17146_ (.A(_05766_),
    .B(_05772_),
    .Y(_05773_));
 NOR2x1_ASAP7_75t_R _17147_ (.A(_01229_),
    .B(_05773_),
    .Y(_03733_));
 INVx1_ASAP7_75t_R _17148_ (.A(_05773_),
    .Y(_03734_));
 NOR2x1_ASAP7_75t_R _17149_ (.A(_01232_),
    .B(_05773_),
    .Y(_03735_));
 NOR2x1_ASAP7_75t_R _17150_ (.A(_01231_),
    .B(_05773_),
    .Y(_03736_));
 NOR2x1_ASAP7_75t_R _17151_ (.A(_01230_),
    .B(_05773_),
    .Y(_03737_));
 NOR2x1_ASAP7_75t_R _17152_ (.A(_01228_),
    .B(_05773_),
    .Y(_03738_));
 NOR2x1_ASAP7_75t_R _17153_ (.A(_01227_),
    .B(_05773_),
    .Y(_03739_));
 INVx1_ASAP7_75t_R _17154_ (.A(_05773_),
    .Y(_03740_));
 AND2x2_ASAP7_75t_R _17155_ (.A(_05683_),
    .B(_00039_),
    .Y(_03741_));
 BUFx6f_ASAP7_75t_R _17156_ (.A(_05337_),
    .Y(_05774_));
 OR4x1_ASAP7_75t_R _17157_ (.A(_01277_),
    .B(_01278_),
    .C(_01281_),
    .D(_02645_),
    .Y(_05775_));
 OR4x1_ASAP7_75t_R _17158_ (.A(_01273_),
    .B(_01274_),
    .C(_01275_),
    .D(_01276_),
    .Y(_05776_));
 OR2x6_ASAP7_75t_R _17159_ (.A(_05775_),
    .B(_05776_),
    .Y(_05777_));
 OR3x1_ASAP7_75t_R _17160_ (.A(_05763_),
    .B(_01302_),
    .C(_05777_),
    .Y(_05778_));
 OAI21x1_ASAP7_75t_R _17161_ (.A1(_05763_),
    .A2(_05777_),
    .B(_01302_),
    .Y(_05779_));
 AND3x1_ASAP7_75t_R _17162_ (.A(_05774_),
    .B(_05778_),
    .C(_05779_),
    .Y(_03742_));
 OR5x2_ASAP7_75t_R _17163_ (.A(_01277_),
    .B(_01278_),
    .C(_01281_),
    .D(_01292_),
    .E(_00039_),
    .Y(_05780_));
 OR2x2_ASAP7_75t_R _17164_ (.A(_05776_),
    .B(_05780_),
    .Y(_05781_));
 OR3x1_ASAP7_75t_R _17165_ (.A(_05763_),
    .B(_01302_),
    .C(_05781_),
    .Y(_05782_));
 XOR2x2_ASAP7_75t_R _17166_ (.A(_01301_),
    .B(_05782_),
    .Y(_05783_));
 AND2x2_ASAP7_75t_R _17167_ (.A(_05683_),
    .B(_05783_),
    .Y(_03743_));
 OR4x1_ASAP7_75t_R _17168_ (.A(_05763_),
    .B(_01300_),
    .C(_01301_),
    .D(_01302_),
    .Y(_05784_));
 OR3x2_ASAP7_75t_R _17169_ (.A(_05775_),
    .B(_05776_),
    .C(_05784_),
    .Y(_05785_));
 OR4x1_ASAP7_75t_R _17170_ (.A(_05763_),
    .B(_01301_),
    .C(_01302_),
    .D(_05777_),
    .Y(_05786_));
 NAND2x1_ASAP7_75t_R _17171_ (.A(_01300_),
    .B(_05786_),
    .Y(_05787_));
 AND3x1_ASAP7_75t_R _17172_ (.A(_05774_),
    .B(_05785_),
    .C(_05787_),
    .Y(_03744_));
 OR3x2_ASAP7_75t_R _17173_ (.A(_05776_),
    .B(_05780_),
    .C(_05784_),
    .Y(_05788_));
 XOR2x2_ASAP7_75t_R _17174_ (.A(_05762_),
    .B(_05788_),
    .Y(_05789_));
 AND2x2_ASAP7_75t_R _17175_ (.A(_05683_),
    .B(_05789_),
    .Y(_03745_));
 OR3x1_ASAP7_75t_R _17176_ (.A(_01298_),
    .B(_05762_),
    .C(_05785_),
    .Y(_05790_));
 OAI21x1_ASAP7_75t_R _17177_ (.A1(_05762_),
    .A2(_05785_),
    .B(_01298_),
    .Y(_05791_));
 AND3x1_ASAP7_75t_R _17178_ (.A(_05774_),
    .B(_05790_),
    .C(_05791_),
    .Y(_03746_));
 OR3x1_ASAP7_75t_R _17179_ (.A(_01298_),
    .B(_05762_),
    .C(_05788_),
    .Y(_05792_));
 XOR2x2_ASAP7_75t_R _17180_ (.A(_01297_),
    .B(_05792_),
    .Y(_05793_));
 AND2x2_ASAP7_75t_R _17181_ (.A(_05683_),
    .B(_05793_),
    .Y(_03747_));
 BUFx6f_ASAP7_75t_R _17182_ (.A(_05426_),
    .Y(_05794_));
 OR4x1_ASAP7_75t_R _17183_ (.A(_01297_),
    .B(_01298_),
    .C(_05762_),
    .D(_05785_),
    .Y(_05795_));
 XOR2x2_ASAP7_75t_R _17184_ (.A(_01296_),
    .B(_05795_),
    .Y(_05796_));
 AND2x2_ASAP7_75t_R _17185_ (.A(_05794_),
    .B(_05796_),
    .Y(_03748_));
 OR5x1_ASAP7_75t_R _17186_ (.A(_01296_),
    .B(_01297_),
    .C(_01298_),
    .D(_05762_),
    .E(_05788_),
    .Y(_05797_));
 XOR2x2_ASAP7_75t_R _17187_ (.A(_01295_),
    .B(_05797_),
    .Y(_05798_));
 AND2x2_ASAP7_75t_R _17188_ (.A(_05794_),
    .B(_05798_),
    .Y(_03749_));
 OR5x2_ASAP7_75t_R _17189_ (.A(_01295_),
    .B(_01296_),
    .C(_01297_),
    .D(_01298_),
    .E(_05762_),
    .Y(_05799_));
 OR3x2_ASAP7_75t_R _17190_ (.A(_01294_),
    .B(_05785_),
    .C(_05799_),
    .Y(_05800_));
 OAI21x1_ASAP7_75t_R _17191_ (.A1(_05785_),
    .A2(_05799_),
    .B(_01294_),
    .Y(_05801_));
 AND3x1_ASAP7_75t_R _17192_ (.A(_05774_),
    .B(_05800_),
    .C(_05801_),
    .Y(_03750_));
 OR3x2_ASAP7_75t_R _17193_ (.A(_01294_),
    .B(_05788_),
    .C(_05799_),
    .Y(_05802_));
 XOR2x2_ASAP7_75t_R _17194_ (.A(_01293_),
    .B(_05802_),
    .Y(_05803_));
 AND2x2_ASAP7_75t_R _17195_ (.A(_05794_),
    .B(_05803_),
    .Y(_03751_));
 NOR2x1_ASAP7_75t_R _17196_ (.A(_05300_),
    .B(_02646_),
    .Y(_03752_));
 OR3x1_ASAP7_75t_R _17197_ (.A(_01291_),
    .B(_01293_),
    .C(_05800_),
    .Y(_05804_));
 OAI21x1_ASAP7_75t_R _17198_ (.A1(_01293_),
    .A2(_05800_),
    .B(_01291_),
    .Y(_05805_));
 AND3x1_ASAP7_75t_R _17199_ (.A(_05774_),
    .B(_05804_),
    .C(_05805_),
    .Y(_03753_));
 OR3x1_ASAP7_75t_R _17200_ (.A(_01291_),
    .B(_01293_),
    .C(_05802_),
    .Y(_05806_));
 XOR2x2_ASAP7_75t_R _17201_ (.A(_01290_),
    .B(_05806_),
    .Y(_05807_));
 AND2x2_ASAP7_75t_R _17202_ (.A(_05794_),
    .B(_05807_),
    .Y(_03754_));
 OR4x1_ASAP7_75t_R _17203_ (.A(_01290_),
    .B(_01291_),
    .C(_01293_),
    .D(_05800_),
    .Y(_05808_));
 XOR2x2_ASAP7_75t_R _17204_ (.A(_01289_),
    .B(_05808_),
    .Y(_05809_));
 AND2x2_ASAP7_75t_R _17205_ (.A(_05794_),
    .B(_05809_),
    .Y(_03755_));
 OR4x1_ASAP7_75t_R _17206_ (.A(_01289_),
    .B(_01290_),
    .C(_01291_),
    .D(_01293_),
    .Y(_05810_));
 OR3x2_ASAP7_75t_R _17207_ (.A(_01288_),
    .B(_05802_),
    .C(_05810_),
    .Y(_05811_));
 OAI21x1_ASAP7_75t_R _17208_ (.A1(_05802_),
    .A2(_05810_),
    .B(_01288_),
    .Y(_05812_));
 AND3x1_ASAP7_75t_R _17209_ (.A(_05774_),
    .B(_05811_),
    .C(_05812_),
    .Y(_03756_));
 OR3x2_ASAP7_75t_R _17210_ (.A(_01288_),
    .B(_05800_),
    .C(_05810_),
    .Y(_05813_));
 XOR2x2_ASAP7_75t_R _17211_ (.A(_01287_),
    .B(_05813_),
    .Y(_05814_));
 AND2x2_ASAP7_75t_R _17212_ (.A(_05794_),
    .B(_05814_),
    .Y(_03757_));
 OR3x1_ASAP7_75t_R _17213_ (.A(_01286_),
    .B(_01287_),
    .C(_05811_),
    .Y(_05815_));
 OAI21x1_ASAP7_75t_R _17214_ (.A1(_01287_),
    .A2(_05811_),
    .B(_01286_),
    .Y(_05816_));
 AND3x1_ASAP7_75t_R _17215_ (.A(_05774_),
    .B(_05815_),
    .C(_05816_),
    .Y(_03758_));
 OR3x1_ASAP7_75t_R _17216_ (.A(_01286_),
    .B(_01287_),
    .C(_05813_),
    .Y(_05817_));
 XOR2x2_ASAP7_75t_R _17217_ (.A(_01285_),
    .B(_05817_),
    .Y(_05818_));
 AND2x2_ASAP7_75t_R _17218_ (.A(_05794_),
    .B(_05818_),
    .Y(_03759_));
 OR4x1_ASAP7_75t_R _17219_ (.A(_01285_),
    .B(_01286_),
    .C(_01287_),
    .D(_05811_),
    .Y(_05819_));
 XOR2x2_ASAP7_75t_R _17220_ (.A(_01284_),
    .B(_05819_),
    .Y(_05820_));
 AND2x2_ASAP7_75t_R _17221_ (.A(_05794_),
    .B(_05820_),
    .Y(_03760_));
 OR4x1_ASAP7_75t_R _17222_ (.A(_01284_),
    .B(_01285_),
    .C(_01286_),
    .D(_01287_),
    .Y(_05821_));
 OR3x1_ASAP7_75t_R _17223_ (.A(_01283_),
    .B(_05813_),
    .C(_05821_),
    .Y(_05822_));
 OAI21x1_ASAP7_75t_R _17224_ (.A1(_05813_),
    .A2(_05821_),
    .B(_01283_),
    .Y(_05823_));
 AND3x1_ASAP7_75t_R _17225_ (.A(_05774_),
    .B(_05822_),
    .C(_05823_),
    .Y(_03761_));
 OR3x1_ASAP7_75t_R _17226_ (.A(_01283_),
    .B(_05811_),
    .C(_05821_),
    .Y(_05824_));
 XOR2x2_ASAP7_75t_R _17227_ (.A(_01282_),
    .B(_05824_),
    .Y(_05825_));
 AND2x2_ASAP7_75t_R _17228_ (.A(_05794_),
    .B(_05825_),
    .Y(_03762_));
 XOR2x2_ASAP7_75t_R _17229_ (.A(_01281_),
    .B(_02645_),
    .Y(_05826_));
 AND2x2_ASAP7_75t_R _17230_ (.A(_05794_),
    .B(_05826_),
    .Y(_03763_));
 BUFx6f_ASAP7_75t_R _17231_ (.A(_05426_),
    .Y(_05827_));
 OR4x1_ASAP7_75t_R _17232_ (.A(_01282_),
    .B(_01283_),
    .C(_05813_),
    .D(_05821_),
    .Y(_05828_));
 XOR2x2_ASAP7_75t_R _17233_ (.A(_01280_),
    .B(_05828_),
    .Y(_05829_));
 AND2x2_ASAP7_75t_R _17234_ (.A(_05827_),
    .B(_05829_),
    .Y(_03764_));
 OR5x1_ASAP7_75t_R _17235_ (.A(_01280_),
    .B(_01282_),
    .C(_01283_),
    .D(_05811_),
    .E(_05821_),
    .Y(_05830_));
 XOR2x2_ASAP7_75t_R _17236_ (.A(_01279_),
    .B(_05830_),
    .Y(_05831_));
 AND2x2_ASAP7_75t_R _17237_ (.A(_05827_),
    .B(_05831_),
    .Y(_03765_));
 OR3x1_ASAP7_75t_R _17238_ (.A(_01281_),
    .B(_01292_),
    .C(_00039_),
    .Y(_05832_));
 XOR2x2_ASAP7_75t_R _17239_ (.A(_01278_),
    .B(_05832_),
    .Y(_05833_));
 AND2x2_ASAP7_75t_R _17240_ (.A(_05827_),
    .B(_05833_),
    .Y(_03766_));
 OR3x1_ASAP7_75t_R _17241_ (.A(_01278_),
    .B(_01281_),
    .C(_02645_),
    .Y(_05834_));
 NAND2x1_ASAP7_75t_R _17242_ (.A(_01277_),
    .B(_05834_),
    .Y(_05835_));
 AND3x1_ASAP7_75t_R _17243_ (.A(_05774_),
    .B(_05775_),
    .C(_05835_),
    .Y(_03767_));
 XOR2x2_ASAP7_75t_R _17244_ (.A(_01276_),
    .B(_05780_),
    .Y(_05836_));
 AND2x2_ASAP7_75t_R _17245_ (.A(_05827_),
    .B(_05836_),
    .Y(_03768_));
 OR3x1_ASAP7_75t_R _17246_ (.A(_01275_),
    .B(_01276_),
    .C(_05775_),
    .Y(_05837_));
 OAI21x1_ASAP7_75t_R _17247_ (.A1(_01276_),
    .A2(_05775_),
    .B(_01275_),
    .Y(_05838_));
 AND3x1_ASAP7_75t_R _17248_ (.A(_05774_),
    .B(_05837_),
    .C(_05838_),
    .Y(_03769_));
 OR3x1_ASAP7_75t_R _17249_ (.A(_01275_),
    .B(_01276_),
    .C(_05780_),
    .Y(_05839_));
 XOR2x2_ASAP7_75t_R _17250_ (.A(_01274_),
    .B(_05839_),
    .Y(_05840_));
 AND2x2_ASAP7_75t_R _17251_ (.A(_05827_),
    .B(_05840_),
    .Y(_03770_));
 BUFx6f_ASAP7_75t_R _17252_ (.A(_05337_),
    .Y(_05841_));
 OR4x1_ASAP7_75t_R _17253_ (.A(_01274_),
    .B(_01275_),
    .C(_01276_),
    .D(_05775_),
    .Y(_05842_));
 NAND2x1_ASAP7_75t_R _17254_ (.A(_01273_),
    .B(_05842_),
    .Y(_05843_));
 AND3x1_ASAP7_75t_R _17255_ (.A(_05841_),
    .B(_05777_),
    .C(_05843_),
    .Y(_03771_));
 XOR2x2_ASAP7_75t_R _17256_ (.A(_05763_),
    .B(_05781_),
    .Y(_05844_));
 AND2x2_ASAP7_75t_R _17257_ (.A(_05827_),
    .B(_05844_),
    .Y(_03772_));
 BUFx6f_ASAP7_75t_R _17258_ (.A(_01256_),
    .Y(_05845_));
 BUFx3_ASAP7_75t_R _17259_ (.A(_01233_),
    .Y(_05846_));
 AND4x1_ASAP7_75t_R _17260_ (.A(_05846_),
    .B(_01261_),
    .C(_01262_),
    .D(_01263_),
    .Y(_05847_));
 AND5x1_ASAP7_75t_R _17261_ (.A(_01252_),
    .B(_01257_),
    .C(_01258_),
    .D(_01260_),
    .E(_05847_),
    .Y(_05848_));
 AND5x2_ASAP7_75t_R _17262_ (.A(_01254_),
    .B(_01255_),
    .C(_05845_),
    .D(_11466_),
    .E(_05848_),
    .Y(_05849_));
 BUFx6f_ASAP7_75t_R _17263_ (.A(_01248_),
    .Y(_05850_));
 AND4x1_ASAP7_75t_R _17264_ (.A(_01247_),
    .B(_05850_),
    .C(_01249_),
    .D(_01250_),
    .Y(_05851_));
 AND4x1_ASAP7_75t_R _17265_ (.A(_01241_),
    .B(_01243_),
    .C(_01244_),
    .D(_01251_),
    .Y(_05852_));
 AND5x1_ASAP7_75t_R _17266_ (.A(_01234_),
    .B(_01235_),
    .C(_01240_),
    .D(_01259_),
    .E(_05852_),
    .Y(_05853_));
 AND3x1_ASAP7_75t_R _17267_ (.A(_01238_),
    .B(_01239_),
    .C(_01242_),
    .Y(_05854_));
 OR3x1_ASAP7_75t_R _17268_ (.A(_01236_),
    .B(_01237_),
    .C(_05854_),
    .Y(_05855_));
 AND5x2_ASAP7_75t_R _17269_ (.A(_01245_),
    .B(_01246_),
    .C(_05851_),
    .D(_05853_),
    .E(_05855_),
    .Y(_05856_));
 NAND2x2_ASAP7_75t_R _17270_ (.A(_05849_),
    .B(_05856_),
    .Y(_05857_));
 NOR2x1_ASAP7_75t_R _17271_ (.A(_01223_),
    .B(_05857_),
    .Y(_03773_));
 INVx1_ASAP7_75t_R _17272_ (.A(_05857_),
    .Y(_03774_));
 NOR2x1_ASAP7_75t_R _17273_ (.A(_01226_),
    .B(_05857_),
    .Y(_03775_));
 NOR2x1_ASAP7_75t_R _17274_ (.A(_01225_),
    .B(_05857_),
    .Y(_03776_));
 NOR2x1_ASAP7_75t_R _17275_ (.A(_01224_),
    .B(_05857_),
    .Y(_03777_));
 NOR2x1_ASAP7_75t_R _17276_ (.A(_01222_),
    .B(_05857_),
    .Y(_03778_));
 NOR2x1_ASAP7_75t_R _17277_ (.A(_01221_),
    .B(_05857_),
    .Y(_03779_));
 INVx1_ASAP7_75t_R _17278_ (.A(_05857_),
    .Y(_03780_));
 AND2x2_ASAP7_75t_R _17279_ (.A(_05827_),
    .B(_00040_),
    .Y(_03781_));
 OR4x1_ASAP7_75t_R _17280_ (.A(_01238_),
    .B(_01239_),
    .C(_01242_),
    .D(_02613_),
    .Y(_05858_));
 OR4x1_ASAP7_75t_R _17281_ (.A(_01234_),
    .B(_01235_),
    .C(_01236_),
    .D(_01237_),
    .Y(_05859_));
 OR2x6_ASAP7_75t_R _17282_ (.A(_05858_),
    .B(_05859_),
    .Y(_05860_));
 OR3x1_ASAP7_75t_R _17283_ (.A(_05846_),
    .B(_01263_),
    .C(_05860_),
    .Y(_05861_));
 OAI21x1_ASAP7_75t_R _17284_ (.A1(_05846_),
    .A2(_05860_),
    .B(_01263_),
    .Y(_05862_));
 AND3x1_ASAP7_75t_R _17285_ (.A(_05841_),
    .B(_05861_),
    .C(_05862_),
    .Y(_03782_));
 OR5x2_ASAP7_75t_R _17286_ (.A(_01238_),
    .B(_01239_),
    .C(_01242_),
    .D(_01253_),
    .E(_00040_),
    .Y(_05863_));
 OR2x6_ASAP7_75t_R _17287_ (.A(_05859_),
    .B(_05863_),
    .Y(_05864_));
 OR3x1_ASAP7_75t_R _17288_ (.A(_05846_),
    .B(_01263_),
    .C(_05864_),
    .Y(_05865_));
 XOR2x2_ASAP7_75t_R _17289_ (.A(_01262_),
    .B(_05865_),
    .Y(_05866_));
 AND2x2_ASAP7_75t_R _17290_ (.A(_05827_),
    .B(_05866_),
    .Y(_03783_));
 OR4x1_ASAP7_75t_R _17291_ (.A(_05846_),
    .B(_01262_),
    .C(_01263_),
    .D(_05860_),
    .Y(_05867_));
 XOR2x2_ASAP7_75t_R _17292_ (.A(_01261_),
    .B(_05867_),
    .Y(_05868_));
 AND2x2_ASAP7_75t_R _17293_ (.A(_05827_),
    .B(_05868_),
    .Y(_03784_));
 OR5x2_ASAP7_75t_R _17294_ (.A(_05846_),
    .B(_01260_),
    .C(_01261_),
    .D(_01262_),
    .E(_01263_),
    .Y(_05869_));
 OR5x1_ASAP7_75t_R _17295_ (.A(_05846_),
    .B(_01261_),
    .C(_01262_),
    .D(_01263_),
    .E(_05864_),
    .Y(_05870_));
 NAND2x1_ASAP7_75t_R _17296_ (.A(_01260_),
    .B(_05870_),
    .Y(_05871_));
 OA211x2_ASAP7_75t_R _17297_ (.A1(_05864_),
    .A2(_05869_),
    .B(_05871_),
    .C(_11589_),
    .Y(_03785_));
 OR3x1_ASAP7_75t_R _17298_ (.A(_05858_),
    .B(_05859_),
    .C(_05869_),
    .Y(_05872_));
 XOR2x2_ASAP7_75t_R _17299_ (.A(_01259_),
    .B(_05872_),
    .Y(_05873_));
 AND2x2_ASAP7_75t_R _17300_ (.A(_05827_),
    .B(_05873_),
    .Y(_03786_));
 BUFx6f_ASAP7_75t_R _17301_ (.A(_05426_),
    .Y(_05874_));
 OR3x1_ASAP7_75t_R _17302_ (.A(_01259_),
    .B(_05864_),
    .C(_05869_),
    .Y(_05875_));
 XOR2x2_ASAP7_75t_R _17303_ (.A(_01258_),
    .B(_05875_),
    .Y(_05876_));
 AND2x2_ASAP7_75t_R _17304_ (.A(_05874_),
    .B(_05876_),
    .Y(_03787_));
 OR4x1_ASAP7_75t_R _17305_ (.A(_01257_),
    .B(_01258_),
    .C(_01259_),
    .D(_05872_),
    .Y(_05877_));
 OR3x1_ASAP7_75t_R _17306_ (.A(_01258_),
    .B(_01259_),
    .C(_05872_),
    .Y(_05878_));
 NAND2x1_ASAP7_75t_R _17307_ (.A(_01257_),
    .B(_05878_),
    .Y(_05879_));
 AND3x1_ASAP7_75t_R _17308_ (.A(_05841_),
    .B(_05877_),
    .C(_05879_),
    .Y(_03788_));
 OR5x2_ASAP7_75t_R _17309_ (.A(_01257_),
    .B(_01258_),
    .C(_01259_),
    .D(_05864_),
    .E(_05869_),
    .Y(_05880_));
 XOR2x2_ASAP7_75t_R _17310_ (.A(_05845_),
    .B(_05880_),
    .Y(_05881_));
 AND2x2_ASAP7_75t_R _17311_ (.A(_05874_),
    .B(_05881_),
    .Y(_03789_));
 OR3x1_ASAP7_75t_R _17312_ (.A(_01255_),
    .B(_05845_),
    .C(_05877_),
    .Y(_05882_));
 OAI21x1_ASAP7_75t_R _17313_ (.A1(_05845_),
    .A2(_05877_),
    .B(_01255_),
    .Y(_05883_));
 AND3x1_ASAP7_75t_R _17314_ (.A(_05841_),
    .B(_05882_),
    .C(_05883_),
    .Y(_03790_));
 OR3x1_ASAP7_75t_R _17315_ (.A(_01255_),
    .B(_05845_),
    .C(_05880_),
    .Y(_05884_));
 XOR2x2_ASAP7_75t_R _17316_ (.A(_01254_),
    .B(_05884_),
    .Y(_05885_));
 AND2x2_ASAP7_75t_R _17317_ (.A(_05874_),
    .B(_05885_),
    .Y(_03791_));
 NOR2x1_ASAP7_75t_R _17318_ (.A(_05300_),
    .B(_02614_),
    .Y(_03792_));
 OR4x1_ASAP7_75t_R _17319_ (.A(_01254_),
    .B(_01255_),
    .C(_05845_),
    .D(_05877_),
    .Y(_05886_));
 XOR2x2_ASAP7_75t_R _17320_ (.A(_01252_),
    .B(_05886_),
    .Y(_05887_));
 AND2x2_ASAP7_75t_R _17321_ (.A(_05874_),
    .B(_05887_),
    .Y(_03793_));
 OR5x1_ASAP7_75t_R _17322_ (.A(_01252_),
    .B(_01254_),
    .C(_01255_),
    .D(_05845_),
    .E(_05880_),
    .Y(_05888_));
 XOR2x2_ASAP7_75t_R _17323_ (.A(_01251_),
    .B(_05888_),
    .Y(_05889_));
 AND2x2_ASAP7_75t_R _17324_ (.A(_05874_),
    .B(_05889_),
    .Y(_03794_));
 OR5x2_ASAP7_75t_R _17325_ (.A(_01251_),
    .B(_01252_),
    .C(_01254_),
    .D(_01255_),
    .E(_05845_),
    .Y(_05890_));
 OR3x1_ASAP7_75t_R _17326_ (.A(_01250_),
    .B(_05877_),
    .C(_05890_),
    .Y(_05891_));
 OAI21x1_ASAP7_75t_R _17327_ (.A1(_05877_),
    .A2(_05890_),
    .B(_01250_),
    .Y(_05892_));
 AND3x1_ASAP7_75t_R _17328_ (.A(_05841_),
    .B(_05891_),
    .C(_05892_),
    .Y(_03795_));
 OR4x1_ASAP7_75t_R _17329_ (.A(_01249_),
    .B(_01250_),
    .C(_05880_),
    .D(_05890_),
    .Y(_05893_));
 OR3x1_ASAP7_75t_R _17330_ (.A(_01250_),
    .B(_05880_),
    .C(_05890_),
    .Y(_05894_));
 NAND2x1_ASAP7_75t_R _17331_ (.A(_01249_),
    .B(_05894_),
    .Y(_05895_));
 AND3x1_ASAP7_75t_R _17332_ (.A(_05841_),
    .B(_05893_),
    .C(_05895_),
    .Y(_03796_));
 OR4x1_ASAP7_75t_R _17333_ (.A(_01249_),
    .B(_01250_),
    .C(_05877_),
    .D(_05890_),
    .Y(_05896_));
 XOR2x2_ASAP7_75t_R _17334_ (.A(_05850_),
    .B(_05896_),
    .Y(_05897_));
 AND2x2_ASAP7_75t_R _17335_ (.A(_05874_),
    .B(_05897_),
    .Y(_03797_));
 OR3x1_ASAP7_75t_R _17336_ (.A(_01247_),
    .B(_05850_),
    .C(_05893_),
    .Y(_05898_));
 OAI21x1_ASAP7_75t_R _17337_ (.A1(_05850_),
    .A2(_05893_),
    .B(_01247_),
    .Y(_05899_));
 AND3x1_ASAP7_75t_R _17338_ (.A(_05841_),
    .B(_05898_),
    .C(_05899_),
    .Y(_03798_));
 OR3x1_ASAP7_75t_R _17339_ (.A(_01247_),
    .B(_05850_),
    .C(_05896_),
    .Y(_05900_));
 XOR2x2_ASAP7_75t_R _17340_ (.A(_01246_),
    .B(_05900_),
    .Y(_05901_));
 AND2x2_ASAP7_75t_R _17341_ (.A(_05874_),
    .B(_05901_),
    .Y(_03799_));
 OR4x1_ASAP7_75t_R _17342_ (.A(_01246_),
    .B(_01247_),
    .C(_05850_),
    .D(_05893_),
    .Y(_05902_));
 XOR2x2_ASAP7_75t_R _17343_ (.A(_01245_),
    .B(_05902_),
    .Y(_05903_));
 AND2x2_ASAP7_75t_R _17344_ (.A(_05874_),
    .B(_05903_),
    .Y(_03800_));
 OR5x1_ASAP7_75t_R _17345_ (.A(_01245_),
    .B(_01246_),
    .C(_01247_),
    .D(_05850_),
    .E(_05896_),
    .Y(_05904_));
 XOR2x2_ASAP7_75t_R _17346_ (.A(_01244_),
    .B(_05904_),
    .Y(_05905_));
 AND2x2_ASAP7_75t_R _17347_ (.A(_05874_),
    .B(_05905_),
    .Y(_03801_));
 OR5x2_ASAP7_75t_R _17348_ (.A(_01244_),
    .B(_01245_),
    .C(_01246_),
    .D(_01247_),
    .E(_05850_),
    .Y(_05906_));
 OR3x1_ASAP7_75t_R _17349_ (.A(_01243_),
    .B(_05893_),
    .C(_05906_),
    .Y(_05907_));
 OAI21x1_ASAP7_75t_R _17350_ (.A1(_05893_),
    .A2(_05906_),
    .B(_01243_),
    .Y(_05908_));
 AND3x1_ASAP7_75t_R _17351_ (.A(_05841_),
    .B(_05907_),
    .C(_05908_),
    .Y(_03802_));
 XOR2x2_ASAP7_75t_R _17352_ (.A(_01242_),
    .B(_02613_),
    .Y(_05909_));
 AND2x2_ASAP7_75t_R _17353_ (.A(_05874_),
    .B(_05909_),
    .Y(_03803_));
 BUFx6f_ASAP7_75t_R _17354_ (.A(_05426_),
    .Y(_05910_));
 OR3x1_ASAP7_75t_R _17355_ (.A(_01243_),
    .B(_05896_),
    .C(_05906_),
    .Y(_05911_));
 XOR2x2_ASAP7_75t_R _17356_ (.A(_01241_),
    .B(_05911_),
    .Y(_05912_));
 AND2x2_ASAP7_75t_R _17357_ (.A(_05910_),
    .B(_05912_),
    .Y(_03804_));
 OR4x1_ASAP7_75t_R _17358_ (.A(_01241_),
    .B(_01243_),
    .C(_05893_),
    .D(_05906_),
    .Y(_05913_));
 XOR2x2_ASAP7_75t_R _17359_ (.A(_01240_),
    .B(_05913_),
    .Y(_05914_));
 AND2x2_ASAP7_75t_R _17360_ (.A(_05910_),
    .B(_05914_),
    .Y(_03805_));
 OR3x1_ASAP7_75t_R _17361_ (.A(_01242_),
    .B(_01253_),
    .C(_00040_),
    .Y(_05915_));
 XOR2x2_ASAP7_75t_R _17362_ (.A(_01239_),
    .B(_05915_),
    .Y(_05916_));
 AND2x2_ASAP7_75t_R _17363_ (.A(_05910_),
    .B(_05916_),
    .Y(_03806_));
 OR3x1_ASAP7_75t_R _17364_ (.A(_01239_),
    .B(_01242_),
    .C(_02613_),
    .Y(_05917_));
 NAND2x1_ASAP7_75t_R _17365_ (.A(_01238_),
    .B(_05917_),
    .Y(_05918_));
 AND3x1_ASAP7_75t_R _17366_ (.A(_05841_),
    .B(_05858_),
    .C(_05918_),
    .Y(_03807_));
 XOR2x2_ASAP7_75t_R _17367_ (.A(_01237_),
    .B(_05863_),
    .Y(_05919_));
 AND2x2_ASAP7_75t_R _17368_ (.A(_05910_),
    .B(_05919_),
    .Y(_03808_));
 OR3x1_ASAP7_75t_R _17369_ (.A(_01236_),
    .B(_01237_),
    .C(_05858_),
    .Y(_05920_));
 OAI21x1_ASAP7_75t_R _17370_ (.A1(_01237_),
    .A2(_05858_),
    .B(_01236_),
    .Y(_05921_));
 AND3x1_ASAP7_75t_R _17371_ (.A(_05841_),
    .B(_05920_),
    .C(_05921_),
    .Y(_03809_));
 OR3x1_ASAP7_75t_R _17372_ (.A(_01236_),
    .B(_01237_),
    .C(_05863_),
    .Y(_05922_));
 XOR2x2_ASAP7_75t_R _17373_ (.A(_01235_),
    .B(_05922_),
    .Y(_05923_));
 AND2x2_ASAP7_75t_R _17374_ (.A(_05910_),
    .B(_05923_),
    .Y(_03810_));
 BUFx6f_ASAP7_75t_R _17375_ (.A(_05337_),
    .Y(_05924_));
 OR4x1_ASAP7_75t_R _17376_ (.A(_01235_),
    .B(_01236_),
    .C(_01237_),
    .D(_05858_),
    .Y(_05925_));
 NAND2x1_ASAP7_75t_R _17377_ (.A(_01234_),
    .B(_05925_),
    .Y(_05926_));
 AND3x1_ASAP7_75t_R _17378_ (.A(_05924_),
    .B(_05860_),
    .C(_05926_),
    .Y(_03811_));
 XOR2x2_ASAP7_75t_R _17379_ (.A(_05846_),
    .B(_05864_),
    .Y(_05927_));
 AND2x2_ASAP7_75t_R _17380_ (.A(_05910_),
    .B(_05927_),
    .Y(_03812_));
 AND2x2_ASAP7_75t_R _17381_ (.A(_05910_),
    .B(_00019_),
    .Y(_03813_));
 INVx2_ASAP7_75t_R _17382_ (.A(_02065_),
    .Y(_05928_));
 INVx1_ASAP7_75t_R _17383_ (.A(_02071_),
    .Y(_05929_));
 NOR2x1_ASAP7_75t_R _17384_ (.A(_01265_),
    .B(_01266_),
    .Y(_05930_));
 AND5x2_ASAP7_75t_R _17385_ (.A(\xs[13].cli1.i[39] ),
    .B(_01267_),
    .C(\xs[13].cli1.i[33] ),
    .D(_01269_),
    .E(_05930_),
    .Y(_05931_));
 NOR2x1_ASAP7_75t_R _17386_ (.A(_01304_),
    .B(_01305_),
    .Y(_05932_));
 AND3x4_ASAP7_75t_R _17387_ (.A(_01306_),
    .B(\peo[26][33] ),
    .C(_05932_),
    .Y(_05933_));
 NOR2x1_ASAP7_75t_R _17388_ (.A(_01303_),
    .B(_01308_),
    .Y(_05934_));
 AO31x2_ASAP7_75t_R _17389_ (.A1(_01267_),
    .A2(\xs[13].cli1.i[33] ),
    .A3(_05930_),
    .B(_01264_),
    .Y(_05935_));
 AND5x1_ASAP7_75t_R _17390_ (.A(_01306_),
    .B(\peo[26][33] ),
    .C(_05929_),
    .D(_05932_),
    .E(_05934_),
    .Y(_05936_));
 AO32x1_ASAP7_75t_R _17391_ (.A1(_05931_),
    .A2(_05933_),
    .A3(_05934_),
    .B1(_05935_),
    .B2(_05936_),
    .Y(_05937_));
 OA211x2_ASAP7_75t_R _17392_ (.A1(_01303_),
    .A2(_05933_),
    .B(_05931_),
    .C(_02071_),
    .Y(_05938_));
 OR2x6_ASAP7_75t_R _17393_ (.A(_05937_),
    .B(_05938_),
    .Y(_05939_));
 OR4x1_ASAP7_75t_R _17394_ (.A(_02064_),
    .B(_05928_),
    .C(_05929_),
    .D(_05939_),
    .Y(_05940_));
 NOR2x1_ASAP7_75t_R _17395_ (.A(_02075_),
    .B(_05940_),
    .Y(_05941_));
 OR2x2_ASAP7_75t_R _17396_ (.A(_01265_),
    .B(_01266_),
    .Y(_05942_));
 OR5x1_ASAP7_75t_R _17397_ (.A(_01264_),
    .B(\xs[13].cli1.i[34] ),
    .C(_01268_),
    .D(\peo[27][32] ),
    .E(_05942_),
    .Y(_05943_));
 OA31x2_ASAP7_75t_R _17398_ (.A1(\xs[13].cli1.i[34] ),
    .A2(_01268_),
    .A3(_05942_),
    .B1(\xs[13].cli1.i[39] ),
    .Y(_05944_));
 OA21x2_ASAP7_75t_R _17399_ (.A1(_05931_),
    .A2(_05944_),
    .B(_02071_),
    .Y(_05945_));
 AO21x1_ASAP7_75t_R _17400_ (.A1(_05928_),
    .A2(_05931_),
    .B(_02064_),
    .Y(_05946_));
 INVx2_ASAP7_75t_R _17401_ (.A(_02064_),
    .Y(_05947_));
 AO21x1_ASAP7_75t_R _17402_ (.A1(_00019_),
    .A2(_05944_),
    .B(_05947_),
    .Y(_05948_));
 NOR2x1_ASAP7_75t_R _17403_ (.A(_01303_),
    .B(_05933_),
    .Y(_05949_));
 OA211x2_ASAP7_75t_R _17404_ (.A1(_05945_),
    .A2(_05946_),
    .B(_05948_),
    .C(_05949_),
    .Y(_05950_));
 BUFx6f_ASAP7_75t_R _17405_ (.A(_05950_),
    .Y(_05951_));
 OR3x1_ASAP7_75t_R _17406_ (.A(\peo[27][0] ),
    .B(_05943_),
    .C(_05951_),
    .Y(_05952_));
 OAI21x1_ASAP7_75t_R _17407_ (.A1(_05943_),
    .A2(_05951_),
    .B(_01310_),
    .Y(_05953_));
 AND3x1_ASAP7_75t_R _17408_ (.A(_05940_),
    .B(_05952_),
    .C(_05953_),
    .Y(_05954_));
 OA21x2_ASAP7_75t_R _17409_ (.A1(_05941_),
    .A2(_05954_),
    .B(_11397_),
    .Y(_03814_));
 OR2x2_ASAP7_75t_R _17410_ (.A(_08683_),
    .B(_05940_),
    .Y(_05955_));
 BUFx3_ASAP7_75t_R _17411_ (.A(_05955_),
    .Y(_05956_));
 NOR2x1_ASAP7_75t_R _17412_ (.A(_02074_),
    .B(_05956_),
    .Y(_03815_));
 NOR2x1_ASAP7_75t_R _17413_ (.A(_02073_),
    .B(_05956_),
    .Y(_03816_));
 NOR2x1_ASAP7_75t_R _17414_ (.A(_02072_),
    .B(_05956_),
    .Y(_03817_));
 NOR2x1_ASAP7_75t_R _17415_ (.A(_02063_),
    .B(_05956_),
    .Y(_03818_));
 NOR2x1_ASAP7_75t_R _17416_ (.A(_02062_),
    .B(_05956_),
    .Y(_03819_));
 NOR2x1_ASAP7_75t_R _17417_ (.A(_02064_),
    .B(_02065_),
    .Y(_05957_));
 AOI21x1_ASAP7_75t_R _17418_ (.A1(_05944_),
    .A2(_05957_),
    .B(_05951_),
    .Y(_05958_));
 AND2x2_ASAP7_75t_R _17419_ (.A(_05933_),
    .B(_05934_),
    .Y(_05959_));
 AO21x1_ASAP7_75t_R _17420_ (.A1(_05935_),
    .A2(_05959_),
    .B(_02071_),
    .Y(_05960_));
 OR4x1_ASAP7_75t_R _17421_ (.A(_02064_),
    .B(_05928_),
    .C(_05939_),
    .D(_05960_),
    .Y(_05961_));
 AND3x1_ASAP7_75t_R _17422_ (.A(\peo[26][0] ),
    .B(_05958_),
    .C(_05961_),
    .Y(_05962_));
 OAI22x1_ASAP7_75t_R _17423_ (.A1(_01271_),
    .A2(_05958_),
    .B1(_05961_),
    .B2(_02075_),
    .Y(_05963_));
 OA21x2_ASAP7_75t_R _17424_ (.A1(_05962_),
    .A2(_05963_),
    .B(_11397_),
    .Y(_03820_));
 OR2x2_ASAP7_75t_R _17425_ (.A(_08683_),
    .B(_05961_),
    .Y(_05964_));
 BUFx3_ASAP7_75t_R _17426_ (.A(_05964_),
    .Y(_05965_));
 NOR2x1_ASAP7_75t_R _17427_ (.A(_02074_),
    .B(_05965_),
    .Y(_03821_));
 NOR2x1_ASAP7_75t_R _17428_ (.A(_02073_),
    .B(_05965_),
    .Y(_03822_));
 NOR2x1_ASAP7_75t_R _17429_ (.A(_02072_),
    .B(_05965_),
    .Y(_03823_));
 NOR2x1_ASAP7_75t_R _17430_ (.A(_02063_),
    .B(_05965_),
    .Y(_03824_));
 NOR2x1_ASAP7_75t_R _17431_ (.A(_02062_),
    .B(_05965_),
    .Y(_03825_));
 OAI21x1_ASAP7_75t_R _17432_ (.A1(_05928_),
    .A2(_05939_),
    .B(_05947_),
    .Y(_05966_));
 AND2x4_ASAP7_75t_R _17433_ (.A(_08876_),
    .B(_05966_),
    .Y(_05967_));
 OR2x6_ASAP7_75t_R _17434_ (.A(_05935_),
    .B(_05957_),
    .Y(_05968_));
 OR3x1_ASAP7_75t_R _17435_ (.A(\peo[27][0] ),
    .B(_05951_),
    .C(_05968_),
    .Y(_05969_));
 OR2x2_ASAP7_75t_R _17436_ (.A(_05951_),
    .B(_05968_),
    .Y(_05970_));
 BUFx6f_ASAP7_75t_R _17437_ (.A(_05970_),
    .Y(_05971_));
 NAND2x1_ASAP7_75t_R _17438_ (.A(_01310_),
    .B(_05971_),
    .Y(_05972_));
 NOR2x1_ASAP7_75t_R _17439_ (.A(_08765_),
    .B(_05966_),
    .Y(_05973_));
 INVx1_ASAP7_75t_R _17440_ (.A(_02075_),
    .Y(_05974_));
 AO32x1_ASAP7_75t_R _17441_ (.A1(_05967_),
    .A2(_05969_),
    .A3(_05972_),
    .B1(_05973_),
    .B2(_05974_),
    .Y(_03826_));
 OR2x2_ASAP7_75t_R _17442_ (.A(_09220_),
    .B(_05966_),
    .Y(_05975_));
 BUFx6f_ASAP7_75t_R _17443_ (.A(_05975_),
    .Y(_05976_));
 NOR2x1_ASAP7_75t_R _17444_ (.A(_02074_),
    .B(_05976_),
    .Y(_03827_));
 NOR2x1_ASAP7_75t_R _17445_ (.A(_02073_),
    .B(_05976_),
    .Y(_03828_));
 NOR2x1_ASAP7_75t_R _17446_ (.A(_02072_),
    .B(_05976_),
    .Y(_03829_));
 OR3x1_ASAP7_75t_R _17447_ (.A(\peo[27][32] ),
    .B(_05951_),
    .C(_05968_),
    .Y(_05977_));
 NAND2x1_ASAP7_75t_R _17448_ (.A(_01308_),
    .B(_05971_),
    .Y(_05978_));
 AO32x1_ASAP7_75t_R _17449_ (.A1(_05967_),
    .A2(_05977_),
    .A3(_05978_),
    .B1(_05973_),
    .B2(_05929_),
    .Y(_03830_));
 OR3x1_ASAP7_75t_R _17450_ (.A(\xs[13].cli1.i[33] ),
    .B(_05951_),
    .C(_05968_),
    .Y(_05979_));
 NAND2x1_ASAP7_75t_R _17451_ (.A(_01307_),
    .B(_05971_),
    .Y(_05980_));
 INVx1_ASAP7_75t_R _17452_ (.A(_02070_),
    .Y(_05981_));
 AO32x1_ASAP7_75t_R _17453_ (.A1(_05967_),
    .A2(_05979_),
    .A3(_05980_),
    .B1(_05973_),
    .B2(_05981_),
    .Y(_03831_));
 OR3x1_ASAP7_75t_R _17454_ (.A(\xs[13].cli1.i[34] ),
    .B(_05951_),
    .C(_05968_),
    .Y(_05982_));
 NAND2x1_ASAP7_75t_R _17455_ (.A(_01306_),
    .B(_05971_),
    .Y(_05983_));
 INVx1_ASAP7_75t_R _17456_ (.A(_02069_),
    .Y(_05984_));
 AO32x1_ASAP7_75t_R _17457_ (.A1(_05967_),
    .A2(_05982_),
    .A3(_05983_),
    .B1(_05973_),
    .B2(_05984_),
    .Y(_03832_));
 OR3x1_ASAP7_75t_R _17458_ (.A(\xs[13].cli1.i[35] ),
    .B(_05951_),
    .C(_05968_),
    .Y(_05985_));
 NAND2x1_ASAP7_75t_R _17459_ (.A(_01305_),
    .B(_05971_),
    .Y(_05986_));
 INVx1_ASAP7_75t_R _17460_ (.A(_02068_),
    .Y(_05987_));
 AO32x1_ASAP7_75t_R _17461_ (.A1(_05967_),
    .A2(_05985_),
    .A3(_05986_),
    .B1(_05973_),
    .B2(_05987_),
    .Y(_03833_));
 OR3x1_ASAP7_75t_R _17462_ (.A(\xs[13].cli1.i[36] ),
    .B(_05951_),
    .C(_05968_),
    .Y(_05988_));
 NAND2x1_ASAP7_75t_R _17463_ (.A(_01304_),
    .B(_05971_),
    .Y(_05989_));
 INVx1_ASAP7_75t_R _17464_ (.A(_02067_),
    .Y(_05990_));
 AO32x1_ASAP7_75t_R _17465_ (.A1(_05967_),
    .A2(_05988_),
    .A3(_05989_),
    .B1(_05973_),
    .B2(_05990_),
    .Y(_03834_));
 NOR2x1_ASAP7_75t_R _17466_ (.A(_02066_),
    .B(_05976_),
    .Y(_03835_));
 AND4x1_ASAP7_75t_R _17467_ (.A(_08999_),
    .B(_05947_),
    .C(_02065_),
    .D(_05939_),
    .Y(_03836_));
 OA21x2_ASAP7_75t_R _17468_ (.A1(_02071_),
    .A2(_05935_),
    .B(_02065_),
    .Y(_05991_));
 OR3x1_ASAP7_75t_R _17469_ (.A(_05947_),
    .B(_00019_),
    .C(_05935_),
    .Y(_05992_));
 OA211x2_ASAP7_75t_R _17470_ (.A1(_02064_),
    .A2(_05991_),
    .B(_05992_),
    .C(_05949_),
    .Y(_05993_));
 NAND2x1_ASAP7_75t_R _17471_ (.A(_05966_),
    .B(_05971_),
    .Y(_05994_));
 OA21x2_ASAP7_75t_R _17472_ (.A1(_05993_),
    .A2(_05994_),
    .B(_11397_),
    .Y(_03837_));
 NOR2x1_ASAP7_75t_R _17473_ (.A(_02063_),
    .B(_05976_),
    .Y(_03838_));
 NOR2x1_ASAP7_75t_R _17474_ (.A(_02062_),
    .B(_05976_),
    .Y(_03839_));
 BUFx12f_ASAP7_75t_R _17475_ (.A(_11465_),
    .Y(_05995_));
 BUFx3_ASAP7_75t_R _17476_ (.A(_01195_),
    .Y(_05996_));
 BUFx3_ASAP7_75t_R _17477_ (.A(_01168_),
    .Y(_05997_));
 AND4x1_ASAP7_75t_R _17478_ (.A(_05997_),
    .B(_01196_),
    .C(_01197_),
    .D(_01198_),
    .Y(_05998_));
 AND5x1_ASAP7_75t_R _17479_ (.A(_01187_),
    .B(_01192_),
    .C(_01193_),
    .D(_05996_),
    .E(_05998_),
    .Y(_05999_));
 AND5x2_ASAP7_75t_R _17480_ (.A(_01189_),
    .B(_01190_),
    .C(_01191_),
    .D(_05995_),
    .E(_05999_),
    .Y(_06000_));
 AND4x1_ASAP7_75t_R _17481_ (.A(_01182_),
    .B(_01183_),
    .C(_01184_),
    .D(_01185_),
    .Y(_06001_));
 AND4x1_ASAP7_75t_R _17482_ (.A(_01176_),
    .B(_01178_),
    .C(_01179_),
    .D(_01186_),
    .Y(_06002_));
 AND5x1_ASAP7_75t_R _17483_ (.A(_01169_),
    .B(_01170_),
    .C(_01175_),
    .D(_01194_),
    .E(_06002_),
    .Y(_06003_));
 AND3x1_ASAP7_75t_R _17484_ (.A(_01173_),
    .B(_01174_),
    .C(_01177_),
    .Y(_06004_));
 OR3x1_ASAP7_75t_R _17485_ (.A(_01171_),
    .B(_01172_),
    .C(_06004_),
    .Y(_06005_));
 AND5x2_ASAP7_75t_R _17486_ (.A(_01180_),
    .B(_01181_),
    .C(_06001_),
    .D(_06003_),
    .E(_06005_),
    .Y(_06006_));
 NAND2x2_ASAP7_75t_R _17487_ (.A(_06000_),
    .B(_06006_),
    .Y(_06007_));
 NOR2x1_ASAP7_75t_R _17488_ (.A(_01125_),
    .B(_06007_),
    .Y(_03840_));
 INVx1_ASAP7_75t_R _17489_ (.A(_06007_),
    .Y(_03841_));
 NOR2x1_ASAP7_75t_R _17490_ (.A(_01128_),
    .B(_06007_),
    .Y(_03842_));
 NOR2x1_ASAP7_75t_R _17491_ (.A(_01127_),
    .B(_06007_),
    .Y(_03843_));
 NOR2x1_ASAP7_75t_R _17492_ (.A(_01126_),
    .B(_06007_),
    .Y(_03844_));
 NOR2x1_ASAP7_75t_R _17493_ (.A(_01124_),
    .B(_06007_),
    .Y(_03845_));
 NOR2x1_ASAP7_75t_R _17494_ (.A(_01123_),
    .B(_06007_),
    .Y(_03846_));
 INVx1_ASAP7_75t_R _17495_ (.A(_06007_),
    .Y(_03847_));
 AND2x2_ASAP7_75t_R _17496_ (.A(_05910_),
    .B(_00041_),
    .Y(_03848_));
 OR4x1_ASAP7_75t_R _17497_ (.A(_01173_),
    .B(_01174_),
    .C(_01177_),
    .D(_02663_),
    .Y(_06008_));
 OR4x1_ASAP7_75t_R _17498_ (.A(_01169_),
    .B(_01170_),
    .C(_01171_),
    .D(_01172_),
    .Y(_06009_));
 OR2x6_ASAP7_75t_R _17499_ (.A(_06008_),
    .B(_06009_),
    .Y(_06010_));
 OR3x1_ASAP7_75t_R _17500_ (.A(_05997_),
    .B(_01198_),
    .C(_06010_),
    .Y(_06011_));
 OAI21x1_ASAP7_75t_R _17501_ (.A1(_05997_),
    .A2(_06010_),
    .B(_01198_),
    .Y(_06012_));
 AND3x1_ASAP7_75t_R _17502_ (.A(_05924_),
    .B(_06011_),
    .C(_06012_),
    .Y(_03849_));
 OR5x2_ASAP7_75t_R _17503_ (.A(_01173_),
    .B(_01174_),
    .C(_01177_),
    .D(_01188_),
    .E(_00041_),
    .Y(_06013_));
 OR2x2_ASAP7_75t_R _17504_ (.A(_06009_),
    .B(_06013_),
    .Y(_06014_));
 OR3x1_ASAP7_75t_R _17505_ (.A(_05997_),
    .B(_01198_),
    .C(_06014_),
    .Y(_06015_));
 XOR2x2_ASAP7_75t_R _17506_ (.A(_01197_),
    .B(_06015_),
    .Y(_06016_));
 AND2x2_ASAP7_75t_R _17507_ (.A(_05910_),
    .B(_06016_),
    .Y(_03850_));
 OR4x1_ASAP7_75t_R _17508_ (.A(_05997_),
    .B(_01196_),
    .C(_01197_),
    .D(_01198_),
    .Y(_06017_));
 OR3x2_ASAP7_75t_R _17509_ (.A(_06008_),
    .B(_06009_),
    .C(_06017_),
    .Y(_06018_));
 OR4x1_ASAP7_75t_R _17510_ (.A(_05997_),
    .B(_01197_),
    .C(_01198_),
    .D(_06010_),
    .Y(_06019_));
 NAND2x1_ASAP7_75t_R _17511_ (.A(_01196_),
    .B(_06019_),
    .Y(_06020_));
 AND3x1_ASAP7_75t_R _17512_ (.A(_05924_),
    .B(_06018_),
    .C(_06020_),
    .Y(_03851_));
 OR3x2_ASAP7_75t_R _17513_ (.A(_06009_),
    .B(_06013_),
    .C(_06017_),
    .Y(_06021_));
 XOR2x2_ASAP7_75t_R _17514_ (.A(_05996_),
    .B(_06021_),
    .Y(_06022_));
 AND2x2_ASAP7_75t_R _17515_ (.A(_05910_),
    .B(_06022_),
    .Y(_03852_));
 OR3x1_ASAP7_75t_R _17516_ (.A(_01194_),
    .B(_05996_),
    .C(_06018_),
    .Y(_06023_));
 OAI21x1_ASAP7_75t_R _17517_ (.A1(_05996_),
    .A2(_06018_),
    .B(_01194_),
    .Y(_06024_));
 AND3x1_ASAP7_75t_R _17518_ (.A(_05924_),
    .B(_06023_),
    .C(_06024_),
    .Y(_03853_));
 BUFx12f_ASAP7_75t_R _17519_ (.A(_08598_),
    .Y(_06025_));
 BUFx6f_ASAP7_75t_R _17520_ (.A(_06025_),
    .Y(_06026_));
 OR3x1_ASAP7_75t_R _17521_ (.A(_01194_),
    .B(_05996_),
    .C(_06021_),
    .Y(_06027_));
 XOR2x2_ASAP7_75t_R _17522_ (.A(_01193_),
    .B(_06027_),
    .Y(_06028_));
 AND2x2_ASAP7_75t_R _17523_ (.A(_06026_),
    .B(_06028_),
    .Y(_03854_));
 OR4x1_ASAP7_75t_R _17524_ (.A(_01193_),
    .B(_01194_),
    .C(_05996_),
    .D(_06018_),
    .Y(_06029_));
 XOR2x2_ASAP7_75t_R _17525_ (.A(_01192_),
    .B(_06029_),
    .Y(_06030_));
 AND2x2_ASAP7_75t_R _17526_ (.A(_06026_),
    .B(_06030_),
    .Y(_03855_));
 OR5x1_ASAP7_75t_R _17527_ (.A(_01192_),
    .B(_01193_),
    .C(_01194_),
    .D(_05996_),
    .E(_06021_),
    .Y(_06031_));
 XOR2x2_ASAP7_75t_R _17528_ (.A(_01191_),
    .B(_06031_),
    .Y(_06032_));
 AND2x2_ASAP7_75t_R _17529_ (.A(_06026_),
    .B(_06032_),
    .Y(_03856_));
 OR5x2_ASAP7_75t_R _17530_ (.A(_01191_),
    .B(_01192_),
    .C(_01193_),
    .D(_01194_),
    .E(_05996_),
    .Y(_06033_));
 OR3x2_ASAP7_75t_R _17531_ (.A(_01190_),
    .B(_06018_),
    .C(_06033_),
    .Y(_06034_));
 OAI21x1_ASAP7_75t_R _17532_ (.A1(_06018_),
    .A2(_06033_),
    .B(_01190_),
    .Y(_06035_));
 AND3x1_ASAP7_75t_R _17533_ (.A(_05924_),
    .B(_06034_),
    .C(_06035_),
    .Y(_03857_));
 OR3x2_ASAP7_75t_R _17534_ (.A(_01190_),
    .B(_06021_),
    .C(_06033_),
    .Y(_06036_));
 XOR2x2_ASAP7_75t_R _17535_ (.A(_01189_),
    .B(_06036_),
    .Y(_06037_));
 AND2x2_ASAP7_75t_R _17536_ (.A(_06026_),
    .B(_06037_),
    .Y(_03858_));
 NOR2x1_ASAP7_75t_R _17537_ (.A(_05300_),
    .B(_02664_),
    .Y(_03859_));
 OR3x1_ASAP7_75t_R _17538_ (.A(_01187_),
    .B(_01189_),
    .C(_06034_),
    .Y(_06038_));
 OAI21x1_ASAP7_75t_R _17539_ (.A1(_01189_),
    .A2(_06034_),
    .B(_01187_),
    .Y(_06039_));
 AND3x1_ASAP7_75t_R _17540_ (.A(_05924_),
    .B(_06038_),
    .C(_06039_),
    .Y(_03860_));
 OR3x1_ASAP7_75t_R _17541_ (.A(_01187_),
    .B(_01189_),
    .C(_06036_),
    .Y(_06040_));
 XOR2x2_ASAP7_75t_R _17542_ (.A(_01186_),
    .B(_06040_),
    .Y(_06041_));
 AND2x2_ASAP7_75t_R _17543_ (.A(_06026_),
    .B(_06041_),
    .Y(_03861_));
 OR4x1_ASAP7_75t_R _17544_ (.A(_01186_),
    .B(_01187_),
    .C(_01189_),
    .D(_06034_),
    .Y(_06042_));
 XOR2x2_ASAP7_75t_R _17545_ (.A(_01185_),
    .B(_06042_),
    .Y(_06043_));
 AND2x2_ASAP7_75t_R _17546_ (.A(_06026_),
    .B(_06043_),
    .Y(_03862_));
 OR4x1_ASAP7_75t_R _17547_ (.A(_01185_),
    .B(_01186_),
    .C(_01187_),
    .D(_01189_),
    .Y(_06044_));
 OR3x2_ASAP7_75t_R _17548_ (.A(_01184_),
    .B(_06036_),
    .C(_06044_),
    .Y(_06045_));
 OAI21x1_ASAP7_75t_R _17549_ (.A1(_06036_),
    .A2(_06044_),
    .B(_01184_),
    .Y(_06046_));
 AND3x1_ASAP7_75t_R _17550_ (.A(_05924_),
    .B(_06045_),
    .C(_06046_),
    .Y(_03863_));
 OR3x2_ASAP7_75t_R _17551_ (.A(_01184_),
    .B(_06034_),
    .C(_06044_),
    .Y(_06047_));
 XOR2x2_ASAP7_75t_R _17552_ (.A(_01183_),
    .B(_06047_),
    .Y(_06048_));
 AND2x2_ASAP7_75t_R _17553_ (.A(_06026_),
    .B(_06048_),
    .Y(_03864_));
 OR3x1_ASAP7_75t_R _17554_ (.A(_01182_),
    .B(_01183_),
    .C(_06045_),
    .Y(_06049_));
 OAI21x1_ASAP7_75t_R _17555_ (.A1(_01183_),
    .A2(_06045_),
    .B(_01182_),
    .Y(_06050_));
 AND3x1_ASAP7_75t_R _17556_ (.A(_05924_),
    .B(_06049_),
    .C(_06050_),
    .Y(_03865_));
 OR3x1_ASAP7_75t_R _17557_ (.A(_01182_),
    .B(_01183_),
    .C(_06047_),
    .Y(_06051_));
 XOR2x2_ASAP7_75t_R _17558_ (.A(_01181_),
    .B(_06051_),
    .Y(_06052_));
 AND2x2_ASAP7_75t_R _17559_ (.A(_06026_),
    .B(_06052_),
    .Y(_03866_));
 OR4x1_ASAP7_75t_R _17560_ (.A(_01181_),
    .B(_01182_),
    .C(_01183_),
    .D(_06045_),
    .Y(_06053_));
 XOR2x2_ASAP7_75t_R _17561_ (.A(_01180_),
    .B(_06053_),
    .Y(_06054_));
 AND2x2_ASAP7_75t_R _17562_ (.A(_06026_),
    .B(_06054_),
    .Y(_03867_));
 OR4x1_ASAP7_75t_R _17563_ (.A(_01180_),
    .B(_01181_),
    .C(_01182_),
    .D(_01183_),
    .Y(_06055_));
 OR3x1_ASAP7_75t_R _17564_ (.A(_01179_),
    .B(_06047_),
    .C(_06055_),
    .Y(_06056_));
 OAI21x1_ASAP7_75t_R _17565_ (.A1(_06047_),
    .A2(_06055_),
    .B(_01179_),
    .Y(_06057_));
 AND3x1_ASAP7_75t_R _17566_ (.A(_05924_),
    .B(_06056_),
    .C(_06057_),
    .Y(_03868_));
 OR3x1_ASAP7_75t_R _17567_ (.A(_01179_),
    .B(_06045_),
    .C(_06055_),
    .Y(_06058_));
 XOR2x2_ASAP7_75t_R _17568_ (.A(_01178_),
    .B(_06058_),
    .Y(_06059_));
 AND2x2_ASAP7_75t_R _17569_ (.A(_06026_),
    .B(_06059_),
    .Y(_03869_));
 BUFx6f_ASAP7_75t_R _17570_ (.A(_06025_),
    .Y(_06060_));
 XOR2x2_ASAP7_75t_R _17571_ (.A(_01177_),
    .B(_02663_),
    .Y(_06061_));
 AND2x2_ASAP7_75t_R _17572_ (.A(_06060_),
    .B(_06061_),
    .Y(_03870_));
 OR4x1_ASAP7_75t_R _17573_ (.A(_01178_),
    .B(_01179_),
    .C(_06047_),
    .D(_06055_),
    .Y(_06062_));
 XOR2x2_ASAP7_75t_R _17574_ (.A(_01176_),
    .B(_06062_),
    .Y(_06063_));
 AND2x2_ASAP7_75t_R _17575_ (.A(_06060_),
    .B(_06063_),
    .Y(_03871_));
 OR5x1_ASAP7_75t_R _17576_ (.A(_01176_),
    .B(_01178_),
    .C(_01179_),
    .D(_06045_),
    .E(_06055_),
    .Y(_06064_));
 XOR2x2_ASAP7_75t_R _17577_ (.A(_01175_),
    .B(_06064_),
    .Y(_06065_));
 AND2x2_ASAP7_75t_R _17578_ (.A(_06060_),
    .B(_06065_),
    .Y(_03872_));
 OR3x1_ASAP7_75t_R _17579_ (.A(_01177_),
    .B(_01188_),
    .C(_00041_),
    .Y(_06066_));
 XOR2x2_ASAP7_75t_R _17580_ (.A(_01174_),
    .B(_06066_),
    .Y(_06067_));
 AND2x2_ASAP7_75t_R _17581_ (.A(_06060_),
    .B(_06067_),
    .Y(_03873_));
 OR3x1_ASAP7_75t_R _17582_ (.A(_01174_),
    .B(_01177_),
    .C(_02663_),
    .Y(_06068_));
 NAND2x1_ASAP7_75t_R _17583_ (.A(_01173_),
    .B(_06068_),
    .Y(_06069_));
 AND3x1_ASAP7_75t_R _17584_ (.A(_05924_),
    .B(_06008_),
    .C(_06069_),
    .Y(_03874_));
 XOR2x2_ASAP7_75t_R _17585_ (.A(_01172_),
    .B(_06013_),
    .Y(_06070_));
 AND2x2_ASAP7_75t_R _17586_ (.A(_06060_),
    .B(_06070_),
    .Y(_03875_));
 BUFx6f_ASAP7_75t_R _17587_ (.A(_05337_),
    .Y(_06071_));
 OR3x1_ASAP7_75t_R _17588_ (.A(_01171_),
    .B(_01172_),
    .C(_06008_),
    .Y(_06072_));
 OAI21x1_ASAP7_75t_R _17589_ (.A1(_01172_),
    .A2(_06008_),
    .B(_01171_),
    .Y(_06073_));
 AND3x1_ASAP7_75t_R _17590_ (.A(_06071_),
    .B(_06072_),
    .C(_06073_),
    .Y(_03876_));
 OR3x1_ASAP7_75t_R _17591_ (.A(_01171_),
    .B(_01172_),
    .C(_06013_),
    .Y(_06074_));
 XOR2x2_ASAP7_75t_R _17592_ (.A(_01170_),
    .B(_06074_),
    .Y(_06075_));
 AND2x2_ASAP7_75t_R _17593_ (.A(_06060_),
    .B(_06075_),
    .Y(_03877_));
 OR4x1_ASAP7_75t_R _17594_ (.A(_01170_),
    .B(_01171_),
    .C(_01172_),
    .D(_06008_),
    .Y(_06076_));
 NAND2x1_ASAP7_75t_R _17595_ (.A(_01169_),
    .B(_06076_),
    .Y(_06077_));
 AND3x1_ASAP7_75t_R _17596_ (.A(_06071_),
    .B(_06010_),
    .C(_06077_),
    .Y(_03878_));
 XOR2x2_ASAP7_75t_R _17597_ (.A(_05997_),
    .B(_06014_),
    .Y(_06078_));
 AND2x2_ASAP7_75t_R _17598_ (.A(_06060_),
    .B(_06078_),
    .Y(_03879_));
 BUFx6f_ASAP7_75t_R _17599_ (.A(_01152_),
    .Y(_06079_));
 BUFx6f_ASAP7_75t_R _17600_ (.A(_01129_),
    .Y(_06080_));
 AND4x1_ASAP7_75t_R _17601_ (.A(_06080_),
    .B(_01157_),
    .C(_01158_),
    .D(_01159_),
    .Y(_06081_));
 AND5x1_ASAP7_75t_R _17602_ (.A(_01148_),
    .B(_01153_),
    .C(_01154_),
    .D(_01156_),
    .E(_06081_),
    .Y(_06082_));
 AND5x2_ASAP7_75t_R _17603_ (.A(_01150_),
    .B(_01151_),
    .C(_06079_),
    .D(_05995_),
    .E(_06082_),
    .Y(_06083_));
 BUFx6f_ASAP7_75t_R _17604_ (.A(_01144_),
    .Y(_06084_));
 AND4x1_ASAP7_75t_R _17605_ (.A(_01143_),
    .B(_06084_),
    .C(_01145_),
    .D(_01146_),
    .Y(_06085_));
 AND4x1_ASAP7_75t_R _17606_ (.A(_01137_),
    .B(_01139_),
    .C(_01140_),
    .D(_01147_),
    .Y(_06086_));
 AND5x1_ASAP7_75t_R _17607_ (.A(_01130_),
    .B(_01131_),
    .C(_01136_),
    .D(_01155_),
    .E(_06086_),
    .Y(_06087_));
 AND3x1_ASAP7_75t_R _17608_ (.A(_01134_),
    .B(_01135_),
    .C(_01138_),
    .Y(_06088_));
 OR3x1_ASAP7_75t_R _17609_ (.A(_01132_),
    .B(_01133_),
    .C(_06088_),
    .Y(_06089_));
 AND5x2_ASAP7_75t_R _17610_ (.A(_01141_),
    .B(_01142_),
    .C(_06085_),
    .D(_06087_),
    .E(_06089_),
    .Y(_06090_));
 NAND2x2_ASAP7_75t_R _17611_ (.A(_06083_),
    .B(_06090_),
    .Y(_06091_));
 NOR2x1_ASAP7_75t_R _17612_ (.A(_01119_),
    .B(_06091_),
    .Y(_03880_));
 INVx1_ASAP7_75t_R _17613_ (.A(_06091_),
    .Y(_03881_));
 NOR2x1_ASAP7_75t_R _17614_ (.A(_01122_),
    .B(_06091_),
    .Y(_03882_));
 NOR2x1_ASAP7_75t_R _17615_ (.A(_01121_),
    .B(_06091_),
    .Y(_03883_));
 NOR2x1_ASAP7_75t_R _17616_ (.A(_01120_),
    .B(_06091_),
    .Y(_03884_));
 NOR2x1_ASAP7_75t_R _17617_ (.A(_01118_),
    .B(_06091_),
    .Y(_03885_));
 NOR2x1_ASAP7_75t_R _17618_ (.A(_01117_),
    .B(_06091_),
    .Y(_03886_));
 INVx1_ASAP7_75t_R _17619_ (.A(_06091_),
    .Y(_03887_));
 AND2x2_ASAP7_75t_R _17620_ (.A(_06060_),
    .B(_00042_),
    .Y(_03888_));
 OR4x1_ASAP7_75t_R _17621_ (.A(_01134_),
    .B(_01135_),
    .C(_01138_),
    .D(_02633_),
    .Y(_06092_));
 OR4x1_ASAP7_75t_R _17622_ (.A(_01130_),
    .B(_01131_),
    .C(_01132_),
    .D(_01133_),
    .Y(_06093_));
 OR2x6_ASAP7_75t_R _17623_ (.A(_06092_),
    .B(_06093_),
    .Y(_06094_));
 OR3x1_ASAP7_75t_R _17624_ (.A(_06080_),
    .B(_01159_),
    .C(_06094_),
    .Y(_06095_));
 OAI21x1_ASAP7_75t_R _17625_ (.A1(_06080_),
    .A2(_06094_),
    .B(_01159_),
    .Y(_06096_));
 AND3x1_ASAP7_75t_R _17626_ (.A(_06071_),
    .B(_06095_),
    .C(_06096_),
    .Y(_03889_));
 OR5x2_ASAP7_75t_R _17627_ (.A(_01134_),
    .B(_01135_),
    .C(_01138_),
    .D(_01149_),
    .E(_00042_),
    .Y(_06097_));
 OR2x6_ASAP7_75t_R _17628_ (.A(_06093_),
    .B(_06097_),
    .Y(_06098_));
 OR3x1_ASAP7_75t_R _17629_ (.A(_06080_),
    .B(_01159_),
    .C(_06098_),
    .Y(_06099_));
 XOR2x2_ASAP7_75t_R _17630_ (.A(_01158_),
    .B(_06099_),
    .Y(_06100_));
 AND2x2_ASAP7_75t_R _17631_ (.A(_06060_),
    .B(_06100_),
    .Y(_03890_));
 OR4x1_ASAP7_75t_R _17632_ (.A(_06080_),
    .B(_01158_),
    .C(_01159_),
    .D(_06094_),
    .Y(_06101_));
 XOR2x2_ASAP7_75t_R _17633_ (.A(_01157_),
    .B(_06101_),
    .Y(_06102_));
 AND2x2_ASAP7_75t_R _17634_ (.A(_06060_),
    .B(_06102_),
    .Y(_03891_));
 OR5x2_ASAP7_75t_R _17635_ (.A(_06080_),
    .B(_01156_),
    .C(_01157_),
    .D(_01158_),
    .E(_01159_),
    .Y(_06103_));
 OR5x1_ASAP7_75t_R _17636_ (.A(_06080_),
    .B(_01157_),
    .C(_01158_),
    .D(_01159_),
    .E(_06098_),
    .Y(_06104_));
 NAND2x1_ASAP7_75t_R _17637_ (.A(_01156_),
    .B(_06104_),
    .Y(_06105_));
 OA211x2_ASAP7_75t_R _17638_ (.A1(_06098_),
    .A2(_06103_),
    .B(_06105_),
    .C(_11589_),
    .Y(_03892_));
 BUFx6f_ASAP7_75t_R _17639_ (.A(_06025_),
    .Y(_06106_));
 OR3x2_ASAP7_75t_R _17640_ (.A(_06092_),
    .B(_06093_),
    .C(_06103_),
    .Y(_06107_));
 XOR2x2_ASAP7_75t_R _17641_ (.A(_01155_),
    .B(_06107_),
    .Y(_06108_));
 AND2x2_ASAP7_75t_R _17642_ (.A(_06106_),
    .B(_06108_),
    .Y(_03893_));
 OR3x1_ASAP7_75t_R _17643_ (.A(_01155_),
    .B(_06098_),
    .C(_06103_),
    .Y(_06109_));
 XOR2x2_ASAP7_75t_R _17644_ (.A(_01154_),
    .B(_06109_),
    .Y(_06110_));
 AND2x2_ASAP7_75t_R _17645_ (.A(_06106_),
    .B(_06110_),
    .Y(_03894_));
 OR4x1_ASAP7_75t_R _17646_ (.A(_01153_),
    .B(_01154_),
    .C(_01155_),
    .D(_06107_),
    .Y(_06111_));
 OR3x1_ASAP7_75t_R _17647_ (.A(_01154_),
    .B(_01155_),
    .C(_06107_),
    .Y(_06112_));
 NAND2x1_ASAP7_75t_R _17648_ (.A(_01153_),
    .B(_06112_),
    .Y(_06113_));
 AND3x1_ASAP7_75t_R _17649_ (.A(_06071_),
    .B(_06111_),
    .C(_06113_),
    .Y(_03895_));
 OR5x2_ASAP7_75t_R _17650_ (.A(_01153_),
    .B(_01154_),
    .C(_01155_),
    .D(_06098_),
    .E(_06103_),
    .Y(_06114_));
 XOR2x2_ASAP7_75t_R _17651_ (.A(_06079_),
    .B(_06114_),
    .Y(_06115_));
 AND2x2_ASAP7_75t_R _17652_ (.A(_06106_),
    .B(_06115_),
    .Y(_03896_));
 OR3x1_ASAP7_75t_R _17653_ (.A(_01151_),
    .B(_06079_),
    .C(_06111_),
    .Y(_06116_));
 OAI21x1_ASAP7_75t_R _17654_ (.A1(_06079_),
    .A2(_06111_),
    .B(_01151_),
    .Y(_06117_));
 AND3x1_ASAP7_75t_R _17655_ (.A(_06071_),
    .B(_06116_),
    .C(_06117_),
    .Y(_03897_));
 OR3x1_ASAP7_75t_R _17656_ (.A(_01151_),
    .B(_06079_),
    .C(_06114_),
    .Y(_06118_));
 XOR2x2_ASAP7_75t_R _17657_ (.A(_01150_),
    .B(_06118_),
    .Y(_06119_));
 AND2x2_ASAP7_75t_R _17658_ (.A(_06106_),
    .B(_06119_),
    .Y(_03898_));
 NOR2x1_ASAP7_75t_R _17659_ (.A(_05300_),
    .B(_02634_),
    .Y(_03899_));
 OR4x1_ASAP7_75t_R _17660_ (.A(_01150_),
    .B(_01151_),
    .C(_06079_),
    .D(_06111_),
    .Y(_06120_));
 XOR2x2_ASAP7_75t_R _17661_ (.A(_01148_),
    .B(_06120_),
    .Y(_06121_));
 AND2x2_ASAP7_75t_R _17662_ (.A(_06106_),
    .B(_06121_),
    .Y(_03900_));
 OR5x1_ASAP7_75t_R _17663_ (.A(_01148_),
    .B(_01150_),
    .C(_01151_),
    .D(_06079_),
    .E(_06114_),
    .Y(_06122_));
 XOR2x2_ASAP7_75t_R _17664_ (.A(_01147_),
    .B(_06122_),
    .Y(_06123_));
 AND2x2_ASAP7_75t_R _17665_ (.A(_06106_),
    .B(_06123_),
    .Y(_03901_));
 OR5x2_ASAP7_75t_R _17666_ (.A(_01147_),
    .B(_01148_),
    .C(_01150_),
    .D(_01151_),
    .E(_06079_),
    .Y(_06124_));
 OR3x1_ASAP7_75t_R _17667_ (.A(_01146_),
    .B(_06111_),
    .C(_06124_),
    .Y(_06125_));
 OAI21x1_ASAP7_75t_R _17668_ (.A1(_06111_),
    .A2(_06124_),
    .B(_01146_),
    .Y(_06126_));
 AND3x1_ASAP7_75t_R _17669_ (.A(_06071_),
    .B(_06125_),
    .C(_06126_),
    .Y(_03902_));
 OR4x1_ASAP7_75t_R _17670_ (.A(_01145_),
    .B(_01146_),
    .C(_06114_),
    .D(_06124_),
    .Y(_06127_));
 OR3x1_ASAP7_75t_R _17671_ (.A(_01146_),
    .B(_06114_),
    .C(_06124_),
    .Y(_06128_));
 NAND2x1_ASAP7_75t_R _17672_ (.A(_01145_),
    .B(_06128_),
    .Y(_06129_));
 AND3x1_ASAP7_75t_R _17673_ (.A(_06071_),
    .B(_06127_),
    .C(_06129_),
    .Y(_03903_));
 OR4x1_ASAP7_75t_R _17674_ (.A(_01145_),
    .B(_01146_),
    .C(_06111_),
    .D(_06124_),
    .Y(_06130_));
 XOR2x2_ASAP7_75t_R _17675_ (.A(_06084_),
    .B(_06130_),
    .Y(_06131_));
 AND2x2_ASAP7_75t_R _17676_ (.A(_06106_),
    .B(_06131_),
    .Y(_03904_));
 OR3x1_ASAP7_75t_R _17677_ (.A(_01143_),
    .B(_06084_),
    .C(_06127_),
    .Y(_06132_));
 OAI21x1_ASAP7_75t_R _17678_ (.A1(_06084_),
    .A2(_06127_),
    .B(_01143_),
    .Y(_06133_));
 AND3x1_ASAP7_75t_R _17679_ (.A(_06071_),
    .B(_06132_),
    .C(_06133_),
    .Y(_03905_));
 OR3x1_ASAP7_75t_R _17680_ (.A(_01143_),
    .B(_06084_),
    .C(_06130_),
    .Y(_06134_));
 XOR2x2_ASAP7_75t_R _17681_ (.A(_01142_),
    .B(_06134_),
    .Y(_06135_));
 AND2x2_ASAP7_75t_R _17682_ (.A(_06106_),
    .B(_06135_),
    .Y(_03906_));
 OR4x1_ASAP7_75t_R _17683_ (.A(_01142_),
    .B(_01143_),
    .C(_06084_),
    .D(_06127_),
    .Y(_06136_));
 XOR2x2_ASAP7_75t_R _17684_ (.A(_01141_),
    .B(_06136_),
    .Y(_06137_));
 AND2x2_ASAP7_75t_R _17685_ (.A(_06106_),
    .B(_06137_),
    .Y(_03907_));
 OR5x1_ASAP7_75t_R _17686_ (.A(_01141_),
    .B(_01142_),
    .C(_01143_),
    .D(_06084_),
    .E(_06130_),
    .Y(_06138_));
 XOR2x2_ASAP7_75t_R _17687_ (.A(_01140_),
    .B(_06138_),
    .Y(_06139_));
 AND2x2_ASAP7_75t_R _17688_ (.A(_06106_),
    .B(_06139_),
    .Y(_03908_));
 OR5x2_ASAP7_75t_R _17689_ (.A(_01140_),
    .B(_01141_),
    .C(_01142_),
    .D(_01143_),
    .E(_06084_),
    .Y(_06140_));
 OR3x1_ASAP7_75t_R _17690_ (.A(_01139_),
    .B(_06127_),
    .C(_06140_),
    .Y(_06141_));
 OAI21x1_ASAP7_75t_R _17691_ (.A1(_06127_),
    .A2(_06140_),
    .B(_01139_),
    .Y(_06142_));
 AND3x1_ASAP7_75t_R _17692_ (.A(_06071_),
    .B(_06141_),
    .C(_06142_),
    .Y(_03909_));
 BUFx6f_ASAP7_75t_R _17693_ (.A(_06025_),
    .Y(_06143_));
 XOR2x2_ASAP7_75t_R _17694_ (.A(_01138_),
    .B(_02633_),
    .Y(_06144_));
 AND2x2_ASAP7_75t_R _17695_ (.A(_06143_),
    .B(_06144_),
    .Y(_03910_));
 OR3x1_ASAP7_75t_R _17696_ (.A(_01139_),
    .B(_06130_),
    .C(_06140_),
    .Y(_06145_));
 XOR2x2_ASAP7_75t_R _17697_ (.A(_01137_),
    .B(_06145_),
    .Y(_06146_));
 AND2x2_ASAP7_75t_R _17698_ (.A(_06143_),
    .B(_06146_),
    .Y(_03911_));
 OR4x1_ASAP7_75t_R _17699_ (.A(_01137_),
    .B(_01139_),
    .C(_06127_),
    .D(_06140_),
    .Y(_06147_));
 XOR2x2_ASAP7_75t_R _17700_ (.A(_01136_),
    .B(_06147_),
    .Y(_06148_));
 AND2x2_ASAP7_75t_R _17701_ (.A(_06143_),
    .B(_06148_),
    .Y(_03912_));
 OR3x1_ASAP7_75t_R _17702_ (.A(_01138_),
    .B(_01149_),
    .C(_00042_),
    .Y(_06149_));
 XOR2x2_ASAP7_75t_R _17703_ (.A(_01135_),
    .B(_06149_),
    .Y(_06150_));
 AND2x2_ASAP7_75t_R _17704_ (.A(_06143_),
    .B(_06150_),
    .Y(_03913_));
 OR3x1_ASAP7_75t_R _17705_ (.A(_01135_),
    .B(_01138_),
    .C(_02633_),
    .Y(_06151_));
 NAND2x1_ASAP7_75t_R _17706_ (.A(_01134_),
    .B(_06151_),
    .Y(_06152_));
 AND3x1_ASAP7_75t_R _17707_ (.A(_06071_),
    .B(_06092_),
    .C(_06152_),
    .Y(_03914_));
 XOR2x2_ASAP7_75t_R _17708_ (.A(_01133_),
    .B(_06097_),
    .Y(_06153_));
 AND2x2_ASAP7_75t_R _17709_ (.A(_06143_),
    .B(_06153_),
    .Y(_03915_));
 BUFx6f_ASAP7_75t_R _17710_ (.A(_05337_),
    .Y(_06154_));
 OR3x1_ASAP7_75t_R _17711_ (.A(_01132_),
    .B(_01133_),
    .C(_06092_),
    .Y(_06155_));
 OAI21x1_ASAP7_75t_R _17712_ (.A1(_01133_),
    .A2(_06092_),
    .B(_01132_),
    .Y(_06156_));
 AND3x1_ASAP7_75t_R _17713_ (.A(_06154_),
    .B(_06155_),
    .C(_06156_),
    .Y(_03916_));
 OR3x1_ASAP7_75t_R _17714_ (.A(_01132_),
    .B(_01133_),
    .C(_06097_),
    .Y(_06157_));
 XOR2x2_ASAP7_75t_R _17715_ (.A(_01131_),
    .B(_06157_),
    .Y(_06158_));
 AND2x2_ASAP7_75t_R _17716_ (.A(_06143_),
    .B(_06158_),
    .Y(_03917_));
 OR4x1_ASAP7_75t_R _17717_ (.A(_01131_),
    .B(_01132_),
    .C(_01133_),
    .D(_06092_),
    .Y(_06159_));
 NAND2x1_ASAP7_75t_R _17718_ (.A(_01130_),
    .B(_06159_),
    .Y(_06160_));
 AND3x1_ASAP7_75t_R _17719_ (.A(_06154_),
    .B(_06094_),
    .C(_06160_),
    .Y(_03918_));
 XOR2x2_ASAP7_75t_R _17720_ (.A(_06080_),
    .B(_06098_),
    .Y(_06161_));
 AND2x2_ASAP7_75t_R _17721_ (.A(_06143_),
    .B(_06161_),
    .Y(_03919_));
 AND2x2_ASAP7_75t_R _17722_ (.A(_06143_),
    .B(_00020_),
    .Y(_03920_));
 OR2x6_ASAP7_75t_R _17723_ (.A(_01161_),
    .B(_01163_),
    .Y(_06162_));
 OR5x2_ASAP7_75t_R _17724_ (.A(_01160_),
    .B(_01162_),
    .C(\xs[14].cli1.i[33] ),
    .D(\peo[29][32] ),
    .E(_06162_),
    .Y(_06163_));
 INVx1_ASAP7_75t_R _17725_ (.A(_02037_),
    .Y(_06164_));
 BUFx6f_ASAP7_75t_R _17726_ (.A(_02043_),
    .Y(_06165_));
 OR4x1_ASAP7_75t_R _17727_ (.A(_01200_),
    .B(_01201_),
    .C(_01202_),
    .D(\peo[28][33] ),
    .Y(_06166_));
 AND2x2_ASAP7_75t_R _17728_ (.A(\peo[28][39] ),
    .B(_06166_),
    .Y(_06167_));
 BUFx6f_ASAP7_75t_R _17729_ (.A(_02036_),
    .Y(_06168_));
 INVx2_ASAP7_75t_R _17730_ (.A(_06168_),
    .Y(_06169_));
 OA211x2_ASAP7_75t_R _17731_ (.A1(_06164_),
    .A2(_06165_),
    .B(_06167_),
    .C(_06169_),
    .Y(_06170_));
 NOR2x1_ASAP7_75t_R _17732_ (.A(_06163_),
    .B(_06170_),
    .Y(_06171_));
 OA31x2_ASAP7_75t_R _17733_ (.A1(_01162_),
    .A2(\xs[14].cli1.i[33] ),
    .A3(_06162_),
    .B1(\xs[14].cli1.i[39] ),
    .Y(_06172_));
 OA21x2_ASAP7_75t_R _17734_ (.A1(_06165_),
    .A2(_06172_),
    .B(_06163_),
    .Y(_06173_));
 INVx2_ASAP7_75t_R _17735_ (.A(_06165_),
    .Y(_06174_));
 OA21x2_ASAP7_75t_R _17736_ (.A1(_01199_),
    .A2(_01204_),
    .B(_06174_),
    .Y(_06175_));
 AO21x2_ASAP7_75t_R _17737_ (.A1(\peo[28][39] ),
    .A2(_06166_),
    .B(_06175_),
    .Y(_06176_));
 AND2x2_ASAP7_75t_R _17738_ (.A(_06169_),
    .B(_02037_),
    .Y(_06177_));
 OA21x2_ASAP7_75t_R _17739_ (.A1(_06173_),
    .A2(_06176_),
    .B(_06177_),
    .Y(_06178_));
 AND3x1_ASAP7_75t_R _17740_ (.A(_06165_),
    .B(_02047_),
    .C(_06178_),
    .Y(_06179_));
 OAI21x1_ASAP7_75t_R _17741_ (.A1(_06173_),
    .A2(_06176_),
    .B(_06177_),
    .Y(_06180_));
 OA21x2_ASAP7_75t_R _17742_ (.A1(_06174_),
    .A2(_06180_),
    .B(_01206_),
    .Y(_06181_));
 OR4x1_ASAP7_75t_R _17743_ (.A(_09221_),
    .B(_06171_),
    .C(_06179_),
    .D(_06181_),
    .Y(_06182_));
 OR4x1_ASAP7_75t_R _17744_ (.A(_09223_),
    .B(_01167_),
    .C(_06163_),
    .D(_06170_),
    .Y(_06183_));
 NAND2x1_ASAP7_75t_R _17745_ (.A(_06182_),
    .B(_06183_),
    .Y(_03921_));
 OR3x2_ASAP7_75t_R _17746_ (.A(_10763_),
    .B(_06174_),
    .C(_06180_),
    .Y(_06184_));
 NOR2x1_ASAP7_75t_R _17747_ (.A(_02046_),
    .B(_06184_),
    .Y(_03922_));
 NOR2x1_ASAP7_75t_R _17748_ (.A(_02045_),
    .B(_06184_),
    .Y(_03923_));
 NOR2x1_ASAP7_75t_R _17749_ (.A(_02044_),
    .B(_06184_),
    .Y(_03924_));
 NOR2x1_ASAP7_75t_R _17750_ (.A(_02035_),
    .B(_06184_),
    .Y(_03925_));
 NOR2x1_ASAP7_75t_R _17751_ (.A(_02034_),
    .B(_06184_),
    .Y(_03926_));
 OR3x1_ASAP7_75t_R _17752_ (.A(_01162_),
    .B(\xs[14].cli1.i[33] ),
    .C(_06162_),
    .Y(_06185_));
 AND2x2_ASAP7_75t_R _17753_ (.A(_06168_),
    .B(_00020_),
    .Y(_06186_));
 NOR2x1_ASAP7_75t_R _17754_ (.A(_01200_),
    .B(_01201_),
    .Y(_06187_));
 AO31x2_ASAP7_75t_R _17755_ (.A1(\peo[28][34] ),
    .A2(_01203_),
    .A3(_06187_),
    .B(_01199_),
    .Y(_06188_));
 OAI21x1_ASAP7_75t_R _17756_ (.A1(_06174_),
    .A2(_06188_),
    .B(_02037_),
    .Y(_06189_));
 AO32x1_ASAP7_75t_R _17757_ (.A1(\peo[28][39] ),
    .A2(_06166_),
    .A3(_06186_),
    .B1(_06189_),
    .B2(_06169_),
    .Y(_06190_));
 INVx1_ASAP7_75t_R _17758_ (.A(_06163_),
    .Y(_06191_));
 AO32x2_ASAP7_75t_R _17759_ (.A1(\xs[14].cli1.i[39] ),
    .A2(_06185_),
    .A3(_06190_),
    .B1(_06170_),
    .B2(_06191_),
    .Y(_06192_));
 NAND2x1_ASAP7_75t_R _17760_ (.A(\peo[29][0] ),
    .B(_06192_),
    .Y(_06193_));
 AND3x1_ASAP7_75t_R _17761_ (.A(_06174_),
    .B(_02047_),
    .C(_06178_),
    .Y(_06194_));
 OA21x2_ASAP7_75t_R _17762_ (.A1(_06165_),
    .A2(_06180_),
    .B(_01206_),
    .Y(_06195_));
 OR3x1_ASAP7_75t_R _17763_ (.A(_06192_),
    .B(_06194_),
    .C(_06195_),
    .Y(_06196_));
 AOI21x1_ASAP7_75t_R _17764_ (.A1(_06193_),
    .A2(_06196_),
    .B(_09081_),
    .Y(_03927_));
 OR3x2_ASAP7_75t_R _17765_ (.A(_10763_),
    .B(_06165_),
    .C(_06180_),
    .Y(_06197_));
 NOR2x1_ASAP7_75t_R _17766_ (.A(_02046_),
    .B(_06197_),
    .Y(_03928_));
 NOR2x1_ASAP7_75t_R _17767_ (.A(_02045_),
    .B(_06197_),
    .Y(_03929_));
 NOR2x1_ASAP7_75t_R _17768_ (.A(_02044_),
    .B(_06197_),
    .Y(_03930_));
 NOR2x1_ASAP7_75t_R _17769_ (.A(_02035_),
    .B(_06197_),
    .Y(_03931_));
 NOR2x1_ASAP7_75t_R _17770_ (.A(_02034_),
    .B(_06197_),
    .Y(_03932_));
 NAND2x1_ASAP7_75t_R _17771_ (.A(\xs[14].cli1.i[39] ),
    .B(_06185_),
    .Y(_06198_));
 AO221x1_ASAP7_75t_R _17772_ (.A1(_06169_),
    .A2(_06189_),
    .B1(_06186_),
    .B2(_06167_),
    .C(_06198_),
    .Y(_06199_));
 BUFx6f_ASAP7_75t_R _17773_ (.A(_06199_),
    .Y(_06200_));
 OR2x2_ASAP7_75t_R _17774_ (.A(\peo[29][0] ),
    .B(_06200_),
    .Y(_06201_));
 NAND2x1_ASAP7_75t_R _17775_ (.A(_01206_),
    .B(_06200_),
    .Y(_06202_));
 OA21x2_ASAP7_75t_R _17776_ (.A1(_06173_),
    .A2(_06176_),
    .B(_02037_),
    .Y(_06203_));
 NOR2x2_ASAP7_75t_R _17777_ (.A(_06168_),
    .B(_06203_),
    .Y(_06204_));
 NOR2x1_ASAP7_75t_R _17778_ (.A(_09223_),
    .B(_06204_),
    .Y(_06205_));
 BUFx12f_ASAP7_75t_R _17779_ (.A(_08578_),
    .Y(_06206_));
 NOR2x1_ASAP7_75t_R _17780_ (.A(_06206_),
    .B(_02047_),
    .Y(_06207_));
 AO32x1_ASAP7_75t_R _17781_ (.A1(_06201_),
    .A2(_06202_),
    .A3(_06205_),
    .B1(_06207_),
    .B2(_06204_),
    .Y(_03933_));
 OR3x1_ASAP7_75t_R _17782_ (.A(_08578_),
    .B(_06168_),
    .C(_06203_),
    .Y(_06208_));
 BUFx6f_ASAP7_75t_R _17783_ (.A(_06208_),
    .Y(_06209_));
 NOR2x1_ASAP7_75t_R _17784_ (.A(_02046_),
    .B(_06209_),
    .Y(_03934_));
 NOR2x1_ASAP7_75t_R _17785_ (.A(_02045_),
    .B(_06209_),
    .Y(_03935_));
 NOR2x1_ASAP7_75t_R _17786_ (.A(_02044_),
    .B(_06209_),
    .Y(_03936_));
 OR2x2_ASAP7_75t_R _17787_ (.A(\peo[29][32] ),
    .B(_06200_),
    .Y(_06210_));
 NAND2x1_ASAP7_75t_R _17788_ (.A(_01204_),
    .B(_06200_),
    .Y(_06211_));
 NOR2x1_ASAP7_75t_R _17789_ (.A(_06206_),
    .B(_06165_),
    .Y(_06212_));
 AO32x1_ASAP7_75t_R _17790_ (.A1(_06205_),
    .A2(_06210_),
    .A3(_06211_),
    .B1(_06212_),
    .B2(_06204_),
    .Y(_03937_));
 OR2x2_ASAP7_75t_R _17791_ (.A(\xs[14].cli1.i[33] ),
    .B(_06200_),
    .Y(_06213_));
 NAND2x1_ASAP7_75t_R _17792_ (.A(_01203_),
    .B(_06200_),
    .Y(_06214_));
 NOR2x1_ASAP7_75t_R _17793_ (.A(_06206_),
    .B(_02042_),
    .Y(_06215_));
 AO32x1_ASAP7_75t_R _17794_ (.A1(_06205_),
    .A2(_06213_),
    .A3(_06214_),
    .B1(_06215_),
    .B2(_06204_),
    .Y(_03938_));
 NOR3x1_ASAP7_75t_R _17795_ (.A(_01160_),
    .B(_06192_),
    .C(_06204_),
    .Y(_06216_));
 OA211x2_ASAP7_75t_R _17796_ (.A1(_06168_),
    .A2(_06203_),
    .B(_06200_),
    .C(_01202_),
    .Y(_06217_));
 AO21x1_ASAP7_75t_R _17797_ (.A1(_02041_),
    .A2(_06204_),
    .B(_06217_),
    .Y(_06218_));
 AOI211x1_ASAP7_75t_R _17798_ (.A1(_01163_),
    .A2(_06216_),
    .B(_06218_),
    .C(_09145_),
    .Y(_03939_));
 OA211x2_ASAP7_75t_R _17799_ (.A1(_06168_),
    .A2(_06203_),
    .B(_06200_),
    .C(_01201_),
    .Y(_06219_));
 AO21x1_ASAP7_75t_R _17800_ (.A1(_02040_),
    .A2(_06204_),
    .B(_06219_),
    .Y(_06220_));
 AOI211x1_ASAP7_75t_R _17801_ (.A1(_01162_),
    .A2(_06216_),
    .B(_06220_),
    .C(_09145_),
    .Y(_03940_));
 OA211x2_ASAP7_75t_R _17802_ (.A1(_06168_),
    .A2(_06203_),
    .B(_06200_),
    .C(_01200_),
    .Y(_06221_));
 AO21x1_ASAP7_75t_R _17803_ (.A1(_02039_),
    .A2(_06204_),
    .B(_06221_),
    .Y(_06222_));
 AOI211x1_ASAP7_75t_R _17804_ (.A1(_01161_),
    .A2(_06216_),
    .B(_06222_),
    .C(_09145_),
    .Y(_03941_));
 NOR2x1_ASAP7_75t_R _17805_ (.A(_02038_),
    .B(_06209_),
    .Y(_03942_));
 OR5x1_ASAP7_75t_R _17806_ (.A(_08684_),
    .B(_06168_),
    .C(_06164_),
    .D(_06173_),
    .E(_06176_),
    .Y(_06223_));
 INVx1_ASAP7_75t_R _17807_ (.A(_06223_),
    .Y(_03943_));
 NOR2x1_ASAP7_75t_R _17808_ (.A(\peo[28][32] ),
    .B(_06166_),
    .Y(_06224_));
 OR4x1_ASAP7_75t_R _17809_ (.A(_01199_),
    .B(_06165_),
    .C(_06198_),
    .D(_06224_),
    .Y(_06225_));
 AO21x1_ASAP7_75t_R _17810_ (.A1(_02037_),
    .A2(_06225_),
    .B(_06168_),
    .Y(_06226_));
 OR3x1_ASAP7_75t_R _17811_ (.A(_06169_),
    .B(_00020_),
    .C(_06198_),
    .Y(_06227_));
 AND3x1_ASAP7_75t_R _17812_ (.A(_06167_),
    .B(_06226_),
    .C(_06227_),
    .Y(_06228_));
 NOR2x1_ASAP7_75t_R _17813_ (.A(_06198_),
    .B(_06190_),
    .Y(_06229_));
 OR2x2_ASAP7_75t_R _17814_ (.A(_06204_),
    .B(_06229_),
    .Y(_06230_));
 OA21x2_ASAP7_75t_R _17815_ (.A1(_06228_),
    .A2(_06230_),
    .B(_11397_),
    .Y(_03944_));
 NOR2x1_ASAP7_75t_R _17816_ (.A(_02035_),
    .B(_06209_),
    .Y(_03945_));
 NOR2x1_ASAP7_75t_R _17817_ (.A(_02034_),
    .B(_06209_),
    .Y(_03946_));
 BUFx6f_ASAP7_75t_R _17818_ (.A(_01091_),
    .Y(_06231_));
 BUFx3_ASAP7_75t_R _17819_ (.A(_01064_),
    .Y(_06232_));
 AND4x1_ASAP7_75t_R _17820_ (.A(_06232_),
    .B(_01092_),
    .C(_01093_),
    .D(_01094_),
    .Y(_06233_));
 AND5x1_ASAP7_75t_R _17821_ (.A(_01083_),
    .B(_01088_),
    .C(_01089_),
    .D(_06231_),
    .E(_06233_),
    .Y(_06234_));
 AND5x2_ASAP7_75t_R _17822_ (.A(_01085_),
    .B(_01086_),
    .C(_01087_),
    .D(_05995_),
    .E(_06234_),
    .Y(_06235_));
 AND4x1_ASAP7_75t_R _17823_ (.A(_01078_),
    .B(_01079_),
    .C(_01080_),
    .D(_01081_),
    .Y(_06236_));
 AND4x1_ASAP7_75t_R _17824_ (.A(_01072_),
    .B(_01074_),
    .C(_01075_),
    .D(_01082_),
    .Y(_06237_));
 AND5x1_ASAP7_75t_R _17825_ (.A(_01065_),
    .B(_01066_),
    .C(_01071_),
    .D(_01090_),
    .E(_06237_),
    .Y(_06238_));
 AND3x1_ASAP7_75t_R _17826_ (.A(_01069_),
    .B(_01070_),
    .C(_01073_),
    .Y(_06239_));
 OR3x1_ASAP7_75t_R _17827_ (.A(_01067_),
    .B(_01068_),
    .C(_06239_),
    .Y(_06240_));
 AND5x2_ASAP7_75t_R _17828_ (.A(_01076_),
    .B(_01077_),
    .C(_06236_),
    .D(_06238_),
    .E(_06240_),
    .Y(_06241_));
 NAND2x2_ASAP7_75t_R _17829_ (.A(_06235_),
    .B(_06241_),
    .Y(_06242_));
 NOR2x1_ASAP7_75t_R _17830_ (.A(_01021_),
    .B(_06242_),
    .Y(_03947_));
 INVx1_ASAP7_75t_R _17831_ (.A(_06242_),
    .Y(_03948_));
 NOR2x1_ASAP7_75t_R _17832_ (.A(_01024_),
    .B(_06242_),
    .Y(_03949_));
 NOR2x1_ASAP7_75t_R _17833_ (.A(_01023_),
    .B(_06242_),
    .Y(_03950_));
 NOR2x1_ASAP7_75t_R _17834_ (.A(_01022_),
    .B(_06242_),
    .Y(_03951_));
 NOR2x1_ASAP7_75t_R _17835_ (.A(_01020_),
    .B(_06242_),
    .Y(_03952_));
 NOR2x1_ASAP7_75t_R _17836_ (.A(_01019_),
    .B(_06242_),
    .Y(_03953_));
 INVx1_ASAP7_75t_R _17837_ (.A(_06242_),
    .Y(_03954_));
 AND2x2_ASAP7_75t_R _17838_ (.A(_06143_),
    .B(_00043_),
    .Y(_03955_));
 OR4x1_ASAP7_75t_R _17839_ (.A(_01069_),
    .B(_01070_),
    .C(_01073_),
    .D(_02629_),
    .Y(_06243_));
 OR4x1_ASAP7_75t_R _17840_ (.A(_01065_),
    .B(_01066_),
    .C(_01067_),
    .D(_01068_),
    .Y(_06244_));
 OR2x6_ASAP7_75t_R _17841_ (.A(_06243_),
    .B(_06244_),
    .Y(_06245_));
 OR3x1_ASAP7_75t_R _17842_ (.A(_06232_),
    .B(_01094_),
    .C(_06245_),
    .Y(_06246_));
 OAI21x1_ASAP7_75t_R _17843_ (.A1(_06232_),
    .A2(_06245_),
    .B(_01094_),
    .Y(_06247_));
 AND3x1_ASAP7_75t_R _17844_ (.A(_06154_),
    .B(_06246_),
    .C(_06247_),
    .Y(_03956_));
 OR5x2_ASAP7_75t_R _17845_ (.A(_01069_),
    .B(_01070_),
    .C(_01073_),
    .D(_01084_),
    .E(_00043_),
    .Y(_06248_));
 OR2x2_ASAP7_75t_R _17846_ (.A(_06244_),
    .B(_06248_),
    .Y(_06249_));
 OR3x1_ASAP7_75t_R _17847_ (.A(_06232_),
    .B(_01094_),
    .C(_06249_),
    .Y(_06250_));
 XOR2x2_ASAP7_75t_R _17848_ (.A(_01093_),
    .B(_06250_),
    .Y(_06251_));
 AND2x2_ASAP7_75t_R _17849_ (.A(_06143_),
    .B(_06251_),
    .Y(_03957_));
 OR4x1_ASAP7_75t_R _17850_ (.A(_06232_),
    .B(_01092_),
    .C(_01093_),
    .D(_01094_),
    .Y(_06252_));
 OR3x2_ASAP7_75t_R _17851_ (.A(_06243_),
    .B(_06244_),
    .C(_06252_),
    .Y(_06253_));
 OR4x1_ASAP7_75t_R _17852_ (.A(_06232_),
    .B(_01093_),
    .C(_01094_),
    .D(_06245_),
    .Y(_06254_));
 NAND2x1_ASAP7_75t_R _17853_ (.A(_01092_),
    .B(_06254_),
    .Y(_06255_));
 AND3x1_ASAP7_75t_R _17854_ (.A(_06154_),
    .B(_06253_),
    .C(_06255_),
    .Y(_03958_));
 BUFx6f_ASAP7_75t_R _17855_ (.A(_06025_),
    .Y(_06256_));
 OR3x2_ASAP7_75t_R _17856_ (.A(_06244_),
    .B(_06248_),
    .C(_06252_),
    .Y(_06257_));
 XOR2x2_ASAP7_75t_R _17857_ (.A(_06231_),
    .B(_06257_),
    .Y(_06258_));
 AND2x2_ASAP7_75t_R _17858_ (.A(_06256_),
    .B(_06258_),
    .Y(_03959_));
 OR3x1_ASAP7_75t_R _17859_ (.A(_01090_),
    .B(_06231_),
    .C(_06253_),
    .Y(_06259_));
 OAI21x1_ASAP7_75t_R _17860_ (.A1(_06231_),
    .A2(_06253_),
    .B(_01090_),
    .Y(_06260_));
 AND3x1_ASAP7_75t_R _17861_ (.A(_06154_),
    .B(_06259_),
    .C(_06260_),
    .Y(_03960_));
 OR3x1_ASAP7_75t_R _17862_ (.A(_01090_),
    .B(_06231_),
    .C(_06257_),
    .Y(_06261_));
 XOR2x2_ASAP7_75t_R _17863_ (.A(_01089_),
    .B(_06261_),
    .Y(_06262_));
 AND2x2_ASAP7_75t_R _17864_ (.A(_06256_),
    .B(_06262_),
    .Y(_03961_));
 OR4x1_ASAP7_75t_R _17865_ (.A(_01089_),
    .B(_01090_),
    .C(_06231_),
    .D(_06253_),
    .Y(_06263_));
 XOR2x2_ASAP7_75t_R _17866_ (.A(_01088_),
    .B(_06263_),
    .Y(_06264_));
 AND2x2_ASAP7_75t_R _17867_ (.A(_06256_),
    .B(_06264_),
    .Y(_03962_));
 OR5x1_ASAP7_75t_R _17868_ (.A(_01088_),
    .B(_01089_),
    .C(_01090_),
    .D(_06231_),
    .E(_06257_),
    .Y(_06265_));
 XOR2x2_ASAP7_75t_R _17869_ (.A(_01087_),
    .B(_06265_),
    .Y(_06266_));
 AND2x2_ASAP7_75t_R _17870_ (.A(_06256_),
    .B(_06266_),
    .Y(_03963_));
 OR5x2_ASAP7_75t_R _17871_ (.A(_01087_),
    .B(_01088_),
    .C(_01089_),
    .D(_01090_),
    .E(_06231_),
    .Y(_06267_));
 OR3x2_ASAP7_75t_R _17872_ (.A(_01086_),
    .B(_06253_),
    .C(_06267_),
    .Y(_06268_));
 OAI21x1_ASAP7_75t_R _17873_ (.A1(_06253_),
    .A2(_06267_),
    .B(_01086_),
    .Y(_06269_));
 AND3x1_ASAP7_75t_R _17874_ (.A(_06154_),
    .B(_06268_),
    .C(_06269_),
    .Y(_03964_));
 OR3x2_ASAP7_75t_R _17875_ (.A(_01086_),
    .B(_06257_),
    .C(_06267_),
    .Y(_06270_));
 XOR2x2_ASAP7_75t_R _17876_ (.A(_01085_),
    .B(_06270_),
    .Y(_06271_));
 AND2x2_ASAP7_75t_R _17877_ (.A(_06256_),
    .B(_06271_),
    .Y(_03965_));
 BUFx12f_ASAP7_75t_R _17878_ (.A(_10012_),
    .Y(_06272_));
 NOR2x1_ASAP7_75t_R _17879_ (.A(_06272_),
    .B(_02630_),
    .Y(_03966_));
 OR3x1_ASAP7_75t_R _17880_ (.A(_01083_),
    .B(_01085_),
    .C(_06268_),
    .Y(_06273_));
 OAI21x1_ASAP7_75t_R _17881_ (.A1(_01085_),
    .A2(_06268_),
    .B(_01083_),
    .Y(_06274_));
 AND3x1_ASAP7_75t_R _17882_ (.A(_06154_),
    .B(_06273_),
    .C(_06274_),
    .Y(_03967_));
 OR3x1_ASAP7_75t_R _17883_ (.A(_01083_),
    .B(_01085_),
    .C(_06270_),
    .Y(_06275_));
 XOR2x2_ASAP7_75t_R _17884_ (.A(_01082_),
    .B(_06275_),
    .Y(_06276_));
 AND2x2_ASAP7_75t_R _17885_ (.A(_06256_),
    .B(_06276_),
    .Y(_03968_));
 OR4x1_ASAP7_75t_R _17886_ (.A(_01082_),
    .B(_01083_),
    .C(_01085_),
    .D(_06268_),
    .Y(_06277_));
 XOR2x2_ASAP7_75t_R _17887_ (.A(_01081_),
    .B(_06277_),
    .Y(_06278_));
 AND2x2_ASAP7_75t_R _17888_ (.A(_06256_),
    .B(_06278_),
    .Y(_03969_));
 OR4x1_ASAP7_75t_R _17889_ (.A(_01081_),
    .B(_01082_),
    .C(_01083_),
    .D(_01085_),
    .Y(_06279_));
 OR3x2_ASAP7_75t_R _17890_ (.A(_01080_),
    .B(_06270_),
    .C(_06279_),
    .Y(_06280_));
 OAI21x1_ASAP7_75t_R _17891_ (.A1(_06270_),
    .A2(_06279_),
    .B(_01080_),
    .Y(_06281_));
 AND3x1_ASAP7_75t_R _17892_ (.A(_06154_),
    .B(_06280_),
    .C(_06281_),
    .Y(_03970_));
 OR3x2_ASAP7_75t_R _17893_ (.A(_01080_),
    .B(_06268_),
    .C(_06279_),
    .Y(_06282_));
 XOR2x2_ASAP7_75t_R _17894_ (.A(_01079_),
    .B(_06282_),
    .Y(_06283_));
 AND2x2_ASAP7_75t_R _17895_ (.A(_06256_),
    .B(_06283_),
    .Y(_03971_));
 OR3x1_ASAP7_75t_R _17896_ (.A(_01078_),
    .B(_01079_),
    .C(_06280_),
    .Y(_06284_));
 OAI21x1_ASAP7_75t_R _17897_ (.A1(_01079_),
    .A2(_06280_),
    .B(_01078_),
    .Y(_06285_));
 AND3x1_ASAP7_75t_R _17898_ (.A(_06154_),
    .B(_06284_),
    .C(_06285_),
    .Y(_03972_));
 OR3x1_ASAP7_75t_R _17899_ (.A(_01078_),
    .B(_01079_),
    .C(_06282_),
    .Y(_06286_));
 XOR2x2_ASAP7_75t_R _17900_ (.A(_01077_),
    .B(_06286_),
    .Y(_06287_));
 AND2x2_ASAP7_75t_R _17901_ (.A(_06256_),
    .B(_06287_),
    .Y(_03973_));
 OR4x1_ASAP7_75t_R _17902_ (.A(_01077_),
    .B(_01078_),
    .C(_01079_),
    .D(_06280_),
    .Y(_06288_));
 XOR2x2_ASAP7_75t_R _17903_ (.A(_01076_),
    .B(_06288_),
    .Y(_06289_));
 AND2x2_ASAP7_75t_R _17904_ (.A(_06256_),
    .B(_06289_),
    .Y(_03974_));
 OR4x1_ASAP7_75t_R _17905_ (.A(_01076_),
    .B(_01077_),
    .C(_01078_),
    .D(_01079_),
    .Y(_06290_));
 OR3x1_ASAP7_75t_R _17906_ (.A(_01075_),
    .B(_06282_),
    .C(_06290_),
    .Y(_06291_));
 OAI21x1_ASAP7_75t_R _17907_ (.A1(_06282_),
    .A2(_06290_),
    .B(_01075_),
    .Y(_06292_));
 AND3x1_ASAP7_75t_R _17908_ (.A(_06154_),
    .B(_06291_),
    .C(_06292_),
    .Y(_03975_));
 BUFx6f_ASAP7_75t_R _17909_ (.A(_06025_),
    .Y(_06293_));
 OR3x1_ASAP7_75t_R _17910_ (.A(_01075_),
    .B(_06280_),
    .C(_06290_),
    .Y(_06294_));
 XOR2x2_ASAP7_75t_R _17911_ (.A(_01074_),
    .B(_06294_),
    .Y(_06295_));
 AND2x2_ASAP7_75t_R _17912_ (.A(_06293_),
    .B(_06295_),
    .Y(_03976_));
 XOR2x2_ASAP7_75t_R _17913_ (.A(_01073_),
    .B(_02629_),
    .Y(_06296_));
 AND2x2_ASAP7_75t_R _17914_ (.A(_06293_),
    .B(_06296_),
    .Y(_03977_));
 OR4x1_ASAP7_75t_R _17915_ (.A(_01074_),
    .B(_01075_),
    .C(_06282_),
    .D(_06290_),
    .Y(_06297_));
 XOR2x2_ASAP7_75t_R _17916_ (.A(_01072_),
    .B(_06297_),
    .Y(_06298_));
 AND2x2_ASAP7_75t_R _17917_ (.A(_06293_),
    .B(_06298_),
    .Y(_03978_));
 OR5x1_ASAP7_75t_R _17918_ (.A(_01072_),
    .B(_01074_),
    .C(_01075_),
    .D(_06280_),
    .E(_06290_),
    .Y(_06299_));
 XOR2x2_ASAP7_75t_R _17919_ (.A(_01071_),
    .B(_06299_),
    .Y(_06300_));
 AND2x2_ASAP7_75t_R _17920_ (.A(_06293_),
    .B(_06300_),
    .Y(_03979_));
 OR3x1_ASAP7_75t_R _17921_ (.A(_01073_),
    .B(_01084_),
    .C(_00043_),
    .Y(_06301_));
 XOR2x2_ASAP7_75t_R _17922_ (.A(_01070_),
    .B(_06301_),
    .Y(_06302_));
 AND2x2_ASAP7_75t_R _17923_ (.A(_06293_),
    .B(_06302_),
    .Y(_03980_));
 BUFx6f_ASAP7_75t_R _17924_ (.A(_05337_),
    .Y(_06303_));
 OR3x1_ASAP7_75t_R _17925_ (.A(_01070_),
    .B(_01073_),
    .C(_02629_),
    .Y(_06304_));
 NAND2x1_ASAP7_75t_R _17926_ (.A(_01069_),
    .B(_06304_),
    .Y(_06305_));
 AND3x1_ASAP7_75t_R _17927_ (.A(_06303_),
    .B(_06243_),
    .C(_06305_),
    .Y(_03981_));
 XOR2x2_ASAP7_75t_R _17928_ (.A(_01068_),
    .B(_06248_),
    .Y(_06306_));
 AND2x2_ASAP7_75t_R _17929_ (.A(_06293_),
    .B(_06306_),
    .Y(_03982_));
 OR3x1_ASAP7_75t_R _17930_ (.A(_01067_),
    .B(_01068_),
    .C(_06243_),
    .Y(_06307_));
 OAI21x1_ASAP7_75t_R _17931_ (.A1(_01068_),
    .A2(_06243_),
    .B(_01067_),
    .Y(_06308_));
 AND3x1_ASAP7_75t_R _17932_ (.A(_06303_),
    .B(_06307_),
    .C(_06308_),
    .Y(_03983_));
 OR3x1_ASAP7_75t_R _17933_ (.A(_01067_),
    .B(_01068_),
    .C(_06248_),
    .Y(_06309_));
 XOR2x2_ASAP7_75t_R _17934_ (.A(_01066_),
    .B(_06309_),
    .Y(_06310_));
 AND2x2_ASAP7_75t_R _17935_ (.A(_06293_),
    .B(_06310_),
    .Y(_03984_));
 OR4x1_ASAP7_75t_R _17936_ (.A(_01066_),
    .B(_01067_),
    .C(_01068_),
    .D(_06243_),
    .Y(_06311_));
 NAND2x1_ASAP7_75t_R _17937_ (.A(_01065_),
    .B(_06311_),
    .Y(_06312_));
 AND3x1_ASAP7_75t_R _17938_ (.A(_06303_),
    .B(_06245_),
    .C(_06312_),
    .Y(_03985_));
 XOR2x2_ASAP7_75t_R _17939_ (.A(_06232_),
    .B(_06249_),
    .Y(_06313_));
 AND2x2_ASAP7_75t_R _17940_ (.A(_06293_),
    .B(_06313_),
    .Y(_03986_));
 BUFx6f_ASAP7_75t_R _17941_ (.A(_01048_),
    .Y(_06314_));
 BUFx6f_ASAP7_75t_R _17942_ (.A(_01025_),
    .Y(_06315_));
 AND4x1_ASAP7_75t_R _17943_ (.A(_06315_),
    .B(_01053_),
    .C(_01054_),
    .D(_01055_),
    .Y(_06316_));
 AND5x1_ASAP7_75t_R _17944_ (.A(_01044_),
    .B(_01049_),
    .C(_01050_),
    .D(_01052_),
    .E(_06316_),
    .Y(_06317_));
 AND5x2_ASAP7_75t_R _17945_ (.A(_01046_),
    .B(_01047_),
    .C(_06314_),
    .D(_05995_),
    .E(_06317_),
    .Y(_06318_));
 BUFx6f_ASAP7_75t_R _17946_ (.A(_01040_),
    .Y(_06319_));
 AND4x1_ASAP7_75t_R _17947_ (.A(_01039_),
    .B(_06319_),
    .C(_01041_),
    .D(_01042_),
    .Y(_06320_));
 AND4x1_ASAP7_75t_R _17948_ (.A(_01033_),
    .B(_01035_),
    .C(_01036_),
    .D(_01043_),
    .Y(_06321_));
 AND5x1_ASAP7_75t_R _17949_ (.A(_01026_),
    .B(_01027_),
    .C(_01032_),
    .D(_01051_),
    .E(_06321_),
    .Y(_06322_));
 AND3x1_ASAP7_75t_R _17950_ (.A(_01030_),
    .B(_01031_),
    .C(_01034_),
    .Y(_06323_));
 OR3x1_ASAP7_75t_R _17951_ (.A(_01028_),
    .B(_01029_),
    .C(_06323_),
    .Y(_06324_));
 AND5x2_ASAP7_75t_R _17952_ (.A(_01037_),
    .B(_01038_),
    .C(_06320_),
    .D(_06322_),
    .E(_06324_),
    .Y(_06325_));
 NAND2x2_ASAP7_75t_R _17953_ (.A(_06318_),
    .B(_06325_),
    .Y(_06326_));
 NOR2x1_ASAP7_75t_R _17954_ (.A(_01015_),
    .B(_06326_),
    .Y(_03987_));
 INVx1_ASAP7_75t_R _17955_ (.A(_06326_),
    .Y(_03988_));
 NOR2x1_ASAP7_75t_R _17956_ (.A(_01018_),
    .B(_06326_),
    .Y(_03989_));
 NOR2x1_ASAP7_75t_R _17957_ (.A(_01017_),
    .B(_06326_),
    .Y(_03990_));
 NOR2x1_ASAP7_75t_R _17958_ (.A(_01016_),
    .B(_06326_),
    .Y(_03991_));
 NOR2x1_ASAP7_75t_R _17959_ (.A(_01014_),
    .B(_06326_),
    .Y(_03992_));
 NOR2x1_ASAP7_75t_R _17960_ (.A(_01013_),
    .B(_06326_),
    .Y(_03993_));
 INVx1_ASAP7_75t_R _17961_ (.A(_06326_),
    .Y(_03994_));
 AND2x2_ASAP7_75t_R _17962_ (.A(_06293_),
    .B(_00044_),
    .Y(_03995_));
 OR4x1_ASAP7_75t_R _17963_ (.A(_01030_),
    .B(_01031_),
    .C(_01034_),
    .D(_02617_),
    .Y(_06327_));
 OR4x1_ASAP7_75t_R _17964_ (.A(_01026_),
    .B(_01027_),
    .C(_01028_),
    .D(_01029_),
    .Y(_06328_));
 OR2x6_ASAP7_75t_R _17965_ (.A(_06327_),
    .B(_06328_),
    .Y(_06329_));
 OR3x1_ASAP7_75t_R _17966_ (.A(_06315_),
    .B(_01055_),
    .C(_06329_),
    .Y(_06330_));
 OAI21x1_ASAP7_75t_R _17967_ (.A1(_06315_),
    .A2(_06329_),
    .B(_01055_),
    .Y(_06331_));
 AND3x1_ASAP7_75t_R _17968_ (.A(_06303_),
    .B(_06330_),
    .C(_06331_),
    .Y(_03996_));
 OR5x2_ASAP7_75t_R _17969_ (.A(_01030_),
    .B(_01031_),
    .C(_01034_),
    .D(_01045_),
    .E(_00044_),
    .Y(_06332_));
 OR2x6_ASAP7_75t_R _17970_ (.A(_06328_),
    .B(_06332_),
    .Y(_06333_));
 OR3x1_ASAP7_75t_R _17971_ (.A(_06315_),
    .B(_01055_),
    .C(_06333_),
    .Y(_06334_));
 XOR2x2_ASAP7_75t_R _17972_ (.A(_01054_),
    .B(_06334_),
    .Y(_06335_));
 AND2x2_ASAP7_75t_R _17973_ (.A(_06293_),
    .B(_06335_),
    .Y(_03997_));
 BUFx6f_ASAP7_75t_R _17974_ (.A(_06025_),
    .Y(_06336_));
 OR4x1_ASAP7_75t_R _17975_ (.A(_06315_),
    .B(_01054_),
    .C(_01055_),
    .D(_06329_),
    .Y(_06337_));
 XOR2x2_ASAP7_75t_R _17976_ (.A(_01053_),
    .B(_06337_),
    .Y(_06338_));
 AND2x2_ASAP7_75t_R _17977_ (.A(_06336_),
    .B(_06338_),
    .Y(_03998_));
 OR5x2_ASAP7_75t_R _17978_ (.A(_06315_),
    .B(_01052_),
    .C(_01053_),
    .D(_01054_),
    .E(_01055_),
    .Y(_06339_));
 OR5x1_ASAP7_75t_R _17979_ (.A(_06315_),
    .B(_01053_),
    .C(_01054_),
    .D(_01055_),
    .E(_06333_),
    .Y(_06340_));
 NAND2x1_ASAP7_75t_R _17980_ (.A(_01052_),
    .B(_06340_),
    .Y(_06341_));
 OA211x2_ASAP7_75t_R _17981_ (.A1(_06333_),
    .A2(_06339_),
    .B(_06341_),
    .C(_11589_),
    .Y(_03999_));
 OR3x2_ASAP7_75t_R _17982_ (.A(_06327_),
    .B(_06328_),
    .C(_06339_),
    .Y(_06342_));
 XOR2x2_ASAP7_75t_R _17983_ (.A(_01051_),
    .B(_06342_),
    .Y(_06343_));
 AND2x2_ASAP7_75t_R _17984_ (.A(_06336_),
    .B(_06343_),
    .Y(_04000_));
 OR3x1_ASAP7_75t_R _17985_ (.A(_01051_),
    .B(_06333_),
    .C(_06339_),
    .Y(_06344_));
 XOR2x2_ASAP7_75t_R _17986_ (.A(_01050_),
    .B(_06344_),
    .Y(_06345_));
 AND2x2_ASAP7_75t_R _17987_ (.A(_06336_),
    .B(_06345_),
    .Y(_04001_));
 OR4x1_ASAP7_75t_R _17988_ (.A(_01049_),
    .B(_01050_),
    .C(_01051_),
    .D(_06342_),
    .Y(_06346_));
 OR3x1_ASAP7_75t_R _17989_ (.A(_01050_),
    .B(_01051_),
    .C(_06342_),
    .Y(_06347_));
 NAND2x1_ASAP7_75t_R _17990_ (.A(_01049_),
    .B(_06347_),
    .Y(_06348_));
 AND3x1_ASAP7_75t_R _17991_ (.A(_06303_),
    .B(_06346_),
    .C(_06348_),
    .Y(_04002_));
 OR5x2_ASAP7_75t_R _17992_ (.A(_01049_),
    .B(_01050_),
    .C(_01051_),
    .D(_06333_),
    .E(_06339_),
    .Y(_06349_));
 XOR2x2_ASAP7_75t_R _17993_ (.A(_06314_),
    .B(_06349_),
    .Y(_06350_));
 AND2x2_ASAP7_75t_R _17994_ (.A(_06336_),
    .B(_06350_),
    .Y(_04003_));
 OR3x1_ASAP7_75t_R _17995_ (.A(_01047_),
    .B(_06314_),
    .C(_06346_),
    .Y(_06351_));
 OAI21x1_ASAP7_75t_R _17996_ (.A1(_06314_),
    .A2(_06346_),
    .B(_01047_),
    .Y(_06352_));
 AND3x1_ASAP7_75t_R _17997_ (.A(_06303_),
    .B(_06351_),
    .C(_06352_),
    .Y(_04004_));
 OR3x1_ASAP7_75t_R _17998_ (.A(_01047_),
    .B(_06314_),
    .C(_06349_),
    .Y(_06353_));
 XOR2x2_ASAP7_75t_R _17999_ (.A(_01046_),
    .B(_06353_),
    .Y(_06354_));
 AND2x2_ASAP7_75t_R _18000_ (.A(_06336_),
    .B(_06354_),
    .Y(_04005_));
 NOR2x1_ASAP7_75t_R _18001_ (.A(_06272_),
    .B(_02618_),
    .Y(_04006_));
 OR4x1_ASAP7_75t_R _18002_ (.A(_01046_),
    .B(_01047_),
    .C(_06314_),
    .D(_06346_),
    .Y(_06355_));
 XOR2x2_ASAP7_75t_R _18003_ (.A(_01044_),
    .B(_06355_),
    .Y(_06356_));
 AND2x2_ASAP7_75t_R _18004_ (.A(_06336_),
    .B(_06356_),
    .Y(_04007_));
 OR5x1_ASAP7_75t_R _18005_ (.A(_01044_),
    .B(_01046_),
    .C(_01047_),
    .D(_06314_),
    .E(_06349_),
    .Y(_06357_));
 XOR2x2_ASAP7_75t_R _18006_ (.A(_01043_),
    .B(_06357_),
    .Y(_06358_));
 AND2x2_ASAP7_75t_R _18007_ (.A(_06336_),
    .B(_06358_),
    .Y(_04008_));
 OR5x2_ASAP7_75t_R _18008_ (.A(_01043_),
    .B(_01044_),
    .C(_01046_),
    .D(_01047_),
    .E(_06314_),
    .Y(_06359_));
 OR3x1_ASAP7_75t_R _18009_ (.A(_01042_),
    .B(_06346_),
    .C(_06359_),
    .Y(_06360_));
 OAI21x1_ASAP7_75t_R _18010_ (.A1(_06346_),
    .A2(_06359_),
    .B(_01042_),
    .Y(_06361_));
 AND3x1_ASAP7_75t_R _18011_ (.A(_06303_),
    .B(_06360_),
    .C(_06361_),
    .Y(_04009_));
 OR4x1_ASAP7_75t_R _18012_ (.A(_01041_),
    .B(_01042_),
    .C(_06349_),
    .D(_06359_),
    .Y(_06362_));
 OR3x1_ASAP7_75t_R _18013_ (.A(_01042_),
    .B(_06349_),
    .C(_06359_),
    .Y(_06363_));
 NAND2x1_ASAP7_75t_R _18014_ (.A(_01041_),
    .B(_06363_),
    .Y(_06364_));
 AND3x1_ASAP7_75t_R _18015_ (.A(_06303_),
    .B(_06362_),
    .C(_06364_),
    .Y(_04010_));
 OR4x1_ASAP7_75t_R _18016_ (.A(_01041_),
    .B(_01042_),
    .C(_06346_),
    .D(_06359_),
    .Y(_06365_));
 XOR2x2_ASAP7_75t_R _18017_ (.A(_06319_),
    .B(_06365_),
    .Y(_06366_));
 AND2x2_ASAP7_75t_R _18018_ (.A(_06336_),
    .B(_06366_),
    .Y(_04011_));
 OR3x1_ASAP7_75t_R _18019_ (.A(_01039_),
    .B(_06319_),
    .C(_06362_),
    .Y(_06367_));
 OAI21x1_ASAP7_75t_R _18020_ (.A1(_06319_),
    .A2(_06362_),
    .B(_01039_),
    .Y(_06368_));
 AND3x1_ASAP7_75t_R _18021_ (.A(_06303_),
    .B(_06367_),
    .C(_06368_),
    .Y(_04012_));
 OR3x1_ASAP7_75t_R _18022_ (.A(_01039_),
    .B(_06319_),
    .C(_06365_),
    .Y(_06369_));
 XOR2x2_ASAP7_75t_R _18023_ (.A(_01038_),
    .B(_06369_),
    .Y(_06370_));
 AND2x2_ASAP7_75t_R _18024_ (.A(_06336_),
    .B(_06370_),
    .Y(_04013_));
 OR4x1_ASAP7_75t_R _18025_ (.A(_01038_),
    .B(_01039_),
    .C(_06319_),
    .D(_06362_),
    .Y(_06371_));
 XOR2x2_ASAP7_75t_R _18026_ (.A(_01037_),
    .B(_06371_),
    .Y(_06372_));
 AND2x2_ASAP7_75t_R _18027_ (.A(_06336_),
    .B(_06372_),
    .Y(_04014_));
 BUFx6f_ASAP7_75t_R _18028_ (.A(_06025_),
    .Y(_06373_));
 OR5x1_ASAP7_75t_R _18029_ (.A(_01037_),
    .B(_01038_),
    .C(_01039_),
    .D(_06319_),
    .E(_06365_),
    .Y(_06374_));
 XOR2x2_ASAP7_75t_R _18030_ (.A(_01036_),
    .B(_06374_),
    .Y(_06375_));
 AND2x2_ASAP7_75t_R _18031_ (.A(_06373_),
    .B(_06375_),
    .Y(_04015_));
 OR5x2_ASAP7_75t_R _18032_ (.A(_01036_),
    .B(_01037_),
    .C(_01038_),
    .D(_01039_),
    .E(_06319_),
    .Y(_06376_));
 OR3x1_ASAP7_75t_R _18033_ (.A(_01035_),
    .B(_06362_),
    .C(_06376_),
    .Y(_06377_));
 OAI21x1_ASAP7_75t_R _18034_ (.A1(_06362_),
    .A2(_06376_),
    .B(_01035_),
    .Y(_06378_));
 AND3x1_ASAP7_75t_R _18035_ (.A(_06303_),
    .B(_06377_),
    .C(_06378_),
    .Y(_04016_));
 XOR2x2_ASAP7_75t_R _18036_ (.A(_01034_),
    .B(_02617_),
    .Y(_06379_));
 AND2x2_ASAP7_75t_R _18037_ (.A(_06373_),
    .B(_06379_),
    .Y(_04017_));
 OR3x1_ASAP7_75t_R _18038_ (.A(_01035_),
    .B(_06365_),
    .C(_06376_),
    .Y(_06380_));
 XOR2x2_ASAP7_75t_R _18039_ (.A(_01033_),
    .B(_06380_),
    .Y(_06381_));
 AND2x2_ASAP7_75t_R _18040_ (.A(_06373_),
    .B(_06381_),
    .Y(_04018_));
 OR4x1_ASAP7_75t_R _18041_ (.A(_01033_),
    .B(_01035_),
    .C(_06362_),
    .D(_06376_),
    .Y(_06382_));
 XOR2x2_ASAP7_75t_R _18042_ (.A(_01032_),
    .B(_06382_),
    .Y(_06383_));
 AND2x2_ASAP7_75t_R _18043_ (.A(_06373_),
    .B(_06383_),
    .Y(_04019_));
 OR3x1_ASAP7_75t_R _18044_ (.A(_01034_),
    .B(_01045_),
    .C(_00044_),
    .Y(_06384_));
 XOR2x2_ASAP7_75t_R _18045_ (.A(_01031_),
    .B(_06384_),
    .Y(_06385_));
 AND2x2_ASAP7_75t_R _18046_ (.A(_06373_),
    .B(_06385_),
    .Y(_04020_));
 BUFx12f_ASAP7_75t_R _18047_ (.A(_08527_),
    .Y(_06386_));
 BUFx6f_ASAP7_75t_R _18048_ (.A(_06386_),
    .Y(_06387_));
 OR3x1_ASAP7_75t_R _18049_ (.A(_01031_),
    .B(_01034_),
    .C(_02617_),
    .Y(_06388_));
 NAND2x1_ASAP7_75t_R _18050_ (.A(_01030_),
    .B(_06388_),
    .Y(_06389_));
 AND3x1_ASAP7_75t_R _18051_ (.A(_06387_),
    .B(_06327_),
    .C(_06389_),
    .Y(_04021_));
 XOR2x2_ASAP7_75t_R _18052_ (.A(_01029_),
    .B(_06332_),
    .Y(_06390_));
 AND2x2_ASAP7_75t_R _18053_ (.A(_06373_),
    .B(_06390_),
    .Y(_04022_));
 OR3x1_ASAP7_75t_R _18054_ (.A(_01028_),
    .B(_01029_),
    .C(_06327_),
    .Y(_06391_));
 OAI21x1_ASAP7_75t_R _18055_ (.A1(_01029_),
    .A2(_06327_),
    .B(_01028_),
    .Y(_06392_));
 AND3x1_ASAP7_75t_R _18056_ (.A(_06387_),
    .B(_06391_),
    .C(_06392_),
    .Y(_04023_));
 OR3x1_ASAP7_75t_R _18057_ (.A(_01028_),
    .B(_01029_),
    .C(_06332_),
    .Y(_06393_));
 XOR2x2_ASAP7_75t_R _18058_ (.A(_01027_),
    .B(_06393_),
    .Y(_06394_));
 AND2x2_ASAP7_75t_R _18059_ (.A(_06373_),
    .B(_06394_),
    .Y(_04024_));
 OR4x1_ASAP7_75t_R _18060_ (.A(_01027_),
    .B(_01028_),
    .C(_01029_),
    .D(_06327_),
    .Y(_06395_));
 NAND2x1_ASAP7_75t_R _18061_ (.A(_01026_),
    .B(_06395_),
    .Y(_06396_));
 AND3x1_ASAP7_75t_R _18062_ (.A(_06387_),
    .B(_06329_),
    .C(_06396_),
    .Y(_04025_));
 XOR2x2_ASAP7_75t_R _18063_ (.A(_06315_),
    .B(_06333_),
    .Y(_06397_));
 AND2x2_ASAP7_75t_R _18064_ (.A(_06373_),
    .B(_06397_),
    .Y(_04026_));
 AND2x2_ASAP7_75t_R _18065_ (.A(_06373_),
    .B(_00021_),
    .Y(_04027_));
 INVx1_ASAP7_75t_R _18066_ (.A(_02033_),
    .Y(_06398_));
 BUFx6f_ASAP7_75t_R _18067_ (.A(_02022_),
    .Y(_06399_));
 INVx1_ASAP7_75t_R _18068_ (.A(_02029_),
    .Y(_06400_));
 OR2x2_ASAP7_75t_R _18069_ (.A(_01095_),
    .B(_01100_),
    .Y(_06401_));
 OR4x1_ASAP7_75t_R _18070_ (.A(_01057_),
    .B(_01058_),
    .C(_01059_),
    .D(_01060_),
    .Y(_06402_));
 OR3x2_ASAP7_75t_R _18071_ (.A(_01056_),
    .B(\peo[31][32] ),
    .C(_06402_),
    .Y(_06403_));
 AO21x1_ASAP7_75t_R _18072_ (.A1(\xs[15].cli1.i[39] ),
    .A2(_06402_),
    .B(_02029_),
    .Y(_06404_));
 OR4x1_ASAP7_75t_R _18073_ (.A(_01096_),
    .B(_01097_),
    .C(_01098_),
    .D(_01099_),
    .Y(_06405_));
 AND2x4_ASAP7_75t_R _18074_ (.A(\peo[30][39] ),
    .B(_06405_),
    .Y(_06406_));
 AO221x1_ASAP7_75t_R _18075_ (.A1(_06400_),
    .A2(_06401_),
    .B1(_06403_),
    .B2(_06404_),
    .C(_06406_),
    .Y(_06407_));
 NAND2x1_ASAP7_75t_R _18076_ (.A(_02023_),
    .B(_06407_),
    .Y(_06408_));
 OR4x1_ASAP7_75t_R _18077_ (.A(_08571_),
    .B(_06399_),
    .C(_06400_),
    .D(_06408_),
    .Y(_06409_));
 BUFx6f_ASAP7_75t_R _18078_ (.A(_06409_),
    .Y(_06410_));
 INVx1_ASAP7_75t_R _18079_ (.A(_06410_),
    .Y(_06411_));
 OR3x1_ASAP7_75t_R _18080_ (.A(_06399_),
    .B(_06400_),
    .C(_06408_),
    .Y(_06412_));
 AND2x4_ASAP7_75t_R _18081_ (.A(\xs[15].cli1.i[39] ),
    .B(_06402_),
    .Y(_06413_));
 INVx2_ASAP7_75t_R _18082_ (.A(_06399_),
    .Y(_06414_));
 AO21x1_ASAP7_75t_R _18083_ (.A1(_00021_),
    .A2(_06413_),
    .B(_06414_),
    .Y(_06415_));
 INVx1_ASAP7_75t_R _18084_ (.A(_02023_),
    .Y(_06416_));
 OR3x1_ASAP7_75t_R _18085_ (.A(_06399_),
    .B(_06416_),
    .C(_02029_),
    .Y(_06417_));
 AND3x1_ASAP7_75t_R _18086_ (.A(_06406_),
    .B(_06415_),
    .C(_06417_),
    .Y(_06418_));
 OAI21x1_ASAP7_75t_R _18087_ (.A1(_06403_),
    .A2(_06418_),
    .B(_01102_),
    .Y(_06419_));
 NOR3x1_ASAP7_75t_R _18088_ (.A(_01056_),
    .B(\peo[31][32] ),
    .C(_06402_),
    .Y(_06420_));
 AO21x1_ASAP7_75t_R _18089_ (.A1(_06406_),
    .A2(_06420_),
    .B(_06413_),
    .Y(_06421_));
 AND2x2_ASAP7_75t_R _18090_ (.A(_06414_),
    .B(_02029_),
    .Y(_06422_));
 OA21x2_ASAP7_75t_R _18091_ (.A1(_01061_),
    .A2(_06402_),
    .B(\xs[15].cli1.i[39] ),
    .Y(_06423_));
 AO32x1_ASAP7_75t_R _18092_ (.A1(_06399_),
    .A2(_00021_),
    .A3(_06413_),
    .B1(_06422_),
    .B2(_06423_),
    .Y(_06424_));
 AO32x2_ASAP7_75t_R _18093_ (.A1(_06414_),
    .A2(_06416_),
    .A3(_06421_),
    .B1(_06424_),
    .B2(_06406_),
    .Y(_06425_));
 OR3x1_ASAP7_75t_R _18094_ (.A(\peo[31][0] ),
    .B(_06403_),
    .C(_06425_),
    .Y(_06426_));
 AND4x1_ASAP7_75t_R _18095_ (.A(_08722_),
    .B(_06412_),
    .C(_06419_),
    .D(_06426_),
    .Y(_06427_));
 AO21x1_ASAP7_75t_R _18096_ (.A1(_06398_),
    .A2(_06411_),
    .B(_06427_),
    .Y(_04028_));
 NOR2x1_ASAP7_75t_R _18097_ (.A(_02032_),
    .B(_06410_),
    .Y(_04029_));
 NOR2x1_ASAP7_75t_R _18098_ (.A(_02031_),
    .B(_06410_),
    .Y(_04030_));
 NOR2x1_ASAP7_75t_R _18099_ (.A(_02030_),
    .B(_06410_),
    .Y(_04031_));
 NOR2x1_ASAP7_75t_R _18100_ (.A(_02021_),
    .B(_06410_),
    .Y(_04032_));
 NOR2x1_ASAP7_75t_R _18101_ (.A(_02020_),
    .B(_06410_),
    .Y(_04033_));
 AND3x1_ASAP7_75t_R _18102_ (.A(_06414_),
    .B(_02023_),
    .C(_06400_),
    .Y(_06428_));
 NAND2x1_ASAP7_75t_R _18103_ (.A(_06407_),
    .B(_06428_),
    .Y(_06429_));
 AND3x1_ASAP7_75t_R _18104_ (.A(_06398_),
    .B(_06407_),
    .C(_06428_),
    .Y(_06430_));
 AO21x1_ASAP7_75t_R _18105_ (.A1(\peo[30][0] ),
    .A2(_06429_),
    .B(_06430_),
    .Y(_06431_));
 NAND2x1_ASAP7_75t_R _18106_ (.A(_01063_),
    .B(_06425_),
    .Y(_06432_));
 BUFx12f_ASAP7_75t_R _18107_ (.A(_08876_),
    .Y(_06433_));
 OA211x2_ASAP7_75t_R _18108_ (.A1(_06425_),
    .A2(_06431_),
    .B(_06432_),
    .C(_06433_),
    .Y(_04034_));
 OR4x1_ASAP7_75t_R _18109_ (.A(_11177_),
    .B(_06399_),
    .C(_02029_),
    .D(_06408_),
    .Y(_06434_));
 NOR2x1_ASAP7_75t_R _18110_ (.A(_02032_),
    .B(_06434_),
    .Y(_04035_));
 NOR2x1_ASAP7_75t_R _18111_ (.A(_02031_),
    .B(_06434_),
    .Y(_04036_));
 NOR2x1_ASAP7_75t_R _18112_ (.A(_02030_),
    .B(_06434_),
    .Y(_04037_));
 NOR2x1_ASAP7_75t_R _18113_ (.A(_02021_),
    .B(_06434_),
    .Y(_04038_));
 NOR2x1_ASAP7_75t_R _18114_ (.A(_02020_),
    .B(_06434_),
    .Y(_04039_));
 INVx1_ASAP7_75t_R _18115_ (.A(_06408_),
    .Y(_06435_));
 OR3x2_ASAP7_75t_R _18116_ (.A(_09220_),
    .B(_06399_),
    .C(_06435_),
    .Y(_06436_));
 BUFx12f_ASAP7_75t_R _18117_ (.A(_06436_),
    .Y(_06437_));
 AO21x2_ASAP7_75t_R _18118_ (.A1(_06414_),
    .A2(_06408_),
    .B(_08572_),
    .Y(_06438_));
 OAI21x1_ASAP7_75t_R _18119_ (.A1(_06399_),
    .A2(_02023_),
    .B(_06413_),
    .Y(_06439_));
 AO21x2_ASAP7_75t_R _18120_ (.A1(_06406_),
    .A2(_06424_),
    .B(_06439_),
    .Y(_06440_));
 NAND2x1_ASAP7_75t_R _18121_ (.A(\peo[30][0] ),
    .B(_06440_),
    .Y(_06441_));
 OA21x2_ASAP7_75t_R _18122_ (.A1(_01063_),
    .A2(_06440_),
    .B(_06441_),
    .Y(_06442_));
 OAI22x1_ASAP7_75t_R _18123_ (.A1(_02033_),
    .A2(_06437_),
    .B1(_06438_),
    .B2(_06442_),
    .Y(_04040_));
 NOR2x1_ASAP7_75t_R _18124_ (.A(_02032_),
    .B(_06437_),
    .Y(_04041_));
 NOR2x1_ASAP7_75t_R _18125_ (.A(_02031_),
    .B(_06437_),
    .Y(_04042_));
 NOR2x1_ASAP7_75t_R _18126_ (.A(_02030_),
    .B(_06437_),
    .Y(_04043_));
 NOR2x1_ASAP7_75t_R _18127_ (.A(\peo[31][32] ),
    .B(_06440_),
    .Y(_06443_));
 AO21x1_ASAP7_75t_R _18128_ (.A1(_01100_),
    .A2(_06440_),
    .B(_06443_),
    .Y(_06444_));
 OAI22x1_ASAP7_75t_R _18129_ (.A1(_02029_),
    .A2(_06437_),
    .B1(_06438_),
    .B2(_06444_),
    .Y(_04044_));
 NOR2x1_ASAP7_75t_R _18130_ (.A(_01056_),
    .B(_06425_),
    .Y(_06445_));
 AO221x1_ASAP7_75t_R _18131_ (.A1(_01099_),
    .A2(_06440_),
    .B1(_06445_),
    .B2(_01060_),
    .C(_06438_),
    .Y(_06446_));
 OAI21x1_ASAP7_75t_R _18132_ (.A1(_02028_),
    .A2(_06437_),
    .B(_06446_),
    .Y(_04045_));
 AO221x1_ASAP7_75t_R _18133_ (.A1(_01098_),
    .A2(_06440_),
    .B1(_06445_),
    .B2(_01059_),
    .C(_06438_),
    .Y(_06447_));
 OAI21x1_ASAP7_75t_R _18134_ (.A1(_02027_),
    .A2(_06437_),
    .B(_06447_),
    .Y(_04046_));
 AO221x1_ASAP7_75t_R _18135_ (.A1(_01097_),
    .A2(_06440_),
    .B1(_06445_),
    .B2(_01058_),
    .C(_06438_),
    .Y(_06448_));
 OAI21x1_ASAP7_75t_R _18136_ (.A1(_02026_),
    .A2(_06437_),
    .B(_06448_),
    .Y(_04047_));
 AO221x1_ASAP7_75t_R _18137_ (.A1(_01096_),
    .A2(_06440_),
    .B1(_06445_),
    .B2(_01057_),
    .C(_06438_),
    .Y(_06449_));
 OAI21x1_ASAP7_75t_R _18138_ (.A1(_02025_),
    .A2(_06437_),
    .B(_06449_),
    .Y(_04048_));
 NOR2x1_ASAP7_75t_R _18139_ (.A(_02024_),
    .B(_06437_),
    .Y(_04049_));
 OR4x1_ASAP7_75t_R _18140_ (.A(_08684_),
    .B(_06399_),
    .C(_06416_),
    .D(_06407_),
    .Y(_06450_));
 INVx1_ASAP7_75t_R _18141_ (.A(_06450_),
    .Y(_04050_));
 AO221x1_ASAP7_75t_R _18142_ (.A1(\xs[15].cli1.i[39] ),
    .A2(_06402_),
    .B1(_06408_),
    .B2(_06414_),
    .C(_06406_),
    .Y(_06451_));
 AND2x2_ASAP7_75t_R _18143_ (.A(_06373_),
    .B(_06451_),
    .Y(_04051_));
 NOR2x1_ASAP7_75t_R _18144_ (.A(_02021_),
    .B(_06436_),
    .Y(_04052_));
 NOR2x1_ASAP7_75t_R _18145_ (.A(_02020_),
    .B(_06436_),
    .Y(_04053_));
 BUFx6f_ASAP7_75t_R _18146_ (.A(_00987_),
    .Y(_06452_));
 BUFx3_ASAP7_75t_R _18147_ (.A(_00960_),
    .Y(_06453_));
 AND4x1_ASAP7_75t_R _18148_ (.A(_06453_),
    .B(_00988_),
    .C(_00989_),
    .D(_00990_),
    .Y(_06454_));
 AND5x1_ASAP7_75t_R _18149_ (.A(_00979_),
    .B(_00984_),
    .C(_00985_),
    .D(_06452_),
    .E(_06454_),
    .Y(_06455_));
 AND5x2_ASAP7_75t_R _18150_ (.A(_00981_),
    .B(_00982_),
    .C(_00983_),
    .D(_05995_),
    .E(_06455_),
    .Y(_06456_));
 AND4x1_ASAP7_75t_R _18151_ (.A(_00974_),
    .B(_00975_),
    .C(_00976_),
    .D(_00977_),
    .Y(_06457_));
 AND4x1_ASAP7_75t_R _18152_ (.A(_00968_),
    .B(_00970_),
    .C(_00971_),
    .D(_00978_),
    .Y(_06458_));
 AND5x1_ASAP7_75t_R _18153_ (.A(_00961_),
    .B(_00962_),
    .C(_00967_),
    .D(_00986_),
    .E(_06458_),
    .Y(_06459_));
 AND3x1_ASAP7_75t_R _18154_ (.A(_00965_),
    .B(_00966_),
    .C(_00969_),
    .Y(_06460_));
 OR3x1_ASAP7_75t_R _18155_ (.A(_00963_),
    .B(_00964_),
    .C(_06460_),
    .Y(_06461_));
 AND5x2_ASAP7_75t_R _18156_ (.A(_00972_),
    .B(_00973_),
    .C(_06457_),
    .D(_06459_),
    .E(_06461_),
    .Y(_06462_));
 NAND2x2_ASAP7_75t_R _18157_ (.A(_06456_),
    .B(_06462_),
    .Y(_06463_));
 NOR2x1_ASAP7_75t_R _18158_ (.A(_00917_),
    .B(_06463_),
    .Y(_04054_));
 INVx1_ASAP7_75t_R _18159_ (.A(_06463_),
    .Y(_04055_));
 NOR2x1_ASAP7_75t_R _18160_ (.A(_00920_),
    .B(_06463_),
    .Y(_04056_));
 NOR2x1_ASAP7_75t_R _18161_ (.A(_00919_),
    .B(_06463_),
    .Y(_04057_));
 NOR2x1_ASAP7_75t_R _18162_ (.A(_00918_),
    .B(_06463_),
    .Y(_04058_));
 NOR2x1_ASAP7_75t_R _18163_ (.A(_00916_),
    .B(_06463_),
    .Y(_04059_));
 NOR2x1_ASAP7_75t_R _18164_ (.A(_00915_),
    .B(_06463_),
    .Y(_04060_));
 INVx1_ASAP7_75t_R _18165_ (.A(_06463_),
    .Y(_04061_));
 BUFx6f_ASAP7_75t_R _18166_ (.A(_06025_),
    .Y(_06464_));
 AND2x2_ASAP7_75t_R _18167_ (.A(_06464_),
    .B(_00045_),
    .Y(_04062_));
 OR4x1_ASAP7_75t_R _18168_ (.A(_00965_),
    .B(_00966_),
    .C(_00969_),
    .D(_02615_),
    .Y(_06465_));
 OR4x1_ASAP7_75t_R _18169_ (.A(_00961_),
    .B(_00962_),
    .C(_00963_),
    .D(_00964_),
    .Y(_06466_));
 OR2x6_ASAP7_75t_R _18170_ (.A(_06465_),
    .B(_06466_),
    .Y(_06467_));
 OR3x1_ASAP7_75t_R _18171_ (.A(_06453_),
    .B(_00990_),
    .C(_06467_),
    .Y(_06468_));
 OAI21x1_ASAP7_75t_R _18172_ (.A1(_06453_),
    .A2(_06467_),
    .B(_00990_),
    .Y(_06469_));
 AND3x1_ASAP7_75t_R _18173_ (.A(_06387_),
    .B(_06468_),
    .C(_06469_),
    .Y(_04063_));
 OR5x2_ASAP7_75t_R _18174_ (.A(_00965_),
    .B(_00966_),
    .C(_00969_),
    .D(_00980_),
    .E(_00045_),
    .Y(_06470_));
 OR2x2_ASAP7_75t_R _18175_ (.A(_06466_),
    .B(_06470_),
    .Y(_06471_));
 OR3x1_ASAP7_75t_R _18176_ (.A(_06453_),
    .B(_00990_),
    .C(_06471_),
    .Y(_06472_));
 XOR2x2_ASAP7_75t_R _18177_ (.A(_00989_),
    .B(_06472_),
    .Y(_06473_));
 AND2x2_ASAP7_75t_R _18178_ (.A(_06464_),
    .B(_06473_),
    .Y(_04064_));
 OR4x1_ASAP7_75t_R _18179_ (.A(_06453_),
    .B(_00988_),
    .C(_00989_),
    .D(_00990_),
    .Y(_06474_));
 OR3x2_ASAP7_75t_R _18180_ (.A(_06465_),
    .B(_06466_),
    .C(_06474_),
    .Y(_06475_));
 OR4x1_ASAP7_75t_R _18181_ (.A(_06453_),
    .B(_00989_),
    .C(_00990_),
    .D(_06467_),
    .Y(_06476_));
 NAND2x1_ASAP7_75t_R _18182_ (.A(_00988_),
    .B(_06476_),
    .Y(_06477_));
 AND3x1_ASAP7_75t_R _18183_ (.A(_06387_),
    .B(_06475_),
    .C(_06477_),
    .Y(_04065_));
 OR3x2_ASAP7_75t_R _18184_ (.A(_06466_),
    .B(_06470_),
    .C(_06474_),
    .Y(_06478_));
 XOR2x2_ASAP7_75t_R _18185_ (.A(_06452_),
    .B(_06478_),
    .Y(_06479_));
 AND2x2_ASAP7_75t_R _18186_ (.A(_06464_),
    .B(_06479_),
    .Y(_04066_));
 OR3x1_ASAP7_75t_R _18187_ (.A(_00986_),
    .B(_06452_),
    .C(_06475_),
    .Y(_06480_));
 OAI21x1_ASAP7_75t_R _18188_ (.A1(_06452_),
    .A2(_06475_),
    .B(_00986_),
    .Y(_06481_));
 AND3x1_ASAP7_75t_R _18189_ (.A(_06387_),
    .B(_06480_),
    .C(_06481_),
    .Y(_04067_));
 OR3x1_ASAP7_75t_R _18190_ (.A(_00986_),
    .B(_06452_),
    .C(_06478_),
    .Y(_06482_));
 XOR2x2_ASAP7_75t_R _18191_ (.A(_00985_),
    .B(_06482_),
    .Y(_06483_));
 AND2x2_ASAP7_75t_R _18192_ (.A(_06464_),
    .B(_06483_),
    .Y(_04068_));
 OR4x1_ASAP7_75t_R _18193_ (.A(_00985_),
    .B(_00986_),
    .C(_06452_),
    .D(_06475_),
    .Y(_06484_));
 XOR2x2_ASAP7_75t_R _18194_ (.A(_00984_),
    .B(_06484_),
    .Y(_06485_));
 AND2x2_ASAP7_75t_R _18195_ (.A(_06464_),
    .B(_06485_),
    .Y(_04069_));
 OR5x1_ASAP7_75t_R _18196_ (.A(_00984_),
    .B(_00985_),
    .C(_00986_),
    .D(_06452_),
    .E(_06478_),
    .Y(_06486_));
 XOR2x2_ASAP7_75t_R _18197_ (.A(_00983_),
    .B(_06486_),
    .Y(_06487_));
 AND2x2_ASAP7_75t_R _18198_ (.A(_06464_),
    .B(_06487_),
    .Y(_04070_));
 OR5x2_ASAP7_75t_R _18199_ (.A(_00983_),
    .B(_00984_),
    .C(_00985_),
    .D(_00986_),
    .E(_06452_),
    .Y(_06488_));
 OR3x2_ASAP7_75t_R _18200_ (.A(_00982_),
    .B(_06475_),
    .C(_06488_),
    .Y(_06489_));
 OAI21x1_ASAP7_75t_R _18201_ (.A1(_06475_),
    .A2(_06488_),
    .B(_00982_),
    .Y(_06490_));
 AND3x1_ASAP7_75t_R _18202_ (.A(_06387_),
    .B(_06489_),
    .C(_06490_),
    .Y(_04071_));
 OR3x2_ASAP7_75t_R _18203_ (.A(_00982_),
    .B(_06478_),
    .C(_06488_),
    .Y(_06491_));
 XOR2x2_ASAP7_75t_R _18204_ (.A(_00981_),
    .B(_06491_),
    .Y(_06492_));
 AND2x2_ASAP7_75t_R _18205_ (.A(_06464_),
    .B(_06492_),
    .Y(_04072_));
 NOR2x1_ASAP7_75t_R _18206_ (.A(_06272_),
    .B(_02616_),
    .Y(_04073_));
 OR3x1_ASAP7_75t_R _18207_ (.A(_00979_),
    .B(_00981_),
    .C(_06489_),
    .Y(_06493_));
 OAI21x1_ASAP7_75t_R _18208_ (.A1(_00981_),
    .A2(_06489_),
    .B(_00979_),
    .Y(_06494_));
 AND3x1_ASAP7_75t_R _18209_ (.A(_06387_),
    .B(_06493_),
    .C(_06494_),
    .Y(_04074_));
 OR3x1_ASAP7_75t_R _18210_ (.A(_00979_),
    .B(_00981_),
    .C(_06491_),
    .Y(_06495_));
 XOR2x2_ASAP7_75t_R _18211_ (.A(_00978_),
    .B(_06495_),
    .Y(_06496_));
 AND2x2_ASAP7_75t_R _18212_ (.A(_06464_),
    .B(_06496_),
    .Y(_04075_));
 OR4x1_ASAP7_75t_R _18213_ (.A(_00978_),
    .B(_00979_),
    .C(_00981_),
    .D(_06489_),
    .Y(_06497_));
 XOR2x2_ASAP7_75t_R _18214_ (.A(_00977_),
    .B(_06497_),
    .Y(_06498_));
 AND2x2_ASAP7_75t_R _18215_ (.A(_06464_),
    .B(_06498_),
    .Y(_04076_));
 OR4x1_ASAP7_75t_R _18216_ (.A(_00977_),
    .B(_00978_),
    .C(_00979_),
    .D(_00981_),
    .Y(_06499_));
 OR3x2_ASAP7_75t_R _18217_ (.A(_00976_),
    .B(_06491_),
    .C(_06499_),
    .Y(_06500_));
 OAI21x1_ASAP7_75t_R _18218_ (.A1(_06491_),
    .A2(_06499_),
    .B(_00976_),
    .Y(_06501_));
 AND3x1_ASAP7_75t_R _18219_ (.A(_06387_),
    .B(_06500_),
    .C(_06501_),
    .Y(_04077_));
 OR3x2_ASAP7_75t_R _18220_ (.A(_00976_),
    .B(_06489_),
    .C(_06499_),
    .Y(_06502_));
 XOR2x2_ASAP7_75t_R _18221_ (.A(_00975_),
    .B(_06502_),
    .Y(_06503_));
 AND2x2_ASAP7_75t_R _18222_ (.A(_06464_),
    .B(_06503_),
    .Y(_04078_));
 OR3x1_ASAP7_75t_R _18223_ (.A(_00974_),
    .B(_00975_),
    .C(_06500_),
    .Y(_06504_));
 OAI21x1_ASAP7_75t_R _18224_ (.A1(_00975_),
    .A2(_06500_),
    .B(_00974_),
    .Y(_06505_));
 AND3x1_ASAP7_75t_R _18225_ (.A(_06387_),
    .B(_06504_),
    .C(_06505_),
    .Y(_04079_));
 BUFx6f_ASAP7_75t_R _18226_ (.A(_06025_),
    .Y(_06506_));
 OR3x1_ASAP7_75t_R _18227_ (.A(_00974_),
    .B(_00975_),
    .C(_06502_),
    .Y(_06507_));
 XOR2x2_ASAP7_75t_R _18228_ (.A(_00973_),
    .B(_06507_),
    .Y(_06508_));
 AND2x2_ASAP7_75t_R _18229_ (.A(_06506_),
    .B(_06508_),
    .Y(_04080_));
 OR4x1_ASAP7_75t_R _18230_ (.A(_00973_),
    .B(_00974_),
    .C(_00975_),
    .D(_06500_),
    .Y(_06509_));
 XOR2x2_ASAP7_75t_R _18231_ (.A(_00972_),
    .B(_06509_),
    .Y(_06510_));
 AND2x2_ASAP7_75t_R _18232_ (.A(_06506_),
    .B(_06510_),
    .Y(_04081_));
 BUFx6f_ASAP7_75t_R _18233_ (.A(_06386_),
    .Y(_06511_));
 OR4x1_ASAP7_75t_R _18234_ (.A(_00972_),
    .B(_00973_),
    .C(_00974_),
    .D(_00975_),
    .Y(_06512_));
 OR3x1_ASAP7_75t_R _18235_ (.A(_00971_),
    .B(_06502_),
    .C(_06512_),
    .Y(_06513_));
 OAI21x1_ASAP7_75t_R _18236_ (.A1(_06502_),
    .A2(_06512_),
    .B(_00971_),
    .Y(_06514_));
 AND3x1_ASAP7_75t_R _18237_ (.A(_06511_),
    .B(_06513_),
    .C(_06514_),
    .Y(_04082_));
 OR3x1_ASAP7_75t_R _18238_ (.A(_00971_),
    .B(_06500_),
    .C(_06512_),
    .Y(_06515_));
 XOR2x2_ASAP7_75t_R _18239_ (.A(_00970_),
    .B(_06515_),
    .Y(_06516_));
 AND2x2_ASAP7_75t_R _18240_ (.A(_06506_),
    .B(_06516_),
    .Y(_04083_));
 XOR2x2_ASAP7_75t_R _18241_ (.A(_00969_),
    .B(_02615_),
    .Y(_06517_));
 AND2x2_ASAP7_75t_R _18242_ (.A(_06506_),
    .B(_06517_),
    .Y(_04084_));
 OR4x1_ASAP7_75t_R _18243_ (.A(_00970_),
    .B(_00971_),
    .C(_06502_),
    .D(_06512_),
    .Y(_06518_));
 XOR2x2_ASAP7_75t_R _18244_ (.A(_00968_),
    .B(_06518_),
    .Y(_06519_));
 AND2x2_ASAP7_75t_R _18245_ (.A(_06506_),
    .B(_06519_),
    .Y(_04085_));
 OR5x1_ASAP7_75t_R _18246_ (.A(_00968_),
    .B(_00970_),
    .C(_00971_),
    .D(_06500_),
    .E(_06512_),
    .Y(_06520_));
 XOR2x2_ASAP7_75t_R _18247_ (.A(_00967_),
    .B(_06520_),
    .Y(_06521_));
 AND2x2_ASAP7_75t_R _18248_ (.A(_06506_),
    .B(_06521_),
    .Y(_04086_));
 OR3x1_ASAP7_75t_R _18249_ (.A(_00969_),
    .B(_00980_),
    .C(_00045_),
    .Y(_06522_));
 XOR2x2_ASAP7_75t_R _18250_ (.A(_00966_),
    .B(_06522_),
    .Y(_06523_));
 AND2x2_ASAP7_75t_R _18251_ (.A(_06506_),
    .B(_06523_),
    .Y(_04087_));
 OR3x1_ASAP7_75t_R _18252_ (.A(_00966_),
    .B(_00969_),
    .C(_02615_),
    .Y(_06524_));
 NAND2x1_ASAP7_75t_R _18253_ (.A(_00965_),
    .B(_06524_),
    .Y(_06525_));
 AND3x1_ASAP7_75t_R _18254_ (.A(_06511_),
    .B(_06465_),
    .C(_06525_),
    .Y(_04088_));
 XOR2x2_ASAP7_75t_R _18255_ (.A(_00964_),
    .B(_06470_),
    .Y(_06526_));
 AND2x2_ASAP7_75t_R _18256_ (.A(_06506_),
    .B(_06526_),
    .Y(_04089_));
 OR3x1_ASAP7_75t_R _18257_ (.A(_00963_),
    .B(_00964_),
    .C(_06465_),
    .Y(_06527_));
 OAI21x1_ASAP7_75t_R _18258_ (.A1(_00964_),
    .A2(_06465_),
    .B(_00963_),
    .Y(_06528_));
 AND3x1_ASAP7_75t_R _18259_ (.A(_06511_),
    .B(_06527_),
    .C(_06528_),
    .Y(_04090_));
 OR3x1_ASAP7_75t_R _18260_ (.A(_00963_),
    .B(_00964_),
    .C(_06470_),
    .Y(_06529_));
 XOR2x2_ASAP7_75t_R _18261_ (.A(_00962_),
    .B(_06529_),
    .Y(_06530_));
 AND2x2_ASAP7_75t_R _18262_ (.A(_06506_),
    .B(_06530_),
    .Y(_04091_));
 OR4x1_ASAP7_75t_R _18263_ (.A(_00962_),
    .B(_00963_),
    .C(_00964_),
    .D(_06465_),
    .Y(_06531_));
 NAND2x1_ASAP7_75t_R _18264_ (.A(_00961_),
    .B(_06531_),
    .Y(_06532_));
 AND3x1_ASAP7_75t_R _18265_ (.A(_06511_),
    .B(_06467_),
    .C(_06532_),
    .Y(_04092_));
 XOR2x2_ASAP7_75t_R _18266_ (.A(_06453_),
    .B(_06471_),
    .Y(_06533_));
 AND2x2_ASAP7_75t_R _18267_ (.A(_06506_),
    .B(_06533_),
    .Y(_04093_));
 BUFx6f_ASAP7_75t_R _18268_ (.A(_00944_),
    .Y(_06534_));
 BUFx6f_ASAP7_75t_R _18269_ (.A(_00921_),
    .Y(_06535_));
 AND4x1_ASAP7_75t_R _18270_ (.A(_06535_),
    .B(_00949_),
    .C(_00950_),
    .D(_00951_),
    .Y(_06536_));
 AND5x1_ASAP7_75t_R _18271_ (.A(_00940_),
    .B(_00945_),
    .C(_00946_),
    .D(_00948_),
    .E(_06536_),
    .Y(_06537_));
 AND5x2_ASAP7_75t_R _18272_ (.A(_00942_),
    .B(_00943_),
    .C(_06534_),
    .D(_05995_),
    .E(_06537_),
    .Y(_06538_));
 BUFx3_ASAP7_75t_R _18273_ (.A(_00936_),
    .Y(_06539_));
 AND4x1_ASAP7_75t_R _18274_ (.A(_00935_),
    .B(_06539_),
    .C(_00937_),
    .D(_00938_),
    .Y(_06540_));
 AND4x1_ASAP7_75t_R _18275_ (.A(_00929_),
    .B(_00931_),
    .C(_00932_),
    .D(_00939_),
    .Y(_06541_));
 AND5x1_ASAP7_75t_R _18276_ (.A(_00922_),
    .B(_00923_),
    .C(_00928_),
    .D(_00947_),
    .E(_06541_),
    .Y(_06542_));
 AND3x1_ASAP7_75t_R _18277_ (.A(_00926_),
    .B(_00927_),
    .C(_00930_),
    .Y(_06543_));
 OR3x1_ASAP7_75t_R _18278_ (.A(_00924_),
    .B(_00925_),
    .C(_06543_),
    .Y(_06544_));
 AND5x2_ASAP7_75t_R _18279_ (.A(_00933_),
    .B(_00934_),
    .C(_06540_),
    .D(_06542_),
    .E(_06544_),
    .Y(_06545_));
 NAND2x2_ASAP7_75t_R _18280_ (.A(_06538_),
    .B(_06545_),
    .Y(_06546_));
 NOR2x1_ASAP7_75t_R _18281_ (.A(_00911_),
    .B(_06546_),
    .Y(_04094_));
 INVx1_ASAP7_75t_R _18282_ (.A(_06546_),
    .Y(_04095_));
 NOR2x1_ASAP7_75t_R _18283_ (.A(_00914_),
    .B(_06546_),
    .Y(_04096_));
 NOR2x1_ASAP7_75t_R _18284_ (.A(_00913_),
    .B(_06546_),
    .Y(_04097_));
 NOR2x1_ASAP7_75t_R _18285_ (.A(_00912_),
    .B(_06546_),
    .Y(_04098_));
 NOR2x1_ASAP7_75t_R _18286_ (.A(_00910_),
    .B(_06546_),
    .Y(_04099_));
 NOR2x1_ASAP7_75t_R _18287_ (.A(_00909_),
    .B(_06546_),
    .Y(_04100_));
 INVx1_ASAP7_75t_R _18288_ (.A(_06546_),
    .Y(_04101_));
 BUFx12f_ASAP7_75t_R _18289_ (.A(_08598_),
    .Y(_06547_));
 BUFx6f_ASAP7_75t_R _18290_ (.A(_06547_),
    .Y(_06548_));
 AND2x2_ASAP7_75t_R _18291_ (.A(_06548_),
    .B(_00046_),
    .Y(_04102_));
 OR4x1_ASAP7_75t_R _18292_ (.A(_00926_),
    .B(_00927_),
    .C(_00930_),
    .D(_02659_),
    .Y(_06549_));
 OR4x1_ASAP7_75t_R _18293_ (.A(_00922_),
    .B(_00923_),
    .C(_00924_),
    .D(_00925_),
    .Y(_06550_));
 OR2x6_ASAP7_75t_R _18294_ (.A(_06549_),
    .B(_06550_),
    .Y(_06551_));
 OR3x1_ASAP7_75t_R _18295_ (.A(_06535_),
    .B(_00951_),
    .C(_06551_),
    .Y(_06552_));
 OAI21x1_ASAP7_75t_R _18296_ (.A1(_06535_),
    .A2(_06551_),
    .B(_00951_),
    .Y(_06553_));
 AND3x1_ASAP7_75t_R _18297_ (.A(_06511_),
    .B(_06552_),
    .C(_06553_),
    .Y(_04103_));
 OR5x2_ASAP7_75t_R _18298_ (.A(_00926_),
    .B(_00927_),
    .C(_00930_),
    .D(_00941_),
    .E(_00046_),
    .Y(_06554_));
 OR2x6_ASAP7_75t_R _18299_ (.A(_06550_),
    .B(_06554_),
    .Y(_06555_));
 OR3x1_ASAP7_75t_R _18300_ (.A(_06535_),
    .B(_00951_),
    .C(_06555_),
    .Y(_06556_));
 XOR2x2_ASAP7_75t_R _18301_ (.A(_00950_),
    .B(_06556_),
    .Y(_06557_));
 AND2x2_ASAP7_75t_R _18302_ (.A(_06548_),
    .B(_06557_),
    .Y(_04104_));
 OR4x1_ASAP7_75t_R _18303_ (.A(_06535_),
    .B(_00950_),
    .C(_00951_),
    .D(_06551_),
    .Y(_06558_));
 XOR2x2_ASAP7_75t_R _18304_ (.A(_00949_),
    .B(_06558_),
    .Y(_06559_));
 AND2x2_ASAP7_75t_R _18305_ (.A(_06548_),
    .B(_06559_),
    .Y(_04105_));
 OR5x2_ASAP7_75t_R _18306_ (.A(_06535_),
    .B(_00948_),
    .C(_00949_),
    .D(_00950_),
    .E(_00951_),
    .Y(_06560_));
 OR5x1_ASAP7_75t_R _18307_ (.A(_06535_),
    .B(_00949_),
    .C(_00950_),
    .D(_00951_),
    .E(_06555_),
    .Y(_06561_));
 NAND2x1_ASAP7_75t_R _18308_ (.A(_00948_),
    .B(_06561_),
    .Y(_06562_));
 OA211x2_ASAP7_75t_R _18309_ (.A1(_06555_),
    .A2(_06560_),
    .B(_06562_),
    .C(_06433_),
    .Y(_04106_));
 OR3x1_ASAP7_75t_R _18310_ (.A(_06549_),
    .B(_06550_),
    .C(_06560_),
    .Y(_06563_));
 XOR2x2_ASAP7_75t_R _18311_ (.A(_00947_),
    .B(_06563_),
    .Y(_06564_));
 AND2x2_ASAP7_75t_R _18312_ (.A(_06548_),
    .B(_06564_),
    .Y(_04107_));
 OR3x1_ASAP7_75t_R _18313_ (.A(_00947_),
    .B(_06555_),
    .C(_06560_),
    .Y(_06565_));
 XOR2x2_ASAP7_75t_R _18314_ (.A(_00946_),
    .B(_06565_),
    .Y(_06566_));
 AND2x2_ASAP7_75t_R _18315_ (.A(_06548_),
    .B(_06566_),
    .Y(_04108_));
 OR4x1_ASAP7_75t_R _18316_ (.A(_00945_),
    .B(_00946_),
    .C(_00947_),
    .D(_06563_),
    .Y(_06567_));
 OR3x1_ASAP7_75t_R _18317_ (.A(_00946_),
    .B(_00947_),
    .C(_06563_),
    .Y(_06568_));
 NAND2x1_ASAP7_75t_R _18318_ (.A(_00945_),
    .B(_06568_),
    .Y(_06569_));
 AND3x1_ASAP7_75t_R _18319_ (.A(_06511_),
    .B(_06567_),
    .C(_06569_),
    .Y(_04109_));
 OR5x2_ASAP7_75t_R _18320_ (.A(_00945_),
    .B(_00946_),
    .C(_00947_),
    .D(_06555_),
    .E(_06560_),
    .Y(_06570_));
 XOR2x2_ASAP7_75t_R _18321_ (.A(_06534_),
    .B(_06570_),
    .Y(_06571_));
 AND2x2_ASAP7_75t_R _18322_ (.A(_06548_),
    .B(_06571_),
    .Y(_04110_));
 OR3x1_ASAP7_75t_R _18323_ (.A(_00943_),
    .B(_06534_),
    .C(_06567_),
    .Y(_06572_));
 OAI21x1_ASAP7_75t_R _18324_ (.A1(_06534_),
    .A2(_06567_),
    .B(_00943_),
    .Y(_06573_));
 AND3x1_ASAP7_75t_R _18325_ (.A(_06511_),
    .B(_06572_),
    .C(_06573_),
    .Y(_04111_));
 OR3x1_ASAP7_75t_R _18326_ (.A(_00943_),
    .B(_06534_),
    .C(_06570_),
    .Y(_06574_));
 XOR2x2_ASAP7_75t_R _18327_ (.A(_00942_),
    .B(_06574_),
    .Y(_06575_));
 AND2x2_ASAP7_75t_R _18328_ (.A(_06548_),
    .B(_06575_),
    .Y(_04112_));
 NOR2x1_ASAP7_75t_R _18329_ (.A(_06272_),
    .B(_02660_),
    .Y(_04113_));
 OR4x1_ASAP7_75t_R _18330_ (.A(_00942_),
    .B(_00943_),
    .C(_06534_),
    .D(_06567_),
    .Y(_06576_));
 XOR2x2_ASAP7_75t_R _18331_ (.A(_00940_),
    .B(_06576_),
    .Y(_06577_));
 AND2x2_ASAP7_75t_R _18332_ (.A(_06548_),
    .B(_06577_),
    .Y(_04114_));
 OR5x1_ASAP7_75t_R _18333_ (.A(_00940_),
    .B(_00942_),
    .C(_00943_),
    .D(_06534_),
    .E(_06570_),
    .Y(_06578_));
 XOR2x2_ASAP7_75t_R _18334_ (.A(_00939_),
    .B(_06578_),
    .Y(_06579_));
 AND2x2_ASAP7_75t_R _18335_ (.A(_06548_),
    .B(_06579_),
    .Y(_04115_));
 OR5x2_ASAP7_75t_R _18336_ (.A(_00939_),
    .B(_00940_),
    .C(_00942_),
    .D(_00943_),
    .E(_06534_),
    .Y(_06580_));
 OR3x1_ASAP7_75t_R _18337_ (.A(_00938_),
    .B(_06567_),
    .C(_06580_),
    .Y(_06581_));
 OAI21x1_ASAP7_75t_R _18338_ (.A1(_06567_),
    .A2(_06580_),
    .B(_00938_),
    .Y(_06582_));
 AND3x1_ASAP7_75t_R _18339_ (.A(_06511_),
    .B(_06581_),
    .C(_06582_),
    .Y(_04116_));
 OR4x1_ASAP7_75t_R _18340_ (.A(_00937_),
    .B(_00938_),
    .C(_06570_),
    .D(_06580_),
    .Y(_06583_));
 OR3x1_ASAP7_75t_R _18341_ (.A(_00938_),
    .B(_06570_),
    .C(_06580_),
    .Y(_06584_));
 NAND2x1_ASAP7_75t_R _18342_ (.A(_00937_),
    .B(_06584_),
    .Y(_06585_));
 AND3x1_ASAP7_75t_R _18343_ (.A(_06511_),
    .B(_06583_),
    .C(_06585_),
    .Y(_04117_));
 OR4x1_ASAP7_75t_R _18344_ (.A(_00937_),
    .B(_00938_),
    .C(_06567_),
    .D(_06580_),
    .Y(_06586_));
 XOR2x2_ASAP7_75t_R _18345_ (.A(_06539_),
    .B(_06586_),
    .Y(_06587_));
 AND2x2_ASAP7_75t_R _18346_ (.A(_06548_),
    .B(_06587_),
    .Y(_04118_));
 OR3x1_ASAP7_75t_R _18347_ (.A(_00935_),
    .B(_06539_),
    .C(_06583_),
    .Y(_06588_));
 OAI21x1_ASAP7_75t_R _18348_ (.A1(_06539_),
    .A2(_06583_),
    .B(_00935_),
    .Y(_06589_));
 AND3x1_ASAP7_75t_R _18349_ (.A(_06511_),
    .B(_06588_),
    .C(_06589_),
    .Y(_04119_));
 BUFx6f_ASAP7_75t_R _18350_ (.A(_06547_),
    .Y(_06590_));
 OR3x1_ASAP7_75t_R _18351_ (.A(_00935_),
    .B(_06539_),
    .C(_06586_),
    .Y(_06591_));
 XOR2x2_ASAP7_75t_R _18352_ (.A(_00934_),
    .B(_06591_),
    .Y(_06592_));
 AND2x2_ASAP7_75t_R _18353_ (.A(_06590_),
    .B(_06592_),
    .Y(_04120_));
 OR4x1_ASAP7_75t_R _18354_ (.A(_00934_),
    .B(_00935_),
    .C(_06539_),
    .D(_06583_),
    .Y(_06593_));
 XOR2x2_ASAP7_75t_R _18355_ (.A(_00933_),
    .B(_06593_),
    .Y(_06594_));
 AND2x2_ASAP7_75t_R _18356_ (.A(_06590_),
    .B(_06594_),
    .Y(_04121_));
 OR5x1_ASAP7_75t_R _18357_ (.A(_00933_),
    .B(_00934_),
    .C(_00935_),
    .D(_06539_),
    .E(_06586_),
    .Y(_06595_));
 XOR2x2_ASAP7_75t_R _18358_ (.A(_00932_),
    .B(_06595_),
    .Y(_06596_));
 AND2x2_ASAP7_75t_R _18359_ (.A(_06590_),
    .B(_06596_),
    .Y(_04122_));
 BUFx6f_ASAP7_75t_R _18360_ (.A(_06386_),
    .Y(_06597_));
 OR5x2_ASAP7_75t_R _18361_ (.A(_00932_),
    .B(_00933_),
    .C(_00934_),
    .D(_00935_),
    .E(_06539_),
    .Y(_06598_));
 OR3x1_ASAP7_75t_R _18362_ (.A(_00931_),
    .B(_06583_),
    .C(_06598_),
    .Y(_06599_));
 OAI21x1_ASAP7_75t_R _18363_ (.A1(_06583_),
    .A2(_06598_),
    .B(_00931_),
    .Y(_06600_));
 AND3x1_ASAP7_75t_R _18364_ (.A(_06597_),
    .B(_06599_),
    .C(_06600_),
    .Y(_04123_));
 XOR2x2_ASAP7_75t_R _18365_ (.A(_00930_),
    .B(_02659_),
    .Y(_06601_));
 AND2x2_ASAP7_75t_R _18366_ (.A(_06590_),
    .B(_06601_),
    .Y(_04124_));
 OR3x1_ASAP7_75t_R _18367_ (.A(_00931_),
    .B(_06586_),
    .C(_06598_),
    .Y(_06602_));
 XOR2x2_ASAP7_75t_R _18368_ (.A(_00929_),
    .B(_06602_),
    .Y(_06603_));
 AND2x2_ASAP7_75t_R _18369_ (.A(_06590_),
    .B(_06603_),
    .Y(_04125_));
 OR4x1_ASAP7_75t_R _18370_ (.A(_00929_),
    .B(_00931_),
    .C(_06583_),
    .D(_06598_),
    .Y(_06604_));
 XOR2x2_ASAP7_75t_R _18371_ (.A(_00928_),
    .B(_06604_),
    .Y(_06605_));
 AND2x2_ASAP7_75t_R _18372_ (.A(_06590_),
    .B(_06605_),
    .Y(_04126_));
 OR3x1_ASAP7_75t_R _18373_ (.A(_00930_),
    .B(_00941_),
    .C(_00046_),
    .Y(_06606_));
 XOR2x2_ASAP7_75t_R _18374_ (.A(_00927_),
    .B(_06606_),
    .Y(_06607_));
 AND2x2_ASAP7_75t_R _18375_ (.A(_06590_),
    .B(_06607_),
    .Y(_04127_));
 OR3x1_ASAP7_75t_R _18376_ (.A(_00927_),
    .B(_00930_),
    .C(_02659_),
    .Y(_06608_));
 NAND2x1_ASAP7_75t_R _18377_ (.A(_00926_),
    .B(_06608_),
    .Y(_06609_));
 AND3x1_ASAP7_75t_R _18378_ (.A(_06597_),
    .B(_06549_),
    .C(_06609_),
    .Y(_04128_));
 XOR2x2_ASAP7_75t_R _18379_ (.A(_00925_),
    .B(_06554_),
    .Y(_06610_));
 AND2x2_ASAP7_75t_R _18380_ (.A(_06590_),
    .B(_06610_),
    .Y(_04129_));
 OR3x1_ASAP7_75t_R _18381_ (.A(_00924_),
    .B(_00925_),
    .C(_06549_),
    .Y(_06611_));
 OAI21x1_ASAP7_75t_R _18382_ (.A1(_00925_),
    .A2(_06549_),
    .B(_00924_),
    .Y(_06612_));
 AND3x1_ASAP7_75t_R _18383_ (.A(_06597_),
    .B(_06611_),
    .C(_06612_),
    .Y(_04130_));
 OR3x1_ASAP7_75t_R _18384_ (.A(_00924_),
    .B(_00925_),
    .C(_06554_),
    .Y(_06613_));
 XOR2x2_ASAP7_75t_R _18385_ (.A(_00923_),
    .B(_06613_),
    .Y(_06614_));
 AND2x2_ASAP7_75t_R _18386_ (.A(_06590_),
    .B(_06614_),
    .Y(_04131_));
 OR4x1_ASAP7_75t_R _18387_ (.A(_00923_),
    .B(_00924_),
    .C(_00925_),
    .D(_06549_),
    .Y(_06615_));
 NAND2x1_ASAP7_75t_R _18388_ (.A(_00922_),
    .B(_06615_),
    .Y(_06616_));
 AND3x1_ASAP7_75t_R _18389_ (.A(_06597_),
    .B(_06551_),
    .C(_06616_),
    .Y(_04132_));
 XOR2x2_ASAP7_75t_R _18390_ (.A(_06535_),
    .B(_06555_),
    .Y(_06617_));
 AND2x2_ASAP7_75t_R _18391_ (.A(_06590_),
    .B(_06617_),
    .Y(_04133_));
 BUFx6f_ASAP7_75t_R _18392_ (.A(_06547_),
    .Y(_06618_));
 AND2x2_ASAP7_75t_R _18393_ (.A(_06618_),
    .B(_00022_),
    .Y(_04134_));
 AND2x4_ASAP7_75t_R _18394_ (.A(_00953_),
    .B(_00954_),
    .Y(_06619_));
 AND5x2_ASAP7_75t_R _18395_ (.A(\xs[1].cli1.i[39] ),
    .B(_00955_),
    .C(\xs[1].cli1.i[33] ),
    .D(_00957_),
    .E(_06619_),
    .Y(_06620_));
 INVx1_ASAP7_75t_R _18396_ (.A(_02323_),
    .Y(_06621_));
 NAND2x1_ASAP7_75t_R _18397_ (.A(_00953_),
    .B(_00954_),
    .Y(_06622_));
 OR5x1_ASAP7_75t_R _18398_ (.A(_00952_),
    .B(\xs[1].cli1.i[34] ),
    .C(_00956_),
    .D(\xs[1].cli1.i[32] ),
    .E(_06622_),
    .Y(_06623_));
 AO31x2_ASAP7_75t_R _18399_ (.A1(_00955_),
    .A2(\xs[1].cli1.i[33] ),
    .A3(_06619_),
    .B(_00952_),
    .Y(_06624_));
 AO221x1_ASAP7_75t_R _18400_ (.A1(_02317_),
    .A2(_06621_),
    .B1(_06623_),
    .B2(_06624_),
    .C(_02316_),
    .Y(_06625_));
 AND2x4_ASAP7_75t_R _18401_ (.A(_00992_),
    .B(_00993_),
    .Y(_06626_));
 AND3x4_ASAP7_75t_R _18402_ (.A(_00994_),
    .B(\peo[2][33] ),
    .C(_06626_),
    .Y(_06627_));
 OA22x2_ASAP7_75t_R _18403_ (.A1(_02317_),
    .A2(_06624_),
    .B1(_06627_),
    .B2(_00991_),
    .Y(_06628_));
 INVx2_ASAP7_75t_R _18404_ (.A(_02316_),
    .Y(_06629_));
 INVx1_ASAP7_75t_R _18405_ (.A(_00022_),
    .Y(_06630_));
 OR5x1_ASAP7_75t_R _18406_ (.A(_06629_),
    .B(_06630_),
    .C(_00991_),
    .D(_06624_),
    .E(_06627_),
    .Y(_06631_));
 OA21x2_ASAP7_75t_R _18407_ (.A1(_06625_),
    .A2(_06628_),
    .B(_06631_),
    .Y(_06632_));
 AND2x2_ASAP7_75t_R _18408_ (.A(_06620_),
    .B(_06632_),
    .Y(_06633_));
 NOR2x1_ASAP7_75t_R _18409_ (.A(_00991_),
    .B(_00996_),
    .Y(_06634_));
 AND5x1_ASAP7_75t_R _18410_ (.A(_00994_),
    .B(\peo[2][33] ),
    .C(_06621_),
    .D(_06626_),
    .E(_06634_),
    .Y(_06635_));
 AO32x1_ASAP7_75t_R _18411_ (.A1(_06620_),
    .A2(_06627_),
    .A3(_06634_),
    .B1(_06635_),
    .B2(_06624_),
    .Y(_06636_));
 OA211x2_ASAP7_75t_R _18412_ (.A1(_00991_),
    .A2(_06627_),
    .B(_06620_),
    .C(_02323_),
    .Y(_06637_));
 NOR2x1_ASAP7_75t_R _18413_ (.A(_06636_),
    .B(_06637_),
    .Y(_06638_));
 AND4x1_ASAP7_75t_R _18414_ (.A(_06629_),
    .B(_02317_),
    .C(_02323_),
    .D(_06638_),
    .Y(_06639_));
 OR3x1_ASAP7_75t_R _18415_ (.A(\peo[2][0] ),
    .B(_06633_),
    .C(_06639_),
    .Y(_06640_));
 AOI22x1_ASAP7_75t_R _18416_ (.A1(_00959_),
    .A2(_06633_),
    .B1(_06639_),
    .B2(_02327_),
    .Y(_06641_));
 AND3x1_ASAP7_75t_R _18417_ (.A(_06597_),
    .B(_06640_),
    .C(_06641_),
    .Y(_04135_));
 NAND2x2_ASAP7_75t_R _18418_ (.A(_08528_),
    .B(_06639_),
    .Y(_06642_));
 NOR2x1_ASAP7_75t_R _18419_ (.A(_02326_),
    .B(_06642_),
    .Y(_04136_));
 NOR2x1_ASAP7_75t_R _18420_ (.A(_02325_),
    .B(_06642_),
    .Y(_04137_));
 NOR2x1_ASAP7_75t_R _18421_ (.A(_02324_),
    .B(_06642_),
    .Y(_04138_));
 NOR2x1_ASAP7_75t_R _18422_ (.A(_02315_),
    .B(_06642_),
    .Y(_04139_));
 NOR2x1_ASAP7_75t_R _18423_ (.A(_02314_),
    .B(_06642_),
    .Y(_04140_));
 NOR2x1_ASAP7_75t_R _18424_ (.A(_00959_),
    .B(_06632_),
    .Y(_06643_));
 NAND2x1_ASAP7_75t_R _18425_ (.A(_06629_),
    .B(_02317_),
    .Y(_06644_));
 AND4x1_ASAP7_75t_R _18426_ (.A(_00994_),
    .B(\peo[2][33] ),
    .C(_06626_),
    .D(_06634_),
    .Y(_06645_));
 AO21x1_ASAP7_75t_R _18427_ (.A1(_06624_),
    .A2(_06645_),
    .B(_02323_),
    .Y(_06646_));
 OR4x1_ASAP7_75t_R _18428_ (.A(_06644_),
    .B(_06636_),
    .C(_06637_),
    .D(_06646_),
    .Y(_06647_));
 NOR2x1_ASAP7_75t_R _18429_ (.A(_02327_),
    .B(_06647_),
    .Y(_06648_));
 AND3x1_ASAP7_75t_R _18430_ (.A(\peo[2][0] ),
    .B(_06632_),
    .C(_06647_),
    .Y(_06649_));
 OR3x1_ASAP7_75t_R _18431_ (.A(_06643_),
    .B(_06648_),
    .C(_06649_),
    .Y(_06650_));
 AND2x2_ASAP7_75t_R _18432_ (.A(_06618_),
    .B(_06650_),
    .Y(_04141_));
 OR2x2_ASAP7_75t_R _18433_ (.A(_08683_),
    .B(_06647_),
    .Y(_06651_));
 BUFx3_ASAP7_75t_R _18434_ (.A(_06651_),
    .Y(_06652_));
 NOR2x1_ASAP7_75t_R _18435_ (.A(_02326_),
    .B(_06652_),
    .Y(_04142_));
 NOR2x1_ASAP7_75t_R _18436_ (.A(_02325_),
    .B(_06652_),
    .Y(_04143_));
 NOR2x1_ASAP7_75t_R _18437_ (.A(_02324_),
    .B(_06652_),
    .Y(_04144_));
 NOR2x1_ASAP7_75t_R _18438_ (.A(_02315_),
    .B(_06652_),
    .Y(_04145_));
 NOR2x1_ASAP7_75t_R _18439_ (.A(_02314_),
    .B(_06652_),
    .Y(_04146_));
 AO21x2_ASAP7_75t_R _18440_ (.A1(_02317_),
    .A2(_06638_),
    .B(_02316_),
    .Y(_06653_));
 BUFx6f_ASAP7_75t_R _18441_ (.A(_06653_),
    .Y(_06654_));
 NOR2x1_ASAP7_75t_R _18442_ (.A(_02327_),
    .B(_06654_),
    .Y(_06655_));
 NAND2x1_ASAP7_75t_R _18443_ (.A(_00992_),
    .B(_00993_),
    .Y(_06656_));
 OA31x2_ASAP7_75t_R _18444_ (.A1(\peo[2][34] ),
    .A2(_00995_),
    .A3(_06656_),
    .B1(\peo[2][39] ),
    .Y(_06657_));
 AND2x2_ASAP7_75t_R _18445_ (.A(_02316_),
    .B(_00022_),
    .Y(_06658_));
 INVx1_ASAP7_75t_R _18446_ (.A(_02317_),
    .Y(_06659_));
 AO21x1_ASAP7_75t_R _18447_ (.A1(_02323_),
    .A2(_06657_),
    .B(_06659_),
    .Y(_06660_));
 AO221x1_ASAP7_75t_R _18448_ (.A1(_06657_),
    .A2(_06658_),
    .B1(_06660_),
    .B2(_06629_),
    .C(_06624_),
    .Y(_06661_));
 BUFx6f_ASAP7_75t_R _18449_ (.A(_06661_),
    .Y(_06662_));
 NAND2x1_ASAP7_75t_R _18450_ (.A(_00998_),
    .B(_06662_),
    .Y(_06663_));
 OA211x2_ASAP7_75t_R _18451_ (.A1(\peo[3][0] ),
    .A2(_06662_),
    .B(_06663_),
    .C(_06654_),
    .Y(_06664_));
 OA21x2_ASAP7_75t_R _18452_ (.A1(_06655_),
    .A2(_06664_),
    .B(_11397_),
    .Y(_04147_));
 OR2x2_ASAP7_75t_R _18453_ (.A(_09220_),
    .B(_06653_),
    .Y(_06665_));
 BUFx6f_ASAP7_75t_R _18454_ (.A(_06665_),
    .Y(_06666_));
 NOR2x1_ASAP7_75t_R _18455_ (.A(_02326_),
    .B(_06666_),
    .Y(_04148_));
 NOR2x1_ASAP7_75t_R _18456_ (.A(_02325_),
    .B(_06666_),
    .Y(_04149_));
 NOR2x1_ASAP7_75t_R _18457_ (.A(_02324_),
    .B(_06666_),
    .Y(_04150_));
 NOR2x1_ASAP7_75t_R _18458_ (.A(_02323_),
    .B(_06654_),
    .Y(_06667_));
 NAND2x1_ASAP7_75t_R _18459_ (.A(_00996_),
    .B(_06662_),
    .Y(_06668_));
 OA211x2_ASAP7_75t_R _18460_ (.A1(\xs[1].cli1.i[32] ),
    .A2(_06662_),
    .B(_06668_),
    .C(_06654_),
    .Y(_06669_));
 OA21x2_ASAP7_75t_R _18461_ (.A1(_06667_),
    .A2(_06669_),
    .B(_11397_),
    .Y(_04151_));
 NOR2x1_ASAP7_75t_R _18462_ (.A(_02322_),
    .B(_06654_),
    .Y(_06670_));
 NAND2x1_ASAP7_75t_R _18463_ (.A(_00995_),
    .B(_06662_),
    .Y(_06671_));
 OA211x2_ASAP7_75t_R _18464_ (.A1(\xs[1].cli1.i[33] ),
    .A2(_06662_),
    .B(_06671_),
    .C(_06654_),
    .Y(_06672_));
 OA21x2_ASAP7_75t_R _18465_ (.A1(_06670_),
    .A2(_06672_),
    .B(_11397_),
    .Y(_04152_));
 NOR2x1_ASAP7_75t_R _18466_ (.A(_02321_),
    .B(_06654_),
    .Y(_06673_));
 NAND2x1_ASAP7_75t_R _18467_ (.A(_00994_),
    .B(_06662_),
    .Y(_06674_));
 OA211x2_ASAP7_75t_R _18468_ (.A1(\xs[1].cli1.i[34] ),
    .A2(_06662_),
    .B(_06674_),
    .C(_06653_),
    .Y(_06675_));
 BUFx12f_ASAP7_75t_R _18469_ (.A(_09229_),
    .Y(_06676_));
 OA21x2_ASAP7_75t_R _18470_ (.A1(_06673_),
    .A2(_06675_),
    .B(_06676_),
    .Y(_04153_));
 NOR2x1_ASAP7_75t_R _18471_ (.A(_02320_),
    .B(_06654_),
    .Y(_06677_));
 NAND2x1_ASAP7_75t_R _18472_ (.A(_00993_),
    .B(_06661_),
    .Y(_06678_));
 OA211x2_ASAP7_75t_R _18473_ (.A1(\xs[1].cli1.i[35] ),
    .A2(_06662_),
    .B(_06678_),
    .C(_06653_),
    .Y(_06679_));
 OA21x2_ASAP7_75t_R _18474_ (.A1(_06677_),
    .A2(_06679_),
    .B(_06676_),
    .Y(_04154_));
 NOR2x1_ASAP7_75t_R _18475_ (.A(_02319_),
    .B(_06654_),
    .Y(_06680_));
 NAND2x1_ASAP7_75t_R _18476_ (.A(_00992_),
    .B(_06661_),
    .Y(_06681_));
 OA211x2_ASAP7_75t_R _18477_ (.A1(\xs[1].cli1.i[36] ),
    .A2(_06662_),
    .B(_06681_),
    .C(_06653_),
    .Y(_06682_));
 OA21x2_ASAP7_75t_R _18478_ (.A1(_06680_),
    .A2(_06682_),
    .B(_06676_),
    .Y(_04155_));
 NOR2x1_ASAP7_75t_R _18479_ (.A(_02318_),
    .B(_06666_),
    .Y(_04156_));
 AO21x1_ASAP7_75t_R _18480_ (.A1(_06621_),
    .A2(_06624_),
    .B(_06620_),
    .Y(_06683_));
 AO32x1_ASAP7_75t_R _18481_ (.A1(\peo[2][39] ),
    .A2(\peo[2][32] ),
    .A3(_06683_),
    .B1(_06620_),
    .B2(_02323_),
    .Y(_06684_));
 AO32x1_ASAP7_75t_R _18482_ (.A1(_00991_),
    .A2(_02323_),
    .A3(_06620_),
    .B1(_06627_),
    .B2(_06684_),
    .Y(_06685_));
 AND4x1_ASAP7_75t_R _18483_ (.A(_08999_),
    .B(_06629_),
    .C(_02317_),
    .D(_06685_),
    .Y(_04157_));
 OA211x2_ASAP7_75t_R _18484_ (.A1(_00991_),
    .A2(_06627_),
    .B(_06654_),
    .C(_06624_),
    .Y(_06686_));
 NOR2x1_ASAP7_75t_R _18485_ (.A(_06272_),
    .B(_06686_),
    .Y(_04158_));
 NOR2x1_ASAP7_75t_R _18486_ (.A(_02315_),
    .B(_06666_),
    .Y(_04159_));
 NOR2x1_ASAP7_75t_R _18487_ (.A(_02314_),
    .B(_06666_),
    .Y(_04160_));
 BUFx3_ASAP7_75t_R _18488_ (.A(_00883_),
    .Y(_06687_));
 BUFx3_ASAP7_75t_R _18489_ (.A(_00856_),
    .Y(_06688_));
 AND4x1_ASAP7_75t_R _18490_ (.A(_06688_),
    .B(_00884_),
    .C(_00885_),
    .D(_00886_),
    .Y(_06689_));
 AND5x1_ASAP7_75t_R _18491_ (.A(_00875_),
    .B(_00880_),
    .C(_00881_),
    .D(_06687_),
    .E(_06689_),
    .Y(_06690_));
 AND5x2_ASAP7_75t_R _18492_ (.A(_00877_),
    .B(_00878_),
    .C(_00879_),
    .D(_05995_),
    .E(_06690_),
    .Y(_06691_));
 AND4x1_ASAP7_75t_R _18493_ (.A(_00870_),
    .B(_00871_),
    .C(_00872_),
    .D(_00873_),
    .Y(_06692_));
 AND4x1_ASAP7_75t_R _18494_ (.A(_00864_),
    .B(_00866_),
    .C(_00867_),
    .D(_00874_),
    .Y(_06693_));
 AND5x1_ASAP7_75t_R _18495_ (.A(_00857_),
    .B(_00858_),
    .C(_00863_),
    .D(_00882_),
    .E(_06693_),
    .Y(_06694_));
 AND3x1_ASAP7_75t_R _18496_ (.A(_00861_),
    .B(_00862_),
    .C(_00865_),
    .Y(_06695_));
 OR3x1_ASAP7_75t_R _18497_ (.A(_00859_),
    .B(_00860_),
    .C(_06695_),
    .Y(_06696_));
 AND5x2_ASAP7_75t_R _18498_ (.A(_00868_),
    .B(_00869_),
    .C(_06692_),
    .D(_06694_),
    .E(_06696_),
    .Y(_06697_));
 NAND2x2_ASAP7_75t_R _18499_ (.A(_06691_),
    .B(_06697_),
    .Y(_06698_));
 NOR2x1_ASAP7_75t_R _18500_ (.A(_00813_),
    .B(_06698_),
    .Y(_04161_));
 INVx1_ASAP7_75t_R _18501_ (.A(_06698_),
    .Y(_04162_));
 NOR2x1_ASAP7_75t_R _18502_ (.A(_00816_),
    .B(_06698_),
    .Y(_04163_));
 NOR2x1_ASAP7_75t_R _18503_ (.A(_00815_),
    .B(_06698_),
    .Y(_04164_));
 NOR2x1_ASAP7_75t_R _18504_ (.A(_00814_),
    .B(_06698_),
    .Y(_04165_));
 NOR2x1_ASAP7_75t_R _18505_ (.A(_00812_),
    .B(_06698_),
    .Y(_04166_));
 NOR2x1_ASAP7_75t_R _18506_ (.A(_00811_),
    .B(_06698_),
    .Y(_04167_));
 INVx1_ASAP7_75t_R _18507_ (.A(_06698_),
    .Y(_04168_));
 AND2x2_ASAP7_75t_R _18508_ (.A(_06618_),
    .B(_00047_),
    .Y(_04169_));
 OR4x1_ASAP7_75t_R _18509_ (.A(_00861_),
    .B(_00862_),
    .C(_00865_),
    .D(_02669_),
    .Y(_06699_));
 OR4x1_ASAP7_75t_R _18510_ (.A(_00857_),
    .B(_00858_),
    .C(_00859_),
    .D(_00860_),
    .Y(_06700_));
 OR2x6_ASAP7_75t_R _18511_ (.A(_06699_),
    .B(_06700_),
    .Y(_06701_));
 OR3x1_ASAP7_75t_R _18512_ (.A(_06688_),
    .B(_00886_),
    .C(_06701_),
    .Y(_06702_));
 OAI21x1_ASAP7_75t_R _18513_ (.A1(_06688_),
    .A2(_06701_),
    .B(_00886_),
    .Y(_06703_));
 AND3x1_ASAP7_75t_R _18514_ (.A(_06597_),
    .B(_06702_),
    .C(_06703_),
    .Y(_04170_));
 OR5x2_ASAP7_75t_R _18515_ (.A(_00861_),
    .B(_00862_),
    .C(_00865_),
    .D(_00876_),
    .E(_00047_),
    .Y(_06704_));
 OR2x2_ASAP7_75t_R _18516_ (.A(_06700_),
    .B(_06704_),
    .Y(_06705_));
 OR3x1_ASAP7_75t_R _18517_ (.A(_06688_),
    .B(_00886_),
    .C(_06705_),
    .Y(_06706_));
 XOR2x2_ASAP7_75t_R _18518_ (.A(_00885_),
    .B(_06706_),
    .Y(_06707_));
 AND2x2_ASAP7_75t_R _18519_ (.A(_06618_),
    .B(_06707_),
    .Y(_04171_));
 OR4x1_ASAP7_75t_R _18520_ (.A(_06688_),
    .B(_00884_),
    .C(_00885_),
    .D(_00886_),
    .Y(_06708_));
 OR3x2_ASAP7_75t_R _18521_ (.A(_06699_),
    .B(_06700_),
    .C(_06708_),
    .Y(_06709_));
 OR4x1_ASAP7_75t_R _18522_ (.A(_06688_),
    .B(_00885_),
    .C(_00886_),
    .D(_06701_),
    .Y(_06710_));
 NAND2x1_ASAP7_75t_R _18523_ (.A(_00884_),
    .B(_06710_),
    .Y(_06711_));
 AND3x1_ASAP7_75t_R _18524_ (.A(_06597_),
    .B(_06709_),
    .C(_06711_),
    .Y(_04172_));
 OR3x2_ASAP7_75t_R _18525_ (.A(_06700_),
    .B(_06704_),
    .C(_06708_),
    .Y(_06712_));
 XOR2x2_ASAP7_75t_R _18526_ (.A(_06687_),
    .B(_06712_),
    .Y(_06713_));
 AND2x2_ASAP7_75t_R _18527_ (.A(_06618_),
    .B(_06713_),
    .Y(_04173_));
 OR3x1_ASAP7_75t_R _18528_ (.A(_00882_),
    .B(_06687_),
    .C(_06709_),
    .Y(_06714_));
 OAI21x1_ASAP7_75t_R _18529_ (.A1(_06687_),
    .A2(_06709_),
    .B(_00882_),
    .Y(_06715_));
 AND3x1_ASAP7_75t_R _18530_ (.A(_06597_),
    .B(_06714_),
    .C(_06715_),
    .Y(_04174_));
 OR3x1_ASAP7_75t_R _18531_ (.A(_00882_),
    .B(_06687_),
    .C(_06712_),
    .Y(_06716_));
 XOR2x2_ASAP7_75t_R _18532_ (.A(_00881_),
    .B(_06716_),
    .Y(_06717_));
 AND2x2_ASAP7_75t_R _18533_ (.A(_06618_),
    .B(_06717_),
    .Y(_04175_));
 OR4x1_ASAP7_75t_R _18534_ (.A(_00881_),
    .B(_00882_),
    .C(_06687_),
    .D(_06709_),
    .Y(_06718_));
 XOR2x2_ASAP7_75t_R _18535_ (.A(_00880_),
    .B(_06718_),
    .Y(_06719_));
 AND2x2_ASAP7_75t_R _18536_ (.A(_06618_),
    .B(_06719_),
    .Y(_04176_));
 OR5x1_ASAP7_75t_R _18537_ (.A(_00880_),
    .B(_00881_),
    .C(_00882_),
    .D(_06687_),
    .E(_06712_),
    .Y(_06720_));
 XOR2x2_ASAP7_75t_R _18538_ (.A(_00879_),
    .B(_06720_),
    .Y(_06721_));
 AND2x2_ASAP7_75t_R _18539_ (.A(_06618_),
    .B(_06721_),
    .Y(_04177_));
 OR5x2_ASAP7_75t_R _18540_ (.A(_00879_),
    .B(_00880_),
    .C(_00881_),
    .D(_00882_),
    .E(_06687_),
    .Y(_06722_));
 OR3x2_ASAP7_75t_R _18541_ (.A(_00878_),
    .B(_06709_),
    .C(_06722_),
    .Y(_06723_));
 OAI21x1_ASAP7_75t_R _18542_ (.A1(_06709_),
    .A2(_06722_),
    .B(_00878_),
    .Y(_06724_));
 AND3x1_ASAP7_75t_R _18543_ (.A(_06597_),
    .B(_06723_),
    .C(_06724_),
    .Y(_04178_));
 OR3x2_ASAP7_75t_R _18544_ (.A(_00878_),
    .B(_06712_),
    .C(_06722_),
    .Y(_06725_));
 XOR2x2_ASAP7_75t_R _18545_ (.A(_00877_),
    .B(_06725_),
    .Y(_06726_));
 AND2x2_ASAP7_75t_R _18546_ (.A(_06618_),
    .B(_06726_),
    .Y(_04179_));
 NOR2x1_ASAP7_75t_R _18547_ (.A(_06272_),
    .B(_02670_),
    .Y(_04180_));
 OR3x1_ASAP7_75t_R _18548_ (.A(_00875_),
    .B(_00877_),
    .C(_06723_),
    .Y(_06727_));
 OAI21x1_ASAP7_75t_R _18549_ (.A1(_00877_),
    .A2(_06723_),
    .B(_00875_),
    .Y(_06728_));
 AND3x1_ASAP7_75t_R _18550_ (.A(_06597_),
    .B(_06727_),
    .C(_06728_),
    .Y(_04181_));
 OR3x1_ASAP7_75t_R _18551_ (.A(_00875_),
    .B(_00877_),
    .C(_06725_),
    .Y(_06729_));
 XOR2x2_ASAP7_75t_R _18552_ (.A(_00874_),
    .B(_06729_),
    .Y(_06730_));
 AND2x2_ASAP7_75t_R _18553_ (.A(_06618_),
    .B(_06730_),
    .Y(_04182_));
 BUFx6f_ASAP7_75t_R _18554_ (.A(_06547_),
    .Y(_06731_));
 OR4x1_ASAP7_75t_R _18555_ (.A(_00874_),
    .B(_00875_),
    .C(_00877_),
    .D(_06723_),
    .Y(_06732_));
 XOR2x2_ASAP7_75t_R _18556_ (.A(_00873_),
    .B(_06732_),
    .Y(_06733_));
 AND2x2_ASAP7_75t_R _18557_ (.A(_06731_),
    .B(_06733_),
    .Y(_04183_));
 BUFx6f_ASAP7_75t_R _18558_ (.A(_06386_),
    .Y(_06734_));
 OR4x1_ASAP7_75t_R _18559_ (.A(_00873_),
    .B(_00874_),
    .C(_00875_),
    .D(_00877_),
    .Y(_06735_));
 OR3x2_ASAP7_75t_R _18560_ (.A(_00872_),
    .B(_06725_),
    .C(_06735_),
    .Y(_06736_));
 OAI21x1_ASAP7_75t_R _18561_ (.A1(_06725_),
    .A2(_06735_),
    .B(_00872_),
    .Y(_06737_));
 AND3x1_ASAP7_75t_R _18562_ (.A(_06734_),
    .B(_06736_),
    .C(_06737_),
    .Y(_04184_));
 OR3x2_ASAP7_75t_R _18563_ (.A(_00872_),
    .B(_06723_),
    .C(_06735_),
    .Y(_06738_));
 XOR2x2_ASAP7_75t_R _18564_ (.A(_00871_),
    .B(_06738_),
    .Y(_06739_));
 AND2x2_ASAP7_75t_R _18565_ (.A(_06731_),
    .B(_06739_),
    .Y(_04185_));
 OR3x1_ASAP7_75t_R _18566_ (.A(_00870_),
    .B(_00871_),
    .C(_06736_),
    .Y(_06740_));
 OAI21x1_ASAP7_75t_R _18567_ (.A1(_00871_),
    .A2(_06736_),
    .B(_00870_),
    .Y(_06741_));
 AND3x1_ASAP7_75t_R _18568_ (.A(_06734_),
    .B(_06740_),
    .C(_06741_),
    .Y(_04186_));
 OR3x1_ASAP7_75t_R _18569_ (.A(_00870_),
    .B(_00871_),
    .C(_06738_),
    .Y(_06742_));
 XOR2x2_ASAP7_75t_R _18570_ (.A(_00869_),
    .B(_06742_),
    .Y(_06743_));
 AND2x2_ASAP7_75t_R _18571_ (.A(_06731_),
    .B(_06743_),
    .Y(_04187_));
 OR4x1_ASAP7_75t_R _18572_ (.A(_00869_),
    .B(_00870_),
    .C(_00871_),
    .D(_06736_),
    .Y(_06744_));
 XOR2x2_ASAP7_75t_R _18573_ (.A(_00868_),
    .B(_06744_),
    .Y(_06745_));
 AND2x2_ASAP7_75t_R _18574_ (.A(_06731_),
    .B(_06745_),
    .Y(_04188_));
 OR4x1_ASAP7_75t_R _18575_ (.A(_00868_),
    .B(_00869_),
    .C(_00870_),
    .D(_00871_),
    .Y(_06746_));
 OR3x1_ASAP7_75t_R _18576_ (.A(_00867_),
    .B(_06738_),
    .C(_06746_),
    .Y(_06747_));
 OAI21x1_ASAP7_75t_R _18577_ (.A1(_06738_),
    .A2(_06746_),
    .B(_00867_),
    .Y(_06748_));
 AND3x1_ASAP7_75t_R _18578_ (.A(_06734_),
    .B(_06747_),
    .C(_06748_),
    .Y(_04189_));
 OR3x1_ASAP7_75t_R _18579_ (.A(_00867_),
    .B(_06736_),
    .C(_06746_),
    .Y(_06749_));
 XOR2x2_ASAP7_75t_R _18580_ (.A(_00866_),
    .B(_06749_),
    .Y(_06750_));
 AND2x2_ASAP7_75t_R _18581_ (.A(_06731_),
    .B(_06750_),
    .Y(_04190_));
 XOR2x2_ASAP7_75t_R _18582_ (.A(_00865_),
    .B(_02669_),
    .Y(_06751_));
 AND2x2_ASAP7_75t_R _18583_ (.A(_06731_),
    .B(_06751_),
    .Y(_04191_));
 OR4x1_ASAP7_75t_R _18584_ (.A(_00866_),
    .B(_00867_),
    .C(_06738_),
    .D(_06746_),
    .Y(_06752_));
 XOR2x2_ASAP7_75t_R _18585_ (.A(_00864_),
    .B(_06752_),
    .Y(_06753_));
 AND2x2_ASAP7_75t_R _18586_ (.A(_06731_),
    .B(_06753_),
    .Y(_04192_));
 OR5x1_ASAP7_75t_R _18587_ (.A(_00864_),
    .B(_00866_),
    .C(_00867_),
    .D(_06736_),
    .E(_06746_),
    .Y(_06754_));
 XOR2x2_ASAP7_75t_R _18588_ (.A(_00863_),
    .B(_06754_),
    .Y(_06755_));
 AND2x2_ASAP7_75t_R _18589_ (.A(_06731_),
    .B(_06755_),
    .Y(_04193_));
 OR3x1_ASAP7_75t_R _18590_ (.A(_00865_),
    .B(_00876_),
    .C(_00047_),
    .Y(_06756_));
 XOR2x2_ASAP7_75t_R _18591_ (.A(_00862_),
    .B(_06756_),
    .Y(_06757_));
 AND2x2_ASAP7_75t_R _18592_ (.A(_06731_),
    .B(_06757_),
    .Y(_04194_));
 OR3x1_ASAP7_75t_R _18593_ (.A(_00862_),
    .B(_00865_),
    .C(_02669_),
    .Y(_06758_));
 NAND2x1_ASAP7_75t_R _18594_ (.A(_00861_),
    .B(_06758_),
    .Y(_06759_));
 AND3x1_ASAP7_75t_R _18595_ (.A(_06734_),
    .B(_06699_),
    .C(_06759_),
    .Y(_04195_));
 XOR2x2_ASAP7_75t_R _18596_ (.A(_00860_),
    .B(_06704_),
    .Y(_06760_));
 AND2x2_ASAP7_75t_R _18597_ (.A(_06731_),
    .B(_06760_),
    .Y(_04196_));
 OR3x1_ASAP7_75t_R _18598_ (.A(_00859_),
    .B(_00860_),
    .C(_06699_),
    .Y(_06761_));
 OAI21x1_ASAP7_75t_R _18599_ (.A1(_00860_),
    .A2(_06699_),
    .B(_00859_),
    .Y(_06762_));
 AND3x1_ASAP7_75t_R _18600_ (.A(_06734_),
    .B(_06761_),
    .C(_06762_),
    .Y(_04197_));
 BUFx6f_ASAP7_75t_R _18601_ (.A(_06547_),
    .Y(_06763_));
 OR3x1_ASAP7_75t_R _18602_ (.A(_00859_),
    .B(_00860_),
    .C(_06704_),
    .Y(_06764_));
 XOR2x2_ASAP7_75t_R _18603_ (.A(_00858_),
    .B(_06764_),
    .Y(_06765_));
 AND2x2_ASAP7_75t_R _18604_ (.A(_06763_),
    .B(_06765_),
    .Y(_04198_));
 OR4x1_ASAP7_75t_R _18605_ (.A(_00858_),
    .B(_00859_),
    .C(_00860_),
    .D(_06699_),
    .Y(_06766_));
 NAND2x1_ASAP7_75t_R _18606_ (.A(_00857_),
    .B(_06766_),
    .Y(_06767_));
 AND3x1_ASAP7_75t_R _18607_ (.A(_06734_),
    .B(_06701_),
    .C(_06767_),
    .Y(_04199_));
 XOR2x2_ASAP7_75t_R _18608_ (.A(_06688_),
    .B(_06705_),
    .Y(_06768_));
 AND2x2_ASAP7_75t_R _18609_ (.A(_06763_),
    .B(_06768_),
    .Y(_04200_));
 BUFx6f_ASAP7_75t_R _18610_ (.A(_00840_),
    .Y(_06769_));
 BUFx6f_ASAP7_75t_R _18611_ (.A(_00817_),
    .Y(_06770_));
 AND4x1_ASAP7_75t_R _18612_ (.A(_06770_),
    .B(_00845_),
    .C(_00846_),
    .D(_00847_),
    .Y(_06771_));
 AND5x1_ASAP7_75t_R _18613_ (.A(_00836_),
    .B(_00841_),
    .C(_00842_),
    .D(_00844_),
    .E(_06771_),
    .Y(_06772_));
 AND5x2_ASAP7_75t_R _18614_ (.A(_00838_),
    .B(_00839_),
    .C(_06769_),
    .D(_05995_),
    .E(_06772_),
    .Y(_06773_));
 BUFx6f_ASAP7_75t_R _18615_ (.A(_00832_),
    .Y(_06774_));
 AND4x1_ASAP7_75t_R _18616_ (.A(_00831_),
    .B(_06774_),
    .C(_00833_),
    .D(_00834_),
    .Y(_06775_));
 AND4x1_ASAP7_75t_R _18617_ (.A(_00825_),
    .B(_00827_),
    .C(_00828_),
    .D(_00835_),
    .Y(_06776_));
 AND5x1_ASAP7_75t_R _18618_ (.A(_00818_),
    .B(_00819_),
    .C(_00824_),
    .D(_00843_),
    .E(_06776_),
    .Y(_06777_));
 AND3x1_ASAP7_75t_R _18619_ (.A(_00822_),
    .B(_00823_),
    .C(_00826_),
    .Y(_06778_));
 OR3x1_ASAP7_75t_R _18620_ (.A(_00820_),
    .B(_00821_),
    .C(_06778_),
    .Y(_06779_));
 AND5x2_ASAP7_75t_R _18621_ (.A(_00829_),
    .B(_00830_),
    .C(_06775_),
    .D(_06777_),
    .E(_06779_),
    .Y(_06780_));
 NAND2x2_ASAP7_75t_R _18622_ (.A(_06773_),
    .B(_06780_),
    .Y(_06781_));
 NOR2x1_ASAP7_75t_R _18623_ (.A(_00807_),
    .B(_06781_),
    .Y(_04201_));
 INVx1_ASAP7_75t_R _18624_ (.A(_06781_),
    .Y(_04202_));
 NOR2x1_ASAP7_75t_R _18625_ (.A(_00810_),
    .B(_06781_),
    .Y(_04203_));
 NOR2x1_ASAP7_75t_R _18626_ (.A(_00809_),
    .B(_06781_),
    .Y(_04204_));
 NOR2x1_ASAP7_75t_R _18627_ (.A(_00808_),
    .B(_06781_),
    .Y(_04205_));
 NOR2x1_ASAP7_75t_R _18628_ (.A(_00806_),
    .B(_06781_),
    .Y(_04206_));
 NOR2x1_ASAP7_75t_R _18629_ (.A(_00805_),
    .B(_06781_),
    .Y(_04207_));
 INVx1_ASAP7_75t_R _18630_ (.A(_06781_),
    .Y(_04208_));
 AND2x2_ASAP7_75t_R _18631_ (.A(_06763_),
    .B(_00048_),
    .Y(_04209_));
 OR4x1_ASAP7_75t_R _18632_ (.A(_00822_),
    .B(_00823_),
    .C(_00826_),
    .D(_02673_),
    .Y(_06782_));
 OR4x1_ASAP7_75t_R _18633_ (.A(_00818_),
    .B(_00819_),
    .C(_00820_),
    .D(_00821_),
    .Y(_06783_));
 OR2x6_ASAP7_75t_R _18634_ (.A(_06782_),
    .B(_06783_),
    .Y(_06784_));
 OR3x1_ASAP7_75t_R _18635_ (.A(_06770_),
    .B(_00847_),
    .C(_06784_),
    .Y(_06785_));
 OAI21x1_ASAP7_75t_R _18636_ (.A1(_06770_),
    .A2(_06784_),
    .B(_00847_),
    .Y(_06786_));
 AND3x1_ASAP7_75t_R _18637_ (.A(_06734_),
    .B(_06785_),
    .C(_06786_),
    .Y(_04210_));
 OR5x2_ASAP7_75t_R _18638_ (.A(_00822_),
    .B(_00823_),
    .C(_00826_),
    .D(_00837_),
    .E(_00048_),
    .Y(_06787_));
 OR2x6_ASAP7_75t_R _18639_ (.A(_06783_),
    .B(_06787_),
    .Y(_06788_));
 OR3x1_ASAP7_75t_R _18640_ (.A(_06770_),
    .B(_00847_),
    .C(_06788_),
    .Y(_06789_));
 XOR2x2_ASAP7_75t_R _18641_ (.A(_00846_),
    .B(_06789_),
    .Y(_06790_));
 AND2x2_ASAP7_75t_R _18642_ (.A(_06763_),
    .B(_06790_),
    .Y(_04211_));
 OR4x1_ASAP7_75t_R _18643_ (.A(_06770_),
    .B(_00846_),
    .C(_00847_),
    .D(_06784_),
    .Y(_06791_));
 XOR2x2_ASAP7_75t_R _18644_ (.A(_00845_),
    .B(_06791_),
    .Y(_06792_));
 AND2x2_ASAP7_75t_R _18645_ (.A(_06763_),
    .B(_06792_),
    .Y(_04212_));
 OR5x2_ASAP7_75t_R _18646_ (.A(_06770_),
    .B(_00844_),
    .C(_00845_),
    .D(_00846_),
    .E(_00847_),
    .Y(_06793_));
 OR5x1_ASAP7_75t_R _18647_ (.A(_06770_),
    .B(_00845_),
    .C(_00846_),
    .D(_00847_),
    .E(_06788_),
    .Y(_06794_));
 NAND2x1_ASAP7_75t_R _18648_ (.A(_00844_),
    .B(_06794_),
    .Y(_06795_));
 OA211x2_ASAP7_75t_R _18649_ (.A1(_06788_),
    .A2(_06793_),
    .B(_06795_),
    .C(_06433_),
    .Y(_04213_));
 OR3x1_ASAP7_75t_R _18650_ (.A(_06782_),
    .B(_06783_),
    .C(_06793_),
    .Y(_06796_));
 XOR2x2_ASAP7_75t_R _18651_ (.A(_00843_),
    .B(_06796_),
    .Y(_06797_));
 AND2x2_ASAP7_75t_R _18652_ (.A(_06763_),
    .B(_06797_),
    .Y(_04214_));
 OR3x1_ASAP7_75t_R _18653_ (.A(_00843_),
    .B(_06788_),
    .C(_06793_),
    .Y(_06798_));
 XOR2x2_ASAP7_75t_R _18654_ (.A(_00842_),
    .B(_06798_),
    .Y(_06799_));
 AND2x2_ASAP7_75t_R _18655_ (.A(_06763_),
    .B(_06799_),
    .Y(_04215_));
 OR4x1_ASAP7_75t_R _18656_ (.A(_00841_),
    .B(_00842_),
    .C(_00843_),
    .D(_06796_),
    .Y(_06800_));
 OR3x1_ASAP7_75t_R _18657_ (.A(_00842_),
    .B(_00843_),
    .C(_06796_),
    .Y(_06801_));
 NAND2x1_ASAP7_75t_R _18658_ (.A(_00841_),
    .B(_06801_),
    .Y(_06802_));
 AND3x1_ASAP7_75t_R _18659_ (.A(_06734_),
    .B(_06800_),
    .C(_06802_),
    .Y(_04216_));
 OR5x2_ASAP7_75t_R _18660_ (.A(_00841_),
    .B(_00842_),
    .C(_00843_),
    .D(_06788_),
    .E(_06793_),
    .Y(_06803_));
 XOR2x2_ASAP7_75t_R _18661_ (.A(_06769_),
    .B(_06803_),
    .Y(_06804_));
 AND2x2_ASAP7_75t_R _18662_ (.A(_06763_),
    .B(_06804_),
    .Y(_04217_));
 OR3x1_ASAP7_75t_R _18663_ (.A(_00839_),
    .B(_06769_),
    .C(_06800_),
    .Y(_06805_));
 OAI21x1_ASAP7_75t_R _18664_ (.A1(_06769_),
    .A2(_06800_),
    .B(_00839_),
    .Y(_06806_));
 AND3x1_ASAP7_75t_R _18665_ (.A(_06734_),
    .B(_06805_),
    .C(_06806_),
    .Y(_04218_));
 OR3x1_ASAP7_75t_R _18666_ (.A(_00839_),
    .B(_06769_),
    .C(_06803_),
    .Y(_06807_));
 XOR2x2_ASAP7_75t_R _18667_ (.A(_00838_),
    .B(_06807_),
    .Y(_06808_));
 AND2x2_ASAP7_75t_R _18668_ (.A(_06763_),
    .B(_06808_),
    .Y(_04219_));
 NOR2x1_ASAP7_75t_R _18669_ (.A(_06272_),
    .B(_02674_),
    .Y(_04220_));
 OR4x1_ASAP7_75t_R _18670_ (.A(_00838_),
    .B(_00839_),
    .C(_06769_),
    .D(_06800_),
    .Y(_06809_));
 XOR2x2_ASAP7_75t_R _18671_ (.A(_00836_),
    .B(_06809_),
    .Y(_06810_));
 AND2x2_ASAP7_75t_R _18672_ (.A(_06763_),
    .B(_06810_),
    .Y(_04221_));
 BUFx6f_ASAP7_75t_R _18673_ (.A(_06547_),
    .Y(_06811_));
 OR5x1_ASAP7_75t_R _18674_ (.A(_00836_),
    .B(_00838_),
    .C(_00839_),
    .D(_06769_),
    .E(_06803_),
    .Y(_06812_));
 XOR2x2_ASAP7_75t_R _18675_ (.A(_00835_),
    .B(_06812_),
    .Y(_06813_));
 AND2x2_ASAP7_75t_R _18676_ (.A(_06811_),
    .B(_06813_),
    .Y(_04222_));
 OR5x2_ASAP7_75t_R _18677_ (.A(_00835_),
    .B(_00836_),
    .C(_00838_),
    .D(_00839_),
    .E(_06769_),
    .Y(_06814_));
 OR3x1_ASAP7_75t_R _18678_ (.A(_00834_),
    .B(_06800_),
    .C(_06814_),
    .Y(_06815_));
 OAI21x1_ASAP7_75t_R _18679_ (.A1(_06800_),
    .A2(_06814_),
    .B(_00834_),
    .Y(_06816_));
 AND3x1_ASAP7_75t_R _18680_ (.A(_06734_),
    .B(_06815_),
    .C(_06816_),
    .Y(_04223_));
 BUFx6f_ASAP7_75t_R _18681_ (.A(_06386_),
    .Y(_06817_));
 OR4x1_ASAP7_75t_R _18682_ (.A(_00833_),
    .B(_00834_),
    .C(_06803_),
    .D(_06814_),
    .Y(_06818_));
 OR3x1_ASAP7_75t_R _18683_ (.A(_00834_),
    .B(_06803_),
    .C(_06814_),
    .Y(_06819_));
 NAND2x1_ASAP7_75t_R _18684_ (.A(_00833_),
    .B(_06819_),
    .Y(_06820_));
 AND3x1_ASAP7_75t_R _18685_ (.A(_06817_),
    .B(_06818_),
    .C(_06820_),
    .Y(_04224_));
 OR4x1_ASAP7_75t_R _18686_ (.A(_00833_),
    .B(_00834_),
    .C(_06800_),
    .D(_06814_),
    .Y(_06821_));
 XOR2x2_ASAP7_75t_R _18687_ (.A(_06774_),
    .B(_06821_),
    .Y(_06822_));
 AND2x2_ASAP7_75t_R _18688_ (.A(_06811_),
    .B(_06822_),
    .Y(_04225_));
 OR3x1_ASAP7_75t_R _18689_ (.A(_00831_),
    .B(_06774_),
    .C(_06818_),
    .Y(_06823_));
 OAI21x1_ASAP7_75t_R _18690_ (.A1(_06774_),
    .A2(_06818_),
    .B(_00831_),
    .Y(_06824_));
 AND3x1_ASAP7_75t_R _18691_ (.A(_06817_),
    .B(_06823_),
    .C(_06824_),
    .Y(_04226_));
 OR3x1_ASAP7_75t_R _18692_ (.A(_00831_),
    .B(_06774_),
    .C(_06821_),
    .Y(_06825_));
 XOR2x2_ASAP7_75t_R _18693_ (.A(_00830_),
    .B(_06825_),
    .Y(_06826_));
 AND2x2_ASAP7_75t_R _18694_ (.A(_06811_),
    .B(_06826_),
    .Y(_04227_));
 OR4x1_ASAP7_75t_R _18695_ (.A(_00830_),
    .B(_00831_),
    .C(_06774_),
    .D(_06818_),
    .Y(_06827_));
 XOR2x2_ASAP7_75t_R _18696_ (.A(_00829_),
    .B(_06827_),
    .Y(_06828_));
 AND2x2_ASAP7_75t_R _18697_ (.A(_06811_),
    .B(_06828_),
    .Y(_04228_));
 OR5x1_ASAP7_75t_R _18698_ (.A(_00829_),
    .B(_00830_),
    .C(_00831_),
    .D(_06774_),
    .E(_06821_),
    .Y(_06829_));
 XOR2x2_ASAP7_75t_R _18699_ (.A(_00828_),
    .B(_06829_),
    .Y(_06830_));
 AND2x2_ASAP7_75t_R _18700_ (.A(_06811_),
    .B(_06830_),
    .Y(_04229_));
 OR5x2_ASAP7_75t_R _18701_ (.A(_00828_),
    .B(_00829_),
    .C(_00830_),
    .D(_00831_),
    .E(_06774_),
    .Y(_06831_));
 OR3x1_ASAP7_75t_R _18702_ (.A(_00827_),
    .B(_06818_),
    .C(_06831_),
    .Y(_06832_));
 OAI21x1_ASAP7_75t_R _18703_ (.A1(_06818_),
    .A2(_06831_),
    .B(_00827_),
    .Y(_06833_));
 AND3x1_ASAP7_75t_R _18704_ (.A(_06817_),
    .B(_06832_),
    .C(_06833_),
    .Y(_04230_));
 XOR2x2_ASAP7_75t_R _18705_ (.A(_00826_),
    .B(_02673_),
    .Y(_06834_));
 AND2x2_ASAP7_75t_R _18706_ (.A(_06811_),
    .B(_06834_),
    .Y(_04231_));
 OR3x1_ASAP7_75t_R _18707_ (.A(_00827_),
    .B(_06821_),
    .C(_06831_),
    .Y(_06835_));
 XOR2x2_ASAP7_75t_R _18708_ (.A(_00825_),
    .B(_06835_),
    .Y(_06836_));
 AND2x2_ASAP7_75t_R _18709_ (.A(_06811_),
    .B(_06836_),
    .Y(_04232_));
 OR4x1_ASAP7_75t_R _18710_ (.A(_00825_),
    .B(_00827_),
    .C(_06818_),
    .D(_06831_),
    .Y(_06837_));
 XOR2x2_ASAP7_75t_R _18711_ (.A(_00824_),
    .B(_06837_),
    .Y(_06838_));
 AND2x2_ASAP7_75t_R _18712_ (.A(_06811_),
    .B(_06838_),
    .Y(_04233_));
 OR3x1_ASAP7_75t_R _18713_ (.A(_00826_),
    .B(_00837_),
    .C(_00048_),
    .Y(_06839_));
 XOR2x2_ASAP7_75t_R _18714_ (.A(_00823_),
    .B(_06839_),
    .Y(_06840_));
 AND2x2_ASAP7_75t_R _18715_ (.A(_06811_),
    .B(_06840_),
    .Y(_04234_));
 OR3x1_ASAP7_75t_R _18716_ (.A(_00823_),
    .B(_00826_),
    .C(_02673_),
    .Y(_06841_));
 NAND2x1_ASAP7_75t_R _18717_ (.A(_00822_),
    .B(_06841_),
    .Y(_06842_));
 AND3x1_ASAP7_75t_R _18718_ (.A(_06817_),
    .B(_06782_),
    .C(_06842_),
    .Y(_04235_));
 XOR2x2_ASAP7_75t_R _18719_ (.A(_00821_),
    .B(_06787_),
    .Y(_06843_));
 AND2x2_ASAP7_75t_R _18720_ (.A(_06811_),
    .B(_06843_),
    .Y(_04236_));
 OR3x1_ASAP7_75t_R _18721_ (.A(_00820_),
    .B(_00821_),
    .C(_06782_),
    .Y(_06844_));
 OAI21x1_ASAP7_75t_R _18722_ (.A1(_00821_),
    .A2(_06782_),
    .B(_00820_),
    .Y(_06845_));
 AND3x1_ASAP7_75t_R _18723_ (.A(_06817_),
    .B(_06844_),
    .C(_06845_),
    .Y(_04237_));
 BUFx6f_ASAP7_75t_R _18724_ (.A(_06547_),
    .Y(_06846_));
 OR3x1_ASAP7_75t_R _18725_ (.A(_00820_),
    .B(_00821_),
    .C(_06787_),
    .Y(_06847_));
 XOR2x2_ASAP7_75t_R _18726_ (.A(_00819_),
    .B(_06847_),
    .Y(_06848_));
 AND2x2_ASAP7_75t_R _18727_ (.A(_06846_),
    .B(_06848_),
    .Y(_04238_));
 OR4x1_ASAP7_75t_R _18728_ (.A(_00819_),
    .B(_00820_),
    .C(_00821_),
    .D(_06782_),
    .Y(_06849_));
 NAND2x1_ASAP7_75t_R _18729_ (.A(_00818_),
    .B(_06849_),
    .Y(_06850_));
 AND3x1_ASAP7_75t_R _18730_ (.A(_06817_),
    .B(_06784_),
    .C(_06850_),
    .Y(_04239_));
 XOR2x2_ASAP7_75t_R _18731_ (.A(_06770_),
    .B(_06788_),
    .Y(_06851_));
 AND2x2_ASAP7_75t_R _18732_ (.A(_06846_),
    .B(_06851_),
    .Y(_04240_));
 AND2x2_ASAP7_75t_R _18733_ (.A(_06846_),
    .B(_00023_),
    .Y(_04241_));
 NAND2x1_ASAP7_75t_R _18734_ (.A(_00849_),
    .B(_00850_),
    .Y(_06852_));
 OR5x1_ASAP7_75t_R _18735_ (.A(_00848_),
    .B(_00851_),
    .C(\xs[2].cli1.i[33] ),
    .D(\xs[2].cli1.i[32] ),
    .E(_06852_),
    .Y(_06853_));
 BUFx3_ASAP7_75t_R _18736_ (.A(_06853_),
    .Y(_06854_));
 AND2x2_ASAP7_75t_R _18737_ (.A(_00849_),
    .B(_00850_),
    .Y(_06855_));
 AO31x2_ASAP7_75t_R _18738_ (.A1(\xs[2].cli1.i[34] ),
    .A2(_00852_),
    .A3(_06855_),
    .B(_00848_),
    .Y(_06856_));
 INVx2_ASAP7_75t_R _18739_ (.A(_02295_),
    .Y(_06857_));
 AOI21x1_ASAP7_75t_R _18740_ (.A1(_06854_),
    .A2(_06856_),
    .B(_06857_),
    .Y(_06858_));
 BUFx3_ASAP7_75t_R _18741_ (.A(_02289_),
    .Y(_06859_));
 INVx3_ASAP7_75t_R _18742_ (.A(_02288_),
    .Y(_06860_));
 OAI21x1_ASAP7_75t_R _18743_ (.A1(_06859_),
    .A2(_06854_),
    .B(_06860_),
    .Y(_06861_));
 OA31x2_ASAP7_75t_R _18744_ (.A1(_00851_),
    .A2(\xs[2].cli1.i[33] ),
    .A3(_06852_),
    .B1(\xs[2].cli1.i[39] ),
    .Y(_06862_));
 AO21x1_ASAP7_75t_R _18745_ (.A1(_00023_),
    .A2(_06862_),
    .B(_06860_),
    .Y(_06863_));
 NAND2x1_ASAP7_75t_R _18746_ (.A(_00888_),
    .B(_00889_),
    .Y(_06864_));
 OA31x2_ASAP7_75t_R _18747_ (.A1(_00890_),
    .A2(\peo[4][33] ),
    .A3(_06864_),
    .B1(\peo[4][39] ),
    .Y(_06865_));
 OA211x2_ASAP7_75t_R _18748_ (.A1(_06858_),
    .A2(_06861_),
    .B(_06863_),
    .C(_06865_),
    .Y(_06866_));
 OAI21x1_ASAP7_75t_R _18749_ (.A1(_06854_),
    .A2(_06866_),
    .B(_00894_),
    .Y(_06867_));
 INVx1_ASAP7_75t_R _18750_ (.A(_06859_),
    .Y(_06868_));
 AND3x1_ASAP7_75t_R _18751_ (.A(_06860_),
    .B(_06868_),
    .C(_06862_),
    .Y(_06869_));
 OR4x1_ASAP7_75t_R _18752_ (.A(\peo[5][0] ),
    .B(_06854_),
    .C(_06866_),
    .D(_06869_),
    .Y(_06870_));
 AND2x2_ASAP7_75t_R _18753_ (.A(_00888_),
    .B(_00889_),
    .Y(_06871_));
 AO31x2_ASAP7_75t_R _18754_ (.A1(\peo[4][34] ),
    .A2(_00891_),
    .A3(_06871_),
    .B(_00887_),
    .Y(_06872_));
 AO21x1_ASAP7_75t_R _18755_ (.A1(\peo[4][39] ),
    .A2(\peo[4][32] ),
    .B(_02295_),
    .Y(_06873_));
 AND2x2_ASAP7_75t_R _18756_ (.A(_06872_),
    .B(_06873_),
    .Y(_06874_));
 OAI21x1_ASAP7_75t_R _18757_ (.A1(_02295_),
    .A2(_06862_),
    .B(_06854_),
    .Y(_06875_));
 NAND2x1_ASAP7_75t_R _18758_ (.A(_06860_),
    .B(_06859_),
    .Y(_06876_));
 AO21x2_ASAP7_75t_R _18759_ (.A1(_06874_),
    .A2(_06875_),
    .B(_06876_),
    .Y(_06877_));
 NOR2x1_ASAP7_75t_R _18760_ (.A(_06857_),
    .B(_06877_),
    .Y(_06878_));
 NOR2x1_ASAP7_75t_R _18761_ (.A(_09314_),
    .B(_06878_),
    .Y(_06879_));
 NOR2x1_ASAP7_75t_R _18762_ (.A(_06206_),
    .B(_02299_),
    .Y(_06880_));
 AO32x1_ASAP7_75t_R _18763_ (.A1(_06867_),
    .A2(_06870_),
    .A3(_06879_),
    .B1(_06880_),
    .B2(_06878_),
    .Y(_04242_));
 OR3x2_ASAP7_75t_R _18764_ (.A(_10763_),
    .B(_06857_),
    .C(_06877_),
    .Y(_06881_));
 NOR2x1_ASAP7_75t_R _18765_ (.A(_02298_),
    .B(_06881_),
    .Y(_04243_));
 NOR2x1_ASAP7_75t_R _18766_ (.A(_02297_),
    .B(_06881_),
    .Y(_04244_));
 NOR2x1_ASAP7_75t_R _18767_ (.A(_02296_),
    .B(_06881_),
    .Y(_04245_));
 NOR2x1_ASAP7_75t_R _18768_ (.A(_02287_),
    .B(_06881_),
    .Y(_04246_));
 NOR2x1_ASAP7_75t_R _18769_ (.A(_02286_),
    .B(_06881_),
    .Y(_04247_));
 NOR2x1_ASAP7_75t_R _18770_ (.A(_06866_),
    .B(_06869_),
    .Y(_06882_));
 OR3x1_ASAP7_75t_R _18771_ (.A(_09207_),
    .B(_00855_),
    .C(_06882_),
    .Y(_06883_));
 NAND2x1_ASAP7_75t_R _18772_ (.A(_06874_),
    .B(_06875_),
    .Y(_06884_));
 AND5x1_ASAP7_75t_R _18773_ (.A(_06860_),
    .B(_06859_),
    .C(_06857_),
    .D(_02299_),
    .E(_06884_),
    .Y(_06885_));
 OA21x2_ASAP7_75t_R _18774_ (.A1(_02295_),
    .A2(_06877_),
    .B(_00894_),
    .Y(_06886_));
 OR5x1_ASAP7_75t_R _18775_ (.A(_10826_),
    .B(_06866_),
    .C(_06869_),
    .D(_06885_),
    .E(_06886_),
    .Y(_06887_));
 NAND2x1_ASAP7_75t_R _18776_ (.A(_06883_),
    .B(_06887_),
    .Y(_04248_));
 OR3x2_ASAP7_75t_R _18777_ (.A(_10763_),
    .B(_02295_),
    .C(_06877_),
    .Y(_06888_));
 NOR2x1_ASAP7_75t_R _18778_ (.A(_02298_),
    .B(_06888_),
    .Y(_04249_));
 NOR2x1_ASAP7_75t_R _18779_ (.A(_02297_),
    .B(_06888_),
    .Y(_04250_));
 NOR2x1_ASAP7_75t_R _18780_ (.A(_02296_),
    .B(_06888_),
    .Y(_04251_));
 NOR2x1_ASAP7_75t_R _18781_ (.A(_02287_),
    .B(_06888_),
    .Y(_04252_));
 NOR2x1_ASAP7_75t_R _18782_ (.A(_02286_),
    .B(_06888_),
    .Y(_04253_));
 AO21x1_ASAP7_75t_R _18783_ (.A1(_06859_),
    .A2(_06884_),
    .B(_02288_),
    .Y(_06889_));
 BUFx6f_ASAP7_75t_R _18784_ (.A(_06889_),
    .Y(_06890_));
 NOR2x1_ASAP7_75t_R _18785_ (.A(_02299_),
    .B(_06890_),
    .Y(_06891_));
 AND2x2_ASAP7_75t_R _18786_ (.A(_06860_),
    .B(_06865_),
    .Y(_06892_));
 AND2x2_ASAP7_75t_R _18787_ (.A(_02288_),
    .B(_00023_),
    .Y(_06893_));
 AO221x1_ASAP7_75t_R _18788_ (.A1(_06860_),
    .A2(_06868_),
    .B1(_06865_),
    .B2(_06893_),
    .C(_06856_),
    .Y(_06894_));
 AOI21x1_ASAP7_75t_R _18789_ (.A1(_06858_),
    .A2(_06892_),
    .B(_06894_),
    .Y(_06895_));
 NAND2x1_ASAP7_75t_R _18790_ (.A(_00855_),
    .B(_06895_),
    .Y(_06896_));
 OA211x2_ASAP7_75t_R _18791_ (.A1(\peo[4][0] ),
    .A2(_06895_),
    .B(_06896_),
    .C(_06890_),
    .Y(_06897_));
 OA21x2_ASAP7_75t_R _18792_ (.A1(_06891_),
    .A2(_06897_),
    .B(_06676_),
    .Y(_04254_));
 AOI21x1_ASAP7_75t_R _18793_ (.A1(_06859_),
    .A2(_06884_),
    .B(_02288_),
    .Y(_06898_));
 NAND2x2_ASAP7_75t_R _18794_ (.A(_08581_),
    .B(_06898_),
    .Y(_06899_));
 NOR2x1_ASAP7_75t_R _18795_ (.A(_02298_),
    .B(_06899_),
    .Y(_04255_));
 NOR2x1_ASAP7_75t_R _18796_ (.A(_02297_),
    .B(_06899_),
    .Y(_04256_));
 NOR2x1_ASAP7_75t_R _18797_ (.A(_02296_),
    .B(_06899_),
    .Y(_04257_));
 AND2x2_ASAP7_75t_R _18798_ (.A(_06857_),
    .B(_06898_),
    .Y(_06900_));
 NAND2x1_ASAP7_75t_R _18799_ (.A(_00853_),
    .B(_06895_),
    .Y(_06901_));
 OA211x2_ASAP7_75t_R _18800_ (.A1(\peo[4][32] ),
    .A2(_06895_),
    .B(_06901_),
    .C(_06890_),
    .Y(_06902_));
 OA21x2_ASAP7_75t_R _18801_ (.A1(_06900_),
    .A2(_06902_),
    .B(_06676_),
    .Y(_04258_));
 NOR2x1_ASAP7_75t_R _18802_ (.A(_02294_),
    .B(_06890_),
    .Y(_06903_));
 NAND2x1_ASAP7_75t_R _18803_ (.A(_00852_),
    .B(_06895_),
    .Y(_06904_));
 OA211x2_ASAP7_75t_R _18804_ (.A1(\peo[4][33] ),
    .A2(_06895_),
    .B(_06904_),
    .C(_06890_),
    .Y(_06905_));
 OA21x2_ASAP7_75t_R _18805_ (.A1(_06903_),
    .A2(_06905_),
    .B(_06676_),
    .Y(_04259_));
 INVx1_ASAP7_75t_R _18806_ (.A(_06866_),
    .Y(_06906_));
 OR2x2_ASAP7_75t_R _18807_ (.A(_06856_),
    .B(_06866_),
    .Y(_06907_));
 AO32x1_ASAP7_75t_R _18808_ (.A1(\xs[2].cli1.i[39] ),
    .A2(_00851_),
    .A3(_06906_),
    .B1(_06907_),
    .B2(_00890_),
    .Y(_06908_));
 NAND2x1_ASAP7_75t_R _18809_ (.A(_08599_),
    .B(_06890_),
    .Y(_06909_));
 OAI22x1_ASAP7_75t_R _18810_ (.A1(_02293_),
    .A2(_06899_),
    .B1(_06908_),
    .B2(_06909_),
    .Y(_04260_));
 NOR2x1_ASAP7_75t_R _18811_ (.A(_02292_),
    .B(_06890_),
    .Y(_06910_));
 NAND2x1_ASAP7_75t_R _18812_ (.A(_00850_),
    .B(_06895_),
    .Y(_06911_));
 OA211x2_ASAP7_75t_R _18813_ (.A1(\peo[4][35] ),
    .A2(_06895_),
    .B(_06911_),
    .C(_06890_),
    .Y(_06912_));
 OA21x2_ASAP7_75t_R _18814_ (.A1(_06910_),
    .A2(_06912_),
    .B(_06676_),
    .Y(_04261_));
 NOR2x1_ASAP7_75t_R _18815_ (.A(_02291_),
    .B(_06890_),
    .Y(_06913_));
 NAND2x1_ASAP7_75t_R _18816_ (.A(_00849_),
    .B(_06895_),
    .Y(_06914_));
 OA211x2_ASAP7_75t_R _18817_ (.A1(\peo[4][36] ),
    .A2(_06895_),
    .B(_06914_),
    .C(_06889_),
    .Y(_06915_));
 OA21x2_ASAP7_75t_R _18818_ (.A1(_06913_),
    .A2(_06915_),
    .B(_06676_),
    .Y(_04262_));
 NOR2x1_ASAP7_75t_R _18819_ (.A(_02290_),
    .B(_06899_),
    .Y(_04263_));
 OR3x1_ASAP7_75t_R _18820_ (.A(_08642_),
    .B(_06884_),
    .C(_06876_),
    .Y(_06916_));
 INVx1_ASAP7_75t_R _18821_ (.A(_06916_),
    .Y(_04264_));
 AND3x1_ASAP7_75t_R _18822_ (.A(_06872_),
    .B(_06856_),
    .C(_06890_),
    .Y(_06917_));
 NOR2x1_ASAP7_75t_R _18823_ (.A(_06272_),
    .B(_06917_),
    .Y(_04265_));
 NOR2x1_ASAP7_75t_R _18824_ (.A(_02287_),
    .B(_06899_),
    .Y(_04266_));
 NOR2x1_ASAP7_75t_R _18825_ (.A(_02286_),
    .B(_06899_),
    .Y(_04267_));
 BUFx6f_ASAP7_75t_R _18826_ (.A(_00773_),
    .Y(_06918_));
 BUFx6f_ASAP7_75t_R _18827_ (.A(_00781_),
    .Y(_06919_));
 AND4x1_ASAP7_75t_R _18828_ (.A(_00752_),
    .B(_00780_),
    .C(_06919_),
    .D(_00782_),
    .Y(_06920_));
 AND5x1_ASAP7_75t_R _18829_ (.A(_00771_),
    .B(_00776_),
    .C(_00777_),
    .D(_00779_),
    .E(_06920_),
    .Y(_06921_));
 AND5x2_ASAP7_75t_R _18830_ (.A(_06918_),
    .B(_00774_),
    .C(_00775_),
    .D(_05995_),
    .E(_06921_),
    .Y(_06922_));
 BUFx3_ASAP7_75t_R _18831_ (.A(_00768_),
    .Y(_06923_));
 AND4x1_ASAP7_75t_R _18832_ (.A(_00766_),
    .B(_00767_),
    .C(_06923_),
    .D(_00769_),
    .Y(_06924_));
 AND4x1_ASAP7_75t_R _18833_ (.A(_00760_),
    .B(_00762_),
    .C(_00763_),
    .D(_00770_),
    .Y(_06925_));
 AND5x1_ASAP7_75t_R _18834_ (.A(_00753_),
    .B(_00754_),
    .C(_00759_),
    .D(_00778_),
    .E(_06925_),
    .Y(_06926_));
 BUFx6f_ASAP7_75t_R _18835_ (.A(_00756_),
    .Y(_06927_));
 AND3x1_ASAP7_75t_R _18836_ (.A(_00757_),
    .B(_00758_),
    .C(_00761_),
    .Y(_06928_));
 OR3x1_ASAP7_75t_R _18837_ (.A(_00755_),
    .B(_06927_),
    .C(_06928_),
    .Y(_06929_));
 AND5x2_ASAP7_75t_R _18838_ (.A(_00764_),
    .B(_00765_),
    .C(_06924_),
    .D(_06926_),
    .E(_06929_),
    .Y(_06930_));
 NAND2x2_ASAP7_75t_R _18839_ (.A(_06922_),
    .B(_06930_),
    .Y(_06931_));
 NOR2x1_ASAP7_75t_R _18840_ (.A(_00709_),
    .B(_06931_),
    .Y(_04268_));
 INVx1_ASAP7_75t_R _18841_ (.A(_06931_),
    .Y(_04269_));
 NOR2x1_ASAP7_75t_R _18842_ (.A(_00712_),
    .B(_06931_),
    .Y(_04270_));
 NOR2x1_ASAP7_75t_R _18843_ (.A(_00711_),
    .B(_06931_),
    .Y(_04271_));
 NOR2x1_ASAP7_75t_R _18844_ (.A(_00710_),
    .B(_06931_),
    .Y(_04272_));
 NOR2x1_ASAP7_75t_R _18845_ (.A(_00708_),
    .B(_06931_),
    .Y(_04273_));
 NOR2x1_ASAP7_75t_R _18846_ (.A(_00707_),
    .B(_06931_),
    .Y(_04274_));
 INVx1_ASAP7_75t_R _18847_ (.A(_06931_),
    .Y(_04275_));
 AND2x2_ASAP7_75t_R _18848_ (.A(_06846_),
    .B(_00049_),
    .Y(_04276_));
 OR4x1_ASAP7_75t_R _18849_ (.A(_00757_),
    .B(_00758_),
    .C(_00761_),
    .D(_02657_),
    .Y(_06932_));
 OR5x2_ASAP7_75t_R _18850_ (.A(_00752_),
    .B(_00753_),
    .C(_00754_),
    .D(_00755_),
    .E(_06927_),
    .Y(_06933_));
 OR3x1_ASAP7_75t_R _18851_ (.A(_00782_),
    .B(_06932_),
    .C(_06933_),
    .Y(_06934_));
 BUFx6f_ASAP7_75t_R _18852_ (.A(_06934_),
    .Y(_06935_));
 OAI21x1_ASAP7_75t_R _18853_ (.A1(_06932_),
    .A2(_06933_),
    .B(_00782_),
    .Y(_06936_));
 AND3x1_ASAP7_75t_R _18854_ (.A(_06817_),
    .B(_06935_),
    .C(_06936_),
    .Y(_04277_));
 OR5x2_ASAP7_75t_R _18855_ (.A(_00757_),
    .B(_00758_),
    .C(_00761_),
    .D(_00772_),
    .E(_00049_),
    .Y(_06937_));
 OR3x2_ASAP7_75t_R _18856_ (.A(_00782_),
    .B(_06933_),
    .C(_06937_),
    .Y(_06938_));
 XOR2x2_ASAP7_75t_R _18857_ (.A(_06919_),
    .B(_06938_),
    .Y(_06939_));
 AND2x2_ASAP7_75t_R _18858_ (.A(_06846_),
    .B(_06939_),
    .Y(_04278_));
 OR3x1_ASAP7_75t_R _18859_ (.A(_00780_),
    .B(_06919_),
    .C(_06935_),
    .Y(_06940_));
 OAI21x1_ASAP7_75t_R _18860_ (.A1(_06919_),
    .A2(_06935_),
    .B(_00780_),
    .Y(_06941_));
 AND3x1_ASAP7_75t_R _18861_ (.A(_06817_),
    .B(_06940_),
    .C(_06941_),
    .Y(_04279_));
 OR3x1_ASAP7_75t_R _18862_ (.A(_00780_),
    .B(_06919_),
    .C(_06938_),
    .Y(_06942_));
 XOR2x2_ASAP7_75t_R _18863_ (.A(_00779_),
    .B(_06942_),
    .Y(_06943_));
 AND2x2_ASAP7_75t_R _18864_ (.A(_06846_),
    .B(_06943_),
    .Y(_04280_));
 OR4x1_ASAP7_75t_R _18865_ (.A(_00779_),
    .B(_00780_),
    .C(_06919_),
    .D(_06935_),
    .Y(_06944_));
 XOR2x2_ASAP7_75t_R _18866_ (.A(_00778_),
    .B(_06944_),
    .Y(_06945_));
 AND2x2_ASAP7_75t_R _18867_ (.A(_06846_),
    .B(_06945_),
    .Y(_04281_));
 OR5x1_ASAP7_75t_R _18868_ (.A(_00778_),
    .B(_00779_),
    .C(_00780_),
    .D(_06919_),
    .E(_06938_),
    .Y(_06946_));
 XOR2x2_ASAP7_75t_R _18869_ (.A(_00777_),
    .B(_06946_),
    .Y(_06947_));
 AND2x2_ASAP7_75t_R _18870_ (.A(_06846_),
    .B(_06947_),
    .Y(_04282_));
 OR5x2_ASAP7_75t_R _18871_ (.A(_00777_),
    .B(_00778_),
    .C(_00779_),
    .D(_00780_),
    .E(_06919_),
    .Y(_06948_));
 OR3x1_ASAP7_75t_R _18872_ (.A(_00776_),
    .B(_06935_),
    .C(_06948_),
    .Y(_06949_));
 OAI21x1_ASAP7_75t_R _18873_ (.A1(_06935_),
    .A2(_06948_),
    .B(_00776_),
    .Y(_06950_));
 AND3x1_ASAP7_75t_R _18874_ (.A(_06817_),
    .B(_06949_),
    .C(_06950_),
    .Y(_04283_));
 OR3x2_ASAP7_75t_R _18875_ (.A(_00775_),
    .B(_00776_),
    .C(_06948_),
    .Y(_06951_));
 OR3x1_ASAP7_75t_R _18876_ (.A(_00776_),
    .B(_06938_),
    .C(_06948_),
    .Y(_06952_));
 NAND2x1_ASAP7_75t_R _18877_ (.A(_00775_),
    .B(_06952_),
    .Y(_06953_));
 OA211x2_ASAP7_75t_R _18878_ (.A1(_06938_),
    .A2(_06951_),
    .B(_06953_),
    .C(_06433_),
    .Y(_04284_));
 OR3x2_ASAP7_75t_R _18879_ (.A(_00774_),
    .B(_06935_),
    .C(_06951_),
    .Y(_06954_));
 OAI21x1_ASAP7_75t_R _18880_ (.A1(_06935_),
    .A2(_06951_),
    .B(_00774_),
    .Y(_06955_));
 AND3x1_ASAP7_75t_R _18881_ (.A(_06817_),
    .B(_06954_),
    .C(_06955_),
    .Y(_04285_));
 OR3x2_ASAP7_75t_R _18882_ (.A(_00774_),
    .B(_06938_),
    .C(_06951_),
    .Y(_06956_));
 XOR2x2_ASAP7_75t_R _18883_ (.A(_06918_),
    .B(_06956_),
    .Y(_06957_));
 AND2x2_ASAP7_75t_R _18884_ (.A(_06846_),
    .B(_06957_),
    .Y(_04286_));
 NOR2x1_ASAP7_75t_R _18885_ (.A(_06272_),
    .B(_02658_),
    .Y(_04287_));
 BUFx6f_ASAP7_75t_R _18886_ (.A(_06386_),
    .Y(_06958_));
 OR3x1_ASAP7_75t_R _18887_ (.A(_00771_),
    .B(_06918_),
    .C(_06954_),
    .Y(_06959_));
 OAI21x1_ASAP7_75t_R _18888_ (.A1(_06918_),
    .A2(_06954_),
    .B(_00771_),
    .Y(_06960_));
 AND3x1_ASAP7_75t_R _18889_ (.A(_06958_),
    .B(_06959_),
    .C(_06960_),
    .Y(_04288_));
 OR3x1_ASAP7_75t_R _18890_ (.A(_00771_),
    .B(_06918_),
    .C(_06956_),
    .Y(_06961_));
 XOR2x2_ASAP7_75t_R _18891_ (.A(_00770_),
    .B(_06961_),
    .Y(_06962_));
 AND2x2_ASAP7_75t_R _18892_ (.A(_06846_),
    .B(_06962_),
    .Y(_04289_));
 OR5x1_ASAP7_75t_R _18893_ (.A(_00769_),
    .B(_00770_),
    .C(_00771_),
    .D(_06918_),
    .E(_06954_),
    .Y(_06963_));
 BUFx3_ASAP7_75t_R _18894_ (.A(_06963_),
    .Y(_06964_));
 OR4x1_ASAP7_75t_R _18895_ (.A(_00770_),
    .B(_00771_),
    .C(_06918_),
    .D(_06954_),
    .Y(_06965_));
 NAND2x1_ASAP7_75t_R _18896_ (.A(_00769_),
    .B(_06965_),
    .Y(_06966_));
 AND3x1_ASAP7_75t_R _18897_ (.A(_06958_),
    .B(_06964_),
    .C(_06966_),
    .Y(_04290_));
 BUFx6f_ASAP7_75t_R _18898_ (.A(_06547_),
    .Y(_06967_));
 OR5x2_ASAP7_75t_R _18899_ (.A(_00769_),
    .B(_00770_),
    .C(_00771_),
    .D(_06918_),
    .E(_06956_),
    .Y(_06968_));
 XOR2x2_ASAP7_75t_R _18900_ (.A(_06923_),
    .B(_06968_),
    .Y(_06969_));
 AND2x2_ASAP7_75t_R _18901_ (.A(_06967_),
    .B(_06969_),
    .Y(_04291_));
 OR3x1_ASAP7_75t_R _18902_ (.A(_00767_),
    .B(_06923_),
    .C(_06964_),
    .Y(_06970_));
 OAI21x1_ASAP7_75t_R _18903_ (.A1(_06923_),
    .A2(_06964_),
    .B(_00767_),
    .Y(_06971_));
 AND3x1_ASAP7_75t_R _18904_ (.A(_06958_),
    .B(_06970_),
    .C(_06971_),
    .Y(_04292_));
 OR3x1_ASAP7_75t_R _18905_ (.A(_00767_),
    .B(_06923_),
    .C(_06968_),
    .Y(_06972_));
 XOR2x2_ASAP7_75t_R _18906_ (.A(_00766_),
    .B(_06972_),
    .Y(_06973_));
 AND2x2_ASAP7_75t_R _18907_ (.A(_06967_),
    .B(_06973_),
    .Y(_04293_));
 OR4x1_ASAP7_75t_R _18908_ (.A(_00766_),
    .B(_00767_),
    .C(_06923_),
    .D(_06964_),
    .Y(_06974_));
 XOR2x2_ASAP7_75t_R _18909_ (.A(_00765_),
    .B(_06974_),
    .Y(_06975_));
 AND2x2_ASAP7_75t_R _18910_ (.A(_06967_),
    .B(_06975_),
    .Y(_04294_));
 OR5x1_ASAP7_75t_R _18911_ (.A(_00765_),
    .B(_00766_),
    .C(_00767_),
    .D(_06923_),
    .E(_06968_),
    .Y(_06976_));
 XOR2x2_ASAP7_75t_R _18912_ (.A(_00764_),
    .B(_06976_),
    .Y(_06977_));
 AND2x2_ASAP7_75t_R _18913_ (.A(_06967_),
    .B(_06977_),
    .Y(_04295_));
 OR5x2_ASAP7_75t_R _18914_ (.A(_00764_),
    .B(_00765_),
    .C(_00766_),
    .D(_00767_),
    .E(_06923_),
    .Y(_06978_));
 OR3x1_ASAP7_75t_R _18915_ (.A(_00763_),
    .B(_06964_),
    .C(_06978_),
    .Y(_06979_));
 OAI21x1_ASAP7_75t_R _18916_ (.A1(_06964_),
    .A2(_06978_),
    .B(_00763_),
    .Y(_06980_));
 AND3x1_ASAP7_75t_R _18917_ (.A(_06958_),
    .B(_06979_),
    .C(_06980_),
    .Y(_04296_));
 OR3x1_ASAP7_75t_R _18918_ (.A(_00763_),
    .B(_06968_),
    .C(_06978_),
    .Y(_06981_));
 XOR2x2_ASAP7_75t_R _18919_ (.A(_00762_),
    .B(_06981_),
    .Y(_06982_));
 AND2x2_ASAP7_75t_R _18920_ (.A(_06967_),
    .B(_06982_),
    .Y(_04297_));
 XOR2x2_ASAP7_75t_R _18921_ (.A(_00761_),
    .B(_02657_),
    .Y(_06983_));
 AND2x2_ASAP7_75t_R _18922_ (.A(_06967_),
    .B(_06983_),
    .Y(_04298_));
 OR4x1_ASAP7_75t_R _18923_ (.A(_00762_),
    .B(_00763_),
    .C(_06964_),
    .D(_06978_),
    .Y(_06984_));
 XOR2x2_ASAP7_75t_R _18924_ (.A(_00760_),
    .B(_06984_),
    .Y(_06985_));
 AND2x2_ASAP7_75t_R _18925_ (.A(_06967_),
    .B(_06985_),
    .Y(_04299_));
 OR5x1_ASAP7_75t_R _18926_ (.A(_00760_),
    .B(_00762_),
    .C(_00763_),
    .D(_06968_),
    .E(_06978_),
    .Y(_06986_));
 XOR2x2_ASAP7_75t_R _18927_ (.A(_00759_),
    .B(_06986_),
    .Y(_06987_));
 AND2x2_ASAP7_75t_R _18928_ (.A(_06967_),
    .B(_06987_),
    .Y(_04300_));
 OR3x1_ASAP7_75t_R _18929_ (.A(_00761_),
    .B(_00772_),
    .C(_00049_),
    .Y(_06988_));
 XOR2x2_ASAP7_75t_R _18930_ (.A(_00758_),
    .B(_06988_),
    .Y(_06989_));
 AND2x2_ASAP7_75t_R _18931_ (.A(_06967_),
    .B(_06989_),
    .Y(_04301_));
 OR3x1_ASAP7_75t_R _18932_ (.A(_00758_),
    .B(_00761_),
    .C(_02657_),
    .Y(_06990_));
 NAND2x1_ASAP7_75t_R _18933_ (.A(_00757_),
    .B(_06990_),
    .Y(_06991_));
 AND3x1_ASAP7_75t_R _18934_ (.A(_06958_),
    .B(_06932_),
    .C(_06991_),
    .Y(_04302_));
 XOR2x2_ASAP7_75t_R _18935_ (.A(_06927_),
    .B(_06937_),
    .Y(_06992_));
 AND2x2_ASAP7_75t_R _18936_ (.A(_06967_),
    .B(_06992_),
    .Y(_04303_));
 OR3x1_ASAP7_75t_R _18937_ (.A(_00755_),
    .B(_06927_),
    .C(_06932_),
    .Y(_06993_));
 OAI21x1_ASAP7_75t_R _18938_ (.A1(_06927_),
    .A2(_06932_),
    .B(_00755_),
    .Y(_06994_));
 AND3x1_ASAP7_75t_R _18939_ (.A(_06958_),
    .B(_06993_),
    .C(_06994_),
    .Y(_04304_));
 BUFx6f_ASAP7_75t_R _18940_ (.A(_06547_),
    .Y(_06995_));
 OR3x1_ASAP7_75t_R _18941_ (.A(_00755_),
    .B(_06927_),
    .C(_06937_),
    .Y(_06996_));
 XOR2x2_ASAP7_75t_R _18942_ (.A(_00754_),
    .B(_06996_),
    .Y(_06997_));
 AND2x2_ASAP7_75t_R _18943_ (.A(_06995_),
    .B(_06997_),
    .Y(_04305_));
 OR4x1_ASAP7_75t_R _18944_ (.A(_00754_),
    .B(_00755_),
    .C(_06927_),
    .D(_06932_),
    .Y(_06998_));
 XOR2x2_ASAP7_75t_R _18945_ (.A(_00753_),
    .B(_06998_),
    .Y(_06999_));
 AND2x2_ASAP7_75t_R _18946_ (.A(_06995_),
    .B(_06999_),
    .Y(_04306_));
 OR5x1_ASAP7_75t_R _18947_ (.A(_00753_),
    .B(_00754_),
    .C(_00755_),
    .D(_06927_),
    .E(_06937_),
    .Y(_07000_));
 NAND2x1_ASAP7_75t_R _18948_ (.A(_00752_),
    .B(_07000_),
    .Y(_07001_));
 OA211x2_ASAP7_75t_R _18949_ (.A1(_06933_),
    .A2(_06937_),
    .B(_07001_),
    .C(_06433_),
    .Y(_04307_));
 BUFx6f_ASAP7_75t_R _18950_ (.A(_00734_),
    .Y(_07002_));
 BUFx3_ASAP7_75t_R _18951_ (.A(_00738_),
    .Y(_07003_));
 BUFx6f_ASAP7_75t_R _18952_ (.A(_00713_),
    .Y(_07004_));
 AND4x1_ASAP7_75t_R _18953_ (.A(_07004_),
    .B(_00741_),
    .C(_00742_),
    .D(_00743_),
    .Y(_07005_));
 AND5x1_ASAP7_75t_R _18954_ (.A(_00732_),
    .B(_00737_),
    .C(_07003_),
    .D(_00740_),
    .E(_07005_),
    .Y(_07006_));
 AND5x2_ASAP7_75t_R _18955_ (.A(_07002_),
    .B(_00735_),
    .C(_00736_),
    .D(_05995_),
    .E(_07006_),
    .Y(_07007_));
 BUFx3_ASAP7_75t_R _18956_ (.A(_00729_),
    .Y(_07008_));
 AND4x1_ASAP7_75t_R _18957_ (.A(_00727_),
    .B(_00728_),
    .C(_07008_),
    .D(_00730_),
    .Y(_07009_));
 AND4x1_ASAP7_75t_R _18958_ (.A(_00721_),
    .B(_00723_),
    .C(_00724_),
    .D(_00731_),
    .Y(_07010_));
 AND5x1_ASAP7_75t_R _18959_ (.A(_00714_),
    .B(_00715_),
    .C(_00720_),
    .D(_00739_),
    .E(_07010_),
    .Y(_07011_));
 AND3x1_ASAP7_75t_R _18960_ (.A(_00718_),
    .B(_00719_),
    .C(_00722_),
    .Y(_07012_));
 OR3x1_ASAP7_75t_R _18961_ (.A(_00716_),
    .B(_00717_),
    .C(_07012_),
    .Y(_07013_));
 AND5x2_ASAP7_75t_R _18962_ (.A(_00725_),
    .B(_00726_),
    .C(_07009_),
    .D(_07011_),
    .E(_07013_),
    .Y(_07014_));
 NAND2x2_ASAP7_75t_R _18963_ (.A(_07007_),
    .B(_07014_),
    .Y(_07015_));
 NOR2x1_ASAP7_75t_R _18964_ (.A(_00703_),
    .B(_07015_),
    .Y(_04308_));
 INVx1_ASAP7_75t_R _18965_ (.A(_07015_),
    .Y(_04309_));
 NOR2x1_ASAP7_75t_R _18966_ (.A(_00706_),
    .B(_07015_),
    .Y(_04310_));
 NOR2x1_ASAP7_75t_R _18967_ (.A(_00705_),
    .B(_07015_),
    .Y(_04311_));
 NOR2x1_ASAP7_75t_R _18968_ (.A(_00704_),
    .B(_07015_),
    .Y(_04312_));
 NOR2x1_ASAP7_75t_R _18969_ (.A(_00702_),
    .B(_07015_),
    .Y(_04313_));
 NOR2x1_ASAP7_75t_R _18970_ (.A(_00701_),
    .B(_07015_),
    .Y(_04314_));
 INVx1_ASAP7_75t_R _18971_ (.A(_07015_),
    .Y(_04315_));
 AND2x2_ASAP7_75t_R _18972_ (.A(_06995_),
    .B(_00050_),
    .Y(_04316_));
 OR4x1_ASAP7_75t_R _18973_ (.A(_00718_),
    .B(_00719_),
    .C(_00722_),
    .D(_02667_),
    .Y(_07016_));
 OR4x1_ASAP7_75t_R _18974_ (.A(_00714_),
    .B(_00715_),
    .C(_00716_),
    .D(_00717_),
    .Y(_07017_));
 OR2x6_ASAP7_75t_R _18975_ (.A(_07016_),
    .B(_07017_),
    .Y(_07018_));
 OR3x1_ASAP7_75t_R _18976_ (.A(_07004_),
    .B(_00743_),
    .C(_07018_),
    .Y(_07019_));
 OAI21x1_ASAP7_75t_R _18977_ (.A1(_07004_),
    .A2(_07018_),
    .B(_00743_),
    .Y(_07020_));
 AND3x1_ASAP7_75t_R _18978_ (.A(_06958_),
    .B(_07019_),
    .C(_07020_),
    .Y(_04317_));
 OR5x2_ASAP7_75t_R _18979_ (.A(_00718_),
    .B(_00719_),
    .C(_00722_),
    .D(_00733_),
    .E(_00050_),
    .Y(_07021_));
 OR2x6_ASAP7_75t_R _18980_ (.A(_07017_),
    .B(_07021_),
    .Y(_07022_));
 OR3x1_ASAP7_75t_R _18981_ (.A(_07004_),
    .B(_00743_),
    .C(_07022_),
    .Y(_07023_));
 XOR2x2_ASAP7_75t_R _18982_ (.A(_00742_),
    .B(_07023_),
    .Y(_07024_));
 AND2x2_ASAP7_75t_R _18983_ (.A(_06995_),
    .B(_07024_),
    .Y(_04318_));
 OR4x1_ASAP7_75t_R _18984_ (.A(_07004_),
    .B(_00742_),
    .C(_00743_),
    .D(_07018_),
    .Y(_07025_));
 XOR2x2_ASAP7_75t_R _18985_ (.A(_00741_),
    .B(_07025_),
    .Y(_07026_));
 AND2x2_ASAP7_75t_R _18986_ (.A(_06995_),
    .B(_07026_),
    .Y(_04319_));
 OR5x2_ASAP7_75t_R _18987_ (.A(_07004_),
    .B(_00740_),
    .C(_00741_),
    .D(_00742_),
    .E(_00743_),
    .Y(_07027_));
 OR5x1_ASAP7_75t_R _18988_ (.A(_07004_),
    .B(_00741_),
    .C(_00742_),
    .D(_00743_),
    .E(_07022_),
    .Y(_07028_));
 NAND2x1_ASAP7_75t_R _18989_ (.A(_00740_),
    .B(_07028_),
    .Y(_07029_));
 OA211x2_ASAP7_75t_R _18990_ (.A1(_07022_),
    .A2(_07027_),
    .B(_07029_),
    .C(_06433_),
    .Y(_04320_));
 OR4x1_ASAP7_75t_R _18991_ (.A(_00739_),
    .B(_07016_),
    .C(_07017_),
    .D(_07027_),
    .Y(_07030_));
 OAI21x1_ASAP7_75t_R _18992_ (.A1(_07018_),
    .A2(_07027_),
    .B(_00739_),
    .Y(_07031_));
 AND3x1_ASAP7_75t_R _18993_ (.A(_06958_),
    .B(_07030_),
    .C(_07031_),
    .Y(_04321_));
 OR4x1_ASAP7_75t_R _18994_ (.A(_00739_),
    .B(_07017_),
    .C(_07021_),
    .D(_07027_),
    .Y(_07032_));
 XOR2x2_ASAP7_75t_R _18995_ (.A(_07003_),
    .B(_07032_),
    .Y(_07033_));
 AND2x2_ASAP7_75t_R _18996_ (.A(_06995_),
    .B(_07033_),
    .Y(_04322_));
 OR3x1_ASAP7_75t_R _18997_ (.A(_00737_),
    .B(_07003_),
    .C(_07030_),
    .Y(_07034_));
 OAI21x1_ASAP7_75t_R _18998_ (.A1(_07003_),
    .A2(_07030_),
    .B(_00737_),
    .Y(_07035_));
 AND3x1_ASAP7_75t_R _18999_ (.A(_06958_),
    .B(_07034_),
    .C(_07035_),
    .Y(_04323_));
 OR3x1_ASAP7_75t_R _19000_ (.A(_00737_),
    .B(_07003_),
    .C(_07032_),
    .Y(_07036_));
 XOR2x2_ASAP7_75t_R _19001_ (.A(_00736_),
    .B(_07036_),
    .Y(_07037_));
 AND2x2_ASAP7_75t_R _19002_ (.A(_06995_),
    .B(_07037_),
    .Y(_04324_));
 OR5x2_ASAP7_75t_R _19003_ (.A(_00735_),
    .B(_00736_),
    .C(_00737_),
    .D(_07003_),
    .E(_07030_),
    .Y(_07038_));
 OR4x1_ASAP7_75t_R _19004_ (.A(_00736_),
    .B(_00737_),
    .C(_07003_),
    .D(_07030_),
    .Y(_07039_));
 NAND2x1_ASAP7_75t_R _19005_ (.A(_00735_),
    .B(_07039_),
    .Y(_07040_));
 AND3x1_ASAP7_75t_R _19006_ (.A(_06958_),
    .B(_07038_),
    .C(_07040_),
    .Y(_04325_));
 OR5x2_ASAP7_75t_R _19007_ (.A(_00735_),
    .B(_00736_),
    .C(_00737_),
    .D(_07003_),
    .E(_07032_),
    .Y(_07041_));
 XOR2x2_ASAP7_75t_R _19008_ (.A(_07002_),
    .B(_07041_),
    .Y(_07042_));
 AND2x2_ASAP7_75t_R _19009_ (.A(_06995_),
    .B(_07042_),
    .Y(_04326_));
 NOR2x1_ASAP7_75t_R _19010_ (.A(_06272_),
    .B(_02668_),
    .Y(_04327_));
 BUFx6f_ASAP7_75t_R _19011_ (.A(_06386_),
    .Y(_07043_));
 OR3x1_ASAP7_75t_R _19012_ (.A(_00732_),
    .B(_07002_),
    .C(_07038_),
    .Y(_07044_));
 OAI21x1_ASAP7_75t_R _19013_ (.A1(_07002_),
    .A2(_07038_),
    .B(_00732_),
    .Y(_07045_));
 AND3x1_ASAP7_75t_R _19014_ (.A(_07043_),
    .B(_07044_),
    .C(_07045_),
    .Y(_04328_));
 OR3x1_ASAP7_75t_R _19015_ (.A(_00732_),
    .B(_07002_),
    .C(_07041_),
    .Y(_07046_));
 XOR2x2_ASAP7_75t_R _19016_ (.A(_00731_),
    .B(_07046_),
    .Y(_07047_));
 AND2x2_ASAP7_75t_R _19017_ (.A(_06995_),
    .B(_07047_),
    .Y(_04329_));
 OR5x1_ASAP7_75t_R _19018_ (.A(_00730_),
    .B(_00731_),
    .C(_00732_),
    .D(_07002_),
    .E(_07038_),
    .Y(_07048_));
 BUFx3_ASAP7_75t_R _19019_ (.A(_07048_),
    .Y(_07049_));
 OR4x1_ASAP7_75t_R _19020_ (.A(_00731_),
    .B(_00732_),
    .C(_07002_),
    .D(_07038_),
    .Y(_07050_));
 NAND2x1_ASAP7_75t_R _19021_ (.A(_00730_),
    .B(_07050_),
    .Y(_07051_));
 AND3x1_ASAP7_75t_R _19022_ (.A(_07043_),
    .B(_07049_),
    .C(_07051_),
    .Y(_04330_));
 OR5x2_ASAP7_75t_R _19023_ (.A(_00730_),
    .B(_00731_),
    .C(_00732_),
    .D(_07002_),
    .E(_07041_),
    .Y(_07052_));
 XOR2x2_ASAP7_75t_R _19024_ (.A(_07008_),
    .B(_07052_),
    .Y(_07053_));
 AND2x2_ASAP7_75t_R _19025_ (.A(_06995_),
    .B(_07053_),
    .Y(_04331_));
 OR3x1_ASAP7_75t_R _19026_ (.A(_00728_),
    .B(_07008_),
    .C(_07049_),
    .Y(_07054_));
 OAI21x1_ASAP7_75t_R _19027_ (.A1(_07008_),
    .A2(_07049_),
    .B(_00728_),
    .Y(_07055_));
 AND3x1_ASAP7_75t_R _19028_ (.A(_07043_),
    .B(_07054_),
    .C(_07055_),
    .Y(_04332_));
 BUFx6f_ASAP7_75t_R _19029_ (.A(_06547_),
    .Y(_07056_));
 OR3x1_ASAP7_75t_R _19030_ (.A(_00728_),
    .B(_07008_),
    .C(_07052_),
    .Y(_07057_));
 XOR2x2_ASAP7_75t_R _19031_ (.A(_00727_),
    .B(_07057_),
    .Y(_07058_));
 AND2x2_ASAP7_75t_R _19032_ (.A(_07056_),
    .B(_07058_),
    .Y(_04333_));
 OR4x1_ASAP7_75t_R _19033_ (.A(_00727_),
    .B(_00728_),
    .C(_07008_),
    .D(_07049_),
    .Y(_07059_));
 XOR2x2_ASAP7_75t_R _19034_ (.A(_00726_),
    .B(_07059_),
    .Y(_07060_));
 AND2x2_ASAP7_75t_R _19035_ (.A(_07056_),
    .B(_07060_),
    .Y(_04334_));
 OR5x1_ASAP7_75t_R _19036_ (.A(_00726_),
    .B(_00727_),
    .C(_00728_),
    .D(_07008_),
    .E(_07052_),
    .Y(_07061_));
 XOR2x2_ASAP7_75t_R _19037_ (.A(_00725_),
    .B(_07061_),
    .Y(_07062_));
 AND2x2_ASAP7_75t_R _19038_ (.A(_07056_),
    .B(_07062_),
    .Y(_04335_));
 OR5x2_ASAP7_75t_R _19039_ (.A(_00725_),
    .B(_00726_),
    .C(_00727_),
    .D(_00728_),
    .E(_07008_),
    .Y(_07063_));
 OR3x1_ASAP7_75t_R _19040_ (.A(_00724_),
    .B(_07049_),
    .C(_07063_),
    .Y(_07064_));
 OAI21x1_ASAP7_75t_R _19041_ (.A1(_07049_),
    .A2(_07063_),
    .B(_00724_),
    .Y(_07065_));
 AND3x1_ASAP7_75t_R _19042_ (.A(_07043_),
    .B(_07064_),
    .C(_07065_),
    .Y(_04336_));
 OR3x1_ASAP7_75t_R _19043_ (.A(_00724_),
    .B(_07052_),
    .C(_07063_),
    .Y(_07066_));
 XOR2x2_ASAP7_75t_R _19044_ (.A(_00723_),
    .B(_07066_),
    .Y(_07067_));
 AND2x2_ASAP7_75t_R _19045_ (.A(_07056_),
    .B(_07067_),
    .Y(_04337_));
 XOR2x2_ASAP7_75t_R _19046_ (.A(_00722_),
    .B(_02667_),
    .Y(_07068_));
 AND2x2_ASAP7_75t_R _19047_ (.A(_07056_),
    .B(_07068_),
    .Y(_04338_));
 OR4x1_ASAP7_75t_R _19048_ (.A(_00723_),
    .B(_00724_),
    .C(_07049_),
    .D(_07063_),
    .Y(_07069_));
 XOR2x2_ASAP7_75t_R _19049_ (.A(_00721_),
    .B(_07069_),
    .Y(_07070_));
 AND2x2_ASAP7_75t_R _19050_ (.A(_07056_),
    .B(_07070_),
    .Y(_04339_));
 OR5x1_ASAP7_75t_R _19051_ (.A(_00721_),
    .B(_00723_),
    .C(_00724_),
    .D(_07052_),
    .E(_07063_),
    .Y(_07071_));
 XOR2x2_ASAP7_75t_R _19052_ (.A(_00720_),
    .B(_07071_),
    .Y(_07072_));
 AND2x2_ASAP7_75t_R _19053_ (.A(_07056_),
    .B(_07072_),
    .Y(_04340_));
 OR3x1_ASAP7_75t_R _19054_ (.A(_00722_),
    .B(_00733_),
    .C(_00050_),
    .Y(_07073_));
 XOR2x2_ASAP7_75t_R _19055_ (.A(_00719_),
    .B(_07073_),
    .Y(_07074_));
 AND2x2_ASAP7_75t_R _19056_ (.A(_07056_),
    .B(_07074_),
    .Y(_04341_));
 OR3x1_ASAP7_75t_R _19057_ (.A(_00719_),
    .B(_00722_),
    .C(_02667_),
    .Y(_07075_));
 NAND2x1_ASAP7_75t_R _19058_ (.A(_00718_),
    .B(_07075_),
    .Y(_07076_));
 AND3x1_ASAP7_75t_R _19059_ (.A(_07043_),
    .B(_07016_),
    .C(_07076_),
    .Y(_04342_));
 XOR2x2_ASAP7_75t_R _19060_ (.A(_00717_),
    .B(_07021_),
    .Y(_07077_));
 AND2x2_ASAP7_75t_R _19061_ (.A(_07056_),
    .B(_07077_),
    .Y(_04343_));
 OR3x1_ASAP7_75t_R _19062_ (.A(_00716_),
    .B(_00717_),
    .C(_07016_),
    .Y(_07078_));
 OAI21x1_ASAP7_75t_R _19063_ (.A1(_00717_),
    .A2(_07016_),
    .B(_00716_),
    .Y(_07079_));
 AND3x1_ASAP7_75t_R _19064_ (.A(_07043_),
    .B(_07078_),
    .C(_07079_),
    .Y(_04344_));
 OR3x1_ASAP7_75t_R _19065_ (.A(_00716_),
    .B(_00717_),
    .C(_07021_),
    .Y(_07080_));
 XOR2x2_ASAP7_75t_R _19066_ (.A(_00715_),
    .B(_07080_),
    .Y(_07081_));
 AND2x2_ASAP7_75t_R _19067_ (.A(_07056_),
    .B(_07081_),
    .Y(_04345_));
 OR4x1_ASAP7_75t_R _19068_ (.A(_00715_),
    .B(_00716_),
    .C(_00717_),
    .D(_07016_),
    .Y(_07082_));
 NAND2x1_ASAP7_75t_R _19069_ (.A(_00714_),
    .B(_07082_),
    .Y(_07083_));
 AND3x1_ASAP7_75t_R _19070_ (.A(_07043_),
    .B(_07018_),
    .C(_07083_),
    .Y(_04346_));
 BUFx12f_ASAP7_75t_R _19071_ (.A(_08598_),
    .Y(_07084_));
 BUFx6f_ASAP7_75t_R _19072_ (.A(_07084_),
    .Y(_07085_));
 XOR2x2_ASAP7_75t_R _19073_ (.A(_07004_),
    .B(_07022_),
    .Y(_07086_));
 AND2x2_ASAP7_75t_R _19074_ (.A(_07085_),
    .B(_07086_),
    .Y(_04347_));
 AND2x2_ASAP7_75t_R _19075_ (.A(_07085_),
    .B(_00024_),
    .Y(_04348_));
 INVx1_ASAP7_75t_R _19076_ (.A(_02274_),
    .Y(_07087_));
 OR2x2_ASAP7_75t_R _19077_ (.A(_00786_),
    .B(_00787_),
    .Y(_07088_));
 NAND2x1_ASAP7_75t_R _19078_ (.A(_00784_),
    .B(_00785_),
    .Y(_07089_));
 OR4x1_ASAP7_75t_R _19079_ (.A(_00783_),
    .B(_00788_),
    .C(_07088_),
    .D(_07089_),
    .Y(_07090_));
 OR2x6_ASAP7_75t_R _19080_ (.A(_00747_),
    .B(_00748_),
    .Y(_07091_));
 NAND2x1_ASAP7_75t_R _19081_ (.A(_00745_),
    .B(_00746_),
    .Y(_07092_));
 OA21x2_ASAP7_75t_R _19082_ (.A1(_07091_),
    .A2(_07092_),
    .B(\xs[3].cli1.i[39] ),
    .Y(_07093_));
 OR4x1_ASAP7_75t_R _19083_ (.A(_00744_),
    .B(\xs[3].cli1.i[32] ),
    .C(_07091_),
    .D(_07092_),
    .Y(_07094_));
 OA21x2_ASAP7_75t_R _19084_ (.A1(_02281_),
    .A2(_07093_),
    .B(_07094_),
    .Y(_07095_));
 INVx1_ASAP7_75t_R _19085_ (.A(_02281_),
    .Y(_07096_));
 OA21x2_ASAP7_75t_R _19086_ (.A1(_07088_),
    .A2(_07089_),
    .B(\peo[6][39] ),
    .Y(_07097_));
 OR3x1_ASAP7_75t_R _19087_ (.A(_07096_),
    .B(_07094_),
    .C(_07097_),
    .Y(_07098_));
 OA21x2_ASAP7_75t_R _19088_ (.A1(_07090_),
    .A2(_07095_),
    .B(_07098_),
    .Y(_07099_));
 AND4x1_ASAP7_75t_R _19089_ (.A(_07087_),
    .B(_02275_),
    .C(_02281_),
    .D(_07099_),
    .Y(_07100_));
 NAND2x1_ASAP7_75t_R _19090_ (.A(_02285_),
    .B(_07100_),
    .Y(_07101_));
 INVx1_ASAP7_75t_R _19091_ (.A(_02275_),
    .Y(_07102_));
 AND2x2_ASAP7_75t_R _19092_ (.A(_00745_),
    .B(_00746_),
    .Y(_07103_));
 AND5x1_ASAP7_75t_R _19093_ (.A(\xs[3].cli1.i[39] ),
    .B(\xs[3].cli1.i[34] ),
    .C(\xs[3].cli1.i[33] ),
    .D(_00749_),
    .E(_07103_),
    .Y(_07104_));
 AO21x1_ASAP7_75t_R _19094_ (.A1(_07104_),
    .A2(_07097_),
    .B(_07093_),
    .Y(_07105_));
 OA31x2_ASAP7_75t_R _19095_ (.A1(_00749_),
    .A2(_07091_),
    .A3(_07092_),
    .B1(\xs[3].cli1.i[39] ),
    .Y(_07106_));
 AND2x2_ASAP7_75t_R _19096_ (.A(_02274_),
    .B(_00024_),
    .Y(_07107_));
 AO32x1_ASAP7_75t_R _19097_ (.A1(_07087_),
    .A2(_02281_),
    .A3(_07106_),
    .B1(_07107_),
    .B2(_07093_),
    .Y(_07108_));
 AO32x2_ASAP7_75t_R _19098_ (.A1(_07087_),
    .A2(_07102_),
    .A3(_07105_),
    .B1(_07108_),
    .B2(_07097_),
    .Y(_07109_));
 NOR2x1_ASAP7_75t_R _19099_ (.A(_07094_),
    .B(_07109_),
    .Y(_07110_));
 OR3x1_ASAP7_75t_R _19100_ (.A(\peo[6][0] ),
    .B(_07100_),
    .C(_07110_),
    .Y(_07111_));
 OR3x1_ASAP7_75t_R _19101_ (.A(\peo[7][0] ),
    .B(_07094_),
    .C(_07109_),
    .Y(_07112_));
 AND4x1_ASAP7_75t_R _19102_ (.A(_08999_),
    .B(_07101_),
    .C(_07111_),
    .D(_07112_),
    .Y(_04349_));
 NAND2x2_ASAP7_75t_R _19103_ (.A(_08528_),
    .B(_07100_),
    .Y(_07113_));
 NOR2x1_ASAP7_75t_R _19104_ (.A(_02284_),
    .B(_07113_),
    .Y(_04350_));
 NOR2x1_ASAP7_75t_R _19105_ (.A(_02283_),
    .B(_07113_),
    .Y(_04351_));
 NOR2x1_ASAP7_75t_R _19106_ (.A(_02282_),
    .B(_07113_),
    .Y(_04352_));
 NOR2x1_ASAP7_75t_R _19107_ (.A(_02273_),
    .B(_07113_),
    .Y(_04353_));
 NOR2x1_ASAP7_75t_R _19108_ (.A(_02272_),
    .B(_07113_),
    .Y(_04354_));
 NOR2x1_ASAP7_75t_R _19109_ (.A(_07090_),
    .B(_07093_),
    .Y(_07114_));
 OR4x1_ASAP7_75t_R _19110_ (.A(_02274_),
    .B(_07102_),
    .C(_02281_),
    .D(_07114_),
    .Y(_07115_));
 NOR2x1_ASAP7_75t_R _19111_ (.A(_02285_),
    .B(_07115_),
    .Y(_07116_));
 AO21x1_ASAP7_75t_R _19112_ (.A1(\peo[6][0] ),
    .A2(_07115_),
    .B(_07116_),
    .Y(_07117_));
 NAND2x1_ASAP7_75t_R _19113_ (.A(_00751_),
    .B(_07109_),
    .Y(_07118_));
 OA211x2_ASAP7_75t_R _19114_ (.A1(_07109_),
    .A2(_07117_),
    .B(_07118_),
    .C(_06433_),
    .Y(_04355_));
 OR2x2_ASAP7_75t_R _19115_ (.A(_08683_),
    .B(_07115_),
    .Y(_07119_));
 BUFx3_ASAP7_75t_R _19116_ (.A(_07119_),
    .Y(_07120_));
 NOR2x1_ASAP7_75t_R _19117_ (.A(_02284_),
    .B(_07120_),
    .Y(_04356_));
 NOR2x1_ASAP7_75t_R _19118_ (.A(_02283_),
    .B(_07120_),
    .Y(_04357_));
 NOR2x1_ASAP7_75t_R _19119_ (.A(_02282_),
    .B(_07120_),
    .Y(_04358_));
 NOR2x1_ASAP7_75t_R _19120_ (.A(_02273_),
    .B(_07120_),
    .Y(_04359_));
 NOR2x1_ASAP7_75t_R _19121_ (.A(_02272_),
    .B(_07120_),
    .Y(_04360_));
 OAI21x1_ASAP7_75t_R _19122_ (.A1(_02274_),
    .A2(_02275_),
    .B(_07093_),
    .Y(_07121_));
 AO21x1_ASAP7_75t_R _19123_ (.A1(_07097_),
    .A2(_07108_),
    .B(_07121_),
    .Y(_07122_));
 BUFx6f_ASAP7_75t_R _19124_ (.A(_07122_),
    .Y(_07123_));
 OR2x2_ASAP7_75t_R _19125_ (.A(\peo[7][0] ),
    .B(_07123_),
    .Y(_07124_));
 NAND2x1_ASAP7_75t_R _19126_ (.A(_00790_),
    .B(_07123_),
    .Y(_07125_));
 AOI21x1_ASAP7_75t_R _19127_ (.A1(_02275_),
    .A2(_07099_),
    .B(_02274_),
    .Y(_07126_));
 BUFx6f_ASAP7_75t_R _19128_ (.A(_07126_),
    .Y(_07127_));
 NOR2x1_ASAP7_75t_R _19129_ (.A(_10826_),
    .B(_07127_),
    .Y(_07128_));
 NOR2x1_ASAP7_75t_R _19130_ (.A(_06206_),
    .B(_02285_),
    .Y(_07129_));
 AO32x1_ASAP7_75t_R _19131_ (.A1(_07124_),
    .A2(_07125_),
    .A3(_07128_),
    .B1(_07129_),
    .B2(_07127_),
    .Y(_04361_));
 NAND2x2_ASAP7_75t_R _19132_ (.A(_09029_),
    .B(_07126_),
    .Y(_07130_));
 NOR2x1_ASAP7_75t_R _19133_ (.A(_02284_),
    .B(_07130_),
    .Y(_04362_));
 NOR2x1_ASAP7_75t_R _19134_ (.A(_02283_),
    .B(_07130_),
    .Y(_04363_));
 NOR2x1_ASAP7_75t_R _19135_ (.A(_02282_),
    .B(_07130_),
    .Y(_04364_));
 NOR2x1_ASAP7_75t_R _19136_ (.A(_00749_),
    .B(_07123_),
    .Y(_07131_));
 AO21x1_ASAP7_75t_R _19137_ (.A1(\peo[6][32] ),
    .A2(_07123_),
    .B(_07131_),
    .Y(_07132_));
 AND3x1_ASAP7_75t_R _19138_ (.A(_08599_),
    .B(_07096_),
    .C(_07127_),
    .Y(_07133_));
 AO21x1_ASAP7_75t_R _19139_ (.A1(_07128_),
    .A2(_07132_),
    .B(_07133_),
    .Y(_04365_));
 NOR2x1_ASAP7_75t_R _19140_ (.A(_00744_),
    .B(_07109_),
    .Y(_07134_));
 AOI22x1_ASAP7_75t_R _19141_ (.A1(_00787_),
    .A2(_07123_),
    .B1(_07134_),
    .B2(_00748_),
    .Y(_07135_));
 NAND2x1_ASAP7_75t_R _19142_ (.A(_02280_),
    .B(_07127_),
    .Y(_07136_));
 OA211x2_ASAP7_75t_R _19143_ (.A1(_07127_),
    .A2(_07135_),
    .B(_07136_),
    .C(_06433_),
    .Y(_04366_));
 AOI22x1_ASAP7_75t_R _19144_ (.A1(_00786_),
    .A2(_07123_),
    .B1(_07134_),
    .B2(_00747_),
    .Y(_07137_));
 NAND2x1_ASAP7_75t_R _19145_ (.A(_02279_),
    .B(_07127_),
    .Y(_07138_));
 OA211x2_ASAP7_75t_R _19146_ (.A1(_07127_),
    .A2(_07137_),
    .B(_07138_),
    .C(_06433_),
    .Y(_04367_));
 OR2x2_ASAP7_75t_R _19147_ (.A(\xs[3].cli1.i[35] ),
    .B(_07123_),
    .Y(_07139_));
 NAND2x1_ASAP7_75t_R _19148_ (.A(_00785_),
    .B(_07123_),
    .Y(_07140_));
 NOR2x1_ASAP7_75t_R _19149_ (.A(_06206_),
    .B(_02278_),
    .Y(_07141_));
 AO32x1_ASAP7_75t_R _19150_ (.A1(_07128_),
    .A2(_07139_),
    .A3(_07140_),
    .B1(_07141_),
    .B2(_07127_),
    .Y(_04368_));
 OR2x2_ASAP7_75t_R _19151_ (.A(\xs[3].cli1.i[36] ),
    .B(_07123_),
    .Y(_07142_));
 NAND2x1_ASAP7_75t_R _19152_ (.A(_00784_),
    .B(_07123_),
    .Y(_07143_));
 NOR2x1_ASAP7_75t_R _19153_ (.A(_06206_),
    .B(_02277_),
    .Y(_07144_));
 AO32x1_ASAP7_75t_R _19154_ (.A1(_07128_),
    .A2(_07142_),
    .A3(_07143_),
    .B1(_07144_),
    .B2(_07127_),
    .Y(_04369_));
 NOR2x1_ASAP7_75t_R _19155_ (.A(_02276_),
    .B(_07130_),
    .Y(_04370_));
 OR4x1_ASAP7_75t_R _19156_ (.A(_08684_),
    .B(_02274_),
    .C(_07102_),
    .D(_07099_),
    .Y(_07145_));
 INVx1_ASAP7_75t_R _19157_ (.A(_07145_),
    .Y(_04371_));
 OR3x1_ASAP7_75t_R _19158_ (.A(_07093_),
    .B(_07097_),
    .C(_07127_),
    .Y(_07146_));
 AND2x2_ASAP7_75t_R _19159_ (.A(_07085_),
    .B(_07146_),
    .Y(_04372_));
 NOR2x1_ASAP7_75t_R _19160_ (.A(_02273_),
    .B(_07130_),
    .Y(_04373_));
 NOR2x1_ASAP7_75t_R _19161_ (.A(_02272_),
    .B(_07130_),
    .Y(_04374_));
 BUFx12f_ASAP7_75t_R _19162_ (.A(_11465_),
    .Y(_07147_));
 BUFx3_ASAP7_75t_R _19163_ (.A(_00648_),
    .Y(_07148_));
 AND4x1_ASAP7_75t_R _19164_ (.A(_07148_),
    .B(_00676_),
    .C(_00677_),
    .D(_00678_),
    .Y(_07149_));
 AND5x1_ASAP7_75t_R _19165_ (.A(_00667_),
    .B(_00672_),
    .C(_00673_),
    .D(_00675_),
    .E(_07149_),
    .Y(_07150_));
 AND5x2_ASAP7_75t_R _19166_ (.A(_00669_),
    .B(_00670_),
    .C(_00671_),
    .D(_07147_),
    .E(_07150_),
    .Y(_07151_));
 BUFx3_ASAP7_75t_R _19167_ (.A(_00664_),
    .Y(_07152_));
 AND4x1_ASAP7_75t_R _19168_ (.A(_00662_),
    .B(_00663_),
    .C(_07152_),
    .D(_00665_),
    .Y(_07153_));
 AND4x1_ASAP7_75t_R _19169_ (.A(_00656_),
    .B(_00658_),
    .C(_00659_),
    .D(_00666_),
    .Y(_07154_));
 AND5x1_ASAP7_75t_R _19170_ (.A(_00649_),
    .B(_00650_),
    .C(_00655_),
    .D(_00674_),
    .E(_07154_),
    .Y(_07155_));
 AND3x1_ASAP7_75t_R _19171_ (.A(_00653_),
    .B(_00654_),
    .C(_00657_),
    .Y(_07156_));
 OR3x1_ASAP7_75t_R _19172_ (.A(_00651_),
    .B(_00652_),
    .C(_07156_),
    .Y(_07157_));
 AND5x2_ASAP7_75t_R _19173_ (.A(_00660_),
    .B(_00661_),
    .C(_07153_),
    .D(_07155_),
    .E(_07157_),
    .Y(_07158_));
 NAND2x2_ASAP7_75t_R _19174_ (.A(_07151_),
    .B(_07158_),
    .Y(_07159_));
 NOR2x1_ASAP7_75t_R _19175_ (.A(_00605_),
    .B(_07159_),
    .Y(_04375_));
 INVx1_ASAP7_75t_R _19176_ (.A(_07159_),
    .Y(_04376_));
 NOR2x1_ASAP7_75t_R _19177_ (.A(_00608_),
    .B(_07159_),
    .Y(_04377_));
 NOR2x1_ASAP7_75t_R _19178_ (.A(_00607_),
    .B(_07159_),
    .Y(_04378_));
 NOR2x1_ASAP7_75t_R _19179_ (.A(_00606_),
    .B(_07159_),
    .Y(_04379_));
 NOR2x1_ASAP7_75t_R _19180_ (.A(_00604_),
    .B(_07159_),
    .Y(_04380_));
 NOR2x1_ASAP7_75t_R _19181_ (.A(_00603_),
    .B(_07159_),
    .Y(_04381_));
 INVx1_ASAP7_75t_R _19182_ (.A(_07159_),
    .Y(_04382_));
 AND2x2_ASAP7_75t_R _19183_ (.A(_07085_),
    .B(_00051_),
    .Y(_04383_));
 OR4x1_ASAP7_75t_R _19184_ (.A(_00653_),
    .B(_00654_),
    .C(_00657_),
    .D(_02661_),
    .Y(_07160_));
 OR4x1_ASAP7_75t_R _19185_ (.A(_00649_),
    .B(_00650_),
    .C(_00651_),
    .D(_00652_),
    .Y(_07161_));
 OR2x6_ASAP7_75t_R _19186_ (.A(_07160_),
    .B(_07161_),
    .Y(_07162_));
 OR3x1_ASAP7_75t_R _19187_ (.A(_07148_),
    .B(_00678_),
    .C(_07162_),
    .Y(_07163_));
 OAI21x1_ASAP7_75t_R _19188_ (.A1(_07148_),
    .A2(_07162_),
    .B(_00678_),
    .Y(_07164_));
 AND3x1_ASAP7_75t_R _19189_ (.A(_07043_),
    .B(_07163_),
    .C(_07164_),
    .Y(_04384_));
 OR5x2_ASAP7_75t_R _19190_ (.A(_00653_),
    .B(_00654_),
    .C(_00657_),
    .D(_00668_),
    .E(_00051_),
    .Y(_07165_));
 OR2x2_ASAP7_75t_R _19191_ (.A(_07161_),
    .B(_07165_),
    .Y(_07166_));
 OR3x1_ASAP7_75t_R _19192_ (.A(_07148_),
    .B(_00678_),
    .C(_07166_),
    .Y(_07167_));
 XOR2x2_ASAP7_75t_R _19193_ (.A(_00677_),
    .B(_07167_),
    .Y(_07168_));
 AND2x2_ASAP7_75t_R _19194_ (.A(_07085_),
    .B(_07168_),
    .Y(_04385_));
 OR4x1_ASAP7_75t_R _19195_ (.A(_07148_),
    .B(_00676_),
    .C(_00677_),
    .D(_00678_),
    .Y(_07169_));
 OR3x2_ASAP7_75t_R _19196_ (.A(_07160_),
    .B(_07161_),
    .C(_07169_),
    .Y(_07170_));
 OR4x1_ASAP7_75t_R _19197_ (.A(_07148_),
    .B(_00677_),
    .C(_00678_),
    .D(_07162_),
    .Y(_07171_));
 NAND2x1_ASAP7_75t_R _19198_ (.A(_00676_),
    .B(_07171_),
    .Y(_07172_));
 AND3x1_ASAP7_75t_R _19199_ (.A(_07043_),
    .B(_07170_),
    .C(_07172_),
    .Y(_04386_));
 OR3x2_ASAP7_75t_R _19200_ (.A(_07161_),
    .B(_07165_),
    .C(_07169_),
    .Y(_07173_));
 XOR2x2_ASAP7_75t_R _19201_ (.A(_00675_),
    .B(_07173_),
    .Y(_07174_));
 AND2x2_ASAP7_75t_R _19202_ (.A(_07085_),
    .B(_07174_),
    .Y(_04387_));
 OR3x1_ASAP7_75t_R _19203_ (.A(_00674_),
    .B(_00675_),
    .C(_07170_),
    .Y(_07175_));
 OAI21x1_ASAP7_75t_R _19204_ (.A1(_00675_),
    .A2(_07170_),
    .B(_00674_),
    .Y(_07176_));
 AND3x1_ASAP7_75t_R _19205_ (.A(_07043_),
    .B(_07175_),
    .C(_07176_),
    .Y(_04388_));
 OR3x1_ASAP7_75t_R _19206_ (.A(_00674_),
    .B(_00675_),
    .C(_07173_),
    .Y(_07177_));
 XOR2x2_ASAP7_75t_R _19207_ (.A(_00673_),
    .B(_07177_),
    .Y(_07178_));
 AND2x2_ASAP7_75t_R _19208_ (.A(_07085_),
    .B(_07178_),
    .Y(_04389_));
 OR4x1_ASAP7_75t_R _19209_ (.A(_00672_),
    .B(_00673_),
    .C(_00674_),
    .D(_00675_),
    .Y(_07179_));
 OR4x1_ASAP7_75t_R _19210_ (.A(_00673_),
    .B(_00674_),
    .C(_00675_),
    .D(_07170_),
    .Y(_07180_));
 NAND2x1_ASAP7_75t_R _19211_ (.A(_00672_),
    .B(_07180_),
    .Y(_07181_));
 OA211x2_ASAP7_75t_R _19212_ (.A1(_07170_),
    .A2(_07179_),
    .B(_07181_),
    .C(_06433_),
    .Y(_04390_));
 BUFx6f_ASAP7_75t_R _19213_ (.A(_06386_),
    .Y(_07182_));
 OR3x1_ASAP7_75t_R _19214_ (.A(_00671_),
    .B(_07173_),
    .C(_07179_),
    .Y(_07183_));
 OAI21x1_ASAP7_75t_R _19215_ (.A1(_07173_),
    .A2(_07179_),
    .B(_00671_),
    .Y(_07184_));
 AND3x1_ASAP7_75t_R _19216_ (.A(_07182_),
    .B(_07183_),
    .C(_07184_),
    .Y(_04391_));
 OR3x1_ASAP7_75t_R _19217_ (.A(_00671_),
    .B(_07170_),
    .C(_07179_),
    .Y(_07185_));
 XOR2x2_ASAP7_75t_R _19218_ (.A(_00670_),
    .B(_07185_),
    .Y(_07186_));
 AND2x2_ASAP7_75t_R _19219_ (.A(_07085_),
    .B(_07186_),
    .Y(_04392_));
 OR5x2_ASAP7_75t_R _19220_ (.A(_00669_),
    .B(_00670_),
    .C(_00671_),
    .D(_07173_),
    .E(_07179_),
    .Y(_07187_));
 OR4x1_ASAP7_75t_R _19221_ (.A(_00670_),
    .B(_00671_),
    .C(_07173_),
    .D(_07179_),
    .Y(_07188_));
 NAND2x1_ASAP7_75t_R _19222_ (.A(_00669_),
    .B(_07188_),
    .Y(_07189_));
 AND3x1_ASAP7_75t_R _19223_ (.A(_07182_),
    .B(_07187_),
    .C(_07189_),
    .Y(_04393_));
 BUFx12f_ASAP7_75t_R _19224_ (.A(_10012_),
    .Y(_07190_));
 NOR2x1_ASAP7_75t_R _19225_ (.A(_07190_),
    .B(_02662_),
    .Y(_04394_));
 OR5x2_ASAP7_75t_R _19226_ (.A(_00669_),
    .B(_00670_),
    .C(_00671_),
    .D(_07170_),
    .E(_07179_),
    .Y(_07191_));
 XOR2x2_ASAP7_75t_R _19227_ (.A(_00667_),
    .B(_07191_),
    .Y(_07192_));
 AND2x2_ASAP7_75t_R _19228_ (.A(_07085_),
    .B(_07192_),
    .Y(_04395_));
 OR3x1_ASAP7_75t_R _19229_ (.A(_00666_),
    .B(_00667_),
    .C(_07187_),
    .Y(_07193_));
 OAI21x1_ASAP7_75t_R _19230_ (.A1(_00667_),
    .A2(_07187_),
    .B(_00666_),
    .Y(_07194_));
 AND3x1_ASAP7_75t_R _19231_ (.A(_07182_),
    .B(_07193_),
    .C(_07194_),
    .Y(_04396_));
 OR4x1_ASAP7_75t_R _19232_ (.A(_00665_),
    .B(_00666_),
    .C(_00667_),
    .D(_07191_),
    .Y(_07195_));
 OR3x1_ASAP7_75t_R _19233_ (.A(_00666_),
    .B(_00667_),
    .C(_07191_),
    .Y(_07196_));
 NAND2x1_ASAP7_75t_R _19234_ (.A(_00665_),
    .B(_07196_),
    .Y(_07197_));
 AND3x1_ASAP7_75t_R _19235_ (.A(_07182_),
    .B(_07195_),
    .C(_07197_),
    .Y(_04397_));
 OR4x1_ASAP7_75t_R _19236_ (.A(_00665_),
    .B(_00666_),
    .C(_00667_),
    .D(_07187_),
    .Y(_07198_));
 XOR2x2_ASAP7_75t_R _19237_ (.A(_07152_),
    .B(_07198_),
    .Y(_07199_));
 AND2x2_ASAP7_75t_R _19238_ (.A(_07085_),
    .B(_07199_),
    .Y(_04398_));
 OR3x1_ASAP7_75t_R _19239_ (.A(_00663_),
    .B(_07152_),
    .C(_07195_),
    .Y(_07200_));
 OAI21x1_ASAP7_75t_R _19240_ (.A1(_07152_),
    .A2(_07195_),
    .B(_00663_),
    .Y(_07201_));
 AND3x1_ASAP7_75t_R _19241_ (.A(_07182_),
    .B(_07200_),
    .C(_07201_),
    .Y(_04399_));
 BUFx6f_ASAP7_75t_R _19242_ (.A(_07084_),
    .Y(_07202_));
 OR3x1_ASAP7_75t_R _19243_ (.A(_00663_),
    .B(_07152_),
    .C(_07198_),
    .Y(_07203_));
 XOR2x2_ASAP7_75t_R _19244_ (.A(_00662_),
    .B(_07203_),
    .Y(_07204_));
 AND2x2_ASAP7_75t_R _19245_ (.A(_07202_),
    .B(_07204_),
    .Y(_04400_));
 OR4x1_ASAP7_75t_R _19246_ (.A(_00662_),
    .B(_00663_),
    .C(_07152_),
    .D(_07195_),
    .Y(_07205_));
 XOR2x2_ASAP7_75t_R _19247_ (.A(_00661_),
    .B(_07205_),
    .Y(_07206_));
 AND2x2_ASAP7_75t_R _19248_ (.A(_07202_),
    .B(_07206_),
    .Y(_04401_));
 OR5x1_ASAP7_75t_R _19249_ (.A(_00661_),
    .B(_00662_),
    .C(_00663_),
    .D(_07152_),
    .E(_07198_),
    .Y(_07207_));
 XOR2x2_ASAP7_75t_R _19250_ (.A(_00660_),
    .B(_07207_),
    .Y(_07208_));
 AND2x2_ASAP7_75t_R _19251_ (.A(_07202_),
    .B(_07208_),
    .Y(_04402_));
 OR5x2_ASAP7_75t_R _19252_ (.A(_00660_),
    .B(_00661_),
    .C(_00662_),
    .D(_00663_),
    .E(_07152_),
    .Y(_07209_));
 OR3x1_ASAP7_75t_R _19253_ (.A(_00659_),
    .B(_07195_),
    .C(_07209_),
    .Y(_07210_));
 OAI21x1_ASAP7_75t_R _19254_ (.A1(_07195_),
    .A2(_07209_),
    .B(_00659_),
    .Y(_07211_));
 AND3x1_ASAP7_75t_R _19255_ (.A(_07182_),
    .B(_07210_),
    .C(_07211_),
    .Y(_04403_));
 OR3x1_ASAP7_75t_R _19256_ (.A(_00659_),
    .B(_07198_),
    .C(_07209_),
    .Y(_07212_));
 XOR2x2_ASAP7_75t_R _19257_ (.A(_00658_),
    .B(_07212_),
    .Y(_07213_));
 AND2x2_ASAP7_75t_R _19258_ (.A(_07202_),
    .B(_07213_),
    .Y(_04404_));
 XOR2x2_ASAP7_75t_R _19259_ (.A(_00657_),
    .B(_02661_),
    .Y(_07214_));
 AND2x2_ASAP7_75t_R _19260_ (.A(_07202_),
    .B(_07214_),
    .Y(_04405_));
 OR4x1_ASAP7_75t_R _19261_ (.A(_00658_),
    .B(_00659_),
    .C(_07195_),
    .D(_07209_),
    .Y(_07215_));
 XOR2x2_ASAP7_75t_R _19262_ (.A(_00656_),
    .B(_07215_),
    .Y(_07216_));
 AND2x2_ASAP7_75t_R _19263_ (.A(_07202_),
    .B(_07216_),
    .Y(_04406_));
 OR5x1_ASAP7_75t_R _19264_ (.A(_00656_),
    .B(_00658_),
    .C(_00659_),
    .D(_07198_),
    .E(_07209_),
    .Y(_07217_));
 XOR2x2_ASAP7_75t_R _19265_ (.A(_00655_),
    .B(_07217_),
    .Y(_07218_));
 AND2x2_ASAP7_75t_R _19266_ (.A(_07202_),
    .B(_07218_),
    .Y(_04407_));
 OR3x1_ASAP7_75t_R _19267_ (.A(_00657_),
    .B(_00668_),
    .C(_00051_),
    .Y(_07219_));
 XOR2x2_ASAP7_75t_R _19268_ (.A(_00654_),
    .B(_07219_),
    .Y(_07220_));
 AND2x2_ASAP7_75t_R _19269_ (.A(_07202_),
    .B(_07220_),
    .Y(_04408_));
 OR3x1_ASAP7_75t_R _19270_ (.A(_00654_),
    .B(_00657_),
    .C(_02661_),
    .Y(_07221_));
 NAND2x1_ASAP7_75t_R _19271_ (.A(_00653_),
    .B(_07221_),
    .Y(_07222_));
 AND3x1_ASAP7_75t_R _19272_ (.A(_07182_),
    .B(_07160_),
    .C(_07222_),
    .Y(_04409_));
 XOR2x2_ASAP7_75t_R _19273_ (.A(_00652_),
    .B(_07165_),
    .Y(_07223_));
 AND2x2_ASAP7_75t_R _19274_ (.A(_07202_),
    .B(_07223_),
    .Y(_04410_));
 OR3x1_ASAP7_75t_R _19275_ (.A(_00651_),
    .B(_00652_),
    .C(_07160_),
    .Y(_07224_));
 OAI21x1_ASAP7_75t_R _19276_ (.A1(_00652_),
    .A2(_07160_),
    .B(_00651_),
    .Y(_07225_));
 AND3x1_ASAP7_75t_R _19277_ (.A(_07182_),
    .B(_07224_),
    .C(_07225_),
    .Y(_04411_));
 OR3x1_ASAP7_75t_R _19278_ (.A(_00651_),
    .B(_00652_),
    .C(_07165_),
    .Y(_07226_));
 XOR2x2_ASAP7_75t_R _19279_ (.A(_00650_),
    .B(_07226_),
    .Y(_07227_));
 AND2x2_ASAP7_75t_R _19280_ (.A(_07202_),
    .B(_07227_),
    .Y(_04412_));
 OR4x1_ASAP7_75t_R _19281_ (.A(_00650_),
    .B(_00651_),
    .C(_00652_),
    .D(_07160_),
    .Y(_07228_));
 NAND2x1_ASAP7_75t_R _19282_ (.A(_00649_),
    .B(_07228_),
    .Y(_07229_));
 AND3x1_ASAP7_75t_R _19283_ (.A(_07182_),
    .B(_07162_),
    .C(_07229_),
    .Y(_04413_));
 BUFx6f_ASAP7_75t_R _19284_ (.A(_07084_),
    .Y(_07230_));
 XOR2x2_ASAP7_75t_R _19285_ (.A(_07148_),
    .B(_07166_),
    .Y(_07231_));
 AND2x2_ASAP7_75t_R _19286_ (.A(_07230_),
    .B(_07231_),
    .Y(_04414_));
 BUFx3_ASAP7_75t_R _19287_ (.A(_00630_),
    .Y(_07232_));
 BUFx3_ASAP7_75t_R _19288_ (.A(_00634_),
    .Y(_07233_));
 BUFx6f_ASAP7_75t_R _19289_ (.A(_00609_),
    .Y(_07234_));
 AND4x1_ASAP7_75t_R _19290_ (.A(_07234_),
    .B(_00637_),
    .C(_00638_),
    .D(_00639_),
    .Y(_07235_));
 AND5x1_ASAP7_75t_R _19291_ (.A(_00628_),
    .B(_00633_),
    .C(_07233_),
    .D(_00636_),
    .E(_07235_),
    .Y(_07236_));
 AND5x1_ASAP7_75t_R _19292_ (.A(_07232_),
    .B(_00631_),
    .C(_00632_),
    .D(_07147_),
    .E(_07236_),
    .Y(_07237_));
 BUFx3_ASAP7_75t_R _19293_ (.A(_00625_),
    .Y(_07238_));
 AND4x1_ASAP7_75t_R _19294_ (.A(_00623_),
    .B(_00624_),
    .C(_07238_),
    .D(_00626_),
    .Y(_07239_));
 AND4x1_ASAP7_75t_R _19295_ (.A(_00617_),
    .B(_00619_),
    .C(_00620_),
    .D(_00627_),
    .Y(_07240_));
 AND5x1_ASAP7_75t_R _19296_ (.A(_00610_),
    .B(_00611_),
    .C(_00616_),
    .D(_00635_),
    .E(_07240_),
    .Y(_07241_));
 AND3x1_ASAP7_75t_R _19297_ (.A(_00614_),
    .B(_00615_),
    .C(_00618_),
    .Y(_07242_));
 OR3x1_ASAP7_75t_R _19298_ (.A(_00612_),
    .B(_00613_),
    .C(_07242_),
    .Y(_07243_));
 AND5x2_ASAP7_75t_R _19299_ (.A(_00621_),
    .B(_00622_),
    .C(_07239_),
    .D(_07241_),
    .E(_07243_),
    .Y(_07244_));
 NAND2x2_ASAP7_75t_R _19300_ (.A(_07237_),
    .B(_07244_),
    .Y(_07245_));
 NOR2x1_ASAP7_75t_R _19301_ (.A(_00599_),
    .B(_07245_),
    .Y(_04415_));
 INVx1_ASAP7_75t_R _19302_ (.A(_07245_),
    .Y(_04416_));
 NOR2x1_ASAP7_75t_R _19303_ (.A(_00602_),
    .B(_07245_),
    .Y(_04417_));
 NOR2x1_ASAP7_75t_R _19304_ (.A(_00601_),
    .B(_07245_),
    .Y(_04418_));
 NOR2x1_ASAP7_75t_R _19305_ (.A(_00600_),
    .B(_07245_),
    .Y(_04419_));
 NOR2x1_ASAP7_75t_R _19306_ (.A(_00598_),
    .B(_07245_),
    .Y(_04420_));
 NOR2x1_ASAP7_75t_R _19307_ (.A(_00597_),
    .B(_07245_),
    .Y(_04421_));
 INVx1_ASAP7_75t_R _19308_ (.A(_07245_),
    .Y(_04422_));
 AND2x2_ASAP7_75t_R _19309_ (.A(_07230_),
    .B(_00052_),
    .Y(_04423_));
 OR4x1_ASAP7_75t_R _19310_ (.A(_00614_),
    .B(_00615_),
    .C(_00618_),
    .D(_02641_),
    .Y(_07246_));
 OR4x1_ASAP7_75t_R _19311_ (.A(_00610_),
    .B(_00611_),
    .C(_00612_),
    .D(_00613_),
    .Y(_07247_));
 OR2x6_ASAP7_75t_R _19312_ (.A(_07246_),
    .B(_07247_),
    .Y(_07248_));
 OR3x1_ASAP7_75t_R _19313_ (.A(_07234_),
    .B(_00639_),
    .C(_07248_),
    .Y(_07249_));
 OAI21x1_ASAP7_75t_R _19314_ (.A1(_07234_),
    .A2(_07248_),
    .B(_00639_),
    .Y(_07250_));
 AND3x1_ASAP7_75t_R _19315_ (.A(_07182_),
    .B(_07249_),
    .C(_07250_),
    .Y(_04424_));
 OR5x2_ASAP7_75t_R _19316_ (.A(_00614_),
    .B(_00615_),
    .C(_00618_),
    .D(_00629_),
    .E(_00052_),
    .Y(_07251_));
 OR2x6_ASAP7_75t_R _19317_ (.A(_07247_),
    .B(_07251_),
    .Y(_07252_));
 OR3x1_ASAP7_75t_R _19318_ (.A(_07234_),
    .B(_00639_),
    .C(_07252_),
    .Y(_07253_));
 XOR2x2_ASAP7_75t_R _19319_ (.A(_00638_),
    .B(_07253_),
    .Y(_07254_));
 AND2x2_ASAP7_75t_R _19320_ (.A(_07230_),
    .B(_07254_),
    .Y(_04425_));
 OR4x1_ASAP7_75t_R _19321_ (.A(_07234_),
    .B(_00638_),
    .C(_00639_),
    .D(_07248_),
    .Y(_07255_));
 XOR2x2_ASAP7_75t_R _19322_ (.A(_00637_),
    .B(_07255_),
    .Y(_07256_));
 AND2x2_ASAP7_75t_R _19323_ (.A(_07230_),
    .B(_07256_),
    .Y(_04426_));
 OR5x2_ASAP7_75t_R _19324_ (.A(_07234_),
    .B(_00636_),
    .C(_00637_),
    .D(_00638_),
    .E(_00639_),
    .Y(_07257_));
 OR5x1_ASAP7_75t_R _19325_ (.A(_07234_),
    .B(_00637_),
    .C(_00638_),
    .D(_00639_),
    .E(_07252_),
    .Y(_07258_));
 NAND2x1_ASAP7_75t_R _19326_ (.A(_00636_),
    .B(_07258_),
    .Y(_07259_));
 BUFx12f_ASAP7_75t_R _19327_ (.A(_08876_),
    .Y(_07260_));
 OA211x2_ASAP7_75t_R _19328_ (.A1(_07252_),
    .A2(_07257_),
    .B(_07259_),
    .C(_07260_),
    .Y(_04427_));
 BUFx6f_ASAP7_75t_R _19329_ (.A(_06386_),
    .Y(_07261_));
 OR4x1_ASAP7_75t_R _19330_ (.A(_00635_),
    .B(_07246_),
    .C(_07247_),
    .D(_07257_),
    .Y(_07262_));
 OAI21x1_ASAP7_75t_R _19331_ (.A1(_07248_),
    .A2(_07257_),
    .B(_00635_),
    .Y(_07263_));
 AND3x1_ASAP7_75t_R _19332_ (.A(_07261_),
    .B(_07262_),
    .C(_07263_),
    .Y(_04428_));
 OR4x1_ASAP7_75t_R _19333_ (.A(_00635_),
    .B(_07247_),
    .C(_07251_),
    .D(_07257_),
    .Y(_07264_));
 XOR2x2_ASAP7_75t_R _19334_ (.A(_07233_),
    .B(_07264_),
    .Y(_07265_));
 AND2x2_ASAP7_75t_R _19335_ (.A(_07230_),
    .B(_07265_),
    .Y(_04429_));
 OR3x1_ASAP7_75t_R _19336_ (.A(_00633_),
    .B(_07233_),
    .C(_07262_),
    .Y(_07266_));
 OAI21x1_ASAP7_75t_R _19337_ (.A1(_07233_),
    .A2(_07262_),
    .B(_00633_),
    .Y(_07267_));
 AND3x1_ASAP7_75t_R _19338_ (.A(_07261_),
    .B(_07266_),
    .C(_07267_),
    .Y(_04430_));
 OR3x1_ASAP7_75t_R _19339_ (.A(_00633_),
    .B(_07233_),
    .C(_07264_),
    .Y(_07268_));
 XOR2x2_ASAP7_75t_R _19340_ (.A(_00632_),
    .B(_07268_),
    .Y(_07269_));
 AND2x2_ASAP7_75t_R _19341_ (.A(_07230_),
    .B(_07269_),
    .Y(_04431_));
 OR5x2_ASAP7_75t_R _19342_ (.A(_00631_),
    .B(_00632_),
    .C(_00633_),
    .D(_07233_),
    .E(_07262_),
    .Y(_07270_));
 OR4x1_ASAP7_75t_R _19343_ (.A(_00632_),
    .B(_00633_),
    .C(_07233_),
    .D(_07262_),
    .Y(_07271_));
 NAND2x1_ASAP7_75t_R _19344_ (.A(_00631_),
    .B(_07271_),
    .Y(_07272_));
 AND3x1_ASAP7_75t_R _19345_ (.A(_07261_),
    .B(_07270_),
    .C(_07272_),
    .Y(_04432_));
 OR5x2_ASAP7_75t_R _19346_ (.A(_00631_),
    .B(_00632_),
    .C(_00633_),
    .D(_07233_),
    .E(_07264_),
    .Y(_07273_));
 XOR2x2_ASAP7_75t_R _19347_ (.A(_07232_),
    .B(_07273_),
    .Y(_07274_));
 AND2x2_ASAP7_75t_R _19348_ (.A(_07230_),
    .B(_07274_),
    .Y(_04433_));
 NOR2x1_ASAP7_75t_R _19349_ (.A(_07190_),
    .B(_02642_),
    .Y(_04434_));
 OR3x1_ASAP7_75t_R _19350_ (.A(_00628_),
    .B(_07232_),
    .C(_07270_),
    .Y(_07275_));
 OAI21x1_ASAP7_75t_R _19351_ (.A1(_07232_),
    .A2(_07270_),
    .B(_00628_),
    .Y(_07276_));
 AND3x1_ASAP7_75t_R _19352_ (.A(_07261_),
    .B(_07275_),
    .C(_07276_),
    .Y(_04435_));
 OR3x1_ASAP7_75t_R _19353_ (.A(_00628_),
    .B(_07232_),
    .C(_07273_),
    .Y(_07277_));
 XOR2x2_ASAP7_75t_R _19354_ (.A(_00627_),
    .B(_07277_),
    .Y(_07278_));
 AND2x2_ASAP7_75t_R _19355_ (.A(_07230_),
    .B(_07278_),
    .Y(_04436_));
 OR5x1_ASAP7_75t_R _19356_ (.A(_00626_),
    .B(_00627_),
    .C(_00628_),
    .D(_07232_),
    .E(_07270_),
    .Y(_07279_));
 BUFx3_ASAP7_75t_R _19357_ (.A(_07279_),
    .Y(_07280_));
 OR4x1_ASAP7_75t_R _19358_ (.A(_00627_),
    .B(_00628_),
    .C(_07232_),
    .D(_07270_),
    .Y(_07281_));
 NAND2x1_ASAP7_75t_R _19359_ (.A(_00626_),
    .B(_07281_),
    .Y(_07282_));
 AND3x1_ASAP7_75t_R _19360_ (.A(_07261_),
    .B(_07280_),
    .C(_07282_),
    .Y(_04437_));
 OR5x2_ASAP7_75t_R _19361_ (.A(_00626_),
    .B(_00627_),
    .C(_00628_),
    .D(_07232_),
    .E(_07273_),
    .Y(_07283_));
 XOR2x2_ASAP7_75t_R _19362_ (.A(_07238_),
    .B(_07283_),
    .Y(_07284_));
 AND2x2_ASAP7_75t_R _19363_ (.A(_07230_),
    .B(_07284_),
    .Y(_04438_));
 OR3x1_ASAP7_75t_R _19364_ (.A(_00624_),
    .B(_07238_),
    .C(_07280_),
    .Y(_07285_));
 OAI21x1_ASAP7_75t_R _19365_ (.A1(_07238_),
    .A2(_07280_),
    .B(_00624_),
    .Y(_07286_));
 AND3x1_ASAP7_75t_R _19366_ (.A(_07261_),
    .B(_07285_),
    .C(_07286_),
    .Y(_04439_));
 OR3x1_ASAP7_75t_R _19367_ (.A(_00624_),
    .B(_07238_),
    .C(_07283_),
    .Y(_07287_));
 XOR2x2_ASAP7_75t_R _19368_ (.A(_00623_),
    .B(_07287_),
    .Y(_07288_));
 AND2x2_ASAP7_75t_R _19369_ (.A(_07230_),
    .B(_07288_),
    .Y(_04440_));
 BUFx6f_ASAP7_75t_R _19370_ (.A(_07084_),
    .Y(_07289_));
 OR4x1_ASAP7_75t_R _19371_ (.A(_00623_),
    .B(_00624_),
    .C(_07238_),
    .D(_07280_),
    .Y(_07290_));
 XOR2x2_ASAP7_75t_R _19372_ (.A(_00622_),
    .B(_07290_),
    .Y(_07291_));
 AND2x2_ASAP7_75t_R _19373_ (.A(_07289_),
    .B(_07291_),
    .Y(_04441_));
 OR5x1_ASAP7_75t_R _19374_ (.A(_00622_),
    .B(_00623_),
    .C(_00624_),
    .D(_07238_),
    .E(_07283_),
    .Y(_07292_));
 XOR2x2_ASAP7_75t_R _19375_ (.A(_00621_),
    .B(_07292_),
    .Y(_07293_));
 AND2x2_ASAP7_75t_R _19376_ (.A(_07289_),
    .B(_07293_),
    .Y(_04442_));
 OR5x2_ASAP7_75t_R _19377_ (.A(_00621_),
    .B(_00622_),
    .C(_00623_),
    .D(_00624_),
    .E(_07238_),
    .Y(_07294_));
 OR3x1_ASAP7_75t_R _19378_ (.A(_00620_),
    .B(_07280_),
    .C(_07294_),
    .Y(_07295_));
 OAI21x1_ASAP7_75t_R _19379_ (.A1(_07280_),
    .A2(_07294_),
    .B(_00620_),
    .Y(_07296_));
 AND3x1_ASAP7_75t_R _19380_ (.A(_07261_),
    .B(_07295_),
    .C(_07296_),
    .Y(_04443_));
 OR3x1_ASAP7_75t_R _19381_ (.A(_00620_),
    .B(_07283_),
    .C(_07294_),
    .Y(_07297_));
 XOR2x2_ASAP7_75t_R _19382_ (.A(_00619_),
    .B(_07297_),
    .Y(_07298_));
 AND2x2_ASAP7_75t_R _19383_ (.A(_07289_),
    .B(_07298_),
    .Y(_04444_));
 XOR2x2_ASAP7_75t_R _19384_ (.A(_00618_),
    .B(_02641_),
    .Y(_07299_));
 AND2x2_ASAP7_75t_R _19385_ (.A(_07289_),
    .B(_07299_),
    .Y(_04445_));
 OR4x1_ASAP7_75t_R _19386_ (.A(_00619_),
    .B(_00620_),
    .C(_07280_),
    .D(_07294_),
    .Y(_07300_));
 XOR2x2_ASAP7_75t_R _19387_ (.A(_00617_),
    .B(_07300_),
    .Y(_07301_));
 AND2x2_ASAP7_75t_R _19388_ (.A(_07289_),
    .B(_07301_),
    .Y(_04446_));
 OR5x1_ASAP7_75t_R _19389_ (.A(_00617_),
    .B(_00619_),
    .C(_00620_),
    .D(_07283_),
    .E(_07294_),
    .Y(_07302_));
 XOR2x2_ASAP7_75t_R _19390_ (.A(_00616_),
    .B(_07302_),
    .Y(_07303_));
 AND2x2_ASAP7_75t_R _19391_ (.A(_07289_),
    .B(_07303_),
    .Y(_04447_));
 OR3x1_ASAP7_75t_R _19392_ (.A(_00618_),
    .B(_00629_),
    .C(_00052_),
    .Y(_07304_));
 XOR2x2_ASAP7_75t_R _19393_ (.A(_00615_),
    .B(_07304_),
    .Y(_07305_));
 AND2x2_ASAP7_75t_R _19394_ (.A(_07289_),
    .B(_07305_),
    .Y(_04448_));
 OR3x1_ASAP7_75t_R _19395_ (.A(_00615_),
    .B(_00618_),
    .C(_02641_),
    .Y(_07306_));
 NAND2x1_ASAP7_75t_R _19396_ (.A(_00614_),
    .B(_07306_),
    .Y(_07307_));
 AND3x1_ASAP7_75t_R _19397_ (.A(_07261_),
    .B(_07246_),
    .C(_07307_),
    .Y(_04449_));
 XOR2x2_ASAP7_75t_R _19398_ (.A(_00613_),
    .B(_07251_),
    .Y(_07308_));
 AND2x2_ASAP7_75t_R _19399_ (.A(_07289_),
    .B(_07308_),
    .Y(_04450_));
 OR3x1_ASAP7_75t_R _19400_ (.A(_00612_),
    .B(_00613_),
    .C(_07246_),
    .Y(_07309_));
 OAI21x1_ASAP7_75t_R _19401_ (.A1(_00613_),
    .A2(_07246_),
    .B(_00612_),
    .Y(_07310_));
 AND3x1_ASAP7_75t_R _19402_ (.A(_07261_),
    .B(_07309_),
    .C(_07310_),
    .Y(_04451_));
 OR3x1_ASAP7_75t_R _19403_ (.A(_00612_),
    .B(_00613_),
    .C(_07251_),
    .Y(_07311_));
 XOR2x2_ASAP7_75t_R _19404_ (.A(_00611_),
    .B(_07311_),
    .Y(_07312_));
 AND2x2_ASAP7_75t_R _19405_ (.A(_07289_),
    .B(_07312_),
    .Y(_04452_));
 OR4x1_ASAP7_75t_R _19406_ (.A(_00611_),
    .B(_00612_),
    .C(_00613_),
    .D(_07246_),
    .Y(_07313_));
 NAND2x1_ASAP7_75t_R _19407_ (.A(_00610_),
    .B(_07313_),
    .Y(_07314_));
 AND3x1_ASAP7_75t_R _19408_ (.A(_07261_),
    .B(_07248_),
    .C(_07314_),
    .Y(_04453_));
 XOR2x2_ASAP7_75t_R _19409_ (.A(_07234_),
    .B(_07252_),
    .Y(_07315_));
 AND2x2_ASAP7_75t_R _19410_ (.A(_07289_),
    .B(_07315_),
    .Y(_04454_));
 BUFx6f_ASAP7_75t_R _19411_ (.A(_07084_),
    .Y(_07316_));
 AND2x2_ASAP7_75t_R _19412_ (.A(_07316_),
    .B(_00025_),
    .Y(_04455_));
 NAND2x1_ASAP7_75t_R _19413_ (.A(_00643_),
    .B(_00644_),
    .Y(_07317_));
 OR5x1_ASAP7_75t_R _19414_ (.A(_00640_),
    .B(\xs[4].cli1.i[36] ),
    .C(_00642_),
    .D(\xs[4].cli1.i[32] ),
    .E(_07317_),
    .Y(_07318_));
 BUFx3_ASAP7_75t_R _19415_ (.A(_07318_),
    .Y(_07319_));
 AND2x2_ASAP7_75t_R _19416_ (.A(_00643_),
    .B(_00644_),
    .Y(_07320_));
 AO31x2_ASAP7_75t_R _19417_ (.A1(_00641_),
    .A2(\xs[4].cli1.i[35] ),
    .A3(_07320_),
    .B(_00640_),
    .Y(_07321_));
 INVx2_ASAP7_75t_R _19418_ (.A(_02253_),
    .Y(_07322_));
 AOI21x1_ASAP7_75t_R _19419_ (.A1(_07319_),
    .A2(_07321_),
    .B(_07322_),
    .Y(_07323_));
 BUFx3_ASAP7_75t_R _19420_ (.A(_02247_),
    .Y(_07324_));
 INVx3_ASAP7_75t_R _19421_ (.A(_02246_),
    .Y(_07325_));
 OAI21x1_ASAP7_75t_R _19422_ (.A1(_07324_),
    .A2(_07319_),
    .B(_07325_),
    .Y(_07326_));
 OA31x2_ASAP7_75t_R _19423_ (.A1(\xs[4].cli1.i[36] ),
    .A2(_00642_),
    .A3(_07317_),
    .B1(\xs[4].cli1.i[39] ),
    .Y(_07327_));
 AO21x1_ASAP7_75t_R _19424_ (.A1(_00025_),
    .A2(_07327_),
    .B(_07325_),
    .Y(_07328_));
 NAND2x1_ASAP7_75t_R _19425_ (.A(_00682_),
    .B(_00683_),
    .Y(_07329_));
 OA31x2_ASAP7_75t_R _19426_ (.A1(\peo[8][36] ),
    .A2(_00681_),
    .A3(_07329_),
    .B1(\peo[8][39] ),
    .Y(_07330_));
 OA211x2_ASAP7_75t_R _19427_ (.A1(_07323_),
    .A2(_07326_),
    .B(_07328_),
    .C(_07330_),
    .Y(_07331_));
 OAI21x1_ASAP7_75t_R _19428_ (.A1(_07319_),
    .A2(_07331_),
    .B(_00686_),
    .Y(_07332_));
 INVx1_ASAP7_75t_R _19429_ (.A(_07324_),
    .Y(_07333_));
 AND3x1_ASAP7_75t_R _19430_ (.A(_07325_),
    .B(_07333_),
    .C(_07327_),
    .Y(_07334_));
 OR4x1_ASAP7_75t_R _19431_ (.A(\peo[9][0] ),
    .B(_07319_),
    .C(_07331_),
    .D(_07334_),
    .Y(_07335_));
 AND2x2_ASAP7_75t_R _19432_ (.A(_00682_),
    .B(_00683_),
    .Y(_07336_));
 AO31x2_ASAP7_75t_R _19433_ (.A1(_00680_),
    .A2(\peo[8][35] ),
    .A3(_07336_),
    .B(_00679_),
    .Y(_07337_));
 AO21x1_ASAP7_75t_R _19434_ (.A1(\peo[8][39] ),
    .A2(\peo[8][32] ),
    .B(_02253_),
    .Y(_07338_));
 AND2x2_ASAP7_75t_R _19435_ (.A(_07337_),
    .B(_07338_),
    .Y(_07339_));
 OAI21x1_ASAP7_75t_R _19436_ (.A1(_02253_),
    .A2(_07327_),
    .B(_07319_),
    .Y(_07340_));
 NAND2x1_ASAP7_75t_R _19437_ (.A(_07325_),
    .B(_07324_),
    .Y(_07341_));
 AO21x2_ASAP7_75t_R _19438_ (.A1(_07339_),
    .A2(_07340_),
    .B(_07341_),
    .Y(_07342_));
 NOR2x1_ASAP7_75t_R _19439_ (.A(_07322_),
    .B(_07342_),
    .Y(_07343_));
 NOR2x1_ASAP7_75t_R _19440_ (.A(_09314_),
    .B(_07343_),
    .Y(_07344_));
 NOR2x1_ASAP7_75t_R _19441_ (.A(_06206_),
    .B(_02257_),
    .Y(_07345_));
 AO32x1_ASAP7_75t_R _19442_ (.A1(_07332_),
    .A2(_07335_),
    .A3(_07344_),
    .B1(_07345_),
    .B2(_07343_),
    .Y(_04456_));
 OR3x2_ASAP7_75t_R _19443_ (.A(_10763_),
    .B(_07322_),
    .C(_07342_),
    .Y(_07346_));
 NOR2x1_ASAP7_75t_R _19444_ (.A(_02256_),
    .B(_07346_),
    .Y(_04457_));
 NOR2x1_ASAP7_75t_R _19445_ (.A(_02255_),
    .B(_07346_),
    .Y(_04458_));
 NOR2x1_ASAP7_75t_R _19446_ (.A(_02254_),
    .B(_07346_),
    .Y(_04459_));
 NOR2x1_ASAP7_75t_R _19447_ (.A(_02245_),
    .B(_07346_),
    .Y(_04460_));
 NOR2x1_ASAP7_75t_R _19448_ (.A(_02244_),
    .B(_07346_),
    .Y(_04461_));
 NOR2x1_ASAP7_75t_R _19449_ (.A(_07331_),
    .B(_07334_),
    .Y(_07347_));
 OR3x1_ASAP7_75t_R _19450_ (.A(_09207_),
    .B(_00647_),
    .C(_07347_),
    .Y(_07348_));
 NAND2x1_ASAP7_75t_R _19451_ (.A(_07339_),
    .B(_07340_),
    .Y(_07349_));
 AND5x1_ASAP7_75t_R _19452_ (.A(_07325_),
    .B(_07324_),
    .C(_07322_),
    .D(_02257_),
    .E(_07349_),
    .Y(_07350_));
 OA21x2_ASAP7_75t_R _19453_ (.A1(_02253_),
    .A2(_07342_),
    .B(_00686_),
    .Y(_07351_));
 OR5x1_ASAP7_75t_R _19454_ (.A(_10826_),
    .B(_07331_),
    .C(_07334_),
    .D(_07350_),
    .E(_07351_),
    .Y(_07352_));
 NAND2x1_ASAP7_75t_R _19455_ (.A(_07348_),
    .B(_07352_),
    .Y(_04462_));
 OR3x2_ASAP7_75t_R _19456_ (.A(_11177_),
    .B(_02253_),
    .C(_07342_),
    .Y(_07353_));
 NOR2x1_ASAP7_75t_R _19457_ (.A(_02256_),
    .B(_07353_),
    .Y(_04463_));
 NOR2x1_ASAP7_75t_R _19458_ (.A(_02255_),
    .B(_07353_),
    .Y(_04464_));
 NOR2x1_ASAP7_75t_R _19459_ (.A(_02254_),
    .B(_07353_),
    .Y(_04465_));
 NOR2x1_ASAP7_75t_R _19460_ (.A(_02245_),
    .B(_07353_),
    .Y(_04466_));
 NOR2x1_ASAP7_75t_R _19461_ (.A(_02244_),
    .B(_07353_),
    .Y(_04467_));
 AO21x1_ASAP7_75t_R _19462_ (.A1(_07324_),
    .A2(_07349_),
    .B(_02246_),
    .Y(_07354_));
 BUFx6f_ASAP7_75t_R _19463_ (.A(_07354_),
    .Y(_07355_));
 NOR2x1_ASAP7_75t_R _19464_ (.A(_02257_),
    .B(_07355_),
    .Y(_07356_));
 AND2x2_ASAP7_75t_R _19465_ (.A(_07325_),
    .B(_07330_),
    .Y(_07357_));
 AND2x2_ASAP7_75t_R _19466_ (.A(_02246_),
    .B(_00025_),
    .Y(_07358_));
 AO221x1_ASAP7_75t_R _19467_ (.A1(_07325_),
    .A2(_07333_),
    .B1(_07330_),
    .B2(_07358_),
    .C(_07321_),
    .Y(_07359_));
 AOI21x1_ASAP7_75t_R _19468_ (.A1(_07323_),
    .A2(_07357_),
    .B(_07359_),
    .Y(_07360_));
 NAND2x1_ASAP7_75t_R _19469_ (.A(_00647_),
    .B(_07360_),
    .Y(_07361_));
 OA211x2_ASAP7_75t_R _19470_ (.A1(\peo[8][0] ),
    .A2(_07360_),
    .B(_07361_),
    .C(_07355_),
    .Y(_07362_));
 OA21x2_ASAP7_75t_R _19471_ (.A1(_07356_),
    .A2(_07362_),
    .B(_06676_),
    .Y(_04468_));
 AOI21x1_ASAP7_75t_R _19472_ (.A1(_07324_),
    .A2(_07349_),
    .B(_02246_),
    .Y(_07363_));
 NAND2x2_ASAP7_75t_R _19473_ (.A(_08581_),
    .B(_07363_),
    .Y(_07364_));
 NOR2x1_ASAP7_75t_R _19474_ (.A(_02256_),
    .B(_07364_),
    .Y(_04469_));
 NOR2x1_ASAP7_75t_R _19475_ (.A(_02255_),
    .B(_07364_),
    .Y(_04470_));
 NOR2x1_ASAP7_75t_R _19476_ (.A(_02254_),
    .B(_07364_),
    .Y(_04471_));
 AND2x2_ASAP7_75t_R _19477_ (.A(_07322_),
    .B(_07363_),
    .Y(_07365_));
 NAND2x1_ASAP7_75t_R _19478_ (.A(_00645_),
    .B(_07360_),
    .Y(_07366_));
 OA211x2_ASAP7_75t_R _19479_ (.A1(\peo[8][32] ),
    .A2(_07360_),
    .B(_07366_),
    .C(_07355_),
    .Y(_07367_));
 OA21x2_ASAP7_75t_R _19480_ (.A1(_07365_),
    .A2(_07367_),
    .B(_06676_),
    .Y(_04472_));
 NOR2x1_ASAP7_75t_R _19481_ (.A(_02252_),
    .B(_07355_),
    .Y(_07368_));
 NAND2x1_ASAP7_75t_R _19482_ (.A(_00644_),
    .B(_07360_),
    .Y(_07369_));
 OA211x2_ASAP7_75t_R _19483_ (.A1(\peo[8][33] ),
    .A2(_07360_),
    .B(_07369_),
    .C(_07355_),
    .Y(_07370_));
 OA21x2_ASAP7_75t_R _19484_ (.A1(_07368_),
    .A2(_07370_),
    .B(_08529_),
    .Y(_04473_));
 NOR2x1_ASAP7_75t_R _19485_ (.A(_02251_),
    .B(_07355_),
    .Y(_07371_));
 NAND2x1_ASAP7_75t_R _19486_ (.A(_00643_),
    .B(_07360_),
    .Y(_07372_));
 OA211x2_ASAP7_75t_R _19487_ (.A1(\peo[8][34] ),
    .A2(_07360_),
    .B(_07372_),
    .C(_07355_),
    .Y(_07373_));
 OA21x2_ASAP7_75t_R _19488_ (.A1(_07371_),
    .A2(_07373_),
    .B(_08529_),
    .Y(_04474_));
 INVx1_ASAP7_75t_R _19489_ (.A(_07331_),
    .Y(_07374_));
 OR2x2_ASAP7_75t_R _19490_ (.A(_07321_),
    .B(_07331_),
    .Y(_07375_));
 AO32x1_ASAP7_75t_R _19491_ (.A1(\xs[4].cli1.i[39] ),
    .A2(_00642_),
    .A3(_07374_),
    .B1(_07375_),
    .B2(_00681_),
    .Y(_07376_));
 NAND2x1_ASAP7_75t_R _19492_ (.A(_08599_),
    .B(_07355_),
    .Y(_07377_));
 OAI22x1_ASAP7_75t_R _19493_ (.A1(_02250_),
    .A2(_07364_),
    .B1(_07376_),
    .B2(_07377_),
    .Y(_04475_));
 NOR2x1_ASAP7_75t_R _19494_ (.A(_02249_),
    .B(_07355_),
    .Y(_07378_));
 NAND2x1_ASAP7_75t_R _19495_ (.A(_00641_),
    .B(_07360_),
    .Y(_07379_));
 OA211x2_ASAP7_75t_R _19496_ (.A1(\peo[8][36] ),
    .A2(_07360_),
    .B(_07379_),
    .C(_07354_),
    .Y(_07380_));
 OA21x2_ASAP7_75t_R _19497_ (.A1(_07378_),
    .A2(_07380_),
    .B(_08529_),
    .Y(_04476_));
 NOR2x1_ASAP7_75t_R _19498_ (.A(_02248_),
    .B(_07364_),
    .Y(_04477_));
 OR3x1_ASAP7_75t_R _19499_ (.A(_08642_),
    .B(_07349_),
    .C(_07341_),
    .Y(_07381_));
 INVx1_ASAP7_75t_R _19500_ (.A(_07381_),
    .Y(_04478_));
 AND3x1_ASAP7_75t_R _19501_ (.A(_07337_),
    .B(_07321_),
    .C(_07355_),
    .Y(_07382_));
 NOR2x1_ASAP7_75t_R _19502_ (.A(_07190_),
    .B(_07382_),
    .Y(_04479_));
 NOR2x1_ASAP7_75t_R _19503_ (.A(_02245_),
    .B(_07364_),
    .Y(_04480_));
 NOR2x1_ASAP7_75t_R _19504_ (.A(_02244_),
    .B(_07364_),
    .Y(_04481_));
 BUFx6f_ASAP7_75t_R _19505_ (.A(_00567_),
    .Y(_07383_));
 AND4x1_ASAP7_75t_R _19506_ (.A(_00544_),
    .B(_00572_),
    .C(_00573_),
    .D(_00574_),
    .Y(_07384_));
 AND5x1_ASAP7_75t_R _19507_ (.A(_00563_),
    .B(_00568_),
    .C(_00569_),
    .D(_00571_),
    .E(_07384_),
    .Y(_07385_));
 AND5x1_ASAP7_75t_R _19508_ (.A(_00565_),
    .B(_00566_),
    .C(_07383_),
    .D(_07147_),
    .E(_07385_),
    .Y(_07386_));
 BUFx3_ASAP7_75t_R _19509_ (.A(_00560_),
    .Y(_07387_));
 AND4x1_ASAP7_75t_R _19510_ (.A(_00558_),
    .B(_00559_),
    .C(_07387_),
    .D(_00561_),
    .Y(_07388_));
 AND4x1_ASAP7_75t_R _19511_ (.A(_00552_),
    .B(_00554_),
    .C(_00555_),
    .D(_00562_),
    .Y(_07389_));
 AND5x1_ASAP7_75t_R _19512_ (.A(_00545_),
    .B(_00546_),
    .C(_00551_),
    .D(_00570_),
    .E(_07389_),
    .Y(_07390_));
 AND3x1_ASAP7_75t_R _19513_ (.A(_00549_),
    .B(_00550_),
    .C(_00553_),
    .Y(_07391_));
 OR3x1_ASAP7_75t_R _19514_ (.A(_00547_),
    .B(_00548_),
    .C(_07391_),
    .Y(_07392_));
 AND5x2_ASAP7_75t_R _19515_ (.A(_00556_),
    .B(_00557_),
    .C(_07388_),
    .D(_07390_),
    .E(_07392_),
    .Y(_07393_));
 NAND2x2_ASAP7_75t_R _19516_ (.A(_07386_),
    .B(_07393_),
    .Y(_07394_));
 NOR2x1_ASAP7_75t_R _19517_ (.A(_00501_),
    .B(_07394_),
    .Y(_04482_));
 INVx1_ASAP7_75t_R _19518_ (.A(_07394_),
    .Y(_04483_));
 NOR2x1_ASAP7_75t_R _19519_ (.A(_00504_),
    .B(_07394_),
    .Y(_04484_));
 NOR2x1_ASAP7_75t_R _19520_ (.A(_00503_),
    .B(_07394_),
    .Y(_04485_));
 NOR2x1_ASAP7_75t_R _19521_ (.A(_00502_),
    .B(_07394_),
    .Y(_04486_));
 NOR2x1_ASAP7_75t_R _19522_ (.A(_00500_),
    .B(_07394_),
    .Y(_04487_));
 NOR2x1_ASAP7_75t_R _19523_ (.A(_00499_),
    .B(_07394_),
    .Y(_04488_));
 INVx1_ASAP7_75t_R _19524_ (.A(_07394_),
    .Y(_04489_));
 AND2x2_ASAP7_75t_R _19525_ (.A(_07316_),
    .B(_00053_),
    .Y(_04490_));
 OR4x1_ASAP7_75t_R _19526_ (.A(_00549_),
    .B(_00550_),
    .C(_00553_),
    .D(_02649_),
    .Y(_07395_));
 OR4x1_ASAP7_75t_R _19527_ (.A(_00545_),
    .B(_00546_),
    .C(_00547_),
    .D(_00548_),
    .Y(_07396_));
 OR3x1_ASAP7_75t_R _19528_ (.A(_00544_),
    .B(_07395_),
    .C(_07396_),
    .Y(_07397_));
 XOR2x2_ASAP7_75t_R _19529_ (.A(_00574_),
    .B(_07397_),
    .Y(_07398_));
 AND2x2_ASAP7_75t_R _19530_ (.A(_07316_),
    .B(_07398_),
    .Y(_04491_));
 OR2x2_ASAP7_75t_R _19531_ (.A(_00544_),
    .B(_00574_),
    .Y(_07399_));
 OR5x2_ASAP7_75t_R _19532_ (.A(_00549_),
    .B(_00550_),
    .C(_00553_),
    .D(_00564_),
    .E(_00053_),
    .Y(_07400_));
 OR3x2_ASAP7_75t_R _19533_ (.A(_07396_),
    .B(_07399_),
    .C(_07400_),
    .Y(_07401_));
 XOR2x2_ASAP7_75t_R _19534_ (.A(_00573_),
    .B(_07401_),
    .Y(_07402_));
 AND2x2_ASAP7_75t_R _19535_ (.A(_07316_),
    .B(_07402_),
    .Y(_04492_));
 BUFx6f_ASAP7_75t_R _19536_ (.A(_06386_),
    .Y(_07403_));
 OR5x2_ASAP7_75t_R _19537_ (.A(_00572_),
    .B(_00573_),
    .C(_07395_),
    .D(_07396_),
    .E(_07399_),
    .Y(_07404_));
 OR3x1_ASAP7_75t_R _19538_ (.A(_00573_),
    .B(_00574_),
    .C(_07397_),
    .Y(_07405_));
 NAND2x1_ASAP7_75t_R _19539_ (.A(_00572_),
    .B(_07405_),
    .Y(_07406_));
 AND3x1_ASAP7_75t_R _19540_ (.A(_07403_),
    .B(_07404_),
    .C(_07406_),
    .Y(_04493_));
 OR3x1_ASAP7_75t_R _19541_ (.A(_00572_),
    .B(_00573_),
    .C(_07401_),
    .Y(_07407_));
 XOR2x2_ASAP7_75t_R _19542_ (.A(_00571_),
    .B(_07407_),
    .Y(_07408_));
 AND2x2_ASAP7_75t_R _19543_ (.A(_07316_),
    .B(_07408_),
    .Y(_04494_));
 OR3x1_ASAP7_75t_R _19544_ (.A(_00570_),
    .B(_00571_),
    .C(_07404_),
    .Y(_07409_));
 OAI21x1_ASAP7_75t_R _19545_ (.A1(_00571_),
    .A2(_07404_),
    .B(_00570_),
    .Y(_07410_));
 AND3x1_ASAP7_75t_R _19546_ (.A(_07403_),
    .B(_07409_),
    .C(_07410_),
    .Y(_04495_));
 OR3x1_ASAP7_75t_R _19547_ (.A(_00570_),
    .B(_00571_),
    .C(_07407_),
    .Y(_07411_));
 XOR2x2_ASAP7_75t_R _19548_ (.A(_00569_),
    .B(_07411_),
    .Y(_07412_));
 AND2x2_ASAP7_75t_R _19549_ (.A(_07316_),
    .B(_07412_),
    .Y(_04496_));
 OR4x1_ASAP7_75t_R _19550_ (.A(_00568_),
    .B(_00569_),
    .C(_00570_),
    .D(_00571_),
    .Y(_07413_));
 OR2x6_ASAP7_75t_R _19551_ (.A(_07404_),
    .B(_07413_),
    .Y(_07414_));
 OR4x1_ASAP7_75t_R _19552_ (.A(_00569_),
    .B(_00570_),
    .C(_00571_),
    .D(_07404_),
    .Y(_07415_));
 NAND2x1_ASAP7_75t_R _19553_ (.A(_00568_),
    .B(_07415_),
    .Y(_07416_));
 AND3x1_ASAP7_75t_R _19554_ (.A(_07403_),
    .B(_07414_),
    .C(_07416_),
    .Y(_04497_));
 OR4x1_ASAP7_75t_R _19555_ (.A(_00572_),
    .B(_00573_),
    .C(_07401_),
    .D(_07413_),
    .Y(_07417_));
 XOR2x2_ASAP7_75t_R _19556_ (.A(_07383_),
    .B(_07417_),
    .Y(_07418_));
 AND2x2_ASAP7_75t_R _19557_ (.A(_07316_),
    .B(_07418_),
    .Y(_04498_));
 OR3x1_ASAP7_75t_R _19558_ (.A(_00566_),
    .B(_07383_),
    .C(_07414_),
    .Y(_07419_));
 OAI21x1_ASAP7_75t_R _19559_ (.A1(_07383_),
    .A2(_07414_),
    .B(_00566_),
    .Y(_07420_));
 AND3x1_ASAP7_75t_R _19560_ (.A(_07403_),
    .B(_07419_),
    .C(_07420_),
    .Y(_04499_));
 OR3x1_ASAP7_75t_R _19561_ (.A(_00566_),
    .B(_07383_),
    .C(_07417_),
    .Y(_07421_));
 XOR2x2_ASAP7_75t_R _19562_ (.A(_00565_),
    .B(_07421_),
    .Y(_07422_));
 AND2x2_ASAP7_75t_R _19563_ (.A(_07316_),
    .B(_07422_),
    .Y(_04500_));
 NOR2x1_ASAP7_75t_R _19564_ (.A(_07190_),
    .B(_02650_),
    .Y(_04501_));
 OR4x1_ASAP7_75t_R _19565_ (.A(_00565_),
    .B(_00566_),
    .C(_07383_),
    .D(_07414_),
    .Y(_07423_));
 XOR2x2_ASAP7_75t_R _19566_ (.A(_00563_),
    .B(_07423_),
    .Y(_07424_));
 AND2x2_ASAP7_75t_R _19567_ (.A(_07316_),
    .B(_07424_),
    .Y(_04502_));
 OR5x1_ASAP7_75t_R _19568_ (.A(_00563_),
    .B(_00565_),
    .C(_00566_),
    .D(_07383_),
    .E(_07417_),
    .Y(_07425_));
 XOR2x2_ASAP7_75t_R _19569_ (.A(_00562_),
    .B(_07425_),
    .Y(_07426_));
 AND2x2_ASAP7_75t_R _19570_ (.A(_07316_),
    .B(_07426_),
    .Y(_04503_));
 OR5x2_ASAP7_75t_R _19571_ (.A(_00562_),
    .B(_00563_),
    .C(_00565_),
    .D(_00566_),
    .E(_07383_),
    .Y(_07427_));
 OR3x2_ASAP7_75t_R _19572_ (.A(_00561_),
    .B(_07414_),
    .C(_07427_),
    .Y(_07428_));
 OAI21x1_ASAP7_75t_R _19573_ (.A1(_07414_),
    .A2(_07427_),
    .B(_00561_),
    .Y(_07429_));
 AND3x1_ASAP7_75t_R _19574_ (.A(_07403_),
    .B(_07428_),
    .C(_07429_),
    .Y(_04504_));
 BUFx6f_ASAP7_75t_R _19575_ (.A(_07084_),
    .Y(_07430_));
 OR3x2_ASAP7_75t_R _19576_ (.A(_00561_),
    .B(_07417_),
    .C(_07427_),
    .Y(_07431_));
 XOR2x2_ASAP7_75t_R _19577_ (.A(_07387_),
    .B(_07431_),
    .Y(_07432_));
 AND2x2_ASAP7_75t_R _19578_ (.A(_07430_),
    .B(_07432_),
    .Y(_04505_));
 OR3x1_ASAP7_75t_R _19579_ (.A(_00559_),
    .B(_07387_),
    .C(_07428_),
    .Y(_07433_));
 OAI21x1_ASAP7_75t_R _19580_ (.A1(_07387_),
    .A2(_07428_),
    .B(_00559_),
    .Y(_07434_));
 AND3x1_ASAP7_75t_R _19581_ (.A(_07403_),
    .B(_07433_),
    .C(_07434_),
    .Y(_04506_));
 OR3x1_ASAP7_75t_R _19582_ (.A(_00559_),
    .B(_07387_),
    .C(_07431_),
    .Y(_07435_));
 XOR2x2_ASAP7_75t_R _19583_ (.A(_00558_),
    .B(_07435_),
    .Y(_07436_));
 AND2x2_ASAP7_75t_R _19584_ (.A(_07430_),
    .B(_07436_),
    .Y(_04507_));
 OR4x1_ASAP7_75t_R _19585_ (.A(_00558_),
    .B(_00559_),
    .C(_07387_),
    .D(_07428_),
    .Y(_07437_));
 XOR2x2_ASAP7_75t_R _19586_ (.A(_00557_),
    .B(_07437_),
    .Y(_07438_));
 AND2x2_ASAP7_75t_R _19587_ (.A(_07430_),
    .B(_07438_),
    .Y(_04508_));
 OR5x1_ASAP7_75t_R _19588_ (.A(_00557_),
    .B(_00558_),
    .C(_00559_),
    .D(_07387_),
    .E(_07431_),
    .Y(_07439_));
 XOR2x2_ASAP7_75t_R _19589_ (.A(_00556_),
    .B(_07439_),
    .Y(_07440_));
 AND2x2_ASAP7_75t_R _19590_ (.A(_07430_),
    .B(_07440_),
    .Y(_04509_));
 OR5x2_ASAP7_75t_R _19591_ (.A(_00556_),
    .B(_00557_),
    .C(_00558_),
    .D(_00559_),
    .E(_07387_),
    .Y(_07441_));
 OR3x1_ASAP7_75t_R _19592_ (.A(_00555_),
    .B(_07428_),
    .C(_07441_),
    .Y(_07442_));
 OAI21x1_ASAP7_75t_R _19593_ (.A1(_07428_),
    .A2(_07441_),
    .B(_00555_),
    .Y(_07443_));
 AND3x1_ASAP7_75t_R _19594_ (.A(_07403_),
    .B(_07442_),
    .C(_07443_),
    .Y(_04510_));
 OR3x1_ASAP7_75t_R _19595_ (.A(_00555_),
    .B(_07431_),
    .C(_07441_),
    .Y(_07444_));
 XOR2x2_ASAP7_75t_R _19596_ (.A(_00554_),
    .B(_07444_),
    .Y(_07445_));
 AND2x2_ASAP7_75t_R _19597_ (.A(_07430_),
    .B(_07445_),
    .Y(_04511_));
 XOR2x2_ASAP7_75t_R _19598_ (.A(_00553_),
    .B(_02649_),
    .Y(_07446_));
 AND2x2_ASAP7_75t_R _19599_ (.A(_07430_),
    .B(_07446_),
    .Y(_04512_));
 OR4x1_ASAP7_75t_R _19600_ (.A(_00554_),
    .B(_00555_),
    .C(_07428_),
    .D(_07441_),
    .Y(_07447_));
 XOR2x2_ASAP7_75t_R _19601_ (.A(_00552_),
    .B(_07447_),
    .Y(_07448_));
 AND2x2_ASAP7_75t_R _19602_ (.A(_07430_),
    .B(_07448_),
    .Y(_04513_));
 OR5x1_ASAP7_75t_R _19603_ (.A(_00552_),
    .B(_00554_),
    .C(_00555_),
    .D(_07431_),
    .E(_07441_),
    .Y(_07449_));
 XOR2x2_ASAP7_75t_R _19604_ (.A(_00551_),
    .B(_07449_),
    .Y(_07450_));
 AND2x2_ASAP7_75t_R _19605_ (.A(_07430_),
    .B(_07450_),
    .Y(_04514_));
 OR3x1_ASAP7_75t_R _19606_ (.A(_00553_),
    .B(_00564_),
    .C(_00053_),
    .Y(_07451_));
 XOR2x2_ASAP7_75t_R _19607_ (.A(_00550_),
    .B(_07451_),
    .Y(_07452_));
 AND2x2_ASAP7_75t_R _19608_ (.A(_07430_),
    .B(_07452_),
    .Y(_04515_));
 OR3x1_ASAP7_75t_R _19609_ (.A(_00550_),
    .B(_00553_),
    .C(_02649_),
    .Y(_07453_));
 NAND2x1_ASAP7_75t_R _19610_ (.A(_00549_),
    .B(_07453_),
    .Y(_07454_));
 AND3x1_ASAP7_75t_R _19611_ (.A(_07403_),
    .B(_07395_),
    .C(_07454_),
    .Y(_04516_));
 XOR2x2_ASAP7_75t_R _19612_ (.A(_00548_),
    .B(_07400_),
    .Y(_07455_));
 AND2x2_ASAP7_75t_R _19613_ (.A(_07430_),
    .B(_07455_),
    .Y(_04517_));
 OR3x1_ASAP7_75t_R _19614_ (.A(_00547_),
    .B(_00548_),
    .C(_07395_),
    .Y(_07456_));
 OAI21x1_ASAP7_75t_R _19615_ (.A1(_00548_),
    .A2(_07395_),
    .B(_00547_),
    .Y(_07457_));
 AND3x1_ASAP7_75t_R _19616_ (.A(_07403_),
    .B(_07456_),
    .C(_07457_),
    .Y(_04518_));
 BUFx6f_ASAP7_75t_R _19617_ (.A(_07084_),
    .Y(_07458_));
 OR3x1_ASAP7_75t_R _19618_ (.A(_00547_),
    .B(_00548_),
    .C(_07400_),
    .Y(_07459_));
 XOR2x2_ASAP7_75t_R _19619_ (.A(_00546_),
    .B(_07459_),
    .Y(_07460_));
 AND2x2_ASAP7_75t_R _19620_ (.A(_07458_),
    .B(_07460_),
    .Y(_04519_));
 OR4x1_ASAP7_75t_R _19621_ (.A(_00546_),
    .B(_00547_),
    .C(_00548_),
    .D(_07395_),
    .Y(_07461_));
 XOR2x2_ASAP7_75t_R _19622_ (.A(_00545_),
    .B(_07461_),
    .Y(_07462_));
 AND2x2_ASAP7_75t_R _19623_ (.A(_07458_),
    .B(_07462_),
    .Y(_04520_));
 OR3x1_ASAP7_75t_R _19624_ (.A(_00544_),
    .B(_07396_),
    .C(_07400_),
    .Y(_07463_));
 OAI21x1_ASAP7_75t_R _19625_ (.A1(_07396_),
    .A2(_07400_),
    .B(_00544_),
    .Y(_07464_));
 AND3x1_ASAP7_75t_R _19626_ (.A(_07403_),
    .B(_07463_),
    .C(_07464_),
    .Y(_04521_));
 BUFx6f_ASAP7_75t_R _19627_ (.A(_00534_),
    .Y(_07465_));
 AND4x1_ASAP7_75t_R _19628_ (.A(_00505_),
    .B(_00533_),
    .C(_07465_),
    .D(_00535_),
    .Y(_07466_));
 AND5x1_ASAP7_75t_R _19629_ (.A(_00524_),
    .B(_00529_),
    .C(_00530_),
    .D(_00532_),
    .E(_07466_),
    .Y(_07467_));
 AND5x2_ASAP7_75t_R _19630_ (.A(_00526_),
    .B(_00527_),
    .C(_00528_),
    .D(_07147_),
    .E(_07467_),
    .Y(_07468_));
 AND4x1_ASAP7_75t_R _19631_ (.A(_00519_),
    .B(_00520_),
    .C(_00521_),
    .D(_00522_),
    .Y(_07469_));
 AND4x1_ASAP7_75t_R _19632_ (.A(_00513_),
    .B(_00515_),
    .C(_00516_),
    .D(_00523_),
    .Y(_07470_));
 AND5x1_ASAP7_75t_R _19633_ (.A(_00506_),
    .B(_00507_),
    .C(_00512_),
    .D(_00531_),
    .E(_07470_),
    .Y(_07471_));
 BUFx3_ASAP7_75t_R _19634_ (.A(_00509_),
    .Y(_07472_));
 AND3x1_ASAP7_75t_R _19635_ (.A(_00510_),
    .B(_00511_),
    .C(_00514_),
    .Y(_07473_));
 OR3x1_ASAP7_75t_R _19636_ (.A(_00508_),
    .B(_07472_),
    .C(_07473_),
    .Y(_07474_));
 AND5x2_ASAP7_75t_R _19637_ (.A(_00517_),
    .B(_00518_),
    .C(_07469_),
    .D(_07471_),
    .E(_07474_),
    .Y(_07475_));
 NAND2x2_ASAP7_75t_R _19638_ (.A(_07468_),
    .B(_07475_),
    .Y(_07476_));
 NOR2x1_ASAP7_75t_R _19639_ (.A(_00495_),
    .B(_07476_),
    .Y(_04522_));
 INVx1_ASAP7_75t_R _19640_ (.A(_07476_),
    .Y(_04523_));
 NOR2x1_ASAP7_75t_R _19641_ (.A(_00498_),
    .B(_07476_),
    .Y(_04524_));
 NOR2x1_ASAP7_75t_R _19642_ (.A(_00497_),
    .B(_07476_),
    .Y(_04525_));
 NOR2x1_ASAP7_75t_R _19643_ (.A(_00496_),
    .B(_07476_),
    .Y(_04526_));
 NOR2x1_ASAP7_75t_R _19644_ (.A(_00494_),
    .B(_07476_),
    .Y(_04527_));
 NOR2x1_ASAP7_75t_R _19645_ (.A(_00493_),
    .B(_07476_),
    .Y(_04528_));
 INVx1_ASAP7_75t_R _19646_ (.A(_07476_),
    .Y(_04529_));
 AND2x2_ASAP7_75t_R _19647_ (.A(_07458_),
    .B(_00054_),
    .Y(_04530_));
 BUFx6f_ASAP7_75t_R _19648_ (.A(_08998_),
    .Y(_07477_));
 OR4x1_ASAP7_75t_R _19649_ (.A(_00510_),
    .B(_00511_),
    .C(_00514_),
    .D(_02619_),
    .Y(_07478_));
 OR5x2_ASAP7_75t_R _19650_ (.A(_00505_),
    .B(_00506_),
    .C(_00507_),
    .D(_00508_),
    .E(_07472_),
    .Y(_07479_));
 OR3x1_ASAP7_75t_R _19651_ (.A(_00535_),
    .B(_07478_),
    .C(_07479_),
    .Y(_07480_));
 BUFx6f_ASAP7_75t_R _19652_ (.A(_07480_),
    .Y(_07481_));
 OAI21x1_ASAP7_75t_R _19653_ (.A1(_07478_),
    .A2(_07479_),
    .B(_00535_),
    .Y(_07482_));
 AND3x1_ASAP7_75t_R _19654_ (.A(_07477_),
    .B(_07481_),
    .C(_07482_),
    .Y(_04531_));
 OR5x2_ASAP7_75t_R _19655_ (.A(_00510_),
    .B(_00511_),
    .C(_00514_),
    .D(_00525_),
    .E(_00054_),
    .Y(_07483_));
 OR3x2_ASAP7_75t_R _19656_ (.A(_00535_),
    .B(_07479_),
    .C(_07483_),
    .Y(_07484_));
 XOR2x2_ASAP7_75t_R _19657_ (.A(_07465_),
    .B(_07484_),
    .Y(_07485_));
 AND2x2_ASAP7_75t_R _19658_ (.A(_07458_),
    .B(_07485_),
    .Y(_04532_));
 OR3x1_ASAP7_75t_R _19659_ (.A(_00533_),
    .B(_07465_),
    .C(_07481_),
    .Y(_07486_));
 OAI21x1_ASAP7_75t_R _19660_ (.A1(_07465_),
    .A2(_07481_),
    .B(_00533_),
    .Y(_07487_));
 AND3x1_ASAP7_75t_R _19661_ (.A(_07477_),
    .B(_07486_),
    .C(_07487_),
    .Y(_04533_));
 OR3x1_ASAP7_75t_R _19662_ (.A(_00533_),
    .B(_07465_),
    .C(_07484_),
    .Y(_07488_));
 XOR2x2_ASAP7_75t_R _19663_ (.A(_00532_),
    .B(_07488_),
    .Y(_07489_));
 AND2x2_ASAP7_75t_R _19664_ (.A(_07458_),
    .B(_07489_),
    .Y(_04534_));
 OR4x1_ASAP7_75t_R _19665_ (.A(_00532_),
    .B(_00533_),
    .C(_07465_),
    .D(_07481_),
    .Y(_07490_));
 XOR2x2_ASAP7_75t_R _19666_ (.A(_00531_),
    .B(_07490_),
    .Y(_07491_));
 AND2x2_ASAP7_75t_R _19667_ (.A(_07458_),
    .B(_07491_),
    .Y(_04535_));
 OR5x2_ASAP7_75t_R _19668_ (.A(_00530_),
    .B(_00531_),
    .C(_00532_),
    .D(_00533_),
    .E(_07465_),
    .Y(_07492_));
 OR5x1_ASAP7_75t_R _19669_ (.A(_00531_),
    .B(_00532_),
    .C(_00533_),
    .D(_07465_),
    .E(_07484_),
    .Y(_07493_));
 NAND2x1_ASAP7_75t_R _19670_ (.A(_00530_),
    .B(_07493_),
    .Y(_07494_));
 OA211x2_ASAP7_75t_R _19671_ (.A1(_07484_),
    .A2(_07492_),
    .B(_07494_),
    .C(_07260_),
    .Y(_04536_));
 OR3x1_ASAP7_75t_R _19672_ (.A(_00529_),
    .B(_07481_),
    .C(_07492_),
    .Y(_07495_));
 OAI21x1_ASAP7_75t_R _19673_ (.A1(_07481_),
    .A2(_07492_),
    .B(_00529_),
    .Y(_07496_));
 AND3x1_ASAP7_75t_R _19674_ (.A(_07477_),
    .B(_07495_),
    .C(_07496_),
    .Y(_04537_));
 OR3x1_ASAP7_75t_R _19675_ (.A(_00529_),
    .B(_07484_),
    .C(_07492_),
    .Y(_07497_));
 XOR2x2_ASAP7_75t_R _19676_ (.A(_00528_),
    .B(_07497_),
    .Y(_07498_));
 AND2x2_ASAP7_75t_R _19677_ (.A(_07458_),
    .B(_07498_),
    .Y(_04538_));
 OR5x2_ASAP7_75t_R _19678_ (.A(_00527_),
    .B(_00528_),
    .C(_00529_),
    .D(_07481_),
    .E(_07492_),
    .Y(_07499_));
 OR4x1_ASAP7_75t_R _19679_ (.A(_00528_),
    .B(_00529_),
    .C(_07481_),
    .D(_07492_),
    .Y(_07500_));
 NAND2x1_ASAP7_75t_R _19680_ (.A(_00527_),
    .B(_07500_),
    .Y(_07501_));
 AND3x1_ASAP7_75t_R _19681_ (.A(_07477_),
    .B(_07499_),
    .C(_07501_),
    .Y(_04539_));
 OR5x2_ASAP7_75t_R _19682_ (.A(_00527_),
    .B(_00528_),
    .C(_00529_),
    .D(_07484_),
    .E(_07492_),
    .Y(_07502_));
 XOR2x2_ASAP7_75t_R _19683_ (.A(_00526_),
    .B(_07502_),
    .Y(_07503_));
 AND2x2_ASAP7_75t_R _19684_ (.A(_07458_),
    .B(_07503_),
    .Y(_04540_));
 NOR2x1_ASAP7_75t_R _19685_ (.A(_07190_),
    .B(_02620_),
    .Y(_04541_));
 OR3x1_ASAP7_75t_R _19686_ (.A(_00524_),
    .B(_00526_),
    .C(_07499_),
    .Y(_07504_));
 OAI21x1_ASAP7_75t_R _19687_ (.A1(_00526_),
    .A2(_07499_),
    .B(_00524_),
    .Y(_07505_));
 AND3x1_ASAP7_75t_R _19688_ (.A(_07477_),
    .B(_07504_),
    .C(_07505_),
    .Y(_04542_));
 OR3x1_ASAP7_75t_R _19689_ (.A(_00524_),
    .B(_00526_),
    .C(_07502_),
    .Y(_07506_));
 XOR2x2_ASAP7_75t_R _19690_ (.A(_00523_),
    .B(_07506_),
    .Y(_07507_));
 AND2x2_ASAP7_75t_R _19691_ (.A(_07458_),
    .B(_07507_),
    .Y(_04543_));
 OR4x1_ASAP7_75t_R _19692_ (.A(_00523_),
    .B(_00524_),
    .C(_00526_),
    .D(_07499_),
    .Y(_07508_));
 XOR2x2_ASAP7_75t_R _19693_ (.A(_00522_),
    .B(_07508_),
    .Y(_07509_));
 AND2x2_ASAP7_75t_R _19694_ (.A(_07458_),
    .B(_07509_),
    .Y(_04544_));
 OR4x1_ASAP7_75t_R _19695_ (.A(_00522_),
    .B(_00523_),
    .C(_00524_),
    .D(_00526_),
    .Y(_07510_));
 OR3x2_ASAP7_75t_R _19696_ (.A(_00521_),
    .B(_07502_),
    .C(_07510_),
    .Y(_07511_));
 OAI21x1_ASAP7_75t_R _19697_ (.A1(_07502_),
    .A2(_07510_),
    .B(_00521_),
    .Y(_07512_));
 AND3x1_ASAP7_75t_R _19698_ (.A(_07477_),
    .B(_07511_),
    .C(_07512_),
    .Y(_04545_));
 BUFx6f_ASAP7_75t_R _19699_ (.A(_07084_),
    .Y(_07513_));
 OR3x2_ASAP7_75t_R _19700_ (.A(_00521_),
    .B(_07499_),
    .C(_07510_),
    .Y(_07514_));
 XOR2x2_ASAP7_75t_R _19701_ (.A(_00520_),
    .B(_07514_),
    .Y(_07515_));
 AND2x2_ASAP7_75t_R _19702_ (.A(_07513_),
    .B(_07515_),
    .Y(_04546_));
 OR3x1_ASAP7_75t_R _19703_ (.A(_00519_),
    .B(_00520_),
    .C(_07511_),
    .Y(_07516_));
 OAI21x1_ASAP7_75t_R _19704_ (.A1(_00520_),
    .A2(_07511_),
    .B(_00519_),
    .Y(_07517_));
 AND3x1_ASAP7_75t_R _19705_ (.A(_07477_),
    .B(_07516_),
    .C(_07517_),
    .Y(_04547_));
 OR3x1_ASAP7_75t_R _19706_ (.A(_00519_),
    .B(_00520_),
    .C(_07514_),
    .Y(_07518_));
 XOR2x2_ASAP7_75t_R _19707_ (.A(_00518_),
    .B(_07518_),
    .Y(_07519_));
 AND2x2_ASAP7_75t_R _19708_ (.A(_07513_),
    .B(_07519_),
    .Y(_04548_));
 OR4x1_ASAP7_75t_R _19709_ (.A(_00518_),
    .B(_00519_),
    .C(_00520_),
    .D(_07511_),
    .Y(_07520_));
 XOR2x2_ASAP7_75t_R _19710_ (.A(_00517_),
    .B(_07520_),
    .Y(_07521_));
 AND2x2_ASAP7_75t_R _19711_ (.A(_07513_),
    .B(_07521_),
    .Y(_04549_));
 OR4x1_ASAP7_75t_R _19712_ (.A(_00517_),
    .B(_00518_),
    .C(_00519_),
    .D(_00520_),
    .Y(_07522_));
 OR3x1_ASAP7_75t_R _19713_ (.A(_00516_),
    .B(_07514_),
    .C(_07522_),
    .Y(_07523_));
 OAI21x1_ASAP7_75t_R _19714_ (.A1(_07514_),
    .A2(_07522_),
    .B(_00516_),
    .Y(_07524_));
 AND3x1_ASAP7_75t_R _19715_ (.A(_07477_),
    .B(_07523_),
    .C(_07524_),
    .Y(_04550_));
 OR3x1_ASAP7_75t_R _19716_ (.A(_00516_),
    .B(_07511_),
    .C(_07522_),
    .Y(_07525_));
 XOR2x2_ASAP7_75t_R _19717_ (.A(_00515_),
    .B(_07525_),
    .Y(_07526_));
 AND2x2_ASAP7_75t_R _19718_ (.A(_07513_),
    .B(_07526_),
    .Y(_04551_));
 XOR2x2_ASAP7_75t_R _19719_ (.A(_00514_),
    .B(_02619_),
    .Y(_07527_));
 AND2x2_ASAP7_75t_R _19720_ (.A(_07513_),
    .B(_07527_),
    .Y(_04552_));
 OR4x1_ASAP7_75t_R _19721_ (.A(_00515_),
    .B(_00516_),
    .C(_07514_),
    .D(_07522_),
    .Y(_07528_));
 XOR2x2_ASAP7_75t_R _19722_ (.A(_00513_),
    .B(_07528_),
    .Y(_07529_));
 AND2x2_ASAP7_75t_R _19723_ (.A(_07513_),
    .B(_07529_),
    .Y(_04553_));
 OR5x1_ASAP7_75t_R _19724_ (.A(_00513_),
    .B(_00515_),
    .C(_00516_),
    .D(_07511_),
    .E(_07522_),
    .Y(_07530_));
 XOR2x2_ASAP7_75t_R _19725_ (.A(_00512_),
    .B(_07530_),
    .Y(_07531_));
 AND2x2_ASAP7_75t_R _19726_ (.A(_07513_),
    .B(_07531_),
    .Y(_04554_));
 OR3x1_ASAP7_75t_R _19727_ (.A(_00514_),
    .B(_00525_),
    .C(_00054_),
    .Y(_07532_));
 XOR2x2_ASAP7_75t_R _19728_ (.A(_00511_),
    .B(_07532_),
    .Y(_07533_));
 AND2x2_ASAP7_75t_R _19729_ (.A(_07513_),
    .B(_07533_),
    .Y(_04555_));
 OR3x1_ASAP7_75t_R _19730_ (.A(_00511_),
    .B(_00514_),
    .C(_02619_),
    .Y(_07534_));
 NAND2x1_ASAP7_75t_R _19731_ (.A(_00510_),
    .B(_07534_),
    .Y(_07535_));
 AND3x1_ASAP7_75t_R _19732_ (.A(_07477_),
    .B(_07478_),
    .C(_07535_),
    .Y(_04556_));
 XOR2x2_ASAP7_75t_R _19733_ (.A(_07472_),
    .B(_07483_),
    .Y(_07536_));
 AND2x2_ASAP7_75t_R _19734_ (.A(_07513_),
    .B(_07536_),
    .Y(_04557_));
 OR3x1_ASAP7_75t_R _19735_ (.A(_00508_),
    .B(_07472_),
    .C(_07478_),
    .Y(_07537_));
 OAI21x1_ASAP7_75t_R _19736_ (.A1(_07472_),
    .A2(_07478_),
    .B(_00508_),
    .Y(_07538_));
 AND3x1_ASAP7_75t_R _19737_ (.A(_07477_),
    .B(_07537_),
    .C(_07538_),
    .Y(_04558_));
 OR3x1_ASAP7_75t_R _19738_ (.A(_00508_),
    .B(_07472_),
    .C(_07483_),
    .Y(_07539_));
 XOR2x2_ASAP7_75t_R _19739_ (.A(_00507_),
    .B(_07539_),
    .Y(_07540_));
 AND2x2_ASAP7_75t_R _19740_ (.A(_07513_),
    .B(_07540_),
    .Y(_04559_));
 BUFx6f_ASAP7_75t_R _19741_ (.A(_07084_),
    .Y(_07541_));
 OR4x1_ASAP7_75t_R _19742_ (.A(_00507_),
    .B(_00508_),
    .C(_07472_),
    .D(_07478_),
    .Y(_07542_));
 XOR2x2_ASAP7_75t_R _19743_ (.A(_00506_),
    .B(_07542_),
    .Y(_07543_));
 AND2x2_ASAP7_75t_R _19744_ (.A(_07541_),
    .B(_07543_),
    .Y(_04560_));
 OR5x1_ASAP7_75t_R _19745_ (.A(_00506_),
    .B(_00507_),
    .C(_00508_),
    .D(_07472_),
    .E(_07483_),
    .Y(_07544_));
 XOR2x2_ASAP7_75t_R _19746_ (.A(_00505_),
    .B(_07544_),
    .Y(_07545_));
 AND2x2_ASAP7_75t_R _19747_ (.A(_07541_),
    .B(_07545_),
    .Y(_04561_));
 AND2x2_ASAP7_75t_R _19748_ (.A(_07541_),
    .B(_00026_),
    .Y(_04562_));
 BUFx6f_ASAP7_75t_R _19749_ (.A(_02232_),
    .Y(_07546_));
 INVx2_ASAP7_75t_R _19750_ (.A(_02239_),
    .Y(_07547_));
 OR2x2_ASAP7_75t_R _19751_ (.A(_00575_),
    .B(_00580_),
    .Y(_07548_));
 AND4x1_ASAP7_75t_R _19752_ (.A(_00537_),
    .B(\xs[5].cli1.i[35] ),
    .C(_00539_),
    .D(\xs[5].cli1.i[33] ),
    .Y(_07549_));
 NAND3x1_ASAP7_75t_R _19753_ (.A(\xs[5].cli1.i[39] ),
    .B(_00541_),
    .C(_07549_),
    .Y(_07550_));
 OAI21x1_ASAP7_75t_R _19754_ (.A1(_08525_),
    .A2(_07549_),
    .B(_07547_),
    .Y(_07551_));
 AND4x1_ASAP7_75t_R _19755_ (.A(_00576_),
    .B(\peo[10][35] ),
    .C(_00578_),
    .D(\peo[10][33] ),
    .Y(_07552_));
 NOR2x1_ASAP7_75t_R _19756_ (.A(_00575_),
    .B(_07552_),
    .Y(_07553_));
 AO221x1_ASAP7_75t_R _19757_ (.A1(_07547_),
    .A2(_07548_),
    .B1(_07550_),
    .B2(_07551_),
    .C(_07553_),
    .Y(_07554_));
 NAND2x1_ASAP7_75t_R _19758_ (.A(_02233_),
    .B(_07554_),
    .Y(_07555_));
 OR4x1_ASAP7_75t_R _19759_ (.A(_09220_),
    .B(_07546_),
    .C(_07547_),
    .D(_07555_),
    .Y(_07556_));
 BUFx6f_ASAP7_75t_R _19760_ (.A(_07556_),
    .Y(_07557_));
 AND2x4_ASAP7_75t_R _19761_ (.A(_02233_),
    .B(_07554_),
    .Y(_07558_));
 INVx2_ASAP7_75t_R _19762_ (.A(_07546_),
    .Y(_07559_));
 NAND2x1_ASAP7_75t_R _19763_ (.A(_07559_),
    .B(_02239_),
    .Y(_07560_));
 INVx1_ASAP7_75t_R _19764_ (.A(_07560_),
    .Y(_07561_));
 AND3x1_ASAP7_75t_R _19765_ (.A(\xs[5].cli1.i[39] ),
    .B(_00541_),
    .C(_07549_),
    .Y(_07562_));
 INVx1_ASAP7_75t_R _19766_ (.A(_00026_),
    .Y(_07563_));
 OR4x1_ASAP7_75t_R _19767_ (.A(_07559_),
    .B(_07563_),
    .C(_08525_),
    .D(_07549_),
    .Y(_07564_));
 AO21x1_ASAP7_75t_R _19768_ (.A1(_02233_),
    .A2(_07547_),
    .B(_07546_),
    .Y(_07565_));
 OR2x6_ASAP7_75t_R _19769_ (.A(_00575_),
    .B(_07552_),
    .Y(_07566_));
 AO21x1_ASAP7_75t_R _19770_ (.A1(_07564_),
    .A2(_07565_),
    .B(_07566_),
    .Y(_07567_));
 NAND2x1_ASAP7_75t_R _19771_ (.A(_07562_),
    .B(_07567_),
    .Y(_07568_));
 AO221x1_ASAP7_75t_R _19772_ (.A1(_07558_),
    .A2(_07561_),
    .B1(_07568_),
    .B2(_00582_),
    .C(_09314_),
    .Y(_07569_));
 INVx1_ASAP7_75t_R _19773_ (.A(_02233_),
    .Y(_07570_));
 NOR2x1_ASAP7_75t_R _19774_ (.A(_08525_),
    .B(_07549_),
    .Y(_07571_));
 AO21x1_ASAP7_75t_R _19775_ (.A1(_07553_),
    .A2(_07562_),
    .B(_07571_),
    .Y(_07572_));
 AO21x1_ASAP7_75t_R _19776_ (.A1(\xs[5].cli1.i[32] ),
    .A2(_07549_),
    .B(_08525_),
    .Y(_07573_));
 OAI21x1_ASAP7_75t_R _19777_ (.A1(_07560_),
    .A2(_07573_),
    .B(_07564_),
    .Y(_07574_));
 AO32x2_ASAP7_75t_R _19778_ (.A1(_07559_),
    .A2(_07570_),
    .A3(_07572_),
    .B1(_07574_),
    .B2(_07553_),
    .Y(_07575_));
 NOR3x1_ASAP7_75t_R _19779_ (.A(\peo[11][0] ),
    .B(_07550_),
    .C(_07575_),
    .Y(_07576_));
 OAI22x1_ASAP7_75t_R _19780_ (.A1(_02243_),
    .A2(_07557_),
    .B1(_07569_),
    .B2(_07576_),
    .Y(_04563_));
 NOR2x1_ASAP7_75t_R _19781_ (.A(_02242_),
    .B(_07557_),
    .Y(_04564_));
 NOR2x1_ASAP7_75t_R _19782_ (.A(_02241_),
    .B(_07557_),
    .Y(_04565_));
 NOR2x1_ASAP7_75t_R _19783_ (.A(_02240_),
    .B(_07557_),
    .Y(_04566_));
 NOR2x1_ASAP7_75t_R _19784_ (.A(_02231_),
    .B(_07557_),
    .Y(_04567_));
 NOR2x1_ASAP7_75t_R _19785_ (.A(_02230_),
    .B(_07557_),
    .Y(_04568_));
 AND3x1_ASAP7_75t_R _19786_ (.A(_07559_),
    .B(_02233_),
    .C(_07547_),
    .Y(_07577_));
 NAND2x1_ASAP7_75t_R _19787_ (.A(_07554_),
    .B(_07577_),
    .Y(_07578_));
 INVx1_ASAP7_75t_R _19788_ (.A(_02243_),
    .Y(_07579_));
 AND3x1_ASAP7_75t_R _19789_ (.A(_07579_),
    .B(_07554_),
    .C(_07577_),
    .Y(_07580_));
 AO21x1_ASAP7_75t_R _19790_ (.A1(\peo[10][0] ),
    .A2(_07578_),
    .B(_07580_),
    .Y(_07581_));
 NAND2x1_ASAP7_75t_R _19791_ (.A(_00543_),
    .B(_07575_),
    .Y(_07582_));
 OA211x2_ASAP7_75t_R _19792_ (.A1(_07575_),
    .A2(_07581_),
    .B(_07582_),
    .C(_07260_),
    .Y(_04569_));
 OR4x1_ASAP7_75t_R _19793_ (.A(_11177_),
    .B(_07546_),
    .C(_02239_),
    .D(_07555_),
    .Y(_07583_));
 NOR2x1_ASAP7_75t_R _19794_ (.A(_02242_),
    .B(_07583_),
    .Y(_04570_));
 NOR2x1_ASAP7_75t_R _19795_ (.A(_02241_),
    .B(_07583_),
    .Y(_04571_));
 NOR2x1_ASAP7_75t_R _19796_ (.A(_02240_),
    .B(_07583_),
    .Y(_04572_));
 NOR2x1_ASAP7_75t_R _19797_ (.A(_02231_),
    .B(_07583_),
    .Y(_04573_));
 NOR2x1_ASAP7_75t_R _19798_ (.A(_02230_),
    .B(_07583_),
    .Y(_04574_));
 OA21x2_ASAP7_75t_R _19799_ (.A1(_07546_),
    .A2(_07558_),
    .B(_08584_),
    .Y(_07584_));
 OA21x2_ASAP7_75t_R _19800_ (.A1(_07560_),
    .A2(_07573_),
    .B(_07564_),
    .Y(_07585_));
 OA21x2_ASAP7_75t_R _19801_ (.A1(_07546_),
    .A2(_02233_),
    .B(_07571_),
    .Y(_07586_));
 OA21x2_ASAP7_75t_R _19802_ (.A1(_07566_),
    .A2(_07585_),
    .B(_07586_),
    .Y(_07587_));
 NAND2x1_ASAP7_75t_R _19803_ (.A(_00543_),
    .B(_07587_),
    .Y(_07588_));
 OAI21x1_ASAP7_75t_R _19804_ (.A1(_07566_),
    .A2(_07585_),
    .B(_07586_),
    .Y(_07589_));
 NAND2x1_ASAP7_75t_R _19805_ (.A(_00582_),
    .B(_07589_),
    .Y(_07590_));
 AND3x4_ASAP7_75t_R _19806_ (.A(_08598_),
    .B(_07559_),
    .C(_07555_),
    .Y(_07591_));
 AO32x1_ASAP7_75t_R _19807_ (.A1(_07584_),
    .A2(_07588_),
    .A3(_07590_),
    .B1(_07591_),
    .B2(_07579_),
    .Y(_04575_));
 OR3x1_ASAP7_75t_R _19808_ (.A(_08578_),
    .B(_07546_),
    .C(_07558_),
    .Y(_07592_));
 BUFx6f_ASAP7_75t_R _19809_ (.A(_07592_),
    .Y(_07593_));
 NOR2x1_ASAP7_75t_R _19810_ (.A(_02242_),
    .B(_07593_),
    .Y(_04576_));
 NOR2x1_ASAP7_75t_R _19811_ (.A(_02241_),
    .B(_07593_),
    .Y(_04577_));
 NOR2x1_ASAP7_75t_R _19812_ (.A(_02240_),
    .B(_07593_),
    .Y(_04578_));
 NAND2x1_ASAP7_75t_R _19813_ (.A(_00541_),
    .B(_07587_),
    .Y(_07594_));
 NAND2x1_ASAP7_75t_R _19814_ (.A(_00580_),
    .B(_07589_),
    .Y(_07595_));
 AO32x1_ASAP7_75t_R _19815_ (.A1(_07584_),
    .A2(_07594_),
    .A3(_07595_),
    .B1(_07591_),
    .B2(_07547_),
    .Y(_04579_));
 OAI21x1_ASAP7_75t_R _19816_ (.A1(_00575_),
    .A2(_07585_),
    .B(_07586_),
    .Y(_07596_));
 NAND2x1_ASAP7_75t_R _19817_ (.A(_00579_),
    .B(_07596_),
    .Y(_07597_));
 OR3x1_ASAP7_75t_R _19818_ (.A(_08525_),
    .B(\xs[5].cli1.i[33] ),
    .C(_07575_),
    .Y(_07598_));
 INVx1_ASAP7_75t_R _19819_ (.A(_02238_),
    .Y(_07599_));
 AO32x1_ASAP7_75t_R _19820_ (.A1(_07584_),
    .A2(_07597_),
    .A3(_07598_),
    .B1(_07591_),
    .B2(_07599_),
    .Y(_04580_));
 NAND2x1_ASAP7_75t_R _19821_ (.A(_00539_),
    .B(_07587_),
    .Y(_07600_));
 NAND2x1_ASAP7_75t_R _19822_ (.A(_00578_),
    .B(_07589_),
    .Y(_07601_));
 INVx1_ASAP7_75t_R _19823_ (.A(_02237_),
    .Y(_07602_));
 AO32x1_ASAP7_75t_R _19824_ (.A1(_07584_),
    .A2(_07600_),
    .A3(_07601_),
    .B1(_07591_),
    .B2(_07602_),
    .Y(_04581_));
 NAND2x1_ASAP7_75t_R _19825_ (.A(_00577_),
    .B(_07596_),
    .Y(_07603_));
 OR3x1_ASAP7_75t_R _19826_ (.A(_08525_),
    .B(\xs[5].cli1.i[35] ),
    .C(_07575_),
    .Y(_07604_));
 INVx1_ASAP7_75t_R _19827_ (.A(_02236_),
    .Y(_07605_));
 AO32x1_ASAP7_75t_R _19828_ (.A1(_07584_),
    .A2(_07603_),
    .A3(_07604_),
    .B1(_07591_),
    .B2(_07605_),
    .Y(_04582_));
 NAND2x1_ASAP7_75t_R _19829_ (.A(_00537_),
    .B(_07587_),
    .Y(_07606_));
 NAND2x1_ASAP7_75t_R _19830_ (.A(_00576_),
    .B(_07589_),
    .Y(_07607_));
 INVx1_ASAP7_75t_R _19831_ (.A(_02235_),
    .Y(_07608_));
 AO32x1_ASAP7_75t_R _19832_ (.A1(_07584_),
    .A2(_07606_),
    .A3(_07607_),
    .B1(_07591_),
    .B2(_07608_),
    .Y(_04583_));
 NOR2x1_ASAP7_75t_R _19833_ (.A(_02234_),
    .B(_07593_),
    .Y(_04584_));
 OR4x1_ASAP7_75t_R _19834_ (.A(_08684_),
    .B(_07546_),
    .C(_07570_),
    .D(_07554_),
    .Y(_07609_));
 INVx1_ASAP7_75t_R _19835_ (.A(_07609_),
    .Y(_04585_));
 INVx1_ASAP7_75t_R _19836_ (.A(_07571_),
    .Y(_07610_));
 OA211x2_ASAP7_75t_R _19837_ (.A1(_07546_),
    .A2(_07558_),
    .B(_07610_),
    .C(_07566_),
    .Y(_07611_));
 NOR2x1_ASAP7_75t_R _19838_ (.A(_07190_),
    .B(_07611_),
    .Y(_04586_));
 NOR2x1_ASAP7_75t_R _19839_ (.A(_02231_),
    .B(_07593_),
    .Y(_04587_));
 NOR2x1_ASAP7_75t_R _19840_ (.A(_02230_),
    .B(_07593_),
    .Y(_04588_));
 AND4x1_ASAP7_75t_R _19841_ (.A(_00440_),
    .B(_00468_),
    .C(_00469_),
    .D(_00470_),
    .Y(_07612_));
 AND5x1_ASAP7_75t_R _19842_ (.A(_00459_),
    .B(_00464_),
    .C(_00465_),
    .D(_00467_),
    .E(_07612_),
    .Y(_07613_));
 AND5x2_ASAP7_75t_R _19843_ (.A(_00461_),
    .B(_00462_),
    .C(_00463_),
    .D(_07147_),
    .E(_07613_),
    .Y(_07614_));
 BUFx3_ASAP7_75t_R _19844_ (.A(_00455_),
    .Y(_07615_));
 AND4x1_ASAP7_75t_R _19845_ (.A(_00454_),
    .B(_07615_),
    .C(_00456_),
    .D(_00457_),
    .Y(_07616_));
 AND4x1_ASAP7_75t_R _19846_ (.A(_00448_),
    .B(_00450_),
    .C(_00451_),
    .D(_00458_),
    .Y(_07617_));
 AND5x1_ASAP7_75t_R _19847_ (.A(_00441_),
    .B(_00442_),
    .C(_00447_),
    .D(_00466_),
    .E(_07617_),
    .Y(_07618_));
 BUFx6f_ASAP7_75t_R _19848_ (.A(_00444_),
    .Y(_07619_));
 AND3x1_ASAP7_75t_R _19849_ (.A(_00445_),
    .B(_00446_),
    .C(_00449_),
    .Y(_07620_));
 OR3x1_ASAP7_75t_R _19850_ (.A(_00443_),
    .B(_07619_),
    .C(_07620_),
    .Y(_07621_));
 AND5x2_ASAP7_75t_R _19851_ (.A(_00452_),
    .B(_00453_),
    .C(_07616_),
    .D(_07618_),
    .E(_07621_),
    .Y(_07622_));
 NAND2x2_ASAP7_75t_R _19852_ (.A(_07614_),
    .B(_07622_),
    .Y(_07623_));
 NOR2x1_ASAP7_75t_R _19853_ (.A(_00397_),
    .B(_07623_),
    .Y(_04589_));
 INVx1_ASAP7_75t_R _19854_ (.A(_07623_),
    .Y(_04590_));
 NOR2x1_ASAP7_75t_R _19855_ (.A(_00400_),
    .B(_07623_),
    .Y(_04591_));
 NOR2x1_ASAP7_75t_R _19856_ (.A(_00399_),
    .B(_07623_),
    .Y(_04592_));
 NOR2x1_ASAP7_75t_R _19857_ (.A(_00398_),
    .B(_07623_),
    .Y(_04593_));
 NOR2x1_ASAP7_75t_R _19858_ (.A(_00396_),
    .B(_07623_),
    .Y(_04594_));
 NOR2x1_ASAP7_75t_R _19859_ (.A(_00395_),
    .B(_07623_),
    .Y(_04595_));
 INVx1_ASAP7_75t_R _19860_ (.A(_07623_),
    .Y(_04596_));
 AND2x2_ASAP7_75t_R _19861_ (.A(_07541_),
    .B(_00055_),
    .Y(_04597_));
 BUFx6f_ASAP7_75t_R _19862_ (.A(_08998_),
    .Y(_07624_));
 OR4x1_ASAP7_75t_R _19863_ (.A(_00445_),
    .B(_00446_),
    .C(_00449_),
    .D(_02621_),
    .Y(_07625_));
 OR5x2_ASAP7_75t_R _19864_ (.A(_00440_),
    .B(_00441_),
    .C(_00442_),
    .D(_00443_),
    .E(_07619_),
    .Y(_07626_));
 OR3x1_ASAP7_75t_R _19865_ (.A(_00470_),
    .B(_07625_),
    .C(_07626_),
    .Y(_07627_));
 OAI21x1_ASAP7_75t_R _19866_ (.A1(_07625_),
    .A2(_07626_),
    .B(_00470_),
    .Y(_07628_));
 AND3x1_ASAP7_75t_R _19867_ (.A(_07624_),
    .B(_07627_),
    .C(_07628_),
    .Y(_04598_));
 OR5x2_ASAP7_75t_R _19868_ (.A(_00445_),
    .B(_00446_),
    .C(_00449_),
    .D(_00460_),
    .E(_00055_),
    .Y(_07629_));
 OR4x1_ASAP7_75t_R _19869_ (.A(_00469_),
    .B(_00470_),
    .C(_07626_),
    .D(_07629_),
    .Y(_07630_));
 OR3x1_ASAP7_75t_R _19870_ (.A(_00470_),
    .B(_07626_),
    .C(_07629_),
    .Y(_07631_));
 NAND2x1_ASAP7_75t_R _19871_ (.A(_00469_),
    .B(_07631_),
    .Y(_07632_));
 AND3x1_ASAP7_75t_R _19872_ (.A(_07624_),
    .B(_07630_),
    .C(_07632_),
    .Y(_04599_));
 OR4x1_ASAP7_75t_R _19873_ (.A(_00469_),
    .B(_00470_),
    .C(_07625_),
    .D(_07626_),
    .Y(_07633_));
 XOR2x2_ASAP7_75t_R _19874_ (.A(_00468_),
    .B(_07633_),
    .Y(_07634_));
 AND2x2_ASAP7_75t_R _19875_ (.A(_07541_),
    .B(_07634_),
    .Y(_04600_));
 OR3x1_ASAP7_75t_R _19876_ (.A(_00467_),
    .B(_00468_),
    .C(_07630_),
    .Y(_07635_));
 OAI21x1_ASAP7_75t_R _19877_ (.A1(_00468_),
    .A2(_07630_),
    .B(_00467_),
    .Y(_07636_));
 AND3x1_ASAP7_75t_R _19878_ (.A(_07624_),
    .B(_07635_),
    .C(_07636_),
    .Y(_04601_));
 OR3x1_ASAP7_75t_R _19879_ (.A(_00467_),
    .B(_00468_),
    .C(_07633_),
    .Y(_07637_));
 XOR2x2_ASAP7_75t_R _19880_ (.A(_00466_),
    .B(_07637_),
    .Y(_07638_));
 AND2x2_ASAP7_75t_R _19881_ (.A(_07541_),
    .B(_07638_),
    .Y(_04602_));
 OR4x1_ASAP7_75t_R _19882_ (.A(_00466_),
    .B(_00467_),
    .C(_00468_),
    .D(_07630_),
    .Y(_07639_));
 XOR2x2_ASAP7_75t_R _19883_ (.A(_00465_),
    .B(_07639_),
    .Y(_07640_));
 AND2x2_ASAP7_75t_R _19884_ (.A(_07541_),
    .B(_07640_),
    .Y(_04603_));
 OR4x1_ASAP7_75t_R _19885_ (.A(_00465_),
    .B(_00466_),
    .C(_00467_),
    .D(_00468_),
    .Y(_07641_));
 OR3x1_ASAP7_75t_R _19886_ (.A(_00464_),
    .B(_07633_),
    .C(_07641_),
    .Y(_07642_));
 OAI21x1_ASAP7_75t_R _19887_ (.A1(_07633_),
    .A2(_07641_),
    .B(_00464_),
    .Y(_07643_));
 AND3x1_ASAP7_75t_R _19888_ (.A(_07624_),
    .B(_07642_),
    .C(_07643_),
    .Y(_04604_));
 OR3x2_ASAP7_75t_R _19889_ (.A(_00463_),
    .B(_00464_),
    .C(_07641_),
    .Y(_07644_));
 OR3x1_ASAP7_75t_R _19890_ (.A(_00464_),
    .B(_07630_),
    .C(_07641_),
    .Y(_07645_));
 NAND2x1_ASAP7_75t_R _19891_ (.A(_00463_),
    .B(_07645_),
    .Y(_07646_));
 OA211x2_ASAP7_75t_R _19892_ (.A1(_07630_),
    .A2(_07644_),
    .B(_07646_),
    .C(_07260_),
    .Y(_04605_));
 OR3x2_ASAP7_75t_R _19893_ (.A(_00462_),
    .B(_07633_),
    .C(_07644_),
    .Y(_07647_));
 OAI21x1_ASAP7_75t_R _19894_ (.A1(_07633_),
    .A2(_07644_),
    .B(_00462_),
    .Y(_07648_));
 AND3x1_ASAP7_75t_R _19895_ (.A(_07624_),
    .B(_07647_),
    .C(_07648_),
    .Y(_04606_));
 OR3x2_ASAP7_75t_R _19896_ (.A(_00462_),
    .B(_07630_),
    .C(_07644_),
    .Y(_07649_));
 XOR2x2_ASAP7_75t_R _19897_ (.A(_00461_),
    .B(_07649_),
    .Y(_07650_));
 AND2x2_ASAP7_75t_R _19898_ (.A(_07541_),
    .B(_07650_),
    .Y(_04607_));
 NOR2x1_ASAP7_75t_R _19899_ (.A(_07190_),
    .B(_02622_),
    .Y(_04608_));
 OR3x1_ASAP7_75t_R _19900_ (.A(_00459_),
    .B(_00461_),
    .C(_07647_),
    .Y(_07651_));
 OAI21x1_ASAP7_75t_R _19901_ (.A1(_00461_),
    .A2(_07647_),
    .B(_00459_),
    .Y(_07652_));
 AND3x1_ASAP7_75t_R _19902_ (.A(_07624_),
    .B(_07651_),
    .C(_07652_),
    .Y(_04609_));
 OR3x1_ASAP7_75t_R _19903_ (.A(_00459_),
    .B(_00461_),
    .C(_07649_),
    .Y(_07653_));
 XOR2x2_ASAP7_75t_R _19904_ (.A(_00458_),
    .B(_07653_),
    .Y(_07654_));
 AND2x2_ASAP7_75t_R _19905_ (.A(_07541_),
    .B(_07654_),
    .Y(_04610_));
 OR4x1_ASAP7_75t_R _19906_ (.A(_00458_),
    .B(_00459_),
    .C(_00461_),
    .D(_07647_),
    .Y(_07655_));
 XOR2x2_ASAP7_75t_R _19907_ (.A(_00457_),
    .B(_07655_),
    .Y(_07656_));
 AND2x2_ASAP7_75t_R _19908_ (.A(_07541_),
    .B(_07656_),
    .Y(_04611_));
 OR4x1_ASAP7_75t_R _19909_ (.A(_00457_),
    .B(_00458_),
    .C(_00459_),
    .D(_00461_),
    .Y(_07657_));
 OR3x2_ASAP7_75t_R _19910_ (.A(_00456_),
    .B(_07649_),
    .C(_07657_),
    .Y(_07658_));
 OAI21x1_ASAP7_75t_R _19911_ (.A1(_07649_),
    .A2(_07657_),
    .B(_00456_),
    .Y(_07659_));
 AND3x1_ASAP7_75t_R _19912_ (.A(_07624_),
    .B(_07658_),
    .C(_07659_),
    .Y(_04612_));
 BUFx6f_ASAP7_75t_R _19913_ (.A(_07084_),
    .Y(_07660_));
 OR3x2_ASAP7_75t_R _19914_ (.A(_00456_),
    .B(_07647_),
    .C(_07657_),
    .Y(_07661_));
 XOR2x2_ASAP7_75t_R _19915_ (.A(_07615_),
    .B(_07661_),
    .Y(_07662_));
 AND2x2_ASAP7_75t_R _19916_ (.A(_07660_),
    .B(_07662_),
    .Y(_04613_));
 OR3x1_ASAP7_75t_R _19917_ (.A(_00454_),
    .B(_07615_),
    .C(_07658_),
    .Y(_07663_));
 OAI21x1_ASAP7_75t_R _19918_ (.A1(_07615_),
    .A2(_07658_),
    .B(_00454_),
    .Y(_07664_));
 AND3x1_ASAP7_75t_R _19919_ (.A(_07624_),
    .B(_07663_),
    .C(_07664_),
    .Y(_04614_));
 OR3x1_ASAP7_75t_R _19920_ (.A(_00454_),
    .B(_07615_),
    .C(_07661_),
    .Y(_07665_));
 XOR2x2_ASAP7_75t_R _19921_ (.A(_00453_),
    .B(_07665_),
    .Y(_07666_));
 AND2x2_ASAP7_75t_R _19922_ (.A(_07660_),
    .B(_07666_),
    .Y(_04615_));
 OR4x1_ASAP7_75t_R _19923_ (.A(_00453_),
    .B(_00454_),
    .C(_07615_),
    .D(_07658_),
    .Y(_07667_));
 XOR2x2_ASAP7_75t_R _19924_ (.A(_00452_),
    .B(_07667_),
    .Y(_07668_));
 AND2x2_ASAP7_75t_R _19925_ (.A(_07660_),
    .B(_07668_),
    .Y(_04616_));
 OR5x1_ASAP7_75t_R _19926_ (.A(_00452_),
    .B(_00453_),
    .C(_00454_),
    .D(_07615_),
    .E(_07661_),
    .Y(_07669_));
 XOR2x2_ASAP7_75t_R _19927_ (.A(_00451_),
    .B(_07669_),
    .Y(_07670_));
 AND2x2_ASAP7_75t_R _19928_ (.A(_07660_),
    .B(_07670_),
    .Y(_04617_));
 OR5x2_ASAP7_75t_R _19929_ (.A(_00451_),
    .B(_00452_),
    .C(_00453_),
    .D(_00454_),
    .E(_07615_),
    .Y(_07671_));
 OR3x1_ASAP7_75t_R _19930_ (.A(_00450_),
    .B(_07658_),
    .C(_07671_),
    .Y(_07672_));
 OAI21x1_ASAP7_75t_R _19931_ (.A1(_07658_),
    .A2(_07671_),
    .B(_00450_),
    .Y(_07673_));
 AND3x1_ASAP7_75t_R _19932_ (.A(_07624_),
    .B(_07672_),
    .C(_07673_),
    .Y(_04618_));
 XOR2x2_ASAP7_75t_R _19933_ (.A(_00449_),
    .B(_02621_),
    .Y(_07674_));
 AND2x2_ASAP7_75t_R _19934_ (.A(_07660_),
    .B(_07674_),
    .Y(_04619_));
 OR3x1_ASAP7_75t_R _19935_ (.A(_00450_),
    .B(_07661_),
    .C(_07671_),
    .Y(_07675_));
 XOR2x2_ASAP7_75t_R _19936_ (.A(_00448_),
    .B(_07675_),
    .Y(_07676_));
 AND2x2_ASAP7_75t_R _19937_ (.A(_07660_),
    .B(_07676_),
    .Y(_04620_));
 OR4x1_ASAP7_75t_R _19938_ (.A(_00448_),
    .B(_00450_),
    .C(_07658_),
    .D(_07671_),
    .Y(_07677_));
 XOR2x2_ASAP7_75t_R _19939_ (.A(_00447_),
    .B(_07677_),
    .Y(_07678_));
 AND2x2_ASAP7_75t_R _19940_ (.A(_07660_),
    .B(_07678_),
    .Y(_04621_));
 OR3x1_ASAP7_75t_R _19941_ (.A(_00449_),
    .B(_00460_),
    .C(_00055_),
    .Y(_07679_));
 XOR2x2_ASAP7_75t_R _19942_ (.A(_00446_),
    .B(_07679_),
    .Y(_07680_));
 AND2x2_ASAP7_75t_R _19943_ (.A(_07660_),
    .B(_07680_),
    .Y(_04622_));
 OR3x1_ASAP7_75t_R _19944_ (.A(_00446_),
    .B(_00449_),
    .C(_02621_),
    .Y(_07681_));
 NAND2x1_ASAP7_75t_R _19945_ (.A(_00445_),
    .B(_07681_),
    .Y(_07682_));
 AND3x1_ASAP7_75t_R _19946_ (.A(_07624_),
    .B(_07625_),
    .C(_07682_),
    .Y(_04623_));
 XOR2x2_ASAP7_75t_R _19947_ (.A(_07619_),
    .B(_07629_),
    .Y(_07683_));
 AND2x2_ASAP7_75t_R _19948_ (.A(_07660_),
    .B(_07683_),
    .Y(_04624_));
 BUFx6f_ASAP7_75t_R _19949_ (.A(_08998_),
    .Y(_07684_));
 OR3x1_ASAP7_75t_R _19950_ (.A(_00443_),
    .B(_07619_),
    .C(_07625_),
    .Y(_07685_));
 OAI21x1_ASAP7_75t_R _19951_ (.A1(_07619_),
    .A2(_07625_),
    .B(_00443_),
    .Y(_07686_));
 AND3x1_ASAP7_75t_R _19952_ (.A(_07684_),
    .B(_07685_),
    .C(_07686_),
    .Y(_04625_));
 OR3x1_ASAP7_75t_R _19953_ (.A(_00443_),
    .B(_07619_),
    .C(_07629_),
    .Y(_07687_));
 XOR2x2_ASAP7_75t_R _19954_ (.A(_00442_),
    .B(_07687_),
    .Y(_07688_));
 AND2x2_ASAP7_75t_R _19955_ (.A(_07660_),
    .B(_07688_),
    .Y(_04626_));
 BUFx12f_ASAP7_75t_R _19956_ (.A(_08527_),
    .Y(_07689_));
 BUFx6f_ASAP7_75t_R _19957_ (.A(_07689_),
    .Y(_07690_));
 OR4x1_ASAP7_75t_R _19958_ (.A(_00442_),
    .B(_00443_),
    .C(_07619_),
    .D(_07625_),
    .Y(_07691_));
 XOR2x2_ASAP7_75t_R _19959_ (.A(_00441_),
    .B(_07691_),
    .Y(_07692_));
 AND2x2_ASAP7_75t_R _19960_ (.A(_07690_),
    .B(_07692_),
    .Y(_04627_));
 OR5x1_ASAP7_75t_R _19961_ (.A(_00441_),
    .B(_00442_),
    .C(_00443_),
    .D(_07619_),
    .E(_07629_),
    .Y(_07693_));
 NAND2x1_ASAP7_75t_R _19962_ (.A(_00440_),
    .B(_07693_),
    .Y(_07694_));
 OA211x2_ASAP7_75t_R _19963_ (.A1(_07626_),
    .A2(_07629_),
    .B(_07694_),
    .C(_07260_),
    .Y(_04628_));
 AND4x1_ASAP7_75t_R _19964_ (.A(_00401_),
    .B(_00429_),
    .C(_00430_),
    .D(_00431_),
    .Y(_07695_));
 AND5x1_ASAP7_75t_R _19965_ (.A(_00420_),
    .B(_00425_),
    .C(_00426_),
    .D(_00428_),
    .E(_07695_),
    .Y(_07696_));
 AND5x1_ASAP7_75t_R _19966_ (.A(_00422_),
    .B(_00423_),
    .C(_00424_),
    .D(_07147_),
    .E(_07696_),
    .Y(_07697_));
 BUFx3_ASAP7_75t_R _19967_ (.A(_00417_),
    .Y(_07698_));
 AND4x1_ASAP7_75t_R _19968_ (.A(_00415_),
    .B(_00416_),
    .C(_07698_),
    .D(_00418_),
    .Y(_07699_));
 BUFx6f_ASAP7_75t_R _19969_ (.A(_00427_),
    .Y(_07700_));
 AND4x1_ASAP7_75t_R _19970_ (.A(_00409_),
    .B(_00411_),
    .C(_00412_),
    .D(_00419_),
    .Y(_07701_));
 AND5x1_ASAP7_75t_R _19971_ (.A(_00402_),
    .B(_00403_),
    .C(_00408_),
    .D(_07700_),
    .E(_07701_),
    .Y(_07702_));
 BUFx3_ASAP7_75t_R _19972_ (.A(_00405_),
    .Y(_07703_));
 AND3x1_ASAP7_75t_R _19973_ (.A(_00406_),
    .B(_00407_),
    .C(_00410_),
    .Y(_07704_));
 OR3x1_ASAP7_75t_R _19974_ (.A(_00404_),
    .B(_07703_),
    .C(_07704_),
    .Y(_07705_));
 AND5x2_ASAP7_75t_R _19975_ (.A(_00413_),
    .B(_00414_),
    .C(_07699_),
    .D(_07702_),
    .E(_07705_),
    .Y(_07706_));
 NAND2x2_ASAP7_75t_R _19976_ (.A(_07697_),
    .B(_07706_),
    .Y(_07707_));
 NOR2x1_ASAP7_75t_R _19977_ (.A(_00391_),
    .B(_07707_),
    .Y(_04629_));
 INVx1_ASAP7_75t_R _19978_ (.A(_07707_),
    .Y(_04630_));
 NOR2x1_ASAP7_75t_R _19979_ (.A(_00394_),
    .B(_07707_),
    .Y(_04631_));
 NOR2x1_ASAP7_75t_R _19980_ (.A(_00393_),
    .B(_07707_),
    .Y(_04632_));
 NOR2x1_ASAP7_75t_R _19981_ (.A(_00392_),
    .B(_07707_),
    .Y(_04633_));
 NOR2x1_ASAP7_75t_R _19982_ (.A(_00390_),
    .B(_07707_),
    .Y(_04634_));
 NOR2x1_ASAP7_75t_R _19983_ (.A(_00389_),
    .B(_07707_),
    .Y(_04635_));
 INVx1_ASAP7_75t_R _19984_ (.A(_07707_),
    .Y(_04636_));
 AND2x2_ASAP7_75t_R _19985_ (.A(_07690_),
    .B(_00056_),
    .Y(_04637_));
 OR4x1_ASAP7_75t_R _19986_ (.A(_00406_),
    .B(_00407_),
    .C(_00410_),
    .D(_02639_),
    .Y(_07708_));
 OR5x2_ASAP7_75t_R _19987_ (.A(_00401_),
    .B(_00402_),
    .C(_00403_),
    .D(_00404_),
    .E(_07703_),
    .Y(_07709_));
 OR2x2_ASAP7_75t_R _19988_ (.A(_07708_),
    .B(_07709_),
    .Y(_07710_));
 XNOR2x2_ASAP7_75t_R _19989_ (.A(_00431_),
    .B(_07710_),
    .Y(_07711_));
 NOR2x1_ASAP7_75t_R _19990_ (.A(_07190_),
    .B(_07711_),
    .Y(_04638_));
 OR5x2_ASAP7_75t_R _19991_ (.A(_00406_),
    .B(_00407_),
    .C(_00410_),
    .D(_00421_),
    .E(_00056_),
    .Y(_07712_));
 OR3x1_ASAP7_75t_R _19992_ (.A(_00431_),
    .B(_07709_),
    .C(_07712_),
    .Y(_07713_));
 XOR2x2_ASAP7_75t_R _19993_ (.A(_00430_),
    .B(_07713_),
    .Y(_07714_));
 AND2x2_ASAP7_75t_R _19994_ (.A(_07690_),
    .B(_07714_),
    .Y(_04639_));
 OR3x1_ASAP7_75t_R _19995_ (.A(_00430_),
    .B(_00431_),
    .C(_07710_),
    .Y(_07715_));
 XOR2x2_ASAP7_75t_R _19996_ (.A(_00429_),
    .B(_07715_),
    .Y(_07716_));
 AND2x2_ASAP7_75t_R _19997_ (.A(_07690_),
    .B(_07716_),
    .Y(_04640_));
 OR3x1_ASAP7_75t_R _19998_ (.A(_00428_),
    .B(_00429_),
    .C(_00430_),
    .Y(_07717_));
 OR4x1_ASAP7_75t_R _19999_ (.A(_00431_),
    .B(_07709_),
    .C(_07712_),
    .D(_07717_),
    .Y(_07718_));
 OR3x1_ASAP7_75t_R _20000_ (.A(_00429_),
    .B(_00430_),
    .C(_07713_),
    .Y(_07719_));
 NAND2x1_ASAP7_75t_R _20001_ (.A(_00428_),
    .B(_07719_),
    .Y(_07720_));
 AND3x1_ASAP7_75t_R _20002_ (.A(_07684_),
    .B(_07718_),
    .C(_07720_),
    .Y(_04641_));
 OR4x1_ASAP7_75t_R _20003_ (.A(_00431_),
    .B(_07708_),
    .C(_07709_),
    .D(_07717_),
    .Y(_07721_));
 XOR2x2_ASAP7_75t_R _20004_ (.A(_07700_),
    .B(_07721_),
    .Y(_07722_));
 AND2x2_ASAP7_75t_R _20005_ (.A(_07690_),
    .B(_07722_),
    .Y(_04642_));
 OR3x1_ASAP7_75t_R _20006_ (.A(_00426_),
    .B(_07700_),
    .C(_07718_),
    .Y(_07723_));
 OAI21x1_ASAP7_75t_R _20007_ (.A1(_07700_),
    .A2(_07718_),
    .B(_00426_),
    .Y(_07724_));
 AND3x1_ASAP7_75t_R _20008_ (.A(_07684_),
    .B(_07723_),
    .C(_07724_),
    .Y(_04643_));
 OR3x1_ASAP7_75t_R _20009_ (.A(_00426_),
    .B(_07700_),
    .C(_07721_),
    .Y(_07725_));
 XOR2x2_ASAP7_75t_R _20010_ (.A(_00425_),
    .B(_07725_),
    .Y(_07726_));
 AND2x2_ASAP7_75t_R _20011_ (.A(_07690_),
    .B(_07726_),
    .Y(_04644_));
 OR5x2_ASAP7_75t_R _20012_ (.A(_00424_),
    .B(_00425_),
    .C(_00426_),
    .D(_07700_),
    .E(_07718_),
    .Y(_07727_));
 OR4x1_ASAP7_75t_R _20013_ (.A(_00425_),
    .B(_00426_),
    .C(_07700_),
    .D(_07718_),
    .Y(_07728_));
 NAND2x1_ASAP7_75t_R _20014_ (.A(_00424_),
    .B(_07728_),
    .Y(_07729_));
 AND3x1_ASAP7_75t_R _20015_ (.A(_07684_),
    .B(_07727_),
    .C(_07729_),
    .Y(_04645_));
 OR5x2_ASAP7_75t_R _20016_ (.A(_00424_),
    .B(_00425_),
    .C(_00426_),
    .D(_07700_),
    .E(_07721_),
    .Y(_07730_));
 XOR2x2_ASAP7_75t_R _20017_ (.A(_00423_),
    .B(_07730_),
    .Y(_07731_));
 AND2x2_ASAP7_75t_R _20018_ (.A(_07690_),
    .B(_07731_),
    .Y(_04646_));
 OR3x1_ASAP7_75t_R _20019_ (.A(_00422_),
    .B(_00423_),
    .C(_07727_),
    .Y(_07732_));
 OAI21x1_ASAP7_75t_R _20020_ (.A1(_00423_),
    .A2(_07727_),
    .B(_00422_),
    .Y(_07733_));
 AND3x1_ASAP7_75t_R _20021_ (.A(_07684_),
    .B(_07732_),
    .C(_07733_),
    .Y(_04647_));
 NOR2x1_ASAP7_75t_R _20022_ (.A(_07190_),
    .B(_02640_),
    .Y(_04648_));
 OR3x1_ASAP7_75t_R _20023_ (.A(_00422_),
    .B(_00423_),
    .C(_07730_),
    .Y(_07734_));
 XOR2x2_ASAP7_75t_R _20024_ (.A(_00420_),
    .B(_07734_),
    .Y(_07735_));
 AND2x2_ASAP7_75t_R _20025_ (.A(_07690_),
    .B(_07735_),
    .Y(_04649_));
 OR4x1_ASAP7_75t_R _20026_ (.A(_00420_),
    .B(_00422_),
    .C(_00423_),
    .D(_07727_),
    .Y(_07736_));
 XOR2x2_ASAP7_75t_R _20027_ (.A(_00419_),
    .B(_07736_),
    .Y(_07737_));
 AND2x2_ASAP7_75t_R _20028_ (.A(_07690_),
    .B(_07737_),
    .Y(_04650_));
 OR4x1_ASAP7_75t_R _20029_ (.A(_00419_),
    .B(_00420_),
    .C(_00422_),
    .D(_00423_),
    .Y(_07738_));
 OR3x2_ASAP7_75t_R _20030_ (.A(_00418_),
    .B(_07730_),
    .C(_07738_),
    .Y(_07739_));
 OAI21x1_ASAP7_75t_R _20031_ (.A1(_07730_),
    .A2(_07738_),
    .B(_00418_),
    .Y(_07740_));
 AND3x1_ASAP7_75t_R _20032_ (.A(_07684_),
    .B(_07739_),
    .C(_07740_),
    .Y(_04651_));
 OR3x2_ASAP7_75t_R _20033_ (.A(_00418_),
    .B(_07727_),
    .C(_07738_),
    .Y(_07741_));
 XOR2x2_ASAP7_75t_R _20034_ (.A(_07698_),
    .B(_07741_),
    .Y(_07742_));
 AND2x2_ASAP7_75t_R _20035_ (.A(_07690_),
    .B(_07742_),
    .Y(_04652_));
 OR3x1_ASAP7_75t_R _20036_ (.A(_00416_),
    .B(_07698_),
    .C(_07739_),
    .Y(_07743_));
 OAI21x1_ASAP7_75t_R _20037_ (.A1(_07698_),
    .A2(_07739_),
    .B(_00416_),
    .Y(_07744_));
 AND3x1_ASAP7_75t_R _20038_ (.A(_07684_),
    .B(_07743_),
    .C(_07744_),
    .Y(_04653_));
 BUFx6f_ASAP7_75t_R _20039_ (.A(_07689_),
    .Y(_07745_));
 OR3x1_ASAP7_75t_R _20040_ (.A(_00416_),
    .B(_07698_),
    .C(_07741_),
    .Y(_07746_));
 XOR2x2_ASAP7_75t_R _20041_ (.A(_00415_),
    .B(_07746_),
    .Y(_07747_));
 AND2x2_ASAP7_75t_R _20042_ (.A(_07745_),
    .B(_07747_),
    .Y(_04654_));
 OR4x1_ASAP7_75t_R _20043_ (.A(_00415_),
    .B(_00416_),
    .C(_07698_),
    .D(_07739_),
    .Y(_07748_));
 XOR2x2_ASAP7_75t_R _20044_ (.A(_00414_),
    .B(_07748_),
    .Y(_07749_));
 AND2x2_ASAP7_75t_R _20045_ (.A(_07745_),
    .B(_07749_),
    .Y(_04655_));
 OR5x1_ASAP7_75t_R _20046_ (.A(_00414_),
    .B(_00415_),
    .C(_00416_),
    .D(_07698_),
    .E(_07741_),
    .Y(_07750_));
 XOR2x2_ASAP7_75t_R _20047_ (.A(_00413_),
    .B(_07750_),
    .Y(_07751_));
 AND2x2_ASAP7_75t_R _20048_ (.A(_07745_),
    .B(_07751_),
    .Y(_04656_));
 OR5x2_ASAP7_75t_R _20049_ (.A(_00413_),
    .B(_00414_),
    .C(_00415_),
    .D(_00416_),
    .E(_07698_),
    .Y(_07752_));
 OR3x1_ASAP7_75t_R _20050_ (.A(_00412_),
    .B(_07739_),
    .C(_07752_),
    .Y(_07753_));
 OAI21x1_ASAP7_75t_R _20051_ (.A1(_07739_),
    .A2(_07752_),
    .B(_00412_),
    .Y(_07754_));
 AND3x1_ASAP7_75t_R _20052_ (.A(_07684_),
    .B(_07753_),
    .C(_07754_),
    .Y(_04657_));
 OR3x1_ASAP7_75t_R _20053_ (.A(_00412_),
    .B(_07741_),
    .C(_07752_),
    .Y(_07755_));
 XOR2x2_ASAP7_75t_R _20054_ (.A(_00411_),
    .B(_07755_),
    .Y(_07756_));
 AND2x2_ASAP7_75t_R _20055_ (.A(_07745_),
    .B(_07756_),
    .Y(_04658_));
 XOR2x2_ASAP7_75t_R _20056_ (.A(_00410_),
    .B(_02639_),
    .Y(_07757_));
 AND2x2_ASAP7_75t_R _20057_ (.A(_07745_),
    .B(_07757_),
    .Y(_04659_));
 OR4x1_ASAP7_75t_R _20058_ (.A(_00411_),
    .B(_00412_),
    .C(_07739_),
    .D(_07752_),
    .Y(_07758_));
 XOR2x2_ASAP7_75t_R _20059_ (.A(_00409_),
    .B(_07758_),
    .Y(_07759_));
 AND2x2_ASAP7_75t_R _20060_ (.A(_07745_),
    .B(_07759_),
    .Y(_04660_));
 OR5x1_ASAP7_75t_R _20061_ (.A(_00409_),
    .B(_00411_),
    .C(_00412_),
    .D(_07741_),
    .E(_07752_),
    .Y(_07760_));
 XOR2x2_ASAP7_75t_R _20062_ (.A(_00408_),
    .B(_07760_),
    .Y(_07761_));
 AND2x2_ASAP7_75t_R _20063_ (.A(_07745_),
    .B(_07761_),
    .Y(_04661_));
 OR3x1_ASAP7_75t_R _20064_ (.A(_00410_),
    .B(_00421_),
    .C(_00056_),
    .Y(_07762_));
 XOR2x2_ASAP7_75t_R _20065_ (.A(_00407_),
    .B(_07762_),
    .Y(_07763_));
 AND2x2_ASAP7_75t_R _20066_ (.A(_07745_),
    .B(_07763_),
    .Y(_04662_));
 OR3x1_ASAP7_75t_R _20067_ (.A(_00407_),
    .B(_00410_),
    .C(_02639_),
    .Y(_07764_));
 NAND2x1_ASAP7_75t_R _20068_ (.A(_00406_),
    .B(_07764_),
    .Y(_07765_));
 AND3x1_ASAP7_75t_R _20069_ (.A(_07684_),
    .B(_07708_),
    .C(_07765_),
    .Y(_04663_));
 XOR2x2_ASAP7_75t_R _20070_ (.A(_07703_),
    .B(_07712_),
    .Y(_07766_));
 AND2x2_ASAP7_75t_R _20071_ (.A(_07745_),
    .B(_07766_),
    .Y(_04664_));
 OR3x1_ASAP7_75t_R _20072_ (.A(_00404_),
    .B(_07703_),
    .C(_07708_),
    .Y(_07767_));
 OAI21x1_ASAP7_75t_R _20073_ (.A1(_07703_),
    .A2(_07708_),
    .B(_00404_),
    .Y(_07768_));
 AND3x1_ASAP7_75t_R _20074_ (.A(_07684_),
    .B(_07767_),
    .C(_07768_),
    .Y(_04665_));
 OR3x1_ASAP7_75t_R _20075_ (.A(_00404_),
    .B(_07703_),
    .C(_07712_),
    .Y(_07769_));
 XOR2x2_ASAP7_75t_R _20076_ (.A(_00403_),
    .B(_07769_),
    .Y(_07770_));
 AND2x2_ASAP7_75t_R _20077_ (.A(_07745_),
    .B(_07770_),
    .Y(_04666_));
 BUFx6f_ASAP7_75t_R _20078_ (.A(_07689_),
    .Y(_07771_));
 OR4x1_ASAP7_75t_R _20079_ (.A(_00403_),
    .B(_00404_),
    .C(_07703_),
    .D(_07708_),
    .Y(_07772_));
 XOR2x2_ASAP7_75t_R _20080_ (.A(_00402_),
    .B(_07772_),
    .Y(_07773_));
 AND2x2_ASAP7_75t_R _20081_ (.A(_07771_),
    .B(_07773_),
    .Y(_04667_));
 OR5x1_ASAP7_75t_R _20082_ (.A(_00402_),
    .B(_00403_),
    .C(_00404_),
    .D(_07703_),
    .E(_07712_),
    .Y(_07774_));
 XOR2x2_ASAP7_75t_R _20083_ (.A(_00401_),
    .B(_07774_),
    .Y(_07775_));
 AND2x2_ASAP7_75t_R _20084_ (.A(_07771_),
    .B(_07775_),
    .Y(_04668_));
 AND2x2_ASAP7_75t_R _20085_ (.A(_07771_),
    .B(_00027_),
    .Y(_04669_));
 INVx2_ASAP7_75t_R _20086_ (.A(_02205_),
    .Y(_07776_));
 AND4x1_ASAP7_75t_R _20087_ (.A(_00433_),
    .B(\xs[6].cli1.i[35] ),
    .C(\xs[6].cli1.i[34] ),
    .D(_00436_),
    .Y(_07777_));
 AND3x1_ASAP7_75t_R _20088_ (.A(\xs[6].cli1.i[39] ),
    .B(_00437_),
    .C(_07777_),
    .Y(_07778_));
 INVx1_ASAP7_75t_R _20089_ (.A(_02211_),
    .Y(_07779_));
 OA21x2_ASAP7_75t_R _20090_ (.A1(_00432_),
    .A2(_07777_),
    .B(_07779_),
    .Y(_07780_));
 NOR2x1_ASAP7_75t_R _20091_ (.A(_00473_),
    .B(_00474_),
    .Y(_07781_));
 AND2x2_ASAP7_75t_R _20092_ (.A(_00472_),
    .B(_00475_),
    .Y(_07782_));
 AO21x1_ASAP7_75t_R _20093_ (.A1(_07781_),
    .A2(_07782_),
    .B(_00471_),
    .Y(_07783_));
 AO21x1_ASAP7_75t_R _20094_ (.A1(\peo[12][39] ),
    .A2(\peo[12][32] ),
    .B(_02211_),
    .Y(_07784_));
 OA211x2_ASAP7_75t_R _20095_ (.A1(_07778_),
    .A2(_07780_),
    .B(_07783_),
    .C(_07784_),
    .Y(_07785_));
 NOR2x1_ASAP7_75t_R _20096_ (.A(_07776_),
    .B(_07785_),
    .Y(_07786_));
 BUFx6f_ASAP7_75t_R _20097_ (.A(_02204_),
    .Y(_07787_));
 INVx2_ASAP7_75t_R _20098_ (.A(_07787_),
    .Y(_07788_));
 AND2x2_ASAP7_75t_R _20099_ (.A(_07788_),
    .B(_02211_),
    .Y(_07789_));
 NOR2x2_ASAP7_75t_R _20100_ (.A(_00432_),
    .B(_07777_),
    .Y(_07790_));
 AO21x1_ASAP7_75t_R _20101_ (.A1(_00027_),
    .A2(_07790_),
    .B(_07788_),
    .Y(_07791_));
 AOI21x1_ASAP7_75t_R _20102_ (.A1(_07781_),
    .A2(_07782_),
    .B(_00471_),
    .Y(_07792_));
 OR3x1_ASAP7_75t_R _20103_ (.A(_07787_),
    .B(_07776_),
    .C(_02211_),
    .Y(_07793_));
 AND2x2_ASAP7_75t_R _20104_ (.A(_07792_),
    .B(_07793_),
    .Y(_07794_));
 INVx1_ASAP7_75t_R _20105_ (.A(_07778_),
    .Y(_07795_));
 AO21x1_ASAP7_75t_R _20106_ (.A1(_07791_),
    .A2(_07794_),
    .B(_07795_),
    .Y(_07796_));
 AOI22x1_ASAP7_75t_R _20107_ (.A1(_07786_),
    .A2(_07789_),
    .B1(_07796_),
    .B2(_00478_),
    .Y(_07797_));
 AO21x1_ASAP7_75t_R _20108_ (.A1(_07792_),
    .A2(_07778_),
    .B(_07790_),
    .Y(_07798_));
 AOI21x1_ASAP7_75t_R _20109_ (.A1(\xs[6].cli1.i[32] ),
    .A2(_07777_),
    .B(_00432_),
    .Y(_07799_));
 AO32x2_ASAP7_75t_R _20110_ (.A1(_07787_),
    .A2(_00027_),
    .A3(_07790_),
    .B1(_07789_),
    .B2(_07799_),
    .Y(_07800_));
 AO32x2_ASAP7_75t_R _20111_ (.A1(_07788_),
    .A2(_07776_),
    .A3(_07798_),
    .B1(_07800_),
    .B2(_07792_),
    .Y(_07801_));
 OR3x1_ASAP7_75t_R _20112_ (.A(\peo[13][0] ),
    .B(_07795_),
    .C(_07801_),
    .Y(_07802_));
 INVx1_ASAP7_75t_R _20113_ (.A(_02215_),
    .Y(_07803_));
 NOR2x2_ASAP7_75t_R _20114_ (.A(_08571_),
    .B(_07787_),
    .Y(_07804_));
 AND3x1_ASAP7_75t_R _20115_ (.A(_02211_),
    .B(_07786_),
    .C(_07804_),
    .Y(_07805_));
 AO32x1_ASAP7_75t_R _20116_ (.A1(_09830_),
    .A2(_07797_),
    .A3(_07802_),
    .B1(_07803_),
    .B2(_07805_),
    .Y(_04670_));
 OR2x6_ASAP7_75t_R _20117_ (.A(_07776_),
    .B(_07785_),
    .Y(_07806_));
 OR4x1_ASAP7_75t_R _20118_ (.A(_11177_),
    .B(_07787_),
    .C(_07779_),
    .D(_07806_),
    .Y(_07807_));
 NOR2x1_ASAP7_75t_R _20119_ (.A(_02214_),
    .B(_07807_),
    .Y(_04671_));
 NOR2x1_ASAP7_75t_R _20120_ (.A(_02213_),
    .B(_07807_),
    .Y(_04672_));
 NOR2x1_ASAP7_75t_R _20121_ (.A(_02212_),
    .B(_07807_),
    .Y(_04673_));
 NOR2x1_ASAP7_75t_R _20122_ (.A(_02203_),
    .B(_07807_),
    .Y(_04674_));
 NOR2x1_ASAP7_75t_R _20123_ (.A(_02202_),
    .B(_07807_),
    .Y(_04675_));
 BUFx6f_ASAP7_75t_R _20124_ (.A(_08998_),
    .Y(_07808_));
 OAI21x1_ASAP7_75t_R _20125_ (.A1(_07785_),
    .A2(_07793_),
    .B(_00478_),
    .Y(_07809_));
 OR3x1_ASAP7_75t_R _20126_ (.A(_07803_),
    .B(_07785_),
    .C(_07793_),
    .Y(_07810_));
 AO21x1_ASAP7_75t_R _20127_ (.A1(_07809_),
    .A2(_07810_),
    .B(_07801_),
    .Y(_07811_));
 NAND2x1_ASAP7_75t_R _20128_ (.A(_00439_),
    .B(_07801_),
    .Y(_07812_));
 AND3x1_ASAP7_75t_R _20129_ (.A(_07808_),
    .B(_07811_),
    .C(_07812_),
    .Y(_04676_));
 OR4x1_ASAP7_75t_R _20130_ (.A(_11177_),
    .B(_07787_),
    .C(_02211_),
    .D(_07806_),
    .Y(_07813_));
 NOR2x1_ASAP7_75t_R _20131_ (.A(_02214_),
    .B(_07813_),
    .Y(_04677_));
 NOR2x1_ASAP7_75t_R _20132_ (.A(_02213_),
    .B(_07813_),
    .Y(_04678_));
 NOR2x1_ASAP7_75t_R _20133_ (.A(_02212_),
    .B(_07813_),
    .Y(_04679_));
 NOR2x1_ASAP7_75t_R _20134_ (.A(_02203_),
    .B(_07813_),
    .Y(_04680_));
 NOR2x1_ASAP7_75t_R _20135_ (.A(_02202_),
    .B(_07813_),
    .Y(_04681_));
 OA21x2_ASAP7_75t_R _20136_ (.A1(_07787_),
    .A2(_07786_),
    .B(_08584_),
    .Y(_07814_));
 OAI21x1_ASAP7_75t_R _20137_ (.A1(_07787_),
    .A2(_02205_),
    .B(_07790_),
    .Y(_07815_));
 AOI21x1_ASAP7_75t_R _20138_ (.A1(_07792_),
    .A2(_07800_),
    .B(_07815_),
    .Y(_07816_));
 NAND2x1_ASAP7_75t_R _20139_ (.A(_00439_),
    .B(_07816_),
    .Y(_07817_));
 AO21x2_ASAP7_75t_R _20140_ (.A1(_07792_),
    .A2(_07800_),
    .B(_07815_),
    .Y(_07818_));
 NAND2x1_ASAP7_75t_R _20141_ (.A(_00478_),
    .B(_07818_),
    .Y(_07819_));
 AND2x4_ASAP7_75t_R _20142_ (.A(_07806_),
    .B(_07804_),
    .Y(_07820_));
 AO32x1_ASAP7_75t_R _20143_ (.A1(_07814_),
    .A2(_07817_),
    .A3(_07819_),
    .B1(_07820_),
    .B2(_07803_),
    .Y(_04682_));
 NAND2x2_ASAP7_75t_R _20144_ (.A(_07806_),
    .B(_07804_),
    .Y(_07821_));
 NOR2x1_ASAP7_75t_R _20145_ (.A(_02214_),
    .B(_07821_),
    .Y(_04683_));
 NOR2x1_ASAP7_75t_R _20146_ (.A(_02213_),
    .B(_07821_),
    .Y(_04684_));
 NOR2x1_ASAP7_75t_R _20147_ (.A(_02212_),
    .B(_07821_),
    .Y(_04685_));
 NAND2x1_ASAP7_75t_R _20148_ (.A(_00437_),
    .B(_07816_),
    .Y(_07822_));
 NAND2x1_ASAP7_75t_R _20149_ (.A(_00476_),
    .B(_07818_),
    .Y(_07823_));
 AO32x1_ASAP7_75t_R _20150_ (.A1(_07814_),
    .A2(_07822_),
    .A3(_07823_),
    .B1(_07820_),
    .B2(_07779_),
    .Y(_04686_));
 NAND2x1_ASAP7_75t_R _20151_ (.A(_00436_),
    .B(_07816_),
    .Y(_07824_));
 NAND2x1_ASAP7_75t_R _20152_ (.A(_00475_),
    .B(_07818_),
    .Y(_07825_));
 INVx1_ASAP7_75t_R _20153_ (.A(_02210_),
    .Y(_07826_));
 AO32x1_ASAP7_75t_R _20154_ (.A1(_07814_),
    .A2(_07824_),
    .A3(_07825_),
    .B1(_07820_),
    .B2(_07826_),
    .Y(_04687_));
 AO21x1_ASAP7_75t_R _20155_ (.A1(\peo[12][39] ),
    .A2(_07800_),
    .B(_07815_),
    .Y(_07827_));
 NAND2x1_ASAP7_75t_R _20156_ (.A(_00474_),
    .B(_07827_),
    .Y(_07828_));
 OR3x1_ASAP7_75t_R _20157_ (.A(_00432_),
    .B(\xs[6].cli1.i[34] ),
    .C(_07801_),
    .Y(_07829_));
 INVx1_ASAP7_75t_R _20158_ (.A(_02209_),
    .Y(_07830_));
 AO32x1_ASAP7_75t_R _20159_ (.A1(_07814_),
    .A2(_07828_),
    .A3(_07829_),
    .B1(_07820_),
    .B2(_07830_),
    .Y(_04688_));
 NAND2x1_ASAP7_75t_R _20160_ (.A(_00473_),
    .B(_07827_),
    .Y(_07831_));
 OR3x1_ASAP7_75t_R _20161_ (.A(_00432_),
    .B(\xs[6].cli1.i[35] ),
    .C(_07801_),
    .Y(_07832_));
 INVx1_ASAP7_75t_R _20162_ (.A(_02208_),
    .Y(_07833_));
 AO32x1_ASAP7_75t_R _20163_ (.A1(_07814_),
    .A2(_07831_),
    .A3(_07832_),
    .B1(_07820_),
    .B2(_07833_),
    .Y(_04689_));
 NAND2x1_ASAP7_75t_R _20164_ (.A(_00433_),
    .B(_07816_),
    .Y(_07834_));
 NAND2x1_ASAP7_75t_R _20165_ (.A(_00472_),
    .B(_07818_),
    .Y(_07835_));
 INVx1_ASAP7_75t_R _20166_ (.A(_02207_),
    .Y(_07836_));
 AO32x1_ASAP7_75t_R _20167_ (.A1(_07814_),
    .A2(_07834_),
    .A3(_07835_),
    .B1(_07820_),
    .B2(_07836_),
    .Y(_04690_));
 NOR2x1_ASAP7_75t_R _20168_ (.A(_02206_),
    .B(_07821_),
    .Y(_04691_));
 AND3x1_ASAP7_75t_R _20169_ (.A(_02205_),
    .B(_07785_),
    .C(_07804_),
    .Y(_04692_));
 AOI211x1_ASAP7_75t_R _20170_ (.A1(_07788_),
    .A2(_07806_),
    .B(_07790_),
    .C(_07792_),
    .Y(_07837_));
 NOR2x1_ASAP7_75t_R _20171_ (.A(_07190_),
    .B(_07837_),
    .Y(_04693_));
 NOR2x1_ASAP7_75t_R _20172_ (.A(_02203_),
    .B(_07821_),
    .Y(_04694_));
 NOR2x1_ASAP7_75t_R _20173_ (.A(_02202_),
    .B(_07821_),
    .Y(_04695_));
 BUFx3_ASAP7_75t_R _20174_ (.A(_00361_),
    .Y(_07838_));
 AND4x1_ASAP7_75t_R _20175_ (.A(_00336_),
    .B(_00364_),
    .C(_00365_),
    .D(_00366_),
    .Y(_07839_));
 AND5x1_ASAP7_75t_R _20176_ (.A(_00355_),
    .B(_00360_),
    .C(_07838_),
    .D(_00363_),
    .E(_07839_),
    .Y(_07840_));
 AND5x1_ASAP7_75t_R _20177_ (.A(_00357_),
    .B(_00358_),
    .C(_00359_),
    .D(_07147_),
    .E(_07840_),
    .Y(_07841_));
 BUFx3_ASAP7_75t_R _20178_ (.A(_00352_),
    .Y(_07842_));
 AND4x1_ASAP7_75t_R _20179_ (.A(_00350_),
    .B(_00351_),
    .C(_07842_),
    .D(_00353_),
    .Y(_07843_));
 AND4x1_ASAP7_75t_R _20180_ (.A(_00344_),
    .B(_00346_),
    .C(_00347_),
    .D(_00354_),
    .Y(_07844_));
 AND5x1_ASAP7_75t_R _20181_ (.A(_00337_),
    .B(_00338_),
    .C(_00343_),
    .D(_00362_),
    .E(_07844_),
    .Y(_07845_));
 AND3x1_ASAP7_75t_R _20182_ (.A(_00341_),
    .B(_00342_),
    .C(_00345_),
    .Y(_07846_));
 OR3x1_ASAP7_75t_R _20183_ (.A(_00339_),
    .B(_00340_),
    .C(_07846_),
    .Y(_07847_));
 AND5x2_ASAP7_75t_R _20184_ (.A(_00348_),
    .B(_00349_),
    .C(_07843_),
    .D(_07845_),
    .E(_07847_),
    .Y(_07848_));
 NAND2x2_ASAP7_75t_R _20185_ (.A(_07841_),
    .B(_07848_),
    .Y(_07849_));
 NOR2x1_ASAP7_75t_R _20186_ (.A(_00293_),
    .B(_07849_),
    .Y(_04696_));
 INVx1_ASAP7_75t_R _20187_ (.A(_07849_),
    .Y(_04697_));
 NOR2x1_ASAP7_75t_R _20188_ (.A(_00296_),
    .B(_07849_),
    .Y(_04698_));
 NOR2x1_ASAP7_75t_R _20189_ (.A(_00295_),
    .B(_07849_),
    .Y(_04699_));
 NOR2x1_ASAP7_75t_R _20190_ (.A(_00294_),
    .B(_07849_),
    .Y(_04700_));
 NOR2x1_ASAP7_75t_R _20191_ (.A(_00292_),
    .B(_07849_),
    .Y(_04701_));
 NOR2x1_ASAP7_75t_R _20192_ (.A(_00291_),
    .B(_07849_),
    .Y(_04702_));
 INVx1_ASAP7_75t_R _20193_ (.A(_07849_),
    .Y(_04703_));
 AND2x2_ASAP7_75t_R _20194_ (.A(_07771_),
    .B(_00057_),
    .Y(_04704_));
 OR3x1_ASAP7_75t_R _20195_ (.A(_00342_),
    .B(_00345_),
    .C(_02651_),
    .Y(_07850_));
 OR2x2_ASAP7_75t_R _20196_ (.A(_00341_),
    .B(_07850_),
    .Y(_07851_));
 BUFx3_ASAP7_75t_R _20197_ (.A(_07851_),
    .Y(_07852_));
 OR4x1_ASAP7_75t_R _20198_ (.A(_00337_),
    .B(_00338_),
    .C(_00339_),
    .D(_00340_),
    .Y(_07853_));
 OR3x1_ASAP7_75t_R _20199_ (.A(_00336_),
    .B(_07852_),
    .C(_07853_),
    .Y(_07854_));
 XOR2x2_ASAP7_75t_R _20200_ (.A(_00366_),
    .B(_07854_),
    .Y(_07855_));
 AND2x2_ASAP7_75t_R _20201_ (.A(_07771_),
    .B(_07855_),
    .Y(_04705_));
 OR3x1_ASAP7_75t_R _20202_ (.A(_00345_),
    .B(_00356_),
    .C(_00057_),
    .Y(_07856_));
 OR3x1_ASAP7_75t_R _20203_ (.A(_00341_),
    .B(_00342_),
    .C(_07856_),
    .Y(_07857_));
 BUFx6f_ASAP7_75t_R _20204_ (.A(_07857_),
    .Y(_07858_));
 OR4x1_ASAP7_75t_R _20205_ (.A(_00336_),
    .B(_00366_),
    .C(_07853_),
    .D(_07858_),
    .Y(_07859_));
 XOR2x2_ASAP7_75t_R _20206_ (.A(_00365_),
    .B(_07859_),
    .Y(_07860_));
 AND2x2_ASAP7_75t_R _20207_ (.A(_07771_),
    .B(_07860_),
    .Y(_04706_));
 OR5x1_ASAP7_75t_R _20208_ (.A(_00336_),
    .B(_00365_),
    .C(_00366_),
    .D(_07852_),
    .E(_07853_),
    .Y(_07861_));
 XOR2x2_ASAP7_75t_R _20209_ (.A(_00364_),
    .B(_07861_),
    .Y(_07862_));
 AND2x2_ASAP7_75t_R _20210_ (.A(_07771_),
    .B(_07862_),
    .Y(_04707_));
 OR5x2_ASAP7_75t_R _20211_ (.A(_00336_),
    .B(_00364_),
    .C(_00365_),
    .D(_00366_),
    .E(_07853_),
    .Y(_07863_));
 OR3x1_ASAP7_75t_R _20212_ (.A(_00363_),
    .B(_07858_),
    .C(_07863_),
    .Y(_07864_));
 OAI21x1_ASAP7_75t_R _20213_ (.A1(_07858_),
    .A2(_07863_),
    .B(_00363_),
    .Y(_07865_));
 AND3x1_ASAP7_75t_R _20214_ (.A(_07808_),
    .B(_07864_),
    .C(_07865_),
    .Y(_04708_));
 OR4x1_ASAP7_75t_R _20215_ (.A(_00362_),
    .B(_00363_),
    .C(_07852_),
    .D(_07863_),
    .Y(_07866_));
 BUFx6f_ASAP7_75t_R _20216_ (.A(_07866_),
    .Y(_07867_));
 OR3x1_ASAP7_75t_R _20217_ (.A(_00363_),
    .B(_07852_),
    .C(_07863_),
    .Y(_07868_));
 NAND2x1_ASAP7_75t_R _20218_ (.A(_00362_),
    .B(_07868_),
    .Y(_07869_));
 AND3x1_ASAP7_75t_R _20219_ (.A(_07808_),
    .B(_07867_),
    .C(_07869_),
    .Y(_04709_));
 OR4x1_ASAP7_75t_R _20220_ (.A(_00362_),
    .B(_00363_),
    .C(_07858_),
    .D(_07863_),
    .Y(_07870_));
 XOR2x2_ASAP7_75t_R _20221_ (.A(_07838_),
    .B(_07870_),
    .Y(_07871_));
 AND2x2_ASAP7_75t_R _20222_ (.A(_07771_),
    .B(_07871_),
    .Y(_04710_));
 OR3x1_ASAP7_75t_R _20223_ (.A(_00360_),
    .B(_07838_),
    .C(_07867_),
    .Y(_07872_));
 OAI21x1_ASAP7_75t_R _20224_ (.A1(_07838_),
    .A2(_07867_),
    .B(_00360_),
    .Y(_07873_));
 AND3x1_ASAP7_75t_R _20225_ (.A(_07808_),
    .B(_07872_),
    .C(_07873_),
    .Y(_04711_));
 OR3x1_ASAP7_75t_R _20226_ (.A(_00360_),
    .B(_07838_),
    .C(_07870_),
    .Y(_07874_));
 XOR2x2_ASAP7_75t_R _20227_ (.A(_00359_),
    .B(_07874_),
    .Y(_07875_));
 AND2x2_ASAP7_75t_R _20228_ (.A(_07771_),
    .B(_07875_),
    .Y(_04712_));
 OR4x1_ASAP7_75t_R _20229_ (.A(_00359_),
    .B(_00360_),
    .C(_07838_),
    .D(_07867_),
    .Y(_07876_));
 XOR2x2_ASAP7_75t_R _20230_ (.A(_00358_),
    .B(_07876_),
    .Y(_07877_));
 AND2x2_ASAP7_75t_R _20231_ (.A(_07771_),
    .B(_07877_),
    .Y(_04713_));
 BUFx6f_ASAP7_75t_R _20232_ (.A(_07689_),
    .Y(_07878_));
 OR5x1_ASAP7_75t_R _20233_ (.A(_00358_),
    .B(_00359_),
    .C(_00360_),
    .D(_07838_),
    .E(_07870_),
    .Y(_07879_));
 XOR2x2_ASAP7_75t_R _20234_ (.A(_00357_),
    .B(_07879_),
    .Y(_07880_));
 AND2x2_ASAP7_75t_R _20235_ (.A(_07878_),
    .B(_07880_),
    .Y(_04714_));
 NOR2x1_ASAP7_75t_R _20236_ (.A(_10986_),
    .B(_02652_),
    .Y(_04715_));
 OR5x2_ASAP7_75t_R _20237_ (.A(_00357_),
    .B(_00358_),
    .C(_00359_),
    .D(_00360_),
    .E(_07838_),
    .Y(_07881_));
 OR3x1_ASAP7_75t_R _20238_ (.A(_00355_),
    .B(_07867_),
    .C(_07881_),
    .Y(_07882_));
 OAI21x1_ASAP7_75t_R _20239_ (.A1(_07867_),
    .A2(_07881_),
    .B(_00355_),
    .Y(_07883_));
 AND3x1_ASAP7_75t_R _20240_ (.A(_07808_),
    .B(_07882_),
    .C(_07883_),
    .Y(_04716_));
 OR3x1_ASAP7_75t_R _20241_ (.A(_00355_),
    .B(_07870_),
    .C(_07881_),
    .Y(_07884_));
 XOR2x2_ASAP7_75t_R _20242_ (.A(_00354_),
    .B(_07884_),
    .Y(_07885_));
 AND2x2_ASAP7_75t_R _20243_ (.A(_07878_),
    .B(_07885_),
    .Y(_04717_));
 OR3x1_ASAP7_75t_R _20244_ (.A(_00354_),
    .B(_00355_),
    .C(_07881_),
    .Y(_07886_));
 OR3x2_ASAP7_75t_R _20245_ (.A(_00353_),
    .B(_07867_),
    .C(_07886_),
    .Y(_07887_));
 OAI21x1_ASAP7_75t_R _20246_ (.A1(_07867_),
    .A2(_07886_),
    .B(_00353_),
    .Y(_07888_));
 AND3x1_ASAP7_75t_R _20247_ (.A(_07808_),
    .B(_07887_),
    .C(_07888_),
    .Y(_04718_));
 OR3x2_ASAP7_75t_R _20248_ (.A(_00353_),
    .B(_07870_),
    .C(_07886_),
    .Y(_07889_));
 XOR2x2_ASAP7_75t_R _20249_ (.A(_07842_),
    .B(_07889_),
    .Y(_07890_));
 AND2x2_ASAP7_75t_R _20250_ (.A(_07878_),
    .B(_07890_),
    .Y(_04719_));
 OR3x1_ASAP7_75t_R _20251_ (.A(_00351_),
    .B(_07842_),
    .C(_07887_),
    .Y(_07891_));
 OAI21x1_ASAP7_75t_R _20252_ (.A1(_07842_),
    .A2(_07887_),
    .B(_00351_),
    .Y(_07892_));
 AND3x1_ASAP7_75t_R _20253_ (.A(_07808_),
    .B(_07891_),
    .C(_07892_),
    .Y(_04720_));
 OR3x1_ASAP7_75t_R _20254_ (.A(_00351_),
    .B(_07842_),
    .C(_07889_),
    .Y(_07893_));
 XOR2x2_ASAP7_75t_R _20255_ (.A(_00350_),
    .B(_07893_),
    .Y(_07894_));
 AND2x2_ASAP7_75t_R _20256_ (.A(_07878_),
    .B(_07894_),
    .Y(_04721_));
 OR4x1_ASAP7_75t_R _20257_ (.A(_00350_),
    .B(_00351_),
    .C(_07842_),
    .D(_07887_),
    .Y(_07895_));
 XOR2x2_ASAP7_75t_R _20258_ (.A(_00349_),
    .B(_07895_),
    .Y(_07896_));
 AND2x2_ASAP7_75t_R _20259_ (.A(_07878_),
    .B(_07896_),
    .Y(_04722_));
 OR5x1_ASAP7_75t_R _20260_ (.A(_00349_),
    .B(_00350_),
    .C(_00351_),
    .D(_07842_),
    .E(_07889_),
    .Y(_07897_));
 XOR2x2_ASAP7_75t_R _20261_ (.A(_00348_),
    .B(_07897_),
    .Y(_07898_));
 AND2x2_ASAP7_75t_R _20262_ (.A(_07878_),
    .B(_07898_),
    .Y(_04723_));
 OR5x2_ASAP7_75t_R _20263_ (.A(_00348_),
    .B(_00349_),
    .C(_00350_),
    .D(_00351_),
    .E(_07842_),
    .Y(_07899_));
 OR3x1_ASAP7_75t_R _20264_ (.A(_00347_),
    .B(_07887_),
    .C(_07899_),
    .Y(_07900_));
 OAI21x1_ASAP7_75t_R _20265_ (.A1(_07887_),
    .A2(_07899_),
    .B(_00347_),
    .Y(_07901_));
 AND3x1_ASAP7_75t_R _20266_ (.A(_07808_),
    .B(_07900_),
    .C(_07901_),
    .Y(_04724_));
 OR3x1_ASAP7_75t_R _20267_ (.A(_00347_),
    .B(_07889_),
    .C(_07899_),
    .Y(_07902_));
 XOR2x2_ASAP7_75t_R _20268_ (.A(_00346_),
    .B(_07902_),
    .Y(_07903_));
 AND2x2_ASAP7_75t_R _20269_ (.A(_07878_),
    .B(_07903_),
    .Y(_04725_));
 XOR2x2_ASAP7_75t_R _20270_ (.A(_00345_),
    .B(_02651_),
    .Y(_07904_));
 AND2x2_ASAP7_75t_R _20271_ (.A(_07878_),
    .B(_07904_),
    .Y(_04726_));
 OR4x1_ASAP7_75t_R _20272_ (.A(_00346_),
    .B(_00347_),
    .C(_07887_),
    .D(_07899_),
    .Y(_07905_));
 XOR2x2_ASAP7_75t_R _20273_ (.A(_00344_),
    .B(_07905_),
    .Y(_07906_));
 AND2x2_ASAP7_75t_R _20274_ (.A(_07878_),
    .B(_07906_),
    .Y(_04727_));
 OR5x1_ASAP7_75t_R _20275_ (.A(_00344_),
    .B(_00346_),
    .C(_00347_),
    .D(_07889_),
    .E(_07899_),
    .Y(_07907_));
 XOR2x2_ASAP7_75t_R _20276_ (.A(_00343_),
    .B(_07907_),
    .Y(_07908_));
 AND2x2_ASAP7_75t_R _20277_ (.A(_07878_),
    .B(_07908_),
    .Y(_04728_));
 BUFx6f_ASAP7_75t_R _20278_ (.A(_07689_),
    .Y(_07909_));
 XOR2x2_ASAP7_75t_R _20279_ (.A(_00342_),
    .B(_07856_),
    .Y(_07910_));
 AND2x2_ASAP7_75t_R _20280_ (.A(_07909_),
    .B(_07910_),
    .Y(_04729_));
 NAND2x1_ASAP7_75t_R _20281_ (.A(_00341_),
    .B(_07850_),
    .Y(_07911_));
 AND3x1_ASAP7_75t_R _20282_ (.A(_07808_),
    .B(_07852_),
    .C(_07911_),
    .Y(_04730_));
 XOR2x2_ASAP7_75t_R _20283_ (.A(_00340_),
    .B(_07858_),
    .Y(_07912_));
 AND2x2_ASAP7_75t_R _20284_ (.A(_07909_),
    .B(_07912_),
    .Y(_04731_));
 OR3x1_ASAP7_75t_R _20285_ (.A(_00339_),
    .B(_00340_),
    .C(_07852_),
    .Y(_07913_));
 OAI21x1_ASAP7_75t_R _20286_ (.A1(_00340_),
    .A2(_07852_),
    .B(_00339_),
    .Y(_07914_));
 AND3x1_ASAP7_75t_R _20287_ (.A(_07808_),
    .B(_07913_),
    .C(_07914_),
    .Y(_04732_));
 OR3x1_ASAP7_75t_R _20288_ (.A(_00339_),
    .B(_00340_),
    .C(_07858_),
    .Y(_07915_));
 XOR2x2_ASAP7_75t_R _20289_ (.A(_00338_),
    .B(_07915_),
    .Y(_07916_));
 AND2x2_ASAP7_75t_R _20290_ (.A(_07909_),
    .B(_07916_),
    .Y(_04733_));
 OR4x1_ASAP7_75t_R _20291_ (.A(_00338_),
    .B(_00339_),
    .C(_00340_),
    .D(_07852_),
    .Y(_07917_));
 XOR2x2_ASAP7_75t_R _20292_ (.A(_00337_),
    .B(_07917_),
    .Y(_07918_));
 AND2x2_ASAP7_75t_R _20293_ (.A(_07909_),
    .B(_07918_),
    .Y(_04734_));
 BUFx6f_ASAP7_75t_R _20294_ (.A(_08998_),
    .Y(_07919_));
 OR3x1_ASAP7_75t_R _20295_ (.A(_00336_),
    .B(_07853_),
    .C(_07858_),
    .Y(_07920_));
 OAI21x1_ASAP7_75t_R _20296_ (.A1(_07853_),
    .A2(_07858_),
    .B(_00336_),
    .Y(_07921_));
 AND3x1_ASAP7_75t_R _20297_ (.A(_07919_),
    .B(_07920_),
    .C(_07921_),
    .Y(_04735_));
 BUFx6f_ASAP7_75t_R _20298_ (.A(_00318_),
    .Y(_07922_));
 BUFx6f_ASAP7_75t_R _20299_ (.A(_00326_),
    .Y(_07923_));
 AND4x1_ASAP7_75t_R _20300_ (.A(_00297_),
    .B(_00325_),
    .C(_07923_),
    .D(_00327_),
    .Y(_07924_));
 AND5x1_ASAP7_75t_R _20301_ (.A(_00316_),
    .B(_00321_),
    .C(_00322_),
    .D(_00324_),
    .E(_07924_),
    .Y(_07925_));
 AND5x2_ASAP7_75t_R _20302_ (.A(_07922_),
    .B(_00319_),
    .C(_00320_),
    .D(_07147_),
    .E(_07925_),
    .Y(_07926_));
 AND4x1_ASAP7_75t_R _20303_ (.A(_00311_),
    .B(_00312_),
    .C(_00313_),
    .D(_00314_),
    .Y(_07927_));
 AND4x1_ASAP7_75t_R _20304_ (.A(_00305_),
    .B(_00307_),
    .C(_00308_),
    .D(_00315_),
    .Y(_07928_));
 AND5x1_ASAP7_75t_R _20305_ (.A(_00298_),
    .B(_00299_),
    .C(_00304_),
    .D(_00323_),
    .E(_07928_),
    .Y(_07929_));
 BUFx3_ASAP7_75t_R _20306_ (.A(_00301_),
    .Y(_07930_));
 AND3x1_ASAP7_75t_R _20307_ (.A(_00302_),
    .B(_00303_),
    .C(_00306_),
    .Y(_07931_));
 OR3x1_ASAP7_75t_R _20308_ (.A(_00300_),
    .B(_07930_),
    .C(_07931_),
    .Y(_07932_));
 AND5x2_ASAP7_75t_R _20309_ (.A(_00309_),
    .B(_00310_),
    .C(_07927_),
    .D(_07929_),
    .E(_07932_),
    .Y(_07933_));
 NAND2x2_ASAP7_75t_R _20310_ (.A(_07926_),
    .B(_07933_),
    .Y(_07934_));
 NOR2x1_ASAP7_75t_R _20311_ (.A(_00287_),
    .B(_07934_),
    .Y(_04736_));
 INVx1_ASAP7_75t_R _20312_ (.A(_07934_),
    .Y(_04737_));
 NOR2x1_ASAP7_75t_R _20313_ (.A(_00290_),
    .B(_07934_),
    .Y(_04738_));
 NOR2x1_ASAP7_75t_R _20314_ (.A(_00289_),
    .B(_07934_),
    .Y(_04739_));
 NOR2x1_ASAP7_75t_R _20315_ (.A(_00288_),
    .B(_07934_),
    .Y(_04740_));
 NOR2x1_ASAP7_75t_R _20316_ (.A(_00286_),
    .B(_07934_),
    .Y(_04741_));
 NOR2x1_ASAP7_75t_R _20317_ (.A(_00285_),
    .B(_07934_),
    .Y(_04742_));
 INVx1_ASAP7_75t_R _20318_ (.A(_07934_),
    .Y(_04743_));
 AND2x2_ASAP7_75t_R _20319_ (.A(_07909_),
    .B(_00058_),
    .Y(_04744_));
 OR4x1_ASAP7_75t_R _20320_ (.A(_00302_),
    .B(_00303_),
    .C(_00306_),
    .D(_02665_),
    .Y(_07935_));
 OR5x2_ASAP7_75t_R _20321_ (.A(_00297_),
    .B(_00298_),
    .C(_00299_),
    .D(_00300_),
    .E(_07930_),
    .Y(_07936_));
 OR3x1_ASAP7_75t_R _20322_ (.A(_00327_),
    .B(_07935_),
    .C(_07936_),
    .Y(_07937_));
 BUFx6f_ASAP7_75t_R _20323_ (.A(_07937_),
    .Y(_07938_));
 OAI21x1_ASAP7_75t_R _20324_ (.A1(_07935_),
    .A2(_07936_),
    .B(_00327_),
    .Y(_07939_));
 AND3x1_ASAP7_75t_R _20325_ (.A(_07919_),
    .B(_07938_),
    .C(_07939_),
    .Y(_04745_));
 OR5x2_ASAP7_75t_R _20326_ (.A(_00302_),
    .B(_00303_),
    .C(_00306_),
    .D(_00317_),
    .E(_00058_),
    .Y(_07940_));
 OR3x2_ASAP7_75t_R _20327_ (.A(_00327_),
    .B(_07936_),
    .C(_07940_),
    .Y(_07941_));
 XOR2x2_ASAP7_75t_R _20328_ (.A(_07923_),
    .B(_07941_),
    .Y(_07942_));
 AND2x2_ASAP7_75t_R _20329_ (.A(_07909_),
    .B(_07942_),
    .Y(_04746_));
 OR3x1_ASAP7_75t_R _20330_ (.A(_00325_),
    .B(_07923_),
    .C(_07938_),
    .Y(_07943_));
 OAI21x1_ASAP7_75t_R _20331_ (.A1(_07923_),
    .A2(_07938_),
    .B(_00325_),
    .Y(_07944_));
 AND3x1_ASAP7_75t_R _20332_ (.A(_07919_),
    .B(_07943_),
    .C(_07944_),
    .Y(_04747_));
 OR3x1_ASAP7_75t_R _20333_ (.A(_00325_),
    .B(_07923_),
    .C(_07941_),
    .Y(_07945_));
 XOR2x2_ASAP7_75t_R _20334_ (.A(_00324_),
    .B(_07945_),
    .Y(_07946_));
 AND2x2_ASAP7_75t_R _20335_ (.A(_07909_),
    .B(_07946_),
    .Y(_04748_));
 OR4x1_ASAP7_75t_R _20336_ (.A(_00324_),
    .B(_00325_),
    .C(_07923_),
    .D(_07938_),
    .Y(_07947_));
 XOR2x2_ASAP7_75t_R _20337_ (.A(_00323_),
    .B(_07947_),
    .Y(_07948_));
 AND2x2_ASAP7_75t_R _20338_ (.A(_07909_),
    .B(_07948_),
    .Y(_04749_));
 OR5x1_ASAP7_75t_R _20339_ (.A(_00323_),
    .B(_00324_),
    .C(_00325_),
    .D(_07923_),
    .E(_07941_),
    .Y(_07949_));
 XOR2x2_ASAP7_75t_R _20340_ (.A(_00322_),
    .B(_07949_),
    .Y(_07950_));
 AND2x2_ASAP7_75t_R _20341_ (.A(_07909_),
    .B(_07950_),
    .Y(_04750_));
 OR5x2_ASAP7_75t_R _20342_ (.A(_00322_),
    .B(_00323_),
    .C(_00324_),
    .D(_00325_),
    .E(_07923_),
    .Y(_07951_));
 OR3x1_ASAP7_75t_R _20343_ (.A(_00321_),
    .B(_07938_),
    .C(_07951_),
    .Y(_07952_));
 OAI21x1_ASAP7_75t_R _20344_ (.A1(_07938_),
    .A2(_07951_),
    .B(_00321_),
    .Y(_07953_));
 AND3x1_ASAP7_75t_R _20345_ (.A(_07919_),
    .B(_07952_),
    .C(_07953_),
    .Y(_04751_));
 OR3x1_ASAP7_75t_R _20346_ (.A(_00321_),
    .B(_07941_),
    .C(_07951_),
    .Y(_07954_));
 XOR2x2_ASAP7_75t_R _20347_ (.A(_00320_),
    .B(_07954_),
    .Y(_07955_));
 AND2x2_ASAP7_75t_R _20348_ (.A(_07909_),
    .B(_07955_),
    .Y(_04752_));
 OR3x2_ASAP7_75t_R _20349_ (.A(_00320_),
    .B(_00321_),
    .C(_07951_),
    .Y(_07956_));
 OR3x1_ASAP7_75t_R _20350_ (.A(_00319_),
    .B(_07938_),
    .C(_07956_),
    .Y(_07957_));
 BUFx6f_ASAP7_75t_R _20351_ (.A(_07957_),
    .Y(_07958_));
 OAI21x1_ASAP7_75t_R _20352_ (.A1(_07938_),
    .A2(_07956_),
    .B(_00319_),
    .Y(_07959_));
 AND3x1_ASAP7_75t_R _20353_ (.A(_07919_),
    .B(_07958_),
    .C(_07959_),
    .Y(_04753_));
 BUFx6f_ASAP7_75t_R _20354_ (.A(_07689_),
    .Y(_07960_));
 OR3x2_ASAP7_75t_R _20355_ (.A(_00319_),
    .B(_07941_),
    .C(_07956_),
    .Y(_07961_));
 XOR2x2_ASAP7_75t_R _20356_ (.A(_07922_),
    .B(_07961_),
    .Y(_07962_));
 AND2x2_ASAP7_75t_R _20357_ (.A(_07960_),
    .B(_07962_),
    .Y(_04754_));
 NOR2x1_ASAP7_75t_R _20358_ (.A(_10986_),
    .B(_02666_),
    .Y(_04755_));
 OR3x1_ASAP7_75t_R _20359_ (.A(_00316_),
    .B(_07922_),
    .C(_07958_),
    .Y(_07963_));
 OAI21x1_ASAP7_75t_R _20360_ (.A1(_07922_),
    .A2(_07958_),
    .B(_00316_),
    .Y(_07964_));
 AND3x1_ASAP7_75t_R _20361_ (.A(_07919_),
    .B(_07963_),
    .C(_07964_),
    .Y(_04756_));
 OR3x1_ASAP7_75t_R _20362_ (.A(_00316_),
    .B(_07922_),
    .C(_07961_),
    .Y(_07965_));
 XOR2x2_ASAP7_75t_R _20363_ (.A(_00315_),
    .B(_07965_),
    .Y(_07966_));
 AND2x2_ASAP7_75t_R _20364_ (.A(_07960_),
    .B(_07966_),
    .Y(_04757_));
 OR4x1_ASAP7_75t_R _20365_ (.A(_00315_),
    .B(_00316_),
    .C(_07922_),
    .D(_07958_),
    .Y(_07967_));
 XOR2x2_ASAP7_75t_R _20366_ (.A(_00314_),
    .B(_07967_),
    .Y(_07968_));
 AND2x2_ASAP7_75t_R _20367_ (.A(_07960_),
    .B(_07968_),
    .Y(_04758_));
 OR5x1_ASAP7_75t_R _20368_ (.A(_00314_),
    .B(_00315_),
    .C(_00316_),
    .D(_07922_),
    .E(_07961_),
    .Y(_07969_));
 XOR2x2_ASAP7_75t_R _20369_ (.A(_00313_),
    .B(_07969_),
    .Y(_07970_));
 AND2x2_ASAP7_75t_R _20370_ (.A(_07960_),
    .B(_07970_),
    .Y(_04759_));
 OR5x2_ASAP7_75t_R _20371_ (.A(_00313_),
    .B(_00314_),
    .C(_00315_),
    .D(_00316_),
    .E(_07922_),
    .Y(_07971_));
 OR3x1_ASAP7_75t_R _20372_ (.A(_00312_),
    .B(_07958_),
    .C(_07971_),
    .Y(_07972_));
 OAI21x1_ASAP7_75t_R _20373_ (.A1(_07958_),
    .A2(_07971_),
    .B(_00312_),
    .Y(_07973_));
 AND3x1_ASAP7_75t_R _20374_ (.A(_07919_),
    .B(_07972_),
    .C(_07973_),
    .Y(_04760_));
 OR3x1_ASAP7_75t_R _20375_ (.A(_00312_),
    .B(_07961_),
    .C(_07971_),
    .Y(_07974_));
 XOR2x2_ASAP7_75t_R _20376_ (.A(_00311_),
    .B(_07974_),
    .Y(_07975_));
 AND2x2_ASAP7_75t_R _20377_ (.A(_07960_),
    .B(_07975_),
    .Y(_04761_));
 OR3x2_ASAP7_75t_R _20378_ (.A(_00311_),
    .B(_00312_),
    .C(_07971_),
    .Y(_07976_));
 OR3x2_ASAP7_75t_R _20379_ (.A(_00310_),
    .B(_07958_),
    .C(_07976_),
    .Y(_07977_));
 OAI21x1_ASAP7_75t_R _20380_ (.A1(_07958_),
    .A2(_07976_),
    .B(_00310_),
    .Y(_07978_));
 AND3x1_ASAP7_75t_R _20381_ (.A(_07919_),
    .B(_07977_),
    .C(_07978_),
    .Y(_04762_));
 OR3x2_ASAP7_75t_R _20382_ (.A(_00310_),
    .B(_07961_),
    .C(_07976_),
    .Y(_07979_));
 XOR2x2_ASAP7_75t_R _20383_ (.A(_00309_),
    .B(_07979_),
    .Y(_07980_));
 AND2x2_ASAP7_75t_R _20384_ (.A(_07960_),
    .B(_07980_),
    .Y(_04763_));
 NOR2x1_ASAP7_75t_R _20385_ (.A(_00309_),
    .B(_07977_),
    .Y(_07981_));
 XNOR2x2_ASAP7_75t_R _20386_ (.A(_00308_),
    .B(_07981_),
    .Y(_07982_));
 AND2x2_ASAP7_75t_R _20387_ (.A(_07960_),
    .B(_07982_),
    .Y(_04764_));
 OR3x1_ASAP7_75t_R _20388_ (.A(_00308_),
    .B(_00309_),
    .C(_07979_),
    .Y(_07983_));
 XOR2x2_ASAP7_75t_R _20389_ (.A(_00307_),
    .B(_07983_),
    .Y(_07984_));
 AND2x2_ASAP7_75t_R _20390_ (.A(_07960_),
    .B(_07984_),
    .Y(_04765_));
 XOR2x2_ASAP7_75t_R _20391_ (.A(_00306_),
    .B(_02665_),
    .Y(_07985_));
 AND2x2_ASAP7_75t_R _20392_ (.A(_07960_),
    .B(_07985_),
    .Y(_04766_));
 OR4x1_ASAP7_75t_R _20393_ (.A(_00307_),
    .B(_00308_),
    .C(_00309_),
    .D(_07977_),
    .Y(_07986_));
 XOR2x2_ASAP7_75t_R _20394_ (.A(_00305_),
    .B(_07986_),
    .Y(_07987_));
 AND2x2_ASAP7_75t_R _20395_ (.A(_07960_),
    .B(_07987_),
    .Y(_04767_));
 BUFx6f_ASAP7_75t_R _20396_ (.A(_07689_),
    .Y(_07988_));
 OR5x1_ASAP7_75t_R _20397_ (.A(_00305_),
    .B(_00307_),
    .C(_00308_),
    .D(_00309_),
    .E(_07979_),
    .Y(_07989_));
 XOR2x2_ASAP7_75t_R _20398_ (.A(_00304_),
    .B(_07989_),
    .Y(_07990_));
 AND2x2_ASAP7_75t_R _20399_ (.A(_07988_),
    .B(_07990_),
    .Y(_04768_));
 OR3x1_ASAP7_75t_R _20400_ (.A(_00306_),
    .B(_00317_),
    .C(_00058_),
    .Y(_07991_));
 XOR2x2_ASAP7_75t_R _20401_ (.A(_00303_),
    .B(_07991_),
    .Y(_07992_));
 AND2x2_ASAP7_75t_R _20402_ (.A(_07988_),
    .B(_07992_),
    .Y(_04769_));
 OR3x1_ASAP7_75t_R _20403_ (.A(_00303_),
    .B(_00306_),
    .C(_02665_),
    .Y(_07993_));
 NAND2x1_ASAP7_75t_R _20404_ (.A(_00302_),
    .B(_07993_),
    .Y(_07994_));
 AND3x1_ASAP7_75t_R _20405_ (.A(_07919_),
    .B(_07935_),
    .C(_07994_),
    .Y(_04770_));
 XOR2x2_ASAP7_75t_R _20406_ (.A(_07930_),
    .B(_07940_),
    .Y(_07995_));
 AND2x2_ASAP7_75t_R _20407_ (.A(_07988_),
    .B(_07995_),
    .Y(_04771_));
 OR3x1_ASAP7_75t_R _20408_ (.A(_00300_),
    .B(_07930_),
    .C(_07935_),
    .Y(_07996_));
 OAI21x1_ASAP7_75t_R _20409_ (.A1(_07930_),
    .A2(_07935_),
    .B(_00300_),
    .Y(_07997_));
 AND3x1_ASAP7_75t_R _20410_ (.A(_07919_),
    .B(_07996_),
    .C(_07997_),
    .Y(_04772_));
 OR3x1_ASAP7_75t_R _20411_ (.A(_00300_),
    .B(_07930_),
    .C(_07940_),
    .Y(_07998_));
 XOR2x2_ASAP7_75t_R _20412_ (.A(_00299_),
    .B(_07998_),
    .Y(_07999_));
 AND2x2_ASAP7_75t_R _20413_ (.A(_07988_),
    .B(_07999_),
    .Y(_04773_));
 OR4x1_ASAP7_75t_R _20414_ (.A(_00299_),
    .B(_00300_),
    .C(_07930_),
    .D(_07935_),
    .Y(_08000_));
 XOR2x2_ASAP7_75t_R _20415_ (.A(_00298_),
    .B(_08000_),
    .Y(_08001_));
 AND2x2_ASAP7_75t_R _20416_ (.A(_07988_),
    .B(_08001_),
    .Y(_04774_));
 OR5x1_ASAP7_75t_R _20417_ (.A(_00298_),
    .B(_00299_),
    .C(_00300_),
    .D(_07930_),
    .E(_07940_),
    .Y(_08002_));
 NAND2x1_ASAP7_75t_R _20418_ (.A(_00297_),
    .B(_08002_),
    .Y(_08003_));
 OA211x2_ASAP7_75t_R _20419_ (.A1(_07936_),
    .A2(_07940_),
    .B(_08003_),
    .C(_07260_),
    .Y(_04775_));
 AND2x2_ASAP7_75t_R _20420_ (.A(_07988_),
    .B(_00028_),
    .Y(_04776_));
 BUFx6f_ASAP7_75t_R _20421_ (.A(_02190_),
    .Y(_08004_));
 INVx1_ASAP7_75t_R _20422_ (.A(_02197_),
    .Y(_08005_));
 OR2x2_ASAP7_75t_R _20423_ (.A(_00367_),
    .B(_00372_),
    .Y(_08006_));
 OR2x2_ASAP7_75t_R _20424_ (.A(_00370_),
    .B(_00371_),
    .Y(_08007_));
 OA31x2_ASAP7_75t_R _20425_ (.A1(\peo[14][36] ),
    .A2(_00369_),
    .A3(_08007_),
    .B1(\peo[14][39] ),
    .Y(_08008_));
 AO21x1_ASAP7_75t_R _20426_ (.A1(_08005_),
    .A2(_08006_),
    .B(_08008_),
    .Y(_08009_));
 OR2x2_ASAP7_75t_R _20427_ (.A(_00331_),
    .B(_00332_),
    .Y(_08010_));
 OA31x2_ASAP7_75t_R _20428_ (.A1(\xs[7].cli1.i[36] ),
    .A2(_00330_),
    .A3(_08010_),
    .B1(\xs[7].cli1.i[39] ),
    .Y(_08011_));
 OR5x2_ASAP7_75t_R _20429_ (.A(_00328_),
    .B(\xs[7].cli1.i[36] ),
    .C(_00330_),
    .D(\xs[7].cli1.i[32] ),
    .E(_08010_),
    .Y(_08012_));
 OA21x2_ASAP7_75t_R _20430_ (.A1(_02197_),
    .A2(_08011_),
    .B(_08012_),
    .Y(_08013_));
 OA21x2_ASAP7_75t_R _20431_ (.A1(_08009_),
    .A2(_08013_),
    .B(_02191_),
    .Y(_08014_));
 INVx2_ASAP7_75t_R _20432_ (.A(_08014_),
    .Y(_08015_));
 OR4x1_ASAP7_75t_R _20433_ (.A(_09220_),
    .B(_08004_),
    .C(_08005_),
    .D(_08015_),
    .Y(_08016_));
 BUFx6f_ASAP7_75t_R _20434_ (.A(_08016_),
    .Y(_08017_));
 INVx3_ASAP7_75t_R _20435_ (.A(_08004_),
    .Y(_08018_));
 AND3x1_ASAP7_75t_R _20436_ (.A(_08018_),
    .B(_02197_),
    .C(_08014_),
    .Y(_08019_));
 AO21x1_ASAP7_75t_R _20437_ (.A1(_00028_),
    .A2(_08011_),
    .B(_08018_),
    .Y(_08020_));
 INVx1_ASAP7_75t_R _20438_ (.A(_02191_),
    .Y(_08021_));
 OR3x1_ASAP7_75t_R _20439_ (.A(_08004_),
    .B(_08021_),
    .C(_02197_),
    .Y(_08022_));
 AND3x1_ASAP7_75t_R _20440_ (.A(_08008_),
    .B(_08020_),
    .C(_08022_),
    .Y(_08023_));
 OA21x2_ASAP7_75t_R _20441_ (.A1(_08012_),
    .A2(_08023_),
    .B(_00374_),
    .Y(_08024_));
 OR3x1_ASAP7_75t_R _20442_ (.A(_08941_),
    .B(_08019_),
    .C(_08024_),
    .Y(_08025_));
 NOR2x1_ASAP7_75t_R _20443_ (.A(_00331_),
    .B(_00332_),
    .Y(_08026_));
 AND5x1_ASAP7_75t_R _20444_ (.A(\xs[7].cli1.i[39] ),
    .B(_00329_),
    .C(\xs[7].cli1.i[35] ),
    .D(_00333_),
    .E(_08026_),
    .Y(_08027_));
 AO21x1_ASAP7_75t_R _20445_ (.A1(_08008_),
    .A2(_08027_),
    .B(_08011_),
    .Y(_08028_));
 OA21x2_ASAP7_75t_R _20446_ (.A1(_08027_),
    .A2(_08011_),
    .B(_02197_),
    .Y(_08029_));
 AND3x1_ASAP7_75t_R _20447_ (.A(_08004_),
    .B(_00028_),
    .C(_08011_),
    .Y(_08030_));
 AO21x1_ASAP7_75t_R _20448_ (.A1(_08018_),
    .A2(_08029_),
    .B(_08030_),
    .Y(_08031_));
 AO32x1_ASAP7_75t_R _20449_ (.A1(_08018_),
    .A2(_08021_),
    .A3(_08028_),
    .B1(_08031_),
    .B2(_08008_),
    .Y(_08032_));
 BUFx3_ASAP7_75t_R _20450_ (.A(_08032_),
    .Y(_08033_));
 NOR3x1_ASAP7_75t_R _20451_ (.A(\peo[15][0] ),
    .B(_08012_),
    .C(_08033_),
    .Y(_08034_));
 OAI22x1_ASAP7_75t_R _20452_ (.A1(_02201_),
    .A2(_08017_),
    .B1(_08025_),
    .B2(_08034_),
    .Y(_04777_));
 NOR2x1_ASAP7_75t_R _20453_ (.A(_02200_),
    .B(_08017_),
    .Y(_04778_));
 NOR2x1_ASAP7_75t_R _20454_ (.A(_02199_),
    .B(_08017_),
    .Y(_04779_));
 NOR2x1_ASAP7_75t_R _20455_ (.A(_02198_),
    .B(_08017_),
    .Y(_04780_));
 NOR2x1_ASAP7_75t_R _20456_ (.A(_02189_),
    .B(_08017_),
    .Y(_04781_));
 NOR2x1_ASAP7_75t_R _20457_ (.A(_02188_),
    .B(_08017_),
    .Y(_04782_));
 BUFx6f_ASAP7_75t_R _20458_ (.A(_08998_),
    .Y(_08035_));
 NOR2x1_ASAP7_75t_R _20459_ (.A(_08009_),
    .B(_08013_),
    .Y(_08036_));
 OAI21x1_ASAP7_75t_R _20460_ (.A1(_08036_),
    .A2(_08022_),
    .B(_00374_),
    .Y(_08037_));
 INVx1_ASAP7_75t_R _20461_ (.A(_02201_),
    .Y(_08038_));
 OR3x1_ASAP7_75t_R _20462_ (.A(_08038_),
    .B(_08036_),
    .C(_08022_),
    .Y(_08039_));
 AO21x1_ASAP7_75t_R _20463_ (.A1(_08037_),
    .A2(_08039_),
    .B(_08033_),
    .Y(_08040_));
 NAND2x1_ASAP7_75t_R _20464_ (.A(_00335_),
    .B(_08033_),
    .Y(_08041_));
 AND3x1_ASAP7_75t_R _20465_ (.A(_08035_),
    .B(_08040_),
    .C(_08041_),
    .Y(_04783_));
 OR4x1_ASAP7_75t_R _20466_ (.A(_11177_),
    .B(_08004_),
    .C(_02197_),
    .D(_08015_),
    .Y(_08042_));
 NOR2x1_ASAP7_75t_R _20467_ (.A(_02200_),
    .B(_08042_),
    .Y(_04784_));
 NOR2x1_ASAP7_75t_R _20468_ (.A(_02199_),
    .B(_08042_),
    .Y(_04785_));
 NOR2x1_ASAP7_75t_R _20469_ (.A(_02198_),
    .B(_08042_),
    .Y(_04786_));
 NOR2x1_ASAP7_75t_R _20470_ (.A(_02189_),
    .B(_08042_),
    .Y(_04787_));
 NOR2x1_ASAP7_75t_R _20471_ (.A(_02188_),
    .B(_08042_),
    .Y(_04788_));
 OA21x2_ASAP7_75t_R _20472_ (.A1(_08004_),
    .A2(_08014_),
    .B(_08581_),
    .Y(_08043_));
 OAI21x1_ASAP7_75t_R _20473_ (.A1(_08004_),
    .A2(_02191_),
    .B(_08011_),
    .Y(_08044_));
 AO21x1_ASAP7_75t_R _20474_ (.A1(_08008_),
    .A2(_08031_),
    .B(_08044_),
    .Y(_08045_));
 BUFx6f_ASAP7_75t_R _20475_ (.A(_08045_),
    .Y(_08046_));
 OR2x2_ASAP7_75t_R _20476_ (.A(\peo[15][0] ),
    .B(_08046_),
    .Y(_08047_));
 NAND2x1_ASAP7_75t_R _20477_ (.A(_00374_),
    .B(_08046_),
    .Y(_08048_));
 AND3x4_ASAP7_75t_R _20478_ (.A(_08598_),
    .B(_08018_),
    .C(_08015_),
    .Y(_08049_));
 AO32x1_ASAP7_75t_R _20479_ (.A1(_08043_),
    .A2(_08047_),
    .A3(_08048_),
    .B1(_08049_),
    .B2(_08038_),
    .Y(_04789_));
 OR3x1_ASAP7_75t_R _20480_ (.A(_08578_),
    .B(_08004_),
    .C(_08014_),
    .Y(_08050_));
 BUFx6f_ASAP7_75t_R _20481_ (.A(_08050_),
    .Y(_08051_));
 NOR2x1_ASAP7_75t_R _20482_ (.A(_02200_),
    .B(_08051_),
    .Y(_04790_));
 NOR2x1_ASAP7_75t_R _20483_ (.A(_02199_),
    .B(_08051_),
    .Y(_04791_));
 NOR2x1_ASAP7_75t_R _20484_ (.A(_02198_),
    .B(_08051_),
    .Y(_04792_));
 OR2x2_ASAP7_75t_R _20485_ (.A(\xs[7].cli1.i[32] ),
    .B(_08046_),
    .Y(_08052_));
 NAND2x1_ASAP7_75t_R _20486_ (.A(_00372_),
    .B(_08046_),
    .Y(_08053_));
 AO32x1_ASAP7_75t_R _20487_ (.A1(_08043_),
    .A2(_08052_),
    .A3(_08053_),
    .B1(_08049_),
    .B2(_08005_),
    .Y(_04793_));
 NAND2x1_ASAP7_75t_R _20488_ (.A(_00371_),
    .B(_08046_),
    .Y(_08054_));
 OR3x1_ASAP7_75t_R _20489_ (.A(_00328_),
    .B(\xs[7].cli1.i[33] ),
    .C(_08033_),
    .Y(_08055_));
 INVx1_ASAP7_75t_R _20490_ (.A(_02196_),
    .Y(_08056_));
 AO32x1_ASAP7_75t_R _20491_ (.A1(_08043_),
    .A2(_08054_),
    .A3(_08055_),
    .B1(_08049_),
    .B2(_08056_),
    .Y(_04794_));
 NAND2x1_ASAP7_75t_R _20492_ (.A(_00370_),
    .B(_08046_),
    .Y(_08057_));
 OR3x1_ASAP7_75t_R _20493_ (.A(_00328_),
    .B(\xs[7].cli1.i[34] ),
    .C(_08033_),
    .Y(_08058_));
 INVx1_ASAP7_75t_R _20494_ (.A(_02195_),
    .Y(_08059_));
 AO32x1_ASAP7_75t_R _20495_ (.A1(_08043_),
    .A2(_08057_),
    .A3(_08058_),
    .B1(_08049_),
    .B2(_08059_),
    .Y(_04795_));
 NAND2x1_ASAP7_75t_R _20496_ (.A(_00369_),
    .B(_08046_),
    .Y(_08060_));
 OR3x1_ASAP7_75t_R _20497_ (.A(_00328_),
    .B(\xs[7].cli1.i[35] ),
    .C(_08033_),
    .Y(_08061_));
 INVx1_ASAP7_75t_R _20498_ (.A(_02194_),
    .Y(_08062_));
 AO32x1_ASAP7_75t_R _20499_ (.A1(_08043_),
    .A2(_08060_),
    .A3(_08061_),
    .B1(_08049_),
    .B2(_08062_),
    .Y(_04796_));
 OR2x2_ASAP7_75t_R _20500_ (.A(\xs[7].cli1.i[36] ),
    .B(_08046_),
    .Y(_08063_));
 NAND2x1_ASAP7_75t_R _20501_ (.A(_00368_),
    .B(_08046_),
    .Y(_08064_));
 INVx1_ASAP7_75t_R _20502_ (.A(_02193_),
    .Y(_08065_));
 AO32x1_ASAP7_75t_R _20503_ (.A1(_08043_),
    .A2(_08063_),
    .A3(_08064_),
    .B1(_08049_),
    .B2(_08065_),
    .Y(_04797_));
 NOR2x1_ASAP7_75t_R _20504_ (.A(_02192_),
    .B(_08051_),
    .Y(_04798_));
 AND4x1_ASAP7_75t_R _20505_ (.A(_08585_),
    .B(_08018_),
    .C(_02191_),
    .D(_08036_),
    .Y(_04799_));
 AOI211x1_ASAP7_75t_R _20506_ (.A1(_08018_),
    .A2(_08015_),
    .B(_08011_),
    .C(_08008_),
    .Y(_08066_));
 NOR2x1_ASAP7_75t_R _20507_ (.A(_10986_),
    .B(_08066_),
    .Y(_04800_));
 NOR2x1_ASAP7_75t_R _20508_ (.A(_02189_),
    .B(_08051_),
    .Y(_04801_));
 NOR2x1_ASAP7_75t_R _20509_ (.A(_02188_),
    .B(_08051_),
    .Y(_04802_));
 BUFx6f_ASAP7_75t_R _20510_ (.A(_00255_),
    .Y(_08067_));
 BUFx3_ASAP7_75t_R _20511_ (.A(_00232_),
    .Y(_08068_));
 AND4x1_ASAP7_75t_R _20512_ (.A(_08068_),
    .B(_00260_),
    .C(_00261_),
    .D(_00262_),
    .Y(_08069_));
 AND5x1_ASAP7_75t_R _20513_ (.A(_00251_),
    .B(_00256_),
    .C(_00257_),
    .D(_00259_),
    .E(_08069_),
    .Y(_08070_));
 AND5x2_ASAP7_75t_R _20514_ (.A(_00253_),
    .B(_00254_),
    .C(_08067_),
    .D(_07147_),
    .E(_08070_),
    .Y(_08071_));
 BUFx6f_ASAP7_75t_R _20515_ (.A(_00247_),
    .Y(_08072_));
 AND4x1_ASAP7_75t_R _20516_ (.A(_00246_),
    .B(_08072_),
    .C(_00248_),
    .D(_00249_),
    .Y(_08073_));
 AND4x1_ASAP7_75t_R _20517_ (.A(_00240_),
    .B(_00242_),
    .C(_00243_),
    .D(_00250_),
    .Y(_08074_));
 AND5x1_ASAP7_75t_R _20518_ (.A(_00233_),
    .B(_00234_),
    .C(_00239_),
    .D(_00258_),
    .E(_08074_),
    .Y(_08075_));
 AND3x1_ASAP7_75t_R _20519_ (.A(_00237_),
    .B(_00238_),
    .C(_00241_),
    .Y(_08076_));
 OR3x1_ASAP7_75t_R _20520_ (.A(_00235_),
    .B(_00236_),
    .C(_08076_),
    .Y(_08077_));
 AND5x2_ASAP7_75t_R _20521_ (.A(_00244_),
    .B(_00245_),
    .C(_08073_),
    .D(_08075_),
    .E(_08077_),
    .Y(_08078_));
 NAND2x2_ASAP7_75t_R _20522_ (.A(_08071_),
    .B(_08078_),
    .Y(_08079_));
 NOR2x1_ASAP7_75t_R _20523_ (.A(_00189_),
    .B(_08079_),
    .Y(_04803_));
 INVx1_ASAP7_75t_R _20524_ (.A(_08079_),
    .Y(_04804_));
 NOR2x1_ASAP7_75t_R _20525_ (.A(_00192_),
    .B(_08079_),
    .Y(_04805_));
 NOR2x1_ASAP7_75t_R _20526_ (.A(_00191_),
    .B(_08079_),
    .Y(_04806_));
 NOR2x1_ASAP7_75t_R _20527_ (.A(_00190_),
    .B(_08079_),
    .Y(_04807_));
 NOR2x1_ASAP7_75t_R _20528_ (.A(_00188_),
    .B(_08079_),
    .Y(_04808_));
 NOR2x1_ASAP7_75t_R _20529_ (.A(_00187_),
    .B(_08079_),
    .Y(_04809_));
 INVx1_ASAP7_75t_R _20530_ (.A(_08079_),
    .Y(_04810_));
 AND2x2_ASAP7_75t_R _20531_ (.A(_07988_),
    .B(_00059_),
    .Y(_04811_));
 OR4x1_ASAP7_75t_R _20532_ (.A(_00237_),
    .B(_00238_),
    .C(_00241_),
    .D(_02671_),
    .Y(_08080_));
 OR4x1_ASAP7_75t_R _20533_ (.A(_00233_),
    .B(_00234_),
    .C(_00235_),
    .D(_00236_),
    .Y(_08081_));
 OR2x6_ASAP7_75t_R _20534_ (.A(_08080_),
    .B(_08081_),
    .Y(_08082_));
 OR3x1_ASAP7_75t_R _20535_ (.A(_08068_),
    .B(_00262_),
    .C(_08082_),
    .Y(_08083_));
 OAI21x1_ASAP7_75t_R _20536_ (.A1(_08068_),
    .A2(_08082_),
    .B(_00262_),
    .Y(_08084_));
 AND3x1_ASAP7_75t_R _20537_ (.A(_08035_),
    .B(_08083_),
    .C(_08084_),
    .Y(_04812_));
 OR5x2_ASAP7_75t_R _20538_ (.A(_00237_),
    .B(_00238_),
    .C(_00241_),
    .D(_00252_),
    .E(_00059_),
    .Y(_08085_));
 OR2x6_ASAP7_75t_R _20539_ (.A(_08081_),
    .B(_08085_),
    .Y(_08086_));
 OR3x1_ASAP7_75t_R _20540_ (.A(_08068_),
    .B(_00262_),
    .C(_08086_),
    .Y(_08087_));
 XOR2x2_ASAP7_75t_R _20541_ (.A(_00261_),
    .B(_08087_),
    .Y(_08088_));
 AND2x2_ASAP7_75t_R _20542_ (.A(_07988_),
    .B(_08088_),
    .Y(_04813_));
 OR4x1_ASAP7_75t_R _20543_ (.A(_08068_),
    .B(_00261_),
    .C(_00262_),
    .D(_08082_),
    .Y(_08089_));
 XOR2x2_ASAP7_75t_R _20544_ (.A(_00260_),
    .B(_08089_),
    .Y(_08090_));
 AND2x2_ASAP7_75t_R _20545_ (.A(_07988_),
    .B(_08090_),
    .Y(_04814_));
 OR5x2_ASAP7_75t_R _20546_ (.A(_08068_),
    .B(_00259_),
    .C(_00260_),
    .D(_00261_),
    .E(_00262_),
    .Y(_08091_));
 OR5x1_ASAP7_75t_R _20547_ (.A(_08068_),
    .B(_00260_),
    .C(_00261_),
    .D(_00262_),
    .E(_08086_),
    .Y(_08092_));
 NAND2x1_ASAP7_75t_R _20548_ (.A(_00259_),
    .B(_08092_),
    .Y(_08093_));
 OA211x2_ASAP7_75t_R _20549_ (.A1(_08086_),
    .A2(_08091_),
    .B(_08093_),
    .C(_07260_),
    .Y(_04815_));
 OR3x2_ASAP7_75t_R _20550_ (.A(_08080_),
    .B(_08081_),
    .C(_08091_),
    .Y(_08094_));
 XOR2x2_ASAP7_75t_R _20551_ (.A(_00258_),
    .B(_08094_),
    .Y(_08095_));
 AND2x2_ASAP7_75t_R _20552_ (.A(_07988_),
    .B(_08095_),
    .Y(_04816_));
 BUFx6f_ASAP7_75t_R _20553_ (.A(_07689_),
    .Y(_08096_));
 OR3x1_ASAP7_75t_R _20554_ (.A(_00258_),
    .B(_08086_),
    .C(_08091_),
    .Y(_08097_));
 XOR2x2_ASAP7_75t_R _20555_ (.A(_00257_),
    .B(_08097_),
    .Y(_08098_));
 AND2x2_ASAP7_75t_R _20556_ (.A(_08096_),
    .B(_08098_),
    .Y(_04817_));
 OR4x1_ASAP7_75t_R _20557_ (.A(_00256_),
    .B(_00257_),
    .C(_00258_),
    .D(_08094_),
    .Y(_08099_));
 OR3x1_ASAP7_75t_R _20558_ (.A(_00257_),
    .B(_00258_),
    .C(_08094_),
    .Y(_08100_));
 NAND2x1_ASAP7_75t_R _20559_ (.A(_00256_),
    .B(_08100_),
    .Y(_08101_));
 AND3x1_ASAP7_75t_R _20560_ (.A(_08035_),
    .B(_08099_),
    .C(_08101_),
    .Y(_04818_));
 OR5x2_ASAP7_75t_R _20561_ (.A(_00256_),
    .B(_00257_),
    .C(_00258_),
    .D(_08086_),
    .E(_08091_),
    .Y(_08102_));
 XOR2x2_ASAP7_75t_R _20562_ (.A(_08067_),
    .B(_08102_),
    .Y(_08103_));
 AND2x2_ASAP7_75t_R _20563_ (.A(_08096_),
    .B(_08103_),
    .Y(_04819_));
 OR3x1_ASAP7_75t_R _20564_ (.A(_00254_),
    .B(_08067_),
    .C(_08099_),
    .Y(_08104_));
 OAI21x1_ASAP7_75t_R _20565_ (.A1(_08067_),
    .A2(_08099_),
    .B(_00254_),
    .Y(_08105_));
 AND3x1_ASAP7_75t_R _20566_ (.A(_08035_),
    .B(_08104_),
    .C(_08105_),
    .Y(_04820_));
 OR3x1_ASAP7_75t_R _20567_ (.A(_00254_),
    .B(_08067_),
    .C(_08102_),
    .Y(_08106_));
 XOR2x2_ASAP7_75t_R _20568_ (.A(_00253_),
    .B(_08106_),
    .Y(_08107_));
 AND2x2_ASAP7_75t_R _20569_ (.A(_08096_),
    .B(_08107_),
    .Y(_04821_));
 NOR2x1_ASAP7_75t_R _20570_ (.A(_10986_),
    .B(_02672_),
    .Y(_04822_));
 OR4x1_ASAP7_75t_R _20571_ (.A(_00253_),
    .B(_00254_),
    .C(_08067_),
    .D(_08099_),
    .Y(_08108_));
 XOR2x2_ASAP7_75t_R _20572_ (.A(_00251_),
    .B(_08108_),
    .Y(_08109_));
 AND2x2_ASAP7_75t_R _20573_ (.A(_08096_),
    .B(_08109_),
    .Y(_04823_));
 OR5x1_ASAP7_75t_R _20574_ (.A(_00251_),
    .B(_00253_),
    .C(_00254_),
    .D(_08067_),
    .E(_08102_),
    .Y(_08110_));
 XOR2x2_ASAP7_75t_R _20575_ (.A(_00250_),
    .B(_08110_),
    .Y(_08111_));
 AND2x2_ASAP7_75t_R _20576_ (.A(_08096_),
    .B(_08111_),
    .Y(_04824_));
 OR5x2_ASAP7_75t_R _20577_ (.A(_00250_),
    .B(_00251_),
    .C(_00253_),
    .D(_00254_),
    .E(_08067_),
    .Y(_08112_));
 OR3x1_ASAP7_75t_R _20578_ (.A(_00249_),
    .B(_08099_),
    .C(_08112_),
    .Y(_08113_));
 OAI21x1_ASAP7_75t_R _20579_ (.A1(_08099_),
    .A2(_08112_),
    .B(_00249_),
    .Y(_08114_));
 AND3x1_ASAP7_75t_R _20580_ (.A(_08035_),
    .B(_08113_),
    .C(_08114_),
    .Y(_04825_));
 OR4x1_ASAP7_75t_R _20581_ (.A(_00248_),
    .B(_00249_),
    .C(_08102_),
    .D(_08112_),
    .Y(_08115_));
 OR3x1_ASAP7_75t_R _20582_ (.A(_00249_),
    .B(_08102_),
    .C(_08112_),
    .Y(_08116_));
 NAND2x1_ASAP7_75t_R _20583_ (.A(_00248_),
    .B(_08116_),
    .Y(_08117_));
 AND3x1_ASAP7_75t_R _20584_ (.A(_08035_),
    .B(_08115_),
    .C(_08117_),
    .Y(_04826_));
 OR4x1_ASAP7_75t_R _20585_ (.A(_00248_),
    .B(_00249_),
    .C(_08099_),
    .D(_08112_),
    .Y(_08118_));
 XOR2x2_ASAP7_75t_R _20586_ (.A(_08072_),
    .B(_08118_),
    .Y(_08119_));
 AND2x2_ASAP7_75t_R _20587_ (.A(_08096_),
    .B(_08119_),
    .Y(_04827_));
 OR3x1_ASAP7_75t_R _20588_ (.A(_00246_),
    .B(_08072_),
    .C(_08115_),
    .Y(_08120_));
 OAI21x1_ASAP7_75t_R _20589_ (.A1(_08072_),
    .A2(_08115_),
    .B(_00246_),
    .Y(_08121_));
 AND3x1_ASAP7_75t_R _20590_ (.A(_08035_),
    .B(_08120_),
    .C(_08121_),
    .Y(_04828_));
 OR3x1_ASAP7_75t_R _20591_ (.A(_00246_),
    .B(_08072_),
    .C(_08118_),
    .Y(_08122_));
 XOR2x2_ASAP7_75t_R _20592_ (.A(_00245_),
    .B(_08122_),
    .Y(_08123_));
 AND2x2_ASAP7_75t_R _20593_ (.A(_08096_),
    .B(_08123_),
    .Y(_04829_));
 OR4x1_ASAP7_75t_R _20594_ (.A(_00245_),
    .B(_00246_),
    .C(_08072_),
    .D(_08115_),
    .Y(_08124_));
 XOR2x2_ASAP7_75t_R _20595_ (.A(_00244_),
    .B(_08124_),
    .Y(_08125_));
 AND2x2_ASAP7_75t_R _20596_ (.A(_08096_),
    .B(_08125_),
    .Y(_04830_));
 OR5x1_ASAP7_75t_R _20597_ (.A(_00244_),
    .B(_00245_),
    .C(_00246_),
    .D(_08072_),
    .E(_08118_),
    .Y(_08126_));
 XOR2x2_ASAP7_75t_R _20598_ (.A(_00243_),
    .B(_08126_),
    .Y(_08127_));
 AND2x2_ASAP7_75t_R _20599_ (.A(_08096_),
    .B(_08127_),
    .Y(_04831_));
 OR5x2_ASAP7_75t_R _20600_ (.A(_00243_),
    .B(_00244_),
    .C(_00245_),
    .D(_00246_),
    .E(_08072_),
    .Y(_08128_));
 OR3x1_ASAP7_75t_R _20601_ (.A(_00242_),
    .B(_08115_),
    .C(_08128_),
    .Y(_08129_));
 OAI21x1_ASAP7_75t_R _20602_ (.A1(_08115_),
    .A2(_08128_),
    .B(_00242_),
    .Y(_08130_));
 AND3x1_ASAP7_75t_R _20603_ (.A(_08035_),
    .B(_08129_),
    .C(_08130_),
    .Y(_04832_));
 XOR2x2_ASAP7_75t_R _20604_ (.A(_00241_),
    .B(_02671_),
    .Y(_08131_));
 AND2x2_ASAP7_75t_R _20605_ (.A(_08096_),
    .B(_08131_),
    .Y(_04833_));
 BUFx6f_ASAP7_75t_R _20606_ (.A(_07689_),
    .Y(_08132_));
 OR3x1_ASAP7_75t_R _20607_ (.A(_00242_),
    .B(_08118_),
    .C(_08128_),
    .Y(_08133_));
 XOR2x2_ASAP7_75t_R _20608_ (.A(_00240_),
    .B(_08133_),
    .Y(_08134_));
 AND2x2_ASAP7_75t_R _20609_ (.A(_08132_),
    .B(_08134_),
    .Y(_04834_));
 OR4x1_ASAP7_75t_R _20610_ (.A(_00240_),
    .B(_00242_),
    .C(_08115_),
    .D(_08128_),
    .Y(_08135_));
 XOR2x2_ASAP7_75t_R _20611_ (.A(_00239_),
    .B(_08135_),
    .Y(_08136_));
 AND2x2_ASAP7_75t_R _20612_ (.A(_08132_),
    .B(_08136_),
    .Y(_04835_));
 OR3x1_ASAP7_75t_R _20613_ (.A(_00241_),
    .B(_00252_),
    .C(_00059_),
    .Y(_08137_));
 XOR2x2_ASAP7_75t_R _20614_ (.A(_00238_),
    .B(_08137_),
    .Y(_08138_));
 AND2x2_ASAP7_75t_R _20615_ (.A(_08132_),
    .B(_08138_),
    .Y(_04836_));
 OR3x1_ASAP7_75t_R _20616_ (.A(_00238_),
    .B(_00241_),
    .C(_02671_),
    .Y(_08139_));
 NAND2x1_ASAP7_75t_R _20617_ (.A(_00237_),
    .B(_08139_),
    .Y(_08140_));
 AND3x1_ASAP7_75t_R _20618_ (.A(_08035_),
    .B(_08080_),
    .C(_08140_),
    .Y(_04837_));
 XOR2x2_ASAP7_75t_R _20619_ (.A(_00236_),
    .B(_08085_),
    .Y(_08141_));
 AND2x2_ASAP7_75t_R _20620_ (.A(_08132_),
    .B(_08141_),
    .Y(_04838_));
 OR3x1_ASAP7_75t_R _20621_ (.A(_00235_),
    .B(_00236_),
    .C(_08080_),
    .Y(_08142_));
 OAI21x1_ASAP7_75t_R _20622_ (.A1(_00236_),
    .A2(_08080_),
    .B(_00235_),
    .Y(_08143_));
 AND3x1_ASAP7_75t_R _20623_ (.A(_08035_),
    .B(_08142_),
    .C(_08143_),
    .Y(_04839_));
 OR3x1_ASAP7_75t_R _20624_ (.A(_00235_),
    .B(_00236_),
    .C(_08085_),
    .Y(_08144_));
 XOR2x2_ASAP7_75t_R _20625_ (.A(_00234_),
    .B(_08144_),
    .Y(_08145_));
 AND2x2_ASAP7_75t_R _20626_ (.A(_08132_),
    .B(_08145_),
    .Y(_04840_));
 BUFx6f_ASAP7_75t_R _20627_ (.A(_08998_),
    .Y(_08146_));
 OR4x1_ASAP7_75t_R _20628_ (.A(_00234_),
    .B(_00235_),
    .C(_00236_),
    .D(_08080_),
    .Y(_08147_));
 NAND2x1_ASAP7_75t_R _20629_ (.A(_00233_),
    .B(_08147_),
    .Y(_08148_));
 AND3x1_ASAP7_75t_R _20630_ (.A(_08146_),
    .B(_08082_),
    .C(_08148_),
    .Y(_04841_));
 XOR2x2_ASAP7_75t_R _20631_ (.A(_08068_),
    .B(_08086_),
    .Y(_08149_));
 AND2x2_ASAP7_75t_R _20632_ (.A(_08132_),
    .B(_08149_),
    .Y(_04842_));
 BUFx3_ASAP7_75t_R _20633_ (.A(_00222_),
    .Y(_08150_));
 AND4x1_ASAP7_75t_R _20634_ (.A(_00193_),
    .B(_00221_),
    .C(_08150_),
    .D(_00223_),
    .Y(_08151_));
 AND5x1_ASAP7_75t_R _20635_ (.A(_00212_),
    .B(_00217_),
    .C(_00218_),
    .D(_00220_),
    .E(_08151_),
    .Y(_08152_));
 AND5x2_ASAP7_75t_R _20636_ (.A(_00214_),
    .B(_00215_),
    .C(_00216_),
    .D(_07147_),
    .E(_08152_),
    .Y(_08153_));
 BUFx3_ASAP7_75t_R _20637_ (.A(_00209_),
    .Y(_08154_));
 AND4x1_ASAP7_75t_R _20638_ (.A(_00207_),
    .B(_00208_),
    .C(_08154_),
    .D(_00210_),
    .Y(_08155_));
 AND4x1_ASAP7_75t_R _20639_ (.A(_00201_),
    .B(_00203_),
    .C(_00204_),
    .D(_00211_),
    .Y(_08156_));
 AND5x1_ASAP7_75t_R _20640_ (.A(_00194_),
    .B(_00195_),
    .C(_00200_),
    .D(_00219_),
    .E(_08156_),
    .Y(_08157_));
 BUFx6f_ASAP7_75t_R _20641_ (.A(_00197_),
    .Y(_08158_));
 AND3x1_ASAP7_75t_R _20642_ (.A(_00198_),
    .B(_00199_),
    .C(_00202_),
    .Y(_08159_));
 OR3x1_ASAP7_75t_R _20643_ (.A(_00196_),
    .B(_08158_),
    .C(_08159_),
    .Y(_08160_));
 AND5x2_ASAP7_75t_R _20644_ (.A(_00205_),
    .B(_00206_),
    .C(_08155_),
    .D(_08157_),
    .E(_08160_),
    .Y(_08161_));
 NAND2x2_ASAP7_75t_R _20645_ (.A(_08153_),
    .B(_08161_),
    .Y(_08162_));
 NOR2x1_ASAP7_75t_R _20646_ (.A(_00183_),
    .B(_08162_),
    .Y(_04843_));
 INVx1_ASAP7_75t_R _20647_ (.A(_08162_),
    .Y(_04844_));
 NOR2x1_ASAP7_75t_R _20648_ (.A(_00186_),
    .B(_08162_),
    .Y(_04845_));
 NOR2x1_ASAP7_75t_R _20649_ (.A(_00185_),
    .B(_08162_),
    .Y(_04846_));
 NOR2x1_ASAP7_75t_R _20650_ (.A(_00184_),
    .B(_08162_),
    .Y(_04847_));
 NOR2x1_ASAP7_75t_R _20651_ (.A(_00182_),
    .B(_08162_),
    .Y(_04848_));
 NOR2x1_ASAP7_75t_R _20652_ (.A(_00181_),
    .B(_08162_),
    .Y(_04849_));
 INVx1_ASAP7_75t_R _20653_ (.A(_08162_),
    .Y(_04850_));
 AND2x2_ASAP7_75t_R _20654_ (.A(_08132_),
    .B(_00060_),
    .Y(_04851_));
 OR4x1_ASAP7_75t_R _20655_ (.A(_00198_),
    .B(_00199_),
    .C(_00202_),
    .D(_02611_),
    .Y(_08163_));
 OR4x1_ASAP7_75t_R _20656_ (.A(_00194_),
    .B(_00195_),
    .C(_00196_),
    .D(_08158_),
    .Y(_08164_));
 OR4x1_ASAP7_75t_R _20657_ (.A(_00193_),
    .B(_00223_),
    .C(_08163_),
    .D(_08164_),
    .Y(_08165_));
 BUFx6f_ASAP7_75t_R _20658_ (.A(_08165_),
    .Y(_08166_));
 OR3x1_ASAP7_75t_R _20659_ (.A(_00193_),
    .B(_08163_),
    .C(_08164_),
    .Y(_08167_));
 NAND2x1_ASAP7_75t_R _20660_ (.A(_00223_),
    .B(_08167_),
    .Y(_08168_));
 AND3x1_ASAP7_75t_R _20661_ (.A(_08146_),
    .B(_08166_),
    .C(_08168_),
    .Y(_04852_));
 OR4x1_ASAP7_75t_R _20662_ (.A(_00193_),
    .B(_00194_),
    .C(_00196_),
    .D(_08158_),
    .Y(_08169_));
 OR5x2_ASAP7_75t_R _20663_ (.A(_00198_),
    .B(_00199_),
    .C(_00202_),
    .D(_00213_),
    .E(_00060_),
    .Y(_08170_));
 OR4x1_ASAP7_75t_R _20664_ (.A(_00195_),
    .B(_00223_),
    .C(_08169_),
    .D(_08170_),
    .Y(_08171_));
 XOR2x2_ASAP7_75t_R _20665_ (.A(_08150_),
    .B(_08171_),
    .Y(_08172_));
 AND2x2_ASAP7_75t_R _20666_ (.A(_08132_),
    .B(_08172_),
    .Y(_04853_));
 OR3x1_ASAP7_75t_R _20667_ (.A(_00221_),
    .B(_08150_),
    .C(_08166_),
    .Y(_08173_));
 OAI21x1_ASAP7_75t_R _20668_ (.A1(_08150_),
    .A2(_08166_),
    .B(_00221_),
    .Y(_08174_));
 AND3x1_ASAP7_75t_R _20669_ (.A(_08146_),
    .B(_08173_),
    .C(_08174_),
    .Y(_04854_));
 OR3x1_ASAP7_75t_R _20670_ (.A(_00221_),
    .B(_08150_),
    .C(_08171_),
    .Y(_08175_));
 XOR2x2_ASAP7_75t_R _20671_ (.A(_00220_),
    .B(_08175_),
    .Y(_08176_));
 AND2x2_ASAP7_75t_R _20672_ (.A(_08132_),
    .B(_08176_),
    .Y(_04855_));
 OR4x1_ASAP7_75t_R _20673_ (.A(_00220_),
    .B(_00221_),
    .C(_08150_),
    .D(_08166_),
    .Y(_08177_));
 XOR2x2_ASAP7_75t_R _20674_ (.A(_00219_),
    .B(_08177_),
    .Y(_08178_));
 AND2x2_ASAP7_75t_R _20675_ (.A(_08132_),
    .B(_08178_),
    .Y(_04856_));
 BUFx6f_ASAP7_75t_R _20676_ (.A(_07689_),
    .Y(_08179_));
 OR5x1_ASAP7_75t_R _20677_ (.A(_00219_),
    .B(_00220_),
    .C(_00221_),
    .D(_08150_),
    .E(_08171_),
    .Y(_08180_));
 XOR2x2_ASAP7_75t_R _20678_ (.A(_00218_),
    .B(_08180_),
    .Y(_08181_));
 AND2x2_ASAP7_75t_R _20679_ (.A(_08179_),
    .B(_08181_),
    .Y(_04857_));
 OR5x2_ASAP7_75t_R _20680_ (.A(_00218_),
    .B(_00219_),
    .C(_00220_),
    .D(_00221_),
    .E(_08150_),
    .Y(_08182_));
 OR3x1_ASAP7_75t_R _20681_ (.A(_00217_),
    .B(_08166_),
    .C(_08182_),
    .Y(_08183_));
 OAI21x1_ASAP7_75t_R _20682_ (.A1(_08166_),
    .A2(_08182_),
    .B(_00217_),
    .Y(_08184_));
 AND3x1_ASAP7_75t_R _20683_ (.A(_08146_),
    .B(_08183_),
    .C(_08184_),
    .Y(_04858_));
 OR3x2_ASAP7_75t_R _20684_ (.A(_00217_),
    .B(_08171_),
    .C(_08182_),
    .Y(_08185_));
 XOR2x2_ASAP7_75t_R _20685_ (.A(_00216_),
    .B(_08185_),
    .Y(_08186_));
 AND2x2_ASAP7_75t_R _20686_ (.A(_08179_),
    .B(_08186_),
    .Y(_04859_));
 OR4x1_ASAP7_75t_R _20687_ (.A(_00216_),
    .B(_00217_),
    .C(_08166_),
    .D(_08182_),
    .Y(_08187_));
 XOR2x2_ASAP7_75t_R _20688_ (.A(_00215_),
    .B(_08187_),
    .Y(_08188_));
 AND2x2_ASAP7_75t_R _20689_ (.A(_08179_),
    .B(_08188_),
    .Y(_04860_));
 OR3x1_ASAP7_75t_R _20690_ (.A(_00215_),
    .B(_00216_),
    .C(_08185_),
    .Y(_08189_));
 XOR2x2_ASAP7_75t_R _20691_ (.A(_00214_),
    .B(_08189_),
    .Y(_08190_));
 AND2x2_ASAP7_75t_R _20692_ (.A(_08179_),
    .B(_08190_),
    .Y(_04861_));
 NOR2x1_ASAP7_75t_R _20693_ (.A(_10986_),
    .B(_02612_),
    .Y(_04862_));
 OR3x1_ASAP7_75t_R _20694_ (.A(_00214_),
    .B(_00215_),
    .C(_08187_),
    .Y(_08191_));
 XOR2x2_ASAP7_75t_R _20695_ (.A(_00212_),
    .B(_08191_),
    .Y(_08192_));
 AND2x2_ASAP7_75t_R _20696_ (.A(_08179_),
    .B(_08192_),
    .Y(_04863_));
 OR2x2_ASAP7_75t_R _20697_ (.A(_00216_),
    .B(_08185_),
    .Y(_08193_));
 OR4x1_ASAP7_75t_R _20698_ (.A(_00212_),
    .B(_00214_),
    .C(_00215_),
    .D(_08193_),
    .Y(_08194_));
 XOR2x2_ASAP7_75t_R _20699_ (.A(_00211_),
    .B(_08194_),
    .Y(_08195_));
 AND2x2_ASAP7_75t_R _20700_ (.A(_08179_),
    .B(_08195_),
    .Y(_04864_));
 OR5x1_ASAP7_75t_R _20701_ (.A(_00210_),
    .B(_00211_),
    .C(_00212_),
    .D(_00214_),
    .E(_00215_),
    .Y(_08196_));
 OR5x2_ASAP7_75t_R _20702_ (.A(_00216_),
    .B(_00217_),
    .C(_08166_),
    .D(_08182_),
    .E(_08196_),
    .Y(_08197_));
 OR5x1_ASAP7_75t_R _20703_ (.A(_00211_),
    .B(_00212_),
    .C(_00214_),
    .D(_00215_),
    .E(_08187_),
    .Y(_08198_));
 NAND2x1_ASAP7_75t_R _20704_ (.A(_00210_),
    .B(_08198_),
    .Y(_08199_));
 AND3x1_ASAP7_75t_R _20705_ (.A(_08146_),
    .B(_08197_),
    .C(_08199_),
    .Y(_04865_));
 OR5x2_ASAP7_75t_R _20706_ (.A(_00216_),
    .B(_00217_),
    .C(_08171_),
    .D(_08182_),
    .E(_08196_),
    .Y(_08200_));
 XOR2x2_ASAP7_75t_R _20707_ (.A(_08154_),
    .B(_08200_),
    .Y(_08201_));
 AND2x2_ASAP7_75t_R _20708_ (.A(_08179_),
    .B(_08201_),
    .Y(_04866_));
 OR3x1_ASAP7_75t_R _20709_ (.A(_00208_),
    .B(_08154_),
    .C(_08197_),
    .Y(_08202_));
 OAI21x1_ASAP7_75t_R _20710_ (.A1(_08154_),
    .A2(_08197_),
    .B(_00208_),
    .Y(_08203_));
 AND3x1_ASAP7_75t_R _20711_ (.A(_08146_),
    .B(_08202_),
    .C(_08203_),
    .Y(_04867_));
 OR3x1_ASAP7_75t_R _20712_ (.A(_00208_),
    .B(_08154_),
    .C(_08200_),
    .Y(_08204_));
 XOR2x2_ASAP7_75t_R _20713_ (.A(_00207_),
    .B(_08204_),
    .Y(_08205_));
 AND2x2_ASAP7_75t_R _20714_ (.A(_08179_),
    .B(_08205_),
    .Y(_04868_));
 OR5x2_ASAP7_75t_R _20715_ (.A(_00206_),
    .B(_00207_),
    .C(_00208_),
    .D(_08154_),
    .E(_08197_),
    .Y(_08206_));
 OR4x1_ASAP7_75t_R _20716_ (.A(_00207_),
    .B(_00208_),
    .C(_08154_),
    .D(_08197_),
    .Y(_08207_));
 NAND2x1_ASAP7_75t_R _20717_ (.A(_00206_),
    .B(_08207_),
    .Y(_08208_));
 AND3x1_ASAP7_75t_R _20718_ (.A(_08146_),
    .B(_08206_),
    .C(_08208_),
    .Y(_04869_));
 OR5x2_ASAP7_75t_R _20719_ (.A(_00206_),
    .B(_00207_),
    .C(_00208_),
    .D(_08154_),
    .E(_08200_),
    .Y(_08209_));
 XOR2x2_ASAP7_75t_R _20720_ (.A(_00205_),
    .B(_08209_),
    .Y(_08210_));
 AND2x2_ASAP7_75t_R _20721_ (.A(_08179_),
    .B(_08210_),
    .Y(_04870_));
 OR3x1_ASAP7_75t_R _20722_ (.A(_00204_),
    .B(_00205_),
    .C(_08206_),
    .Y(_08211_));
 OAI21x1_ASAP7_75t_R _20723_ (.A1(_00205_),
    .A2(_08206_),
    .B(_00204_),
    .Y(_08212_));
 AND3x1_ASAP7_75t_R _20724_ (.A(_08146_),
    .B(_08211_),
    .C(_08212_),
    .Y(_04871_));
 OR3x1_ASAP7_75t_R _20725_ (.A(_00204_),
    .B(_00205_),
    .C(_08209_),
    .Y(_08213_));
 XOR2x2_ASAP7_75t_R _20726_ (.A(_00203_),
    .B(_08213_),
    .Y(_08214_));
 AND2x2_ASAP7_75t_R _20727_ (.A(_08179_),
    .B(_08214_),
    .Y(_04872_));
 BUFx6f_ASAP7_75t_R _20728_ (.A(_09029_),
    .Y(_08215_));
 XOR2x2_ASAP7_75t_R _20729_ (.A(_00202_),
    .B(_02611_),
    .Y(_08216_));
 AND2x2_ASAP7_75t_R _20730_ (.A(_08215_),
    .B(_08216_),
    .Y(_04873_));
 OR4x1_ASAP7_75t_R _20731_ (.A(_00203_),
    .B(_00204_),
    .C(_00205_),
    .D(_08206_),
    .Y(_08217_));
 XOR2x2_ASAP7_75t_R _20732_ (.A(_00201_),
    .B(_08217_),
    .Y(_08218_));
 AND2x2_ASAP7_75t_R _20733_ (.A(_08215_),
    .B(_08218_),
    .Y(_04874_));
 OR5x1_ASAP7_75t_R _20734_ (.A(_00201_),
    .B(_00203_),
    .C(_00204_),
    .D(_00205_),
    .E(_08209_),
    .Y(_08219_));
 XOR2x2_ASAP7_75t_R _20735_ (.A(_00200_),
    .B(_08219_),
    .Y(_08220_));
 AND2x2_ASAP7_75t_R _20736_ (.A(_08215_),
    .B(_08220_),
    .Y(_04875_));
 OR3x1_ASAP7_75t_R _20737_ (.A(_00202_),
    .B(_00213_),
    .C(_00060_),
    .Y(_08221_));
 XOR2x2_ASAP7_75t_R _20738_ (.A(_00199_),
    .B(_08221_),
    .Y(_08222_));
 AND2x2_ASAP7_75t_R _20739_ (.A(_08215_),
    .B(_08222_),
    .Y(_04876_));
 OR3x1_ASAP7_75t_R _20740_ (.A(_00199_),
    .B(_00202_),
    .C(_02611_),
    .Y(_08223_));
 NAND2x1_ASAP7_75t_R _20741_ (.A(_00198_),
    .B(_08223_),
    .Y(_08224_));
 AND3x1_ASAP7_75t_R _20742_ (.A(_08146_),
    .B(_08163_),
    .C(_08224_),
    .Y(_04877_));
 XOR2x2_ASAP7_75t_R _20743_ (.A(_08158_),
    .B(_08170_),
    .Y(_08225_));
 AND2x2_ASAP7_75t_R _20744_ (.A(_08215_),
    .B(_08225_),
    .Y(_04878_));
 OR3x1_ASAP7_75t_R _20745_ (.A(_00196_),
    .B(_08158_),
    .C(_08163_),
    .Y(_08226_));
 OAI21x1_ASAP7_75t_R _20746_ (.A1(_08158_),
    .A2(_08163_),
    .B(_00196_),
    .Y(_08227_));
 AND3x1_ASAP7_75t_R _20747_ (.A(_08146_),
    .B(_08226_),
    .C(_08227_),
    .Y(_04879_));
 OR3x1_ASAP7_75t_R _20748_ (.A(_00196_),
    .B(_08158_),
    .C(_08170_),
    .Y(_08228_));
 XOR2x2_ASAP7_75t_R _20749_ (.A(_00195_),
    .B(_08228_),
    .Y(_08229_));
 AND2x2_ASAP7_75t_R _20750_ (.A(_08215_),
    .B(_08229_),
    .Y(_04880_));
 OR4x1_ASAP7_75t_R _20751_ (.A(_00195_),
    .B(_00196_),
    .C(_08158_),
    .D(_08163_),
    .Y(_08230_));
 NAND2x1_ASAP7_75t_R _20752_ (.A(_00194_),
    .B(_08230_),
    .Y(_08231_));
 OA211x2_ASAP7_75t_R _20753_ (.A1(_08163_),
    .A2(_08164_),
    .B(_08231_),
    .C(_07260_),
    .Y(_04881_));
 BUFx6f_ASAP7_75t_R _20754_ (.A(_08998_),
    .Y(_08232_));
 OR3x1_ASAP7_75t_R _20755_ (.A(_00193_),
    .B(_08164_),
    .C(_08170_),
    .Y(_08233_));
 OAI21x1_ASAP7_75t_R _20756_ (.A1(_08164_),
    .A2(_08170_),
    .B(_00193_),
    .Y(_08234_));
 AND3x1_ASAP7_75t_R _20757_ (.A(_08232_),
    .B(_08233_),
    .C(_08234_),
    .Y(_04882_));
 AND2x2_ASAP7_75t_R _20758_ (.A(_08215_),
    .B(_00029_),
    .Y(_04883_));
 AND2x4_ASAP7_75t_R _20759_ (.A(_00226_),
    .B(_00227_),
    .Y(_08235_));
 AND5x2_ASAP7_75t_R _20760_ (.A(\xs[8].cli1.i[39] ),
    .B(\xs[8].cli1.i[36] ),
    .C(_00228_),
    .D(_00229_),
    .E(_08235_),
    .Y(_08236_));
 NAND2x1_ASAP7_75t_R _20761_ (.A(_00226_),
    .B(_00227_),
    .Y(_08237_));
 OA31x2_ASAP7_75t_R _20762_ (.A1(_00225_),
    .A2(\xs[8].cli1.i[33] ),
    .A3(_08237_),
    .B1(\xs[8].cli1.i[39] ),
    .Y(_08238_));
 BUFx3_ASAP7_75t_R _20763_ (.A(_02163_),
    .Y(_08239_));
 NOR2x1_ASAP7_75t_R _20764_ (.A(_02162_),
    .B(_08239_),
    .Y(_08240_));
 OA21x2_ASAP7_75t_R _20765_ (.A1(_08236_),
    .A2(_08238_),
    .B(_02169_),
    .Y(_08241_));
 INVx1_ASAP7_75t_R _20766_ (.A(_08239_),
    .Y(_08242_));
 AO21x1_ASAP7_75t_R _20767_ (.A1(_08242_),
    .A2(_08236_),
    .B(_02162_),
    .Y(_08243_));
 INVx2_ASAP7_75t_R _20768_ (.A(_02162_),
    .Y(_08244_));
 AO21x1_ASAP7_75t_R _20769_ (.A1(_00029_),
    .A2(_08238_),
    .B(_08244_),
    .Y(_08245_));
 NAND2x1_ASAP7_75t_R _20770_ (.A(_00266_),
    .B(_00267_),
    .Y(_08246_));
 OA31x2_ASAP7_75t_R _20771_ (.A1(_00264_),
    .A2(\peo[16][35] ),
    .A3(_08246_),
    .B1(\peo[16][39] ),
    .Y(_08247_));
 OA211x2_ASAP7_75t_R _20772_ (.A1(_08241_),
    .A2(_08243_),
    .B(_08245_),
    .C(_08247_),
    .Y(_08248_));
 AOI21x1_ASAP7_75t_R _20773_ (.A1(_08238_),
    .A2(_08240_),
    .B(_08248_),
    .Y(_08249_));
 NOR2x1_ASAP7_75t_R _20774_ (.A(_09314_),
    .B(_00231_),
    .Y(_08250_));
 AOI21x1_ASAP7_75t_R _20775_ (.A1(_08236_),
    .A2(_08249_),
    .B(_09818_),
    .Y(_08251_));
 AND2x2_ASAP7_75t_R _20776_ (.A(_00266_),
    .B(_00267_),
    .Y(_08252_));
 AO31x2_ASAP7_75t_R _20777_ (.A1(\peo[16][36] ),
    .A2(_00265_),
    .A3(_08252_),
    .B(_00263_),
    .Y(_08253_));
 AO21x1_ASAP7_75t_R _20778_ (.A1(\peo[16][39] ),
    .A2(\peo[16][32] ),
    .B(_02169_),
    .Y(_08254_));
 AND2x2_ASAP7_75t_R _20779_ (.A(_08253_),
    .B(_08254_),
    .Y(_08255_));
 INVx2_ASAP7_75t_R _20780_ (.A(_02169_),
    .Y(_08256_));
 AO31x2_ASAP7_75t_R _20781_ (.A1(\xs[8].cli1.i[36] ),
    .A2(_00228_),
    .A3(_08235_),
    .B(_00224_),
    .Y(_08257_));
 AO21x1_ASAP7_75t_R _20782_ (.A1(_08256_),
    .A2(_08257_),
    .B(_08236_),
    .Y(_08258_));
 NAND2x1_ASAP7_75t_R _20783_ (.A(_08255_),
    .B(_08258_),
    .Y(_08259_));
 AND2x2_ASAP7_75t_R _20784_ (.A(_08244_),
    .B(_08239_),
    .Y(_08260_));
 AND4x1_ASAP7_75t_R _20785_ (.A(_02169_),
    .B(_02173_),
    .C(_08259_),
    .D(_08260_),
    .Y(_08261_));
 NAND2x1_ASAP7_75t_R _20786_ (.A(_08244_),
    .B(_08239_),
    .Y(_08262_));
 AO21x2_ASAP7_75t_R _20787_ (.A1(_08255_),
    .A2(_08258_),
    .B(_08262_),
    .Y(_08263_));
 OA21x2_ASAP7_75t_R _20788_ (.A1(_08256_),
    .A2(_08263_),
    .B(_00270_),
    .Y(_08264_));
 NOR2x1_ASAP7_75t_R _20789_ (.A(_08261_),
    .B(_08264_),
    .Y(_08265_));
 AO32x1_ASAP7_75t_R _20790_ (.A1(_08236_),
    .A2(_08249_),
    .A3(_08250_),
    .B1(_08251_),
    .B2(_08265_),
    .Y(_04884_));
 OR3x2_ASAP7_75t_R _20791_ (.A(_11177_),
    .B(_08256_),
    .C(_08263_),
    .Y(_08266_));
 NOR2x1_ASAP7_75t_R _20792_ (.A(_02172_),
    .B(_08266_),
    .Y(_04885_));
 NOR2x1_ASAP7_75t_R _20793_ (.A(_02171_),
    .B(_08266_),
    .Y(_04886_));
 NOR2x1_ASAP7_75t_R _20794_ (.A(_02170_),
    .B(_08266_),
    .Y(_04887_));
 NOR2x1_ASAP7_75t_R _20795_ (.A(_02161_),
    .B(_08266_),
    .Y(_04888_));
 NOR2x1_ASAP7_75t_R _20796_ (.A(_02160_),
    .B(_08266_),
    .Y(_04889_));
 AND4x1_ASAP7_75t_R _20797_ (.A(_08256_),
    .B(_02173_),
    .C(_08259_),
    .D(_08260_),
    .Y(_08267_));
 OA21x2_ASAP7_75t_R _20798_ (.A1(_02169_),
    .A2(_08263_),
    .B(_00270_),
    .Y(_08268_));
 OAI21x1_ASAP7_75t_R _20799_ (.A1(_08267_),
    .A2(_08268_),
    .B(_08249_),
    .Y(_08269_));
 OA211x2_ASAP7_75t_R _20800_ (.A1(\peo[17][0] ),
    .A2(_08249_),
    .B(_08269_),
    .C(_07260_),
    .Y(_04890_));
 OR3x2_ASAP7_75t_R _20801_ (.A(_11177_),
    .B(_02169_),
    .C(_08263_),
    .Y(_08270_));
 NOR2x1_ASAP7_75t_R _20802_ (.A(_02172_),
    .B(_08270_),
    .Y(_04891_));
 NOR2x1_ASAP7_75t_R _20803_ (.A(_02171_),
    .B(_08270_),
    .Y(_04892_));
 NOR2x1_ASAP7_75t_R _20804_ (.A(_02170_),
    .B(_08270_),
    .Y(_04893_));
 NOR2x1_ASAP7_75t_R _20805_ (.A(_02161_),
    .B(_08270_),
    .Y(_04894_));
 NOR2x1_ASAP7_75t_R _20806_ (.A(_02160_),
    .B(_08270_),
    .Y(_04895_));
 AO21x1_ASAP7_75t_R _20807_ (.A1(_08239_),
    .A2(_08259_),
    .B(_02162_),
    .Y(_08271_));
 BUFx6f_ASAP7_75t_R _20808_ (.A(_08271_),
    .Y(_08272_));
 NOR2x1_ASAP7_75t_R _20809_ (.A(_02173_),
    .B(_08272_),
    .Y(_08273_));
 AND2x2_ASAP7_75t_R _20810_ (.A(_08244_),
    .B(_08247_),
    .Y(_08274_));
 OR2x2_ASAP7_75t_R _20811_ (.A(_08257_),
    .B(_08240_),
    .Y(_08275_));
 AND3x1_ASAP7_75t_R _20812_ (.A(_02162_),
    .B(_00029_),
    .C(_08247_),
    .Y(_08276_));
 AOI211x1_ASAP7_75t_R _20813_ (.A1(_08241_),
    .A2(_08274_),
    .B(_08275_),
    .C(_08276_),
    .Y(_08277_));
 NAND2x1_ASAP7_75t_R _20814_ (.A(_00231_),
    .B(_08277_),
    .Y(_08278_));
 OA211x2_ASAP7_75t_R _20815_ (.A1(\peo[16][0] ),
    .A2(_08277_),
    .B(_08278_),
    .C(_08272_),
    .Y(_08279_));
 OA21x2_ASAP7_75t_R _20816_ (.A1(_08273_),
    .A2(_08279_),
    .B(_08529_),
    .Y(_04896_));
 AOI21x1_ASAP7_75t_R _20817_ (.A1(_08239_),
    .A2(_08259_),
    .B(_02162_),
    .Y(_08280_));
 NAND2x2_ASAP7_75t_R _20818_ (.A(_08584_),
    .B(_08280_),
    .Y(_08281_));
 NOR2x1_ASAP7_75t_R _20819_ (.A(_02172_),
    .B(_08281_),
    .Y(_04897_));
 NOR2x1_ASAP7_75t_R _20820_ (.A(_02171_),
    .B(_08281_),
    .Y(_04898_));
 NOR2x1_ASAP7_75t_R _20821_ (.A(_02170_),
    .B(_08281_),
    .Y(_04899_));
 AND2x2_ASAP7_75t_R _20822_ (.A(_08256_),
    .B(_08280_),
    .Y(_08282_));
 NAND2x1_ASAP7_75t_R _20823_ (.A(_00229_),
    .B(_08277_),
    .Y(_08283_));
 OA211x2_ASAP7_75t_R _20824_ (.A1(\peo[16][32] ),
    .A2(_08277_),
    .B(_08283_),
    .C(_08272_),
    .Y(_08284_));
 OA21x2_ASAP7_75t_R _20825_ (.A1(_08282_),
    .A2(_08284_),
    .B(_08529_),
    .Y(_04900_));
 NOR2x1_ASAP7_75t_R _20826_ (.A(_02168_),
    .B(_08272_),
    .Y(_08285_));
 NAND2x1_ASAP7_75t_R _20827_ (.A(_00228_),
    .B(_08277_),
    .Y(_08286_));
 OA211x2_ASAP7_75t_R _20828_ (.A1(\peo[16][33] ),
    .A2(_08277_),
    .B(_08286_),
    .C(_08272_),
    .Y(_08287_));
 OA21x2_ASAP7_75t_R _20829_ (.A1(_08285_),
    .A2(_08287_),
    .B(_08529_),
    .Y(_04901_));
 NOR2x1_ASAP7_75t_R _20830_ (.A(_02167_),
    .B(_08272_),
    .Y(_08288_));
 NAND2x1_ASAP7_75t_R _20831_ (.A(_00227_),
    .B(_08277_),
    .Y(_08289_));
 OA211x2_ASAP7_75t_R _20832_ (.A1(\peo[16][34] ),
    .A2(_08277_),
    .B(_08289_),
    .C(_08272_),
    .Y(_08290_));
 OA21x2_ASAP7_75t_R _20833_ (.A1(_08288_),
    .A2(_08290_),
    .B(_08529_),
    .Y(_04902_));
 NOR2x1_ASAP7_75t_R _20834_ (.A(_02166_),
    .B(_08272_),
    .Y(_08291_));
 NAND2x1_ASAP7_75t_R _20835_ (.A(_00226_),
    .B(_08277_),
    .Y(_08292_));
 OA211x2_ASAP7_75t_R _20836_ (.A1(\peo[16][35] ),
    .A2(_08277_),
    .B(_08292_),
    .C(_08272_),
    .Y(_08293_));
 OA21x2_ASAP7_75t_R _20837_ (.A1(_08291_),
    .A2(_08293_),
    .B(_08529_),
    .Y(_04903_));
 OA21x2_ASAP7_75t_R _20838_ (.A1(_08257_),
    .A2(_08248_),
    .B(_00264_),
    .Y(_08294_));
 NOR3x1_ASAP7_75t_R _20839_ (.A(_00224_),
    .B(\xs[8].cli1.i[36] ),
    .C(_08248_),
    .Y(_08295_));
 OR4x1_ASAP7_75t_R _20840_ (.A(_09314_),
    .B(_08280_),
    .C(_08294_),
    .D(_08295_),
    .Y(_08296_));
 OAI21x1_ASAP7_75t_R _20841_ (.A1(_02165_),
    .A2(_08281_),
    .B(_08296_),
    .Y(_04904_));
 NOR2x1_ASAP7_75t_R _20842_ (.A(_02164_),
    .B(_08281_),
    .Y(_04905_));
 OR3x1_ASAP7_75t_R _20843_ (.A(_08642_),
    .B(_08259_),
    .C(_08262_),
    .Y(_08297_));
 INVx1_ASAP7_75t_R _20844_ (.A(_08297_),
    .Y(_04906_));
 AND3x1_ASAP7_75t_R _20845_ (.A(_08253_),
    .B(_08257_),
    .C(_08272_),
    .Y(_08298_));
 NOR2x1_ASAP7_75t_R _20846_ (.A(_10986_),
    .B(_08298_),
    .Y(_04907_));
 NOR2x1_ASAP7_75t_R _20847_ (.A(_02161_),
    .B(_08281_),
    .Y(_04908_));
 NOR2x1_ASAP7_75t_R _20848_ (.A(_02160_),
    .B(_08281_),
    .Y(_04909_));
 BUFx3_ASAP7_75t_R _20849_ (.A(_00155_),
    .Y(_08299_));
 BUFx3_ASAP7_75t_R _20850_ (.A(_00128_),
    .Y(_08300_));
 AND4x1_ASAP7_75t_R _20851_ (.A(_08300_),
    .B(_00156_),
    .C(_00157_),
    .D(_00158_),
    .Y(_08301_));
 AND5x1_ASAP7_75t_R _20852_ (.A(_00147_),
    .B(_00152_),
    .C(_00153_),
    .D(_08299_),
    .E(_08301_),
    .Y(_08302_));
 AND5x2_ASAP7_75t_R _20853_ (.A(_00149_),
    .B(_00150_),
    .C(_00151_),
    .D(_11465_),
    .E(_08302_),
    .Y(_08303_));
 AND4x1_ASAP7_75t_R _20854_ (.A(_00142_),
    .B(_00143_),
    .C(_00144_),
    .D(_00145_),
    .Y(_08304_));
 AND4x1_ASAP7_75t_R _20855_ (.A(_00136_),
    .B(_00138_),
    .C(_00139_),
    .D(_00146_),
    .Y(_08305_));
 AND5x1_ASAP7_75t_R _20856_ (.A(_00129_),
    .B(_00130_),
    .C(_00135_),
    .D(_00154_),
    .E(_08305_),
    .Y(_08306_));
 AND3x1_ASAP7_75t_R _20857_ (.A(_00133_),
    .B(_00134_),
    .C(_00137_),
    .Y(_08307_));
 OR3x1_ASAP7_75t_R _20858_ (.A(_00131_),
    .B(_00132_),
    .C(_08307_),
    .Y(_08308_));
 AND5x2_ASAP7_75t_R _20859_ (.A(_00140_),
    .B(_00141_),
    .C(_08304_),
    .D(_08306_),
    .E(_08308_),
    .Y(_08309_));
 NAND2x2_ASAP7_75t_R _20860_ (.A(_08303_),
    .B(_08309_),
    .Y(_08310_));
 NOR2x1_ASAP7_75t_R _20861_ (.A(_00085_),
    .B(_08310_),
    .Y(_04910_));
 INVx1_ASAP7_75t_R _20862_ (.A(_08310_),
    .Y(_04911_));
 NOR2x1_ASAP7_75t_R _20863_ (.A(_00088_),
    .B(_08310_),
    .Y(_04912_));
 NOR2x1_ASAP7_75t_R _20864_ (.A(_00087_),
    .B(_08310_),
    .Y(_04913_));
 NOR2x1_ASAP7_75t_R _20865_ (.A(_00086_),
    .B(_08310_),
    .Y(_04914_));
 NOR2x1_ASAP7_75t_R _20866_ (.A(_00084_),
    .B(_08310_),
    .Y(_04915_));
 NOR2x1_ASAP7_75t_R _20867_ (.A(_00083_),
    .B(_08310_),
    .Y(_04916_));
 INVx1_ASAP7_75t_R _20868_ (.A(_08310_),
    .Y(_04917_));
 AND2x2_ASAP7_75t_R _20869_ (.A(_08215_),
    .B(_00061_),
    .Y(_04918_));
 OR4x1_ASAP7_75t_R _20870_ (.A(_00133_),
    .B(_00134_),
    .C(_00137_),
    .D(_02647_),
    .Y(_08311_));
 OR4x1_ASAP7_75t_R _20871_ (.A(_00129_),
    .B(_00130_),
    .C(_00131_),
    .D(_00132_),
    .Y(_08312_));
 OR2x6_ASAP7_75t_R _20872_ (.A(_08311_),
    .B(_08312_),
    .Y(_08313_));
 OR3x1_ASAP7_75t_R _20873_ (.A(_08300_),
    .B(_00158_),
    .C(_08313_),
    .Y(_08314_));
 OAI21x1_ASAP7_75t_R _20874_ (.A1(_08300_),
    .A2(_08313_),
    .B(_00158_),
    .Y(_08315_));
 AND3x1_ASAP7_75t_R _20875_ (.A(_08232_),
    .B(_08314_),
    .C(_08315_),
    .Y(_04919_));
 OR5x2_ASAP7_75t_R _20876_ (.A(_00133_),
    .B(_00134_),
    .C(_00137_),
    .D(_00148_),
    .E(_00061_),
    .Y(_08316_));
 OR2x2_ASAP7_75t_R _20877_ (.A(_08312_),
    .B(_08316_),
    .Y(_08317_));
 OR3x1_ASAP7_75t_R _20878_ (.A(_08300_),
    .B(_00158_),
    .C(_08317_),
    .Y(_08318_));
 XOR2x2_ASAP7_75t_R _20879_ (.A(_00157_),
    .B(_08318_),
    .Y(_08319_));
 AND2x2_ASAP7_75t_R _20880_ (.A(_08215_),
    .B(_08319_),
    .Y(_04920_));
 OR4x1_ASAP7_75t_R _20881_ (.A(_08300_),
    .B(_00156_),
    .C(_00157_),
    .D(_00158_),
    .Y(_08320_));
 OR3x2_ASAP7_75t_R _20882_ (.A(_08311_),
    .B(_08312_),
    .C(_08320_),
    .Y(_08321_));
 OR4x1_ASAP7_75t_R _20883_ (.A(_08300_),
    .B(_00157_),
    .C(_00158_),
    .D(_08313_),
    .Y(_08322_));
 NAND2x1_ASAP7_75t_R _20884_ (.A(_00156_),
    .B(_08322_),
    .Y(_08323_));
 AND3x1_ASAP7_75t_R _20885_ (.A(_08232_),
    .B(_08321_),
    .C(_08323_),
    .Y(_04921_));
 OR3x2_ASAP7_75t_R _20886_ (.A(_08312_),
    .B(_08316_),
    .C(_08320_),
    .Y(_08324_));
 XOR2x2_ASAP7_75t_R _20887_ (.A(_08299_),
    .B(_08324_),
    .Y(_08325_));
 AND2x2_ASAP7_75t_R _20888_ (.A(_08215_),
    .B(_08325_),
    .Y(_04922_));
 OR3x1_ASAP7_75t_R _20889_ (.A(_00154_),
    .B(_08299_),
    .C(_08321_),
    .Y(_08326_));
 OAI21x1_ASAP7_75t_R _20890_ (.A1(_08299_),
    .A2(_08321_),
    .B(_00154_),
    .Y(_08327_));
 AND3x1_ASAP7_75t_R _20891_ (.A(_08232_),
    .B(_08326_),
    .C(_08327_),
    .Y(_04923_));
 BUFx6f_ASAP7_75t_R _20892_ (.A(_09029_),
    .Y(_08328_));
 OR3x1_ASAP7_75t_R _20893_ (.A(_00154_),
    .B(_08299_),
    .C(_08324_),
    .Y(_08329_));
 XOR2x2_ASAP7_75t_R _20894_ (.A(_00153_),
    .B(_08329_),
    .Y(_08330_));
 AND2x2_ASAP7_75t_R _20895_ (.A(_08328_),
    .B(_08330_),
    .Y(_04924_));
 OR4x1_ASAP7_75t_R _20896_ (.A(_00153_),
    .B(_00154_),
    .C(_08299_),
    .D(_08321_),
    .Y(_08331_));
 XOR2x2_ASAP7_75t_R _20897_ (.A(_00152_),
    .B(_08331_),
    .Y(_08332_));
 AND2x2_ASAP7_75t_R _20898_ (.A(_08328_),
    .B(_08332_),
    .Y(_04925_));
 OR5x1_ASAP7_75t_R _20899_ (.A(_00152_),
    .B(_00153_),
    .C(_00154_),
    .D(_08299_),
    .E(_08324_),
    .Y(_08333_));
 XOR2x2_ASAP7_75t_R _20900_ (.A(_00151_),
    .B(_08333_),
    .Y(_08334_));
 AND2x2_ASAP7_75t_R _20901_ (.A(_08328_),
    .B(_08334_),
    .Y(_04926_));
 OR5x2_ASAP7_75t_R _20902_ (.A(_00151_),
    .B(_00152_),
    .C(_00153_),
    .D(_00154_),
    .E(_08299_),
    .Y(_08335_));
 OR3x2_ASAP7_75t_R _20903_ (.A(_00150_),
    .B(_08321_),
    .C(_08335_),
    .Y(_08336_));
 OAI21x1_ASAP7_75t_R _20904_ (.A1(_08321_),
    .A2(_08335_),
    .B(_00150_),
    .Y(_08337_));
 AND3x1_ASAP7_75t_R _20905_ (.A(_08232_),
    .B(_08336_),
    .C(_08337_),
    .Y(_04927_));
 OR3x2_ASAP7_75t_R _20906_ (.A(_00150_),
    .B(_08324_),
    .C(_08335_),
    .Y(_08338_));
 XOR2x2_ASAP7_75t_R _20907_ (.A(_00149_),
    .B(_08338_),
    .Y(_08339_));
 AND2x2_ASAP7_75t_R _20908_ (.A(_08328_),
    .B(_08339_),
    .Y(_04928_));
 NOR2x1_ASAP7_75t_R _20909_ (.A(_10986_),
    .B(_02648_),
    .Y(_04929_));
 OR3x1_ASAP7_75t_R _20910_ (.A(_00147_),
    .B(_00149_),
    .C(_08336_),
    .Y(_08340_));
 OAI21x1_ASAP7_75t_R _20911_ (.A1(_00149_),
    .A2(_08336_),
    .B(_00147_),
    .Y(_08341_));
 AND3x1_ASAP7_75t_R _20912_ (.A(_08232_),
    .B(_08340_),
    .C(_08341_),
    .Y(_04930_));
 OR3x1_ASAP7_75t_R _20913_ (.A(_00147_),
    .B(_00149_),
    .C(_08338_),
    .Y(_08342_));
 XOR2x2_ASAP7_75t_R _20914_ (.A(_00146_),
    .B(_08342_),
    .Y(_08343_));
 AND2x2_ASAP7_75t_R _20915_ (.A(_08328_),
    .B(_08343_),
    .Y(_04931_));
 OR4x1_ASAP7_75t_R _20916_ (.A(_00146_),
    .B(_00147_),
    .C(_00149_),
    .D(_08336_),
    .Y(_08344_));
 XOR2x2_ASAP7_75t_R _20917_ (.A(_00145_),
    .B(_08344_),
    .Y(_08345_));
 AND2x2_ASAP7_75t_R _20918_ (.A(_08328_),
    .B(_08345_),
    .Y(_04932_));
 OR4x1_ASAP7_75t_R _20919_ (.A(_00145_),
    .B(_00146_),
    .C(_00147_),
    .D(_00149_),
    .Y(_08346_));
 OR3x2_ASAP7_75t_R _20920_ (.A(_00144_),
    .B(_08338_),
    .C(_08346_),
    .Y(_08347_));
 OAI21x1_ASAP7_75t_R _20921_ (.A1(_08338_),
    .A2(_08346_),
    .B(_00144_),
    .Y(_08348_));
 AND3x1_ASAP7_75t_R _20922_ (.A(_08232_),
    .B(_08347_),
    .C(_08348_),
    .Y(_04933_));
 OR3x2_ASAP7_75t_R _20923_ (.A(_00144_),
    .B(_08336_),
    .C(_08346_),
    .Y(_08349_));
 XOR2x2_ASAP7_75t_R _20924_ (.A(_00143_),
    .B(_08349_),
    .Y(_08350_));
 AND2x2_ASAP7_75t_R _20925_ (.A(_08328_),
    .B(_08350_),
    .Y(_04934_));
 OR3x1_ASAP7_75t_R _20926_ (.A(_00142_),
    .B(_00143_),
    .C(_08347_),
    .Y(_08351_));
 OAI21x1_ASAP7_75t_R _20927_ (.A1(_00143_),
    .A2(_08347_),
    .B(_00142_),
    .Y(_08352_));
 AND3x1_ASAP7_75t_R _20928_ (.A(_08232_),
    .B(_08351_),
    .C(_08352_),
    .Y(_04935_));
 OR3x1_ASAP7_75t_R _20929_ (.A(_00142_),
    .B(_00143_),
    .C(_08349_),
    .Y(_08353_));
 XOR2x2_ASAP7_75t_R _20930_ (.A(_00141_),
    .B(_08353_),
    .Y(_08354_));
 AND2x2_ASAP7_75t_R _20931_ (.A(_08328_),
    .B(_08354_),
    .Y(_04936_));
 OR4x1_ASAP7_75t_R _20932_ (.A(_00141_),
    .B(_00142_),
    .C(_00143_),
    .D(_08347_),
    .Y(_08355_));
 XOR2x2_ASAP7_75t_R _20933_ (.A(_00140_),
    .B(_08355_),
    .Y(_08356_));
 AND2x2_ASAP7_75t_R _20934_ (.A(_08328_),
    .B(_08356_),
    .Y(_04937_));
 OR4x1_ASAP7_75t_R _20935_ (.A(_00140_),
    .B(_00141_),
    .C(_00142_),
    .D(_00143_),
    .Y(_08357_));
 OR3x1_ASAP7_75t_R _20936_ (.A(_00139_),
    .B(_08349_),
    .C(_08357_),
    .Y(_08358_));
 OAI21x1_ASAP7_75t_R _20937_ (.A1(_08349_),
    .A2(_08357_),
    .B(_00139_),
    .Y(_08359_));
 AND3x1_ASAP7_75t_R _20938_ (.A(_08232_),
    .B(_08358_),
    .C(_08359_),
    .Y(_04938_));
 OR3x1_ASAP7_75t_R _20939_ (.A(_00139_),
    .B(_08347_),
    .C(_08357_),
    .Y(_08360_));
 XOR2x2_ASAP7_75t_R _20940_ (.A(_00138_),
    .B(_08360_),
    .Y(_08361_));
 AND2x2_ASAP7_75t_R _20941_ (.A(_08328_),
    .B(_08361_),
    .Y(_04939_));
 BUFx6f_ASAP7_75t_R _20942_ (.A(_09029_),
    .Y(_08362_));
 XOR2x2_ASAP7_75t_R _20943_ (.A(_00137_),
    .B(_02647_),
    .Y(_08363_));
 AND2x2_ASAP7_75t_R _20944_ (.A(_08362_),
    .B(_08363_),
    .Y(_04940_));
 OR4x1_ASAP7_75t_R _20945_ (.A(_00138_),
    .B(_00139_),
    .C(_08349_),
    .D(_08357_),
    .Y(_08364_));
 XOR2x2_ASAP7_75t_R _20946_ (.A(_00136_),
    .B(_08364_),
    .Y(_08365_));
 AND2x2_ASAP7_75t_R _20947_ (.A(_08362_),
    .B(_08365_),
    .Y(_04941_));
 OR5x1_ASAP7_75t_R _20948_ (.A(_00136_),
    .B(_00138_),
    .C(_00139_),
    .D(_08347_),
    .E(_08357_),
    .Y(_08366_));
 XOR2x2_ASAP7_75t_R _20949_ (.A(_00135_),
    .B(_08366_),
    .Y(_08367_));
 AND2x2_ASAP7_75t_R _20950_ (.A(_08362_),
    .B(_08367_),
    .Y(_04942_));
 OR3x1_ASAP7_75t_R _20951_ (.A(_00137_),
    .B(_00148_),
    .C(_00061_),
    .Y(_08368_));
 XOR2x2_ASAP7_75t_R _20952_ (.A(_00134_),
    .B(_08368_),
    .Y(_08369_));
 AND2x2_ASAP7_75t_R _20953_ (.A(_08362_),
    .B(_08369_),
    .Y(_04943_));
 OR3x1_ASAP7_75t_R _20954_ (.A(_00134_),
    .B(_00137_),
    .C(_02647_),
    .Y(_08370_));
 NAND2x1_ASAP7_75t_R _20955_ (.A(_00133_),
    .B(_08370_),
    .Y(_08371_));
 AND3x1_ASAP7_75t_R _20956_ (.A(_08232_),
    .B(_08311_),
    .C(_08371_),
    .Y(_04944_));
 XOR2x2_ASAP7_75t_R _20957_ (.A(_00132_),
    .B(_08316_),
    .Y(_08372_));
 AND2x2_ASAP7_75t_R _20958_ (.A(_08362_),
    .B(_08372_),
    .Y(_04945_));
 BUFx6f_ASAP7_75t_R _20959_ (.A(_08998_),
    .Y(_08373_));
 OR3x1_ASAP7_75t_R _20960_ (.A(_00131_),
    .B(_00132_),
    .C(_08311_),
    .Y(_08374_));
 OAI21x1_ASAP7_75t_R _20961_ (.A1(_00132_),
    .A2(_08311_),
    .B(_00131_),
    .Y(_08375_));
 AND3x1_ASAP7_75t_R _20962_ (.A(_08373_),
    .B(_08374_),
    .C(_08375_),
    .Y(_04946_));
 OR3x1_ASAP7_75t_R _20963_ (.A(_00131_),
    .B(_00132_),
    .C(_08316_),
    .Y(_08376_));
 XOR2x2_ASAP7_75t_R _20964_ (.A(_00130_),
    .B(_08376_),
    .Y(_08377_));
 AND2x2_ASAP7_75t_R _20965_ (.A(_08362_),
    .B(_08377_),
    .Y(_04947_));
 OR4x1_ASAP7_75t_R _20966_ (.A(_00130_),
    .B(_00131_),
    .C(_00132_),
    .D(_08311_),
    .Y(_08378_));
 NAND2x1_ASAP7_75t_R _20967_ (.A(_00129_),
    .B(_08378_),
    .Y(_08379_));
 AND3x1_ASAP7_75t_R _20968_ (.A(_08373_),
    .B(_08313_),
    .C(_08379_),
    .Y(_04948_));
 XOR2x2_ASAP7_75t_R _20969_ (.A(_08300_),
    .B(_08317_),
    .Y(_08380_));
 AND2x2_ASAP7_75t_R _20970_ (.A(_08362_),
    .B(_08380_),
    .Y(_04949_));
 BUFx3_ASAP7_75t_R _20971_ (.A(_00118_),
    .Y(_08381_));
 AND4x1_ASAP7_75t_R _20972_ (.A(_00089_),
    .B(_00117_),
    .C(_08381_),
    .D(_00119_),
    .Y(_08382_));
 AND5x1_ASAP7_75t_R _20973_ (.A(_00108_),
    .B(_00113_),
    .C(_00114_),
    .D(_00116_),
    .E(_08382_),
    .Y(_08383_));
 AND5x2_ASAP7_75t_R _20974_ (.A(_00110_),
    .B(_00111_),
    .C(_00112_),
    .D(_11465_),
    .E(_08383_),
    .Y(_08384_));
 BUFx3_ASAP7_75t_R _20975_ (.A(_00105_),
    .Y(_08385_));
 AND4x1_ASAP7_75t_R _20976_ (.A(_00103_),
    .B(_00104_),
    .C(_08385_),
    .D(_00106_),
    .Y(_08386_));
 AND4x1_ASAP7_75t_R _20977_ (.A(_00097_),
    .B(_00099_),
    .C(_00100_),
    .D(_00107_),
    .Y(_08387_));
 AND5x1_ASAP7_75t_R _20978_ (.A(_00090_),
    .B(_00091_),
    .C(_00096_),
    .D(_00115_),
    .E(_08387_),
    .Y(_08388_));
 BUFx3_ASAP7_75t_R _20979_ (.A(_00093_),
    .Y(_08389_));
 AND3x1_ASAP7_75t_R _20980_ (.A(_00094_),
    .B(_00095_),
    .C(_00098_),
    .Y(_08390_));
 OR3x1_ASAP7_75t_R _20981_ (.A(_00092_),
    .B(_08389_),
    .C(_08390_),
    .Y(_08391_));
 AND5x2_ASAP7_75t_R _20982_ (.A(_00101_),
    .B(_00102_),
    .C(_08386_),
    .D(_08388_),
    .E(_08391_),
    .Y(_08392_));
 NAND2x2_ASAP7_75t_R _20983_ (.A(_08384_),
    .B(_08392_),
    .Y(_08393_));
 NOR2x1_ASAP7_75t_R _20984_ (.A(_00079_),
    .B(_08393_),
    .Y(_04950_));
 INVx1_ASAP7_75t_R _20985_ (.A(_08393_),
    .Y(_04951_));
 NOR2x1_ASAP7_75t_R _20986_ (.A(_00082_),
    .B(_08393_),
    .Y(_04952_));
 NOR2x1_ASAP7_75t_R _20987_ (.A(_00081_),
    .B(_08393_),
    .Y(_04953_));
 NOR2x1_ASAP7_75t_R _20988_ (.A(_00080_),
    .B(_08393_),
    .Y(_04954_));
 NOR2x1_ASAP7_75t_R _20989_ (.A(_00078_),
    .B(_08393_),
    .Y(_04955_));
 NOR2x1_ASAP7_75t_R _20990_ (.A(_00077_),
    .B(_08393_),
    .Y(_04956_));
 INVx1_ASAP7_75t_R _20991_ (.A(_08393_),
    .Y(_04957_));
 AND2x2_ASAP7_75t_R _20992_ (.A(_08362_),
    .B(_00062_),
    .Y(_04958_));
 OR4x1_ASAP7_75t_R _20993_ (.A(_00094_),
    .B(_00095_),
    .C(_00098_),
    .D(_02653_),
    .Y(_08394_));
 OR4x1_ASAP7_75t_R _20994_ (.A(_00090_),
    .B(_00091_),
    .C(_00092_),
    .D(_08389_),
    .Y(_08395_));
 OR4x1_ASAP7_75t_R _20995_ (.A(_00089_),
    .B(_00119_),
    .C(_08394_),
    .D(_08395_),
    .Y(_08396_));
 BUFx6f_ASAP7_75t_R _20996_ (.A(_08396_),
    .Y(_08397_));
 OR3x1_ASAP7_75t_R _20997_ (.A(_00089_),
    .B(_08394_),
    .C(_08395_),
    .Y(_08398_));
 NAND2x1_ASAP7_75t_R _20998_ (.A(_00119_),
    .B(_08398_),
    .Y(_08399_));
 AND3x1_ASAP7_75t_R _20999_ (.A(_08373_),
    .B(_08397_),
    .C(_08399_),
    .Y(_04959_));
 OR4x1_ASAP7_75t_R _21000_ (.A(_00089_),
    .B(_00090_),
    .C(_00092_),
    .D(_08389_),
    .Y(_08400_));
 OR5x2_ASAP7_75t_R _21001_ (.A(_00094_),
    .B(_00095_),
    .C(_00098_),
    .D(_00109_),
    .E(_00062_),
    .Y(_08401_));
 OR4x1_ASAP7_75t_R _21002_ (.A(_00091_),
    .B(_00119_),
    .C(_08400_),
    .D(_08401_),
    .Y(_08402_));
 XOR2x2_ASAP7_75t_R _21003_ (.A(_08381_),
    .B(_08402_),
    .Y(_08403_));
 AND2x2_ASAP7_75t_R _21004_ (.A(_08362_),
    .B(_08403_),
    .Y(_04960_));
 OR3x1_ASAP7_75t_R _21005_ (.A(_00117_),
    .B(_08381_),
    .C(_08397_),
    .Y(_08404_));
 OAI21x1_ASAP7_75t_R _21006_ (.A1(_08381_),
    .A2(_08397_),
    .B(_00117_),
    .Y(_08405_));
 AND3x1_ASAP7_75t_R _21007_ (.A(_08373_),
    .B(_08404_),
    .C(_08405_),
    .Y(_04961_));
 OR3x1_ASAP7_75t_R _21008_ (.A(_00117_),
    .B(_08381_),
    .C(_08402_),
    .Y(_08406_));
 XOR2x2_ASAP7_75t_R _21009_ (.A(_00116_),
    .B(_08406_),
    .Y(_08407_));
 AND2x2_ASAP7_75t_R _21010_ (.A(_08362_),
    .B(_08407_),
    .Y(_04962_));
 BUFx6f_ASAP7_75t_R _21011_ (.A(_09029_),
    .Y(_08408_));
 OR4x1_ASAP7_75t_R _21012_ (.A(_00116_),
    .B(_00117_),
    .C(_08381_),
    .D(_08397_),
    .Y(_08409_));
 XOR2x2_ASAP7_75t_R _21013_ (.A(_00115_),
    .B(_08409_),
    .Y(_08410_));
 AND2x2_ASAP7_75t_R _21014_ (.A(_08408_),
    .B(_08410_),
    .Y(_04963_));
 OR5x1_ASAP7_75t_R _21015_ (.A(_00115_),
    .B(_00116_),
    .C(_00117_),
    .D(_08381_),
    .E(_08402_),
    .Y(_08411_));
 XOR2x2_ASAP7_75t_R _21016_ (.A(_00114_),
    .B(_08411_),
    .Y(_08412_));
 AND2x2_ASAP7_75t_R _21017_ (.A(_08408_),
    .B(_08412_),
    .Y(_04964_));
 OR5x2_ASAP7_75t_R _21018_ (.A(_00114_),
    .B(_00115_),
    .C(_00116_),
    .D(_00117_),
    .E(_08381_),
    .Y(_08413_));
 OR3x1_ASAP7_75t_R _21019_ (.A(_00113_),
    .B(_08397_),
    .C(_08413_),
    .Y(_08414_));
 OAI21x1_ASAP7_75t_R _21020_ (.A1(_08397_),
    .A2(_08413_),
    .B(_00113_),
    .Y(_08415_));
 AND3x1_ASAP7_75t_R _21021_ (.A(_08373_),
    .B(_08414_),
    .C(_08415_),
    .Y(_04965_));
 OR3x1_ASAP7_75t_R _21022_ (.A(_00113_),
    .B(_08402_),
    .C(_08413_),
    .Y(_08416_));
 XOR2x2_ASAP7_75t_R _21023_ (.A(_00112_),
    .B(_08416_),
    .Y(_08417_));
 AND2x2_ASAP7_75t_R _21024_ (.A(_08408_),
    .B(_08417_),
    .Y(_04966_));
 OR4x1_ASAP7_75t_R _21025_ (.A(_00112_),
    .B(_00113_),
    .C(_08397_),
    .D(_08413_),
    .Y(_08418_));
 XOR2x2_ASAP7_75t_R _21026_ (.A(_00111_),
    .B(_08418_),
    .Y(_08419_));
 AND2x2_ASAP7_75t_R _21027_ (.A(_08408_),
    .B(_08419_),
    .Y(_04967_));
 OR3x1_ASAP7_75t_R _21028_ (.A(_00111_),
    .B(_00112_),
    .C(_08416_),
    .Y(_08420_));
 XOR2x2_ASAP7_75t_R _21029_ (.A(_00110_),
    .B(_08420_),
    .Y(_08421_));
 AND2x2_ASAP7_75t_R _21030_ (.A(_08408_),
    .B(_08421_),
    .Y(_04968_));
 NOR2x1_ASAP7_75t_R _21031_ (.A(_10986_),
    .B(_02654_),
    .Y(_04969_));
 OR3x1_ASAP7_75t_R _21032_ (.A(_00110_),
    .B(_00111_),
    .C(_08418_),
    .Y(_08422_));
 XOR2x2_ASAP7_75t_R _21033_ (.A(_00108_),
    .B(_08422_),
    .Y(_08423_));
 AND2x2_ASAP7_75t_R _21034_ (.A(_08408_),
    .B(_08423_),
    .Y(_04970_));
 OR2x2_ASAP7_75t_R _21035_ (.A(_00112_),
    .B(_08416_),
    .Y(_08424_));
 OR4x1_ASAP7_75t_R _21036_ (.A(_00108_),
    .B(_00110_),
    .C(_00111_),
    .D(_08424_),
    .Y(_08425_));
 XOR2x2_ASAP7_75t_R _21037_ (.A(_00107_),
    .B(_08425_),
    .Y(_08426_));
 AND2x2_ASAP7_75t_R _21038_ (.A(_08408_),
    .B(_08426_),
    .Y(_04971_));
 OR5x1_ASAP7_75t_R _21039_ (.A(_00106_),
    .B(_00107_),
    .C(_00108_),
    .D(_00110_),
    .E(_00111_),
    .Y(_08427_));
 OR5x2_ASAP7_75t_R _21040_ (.A(_00112_),
    .B(_00113_),
    .C(_08397_),
    .D(_08413_),
    .E(_08427_),
    .Y(_08428_));
 OR5x1_ASAP7_75t_R _21041_ (.A(_00107_),
    .B(_00108_),
    .C(_00110_),
    .D(_00111_),
    .E(_08418_),
    .Y(_08429_));
 NAND2x1_ASAP7_75t_R _21042_ (.A(_00106_),
    .B(_08429_),
    .Y(_08430_));
 AND3x1_ASAP7_75t_R _21043_ (.A(_08373_),
    .B(_08428_),
    .C(_08430_),
    .Y(_04972_));
 OR5x2_ASAP7_75t_R _21044_ (.A(_00112_),
    .B(_00113_),
    .C(_08402_),
    .D(_08413_),
    .E(_08427_),
    .Y(_08431_));
 XOR2x2_ASAP7_75t_R _21045_ (.A(_08385_),
    .B(_08431_),
    .Y(_08432_));
 AND2x2_ASAP7_75t_R _21046_ (.A(_08408_),
    .B(_08432_),
    .Y(_04973_));
 OR3x1_ASAP7_75t_R _21047_ (.A(_00104_),
    .B(_08385_),
    .C(_08428_),
    .Y(_08433_));
 OAI21x1_ASAP7_75t_R _21048_ (.A1(_08385_),
    .A2(_08428_),
    .B(_00104_),
    .Y(_08434_));
 AND3x1_ASAP7_75t_R _21049_ (.A(_08373_),
    .B(_08433_),
    .C(_08434_),
    .Y(_04974_));
 OR3x1_ASAP7_75t_R _21050_ (.A(_00104_),
    .B(_08385_),
    .C(_08431_),
    .Y(_08435_));
 XOR2x2_ASAP7_75t_R _21051_ (.A(_00103_),
    .B(_08435_),
    .Y(_08436_));
 AND2x2_ASAP7_75t_R _21052_ (.A(_08408_),
    .B(_08436_),
    .Y(_04975_));
 OR5x2_ASAP7_75t_R _21053_ (.A(_00102_),
    .B(_00103_),
    .C(_00104_),
    .D(_08385_),
    .E(_08428_),
    .Y(_08437_));
 OR4x1_ASAP7_75t_R _21054_ (.A(_00103_),
    .B(_00104_),
    .C(_08385_),
    .D(_08428_),
    .Y(_08438_));
 NAND2x1_ASAP7_75t_R _21055_ (.A(_00102_),
    .B(_08438_),
    .Y(_08439_));
 AND3x1_ASAP7_75t_R _21056_ (.A(_08373_),
    .B(_08437_),
    .C(_08439_),
    .Y(_04976_));
 OR5x2_ASAP7_75t_R _21057_ (.A(_00102_),
    .B(_00103_),
    .C(_00104_),
    .D(_08385_),
    .E(_08431_),
    .Y(_08440_));
 XOR2x2_ASAP7_75t_R _21058_ (.A(_00101_),
    .B(_08440_),
    .Y(_08441_));
 AND2x2_ASAP7_75t_R _21059_ (.A(_08408_),
    .B(_08441_),
    .Y(_04977_));
 OR3x1_ASAP7_75t_R _21060_ (.A(_00100_),
    .B(_00101_),
    .C(_08437_),
    .Y(_08442_));
 OAI21x1_ASAP7_75t_R _21061_ (.A1(_00101_),
    .A2(_08437_),
    .B(_00100_),
    .Y(_08443_));
 AND3x1_ASAP7_75t_R _21062_ (.A(_08373_),
    .B(_08442_),
    .C(_08443_),
    .Y(_04978_));
 OR3x1_ASAP7_75t_R _21063_ (.A(_00100_),
    .B(_00101_),
    .C(_08440_),
    .Y(_08444_));
 XOR2x2_ASAP7_75t_R _21064_ (.A(_00099_),
    .B(_08444_),
    .Y(_08445_));
 AND2x2_ASAP7_75t_R _21065_ (.A(_08877_),
    .B(_08445_),
    .Y(_04979_));
 XOR2x2_ASAP7_75t_R _21066_ (.A(_00098_),
    .B(_02653_),
    .Y(_08446_));
 AND2x2_ASAP7_75t_R _21067_ (.A(_08877_),
    .B(_08446_),
    .Y(_04980_));
 OR4x1_ASAP7_75t_R _21068_ (.A(_00099_),
    .B(_00100_),
    .C(_00101_),
    .D(_08437_),
    .Y(_08447_));
 XOR2x2_ASAP7_75t_R _21069_ (.A(_00097_),
    .B(_08447_),
    .Y(_08448_));
 AND2x2_ASAP7_75t_R _21070_ (.A(_08877_),
    .B(_08448_),
    .Y(_04981_));
 OR5x1_ASAP7_75t_R _21071_ (.A(_00097_),
    .B(_00099_),
    .C(_00100_),
    .D(_00101_),
    .E(_08440_),
    .Y(_08449_));
 XOR2x2_ASAP7_75t_R _21072_ (.A(_00096_),
    .B(_08449_),
    .Y(_08450_));
 AND2x2_ASAP7_75t_R _21073_ (.A(_08877_),
    .B(_08450_),
    .Y(_04982_));
 OR3x1_ASAP7_75t_R _21074_ (.A(_00098_),
    .B(_00109_),
    .C(_00062_),
    .Y(_08451_));
 XOR2x2_ASAP7_75t_R _21075_ (.A(_00095_),
    .B(_08451_),
    .Y(_08452_));
 AND2x2_ASAP7_75t_R _21076_ (.A(_08877_),
    .B(_08452_),
    .Y(_04983_));
 OR3x1_ASAP7_75t_R _21077_ (.A(_00095_),
    .B(_00098_),
    .C(_02653_),
    .Y(_08453_));
 NAND2x1_ASAP7_75t_R _21078_ (.A(_00094_),
    .B(_08453_),
    .Y(_08454_));
 AND3x1_ASAP7_75t_R _21079_ (.A(_08373_),
    .B(_08394_),
    .C(_08454_),
    .Y(_04984_));
 XOR2x2_ASAP7_75t_R _21080_ (.A(_08389_),
    .B(_08401_),
    .Y(_08455_));
 AND2x2_ASAP7_75t_R _21081_ (.A(_08877_),
    .B(_08455_),
    .Y(_04985_));
 OR3x1_ASAP7_75t_R _21082_ (.A(_00092_),
    .B(_08389_),
    .C(_08394_),
    .Y(_08456_));
 OAI21x1_ASAP7_75t_R _21083_ (.A1(_08389_),
    .A2(_08394_),
    .B(_00092_),
    .Y(_08457_));
 AND3x1_ASAP7_75t_R _21084_ (.A(_08999_),
    .B(_08456_),
    .C(_08457_),
    .Y(_04986_));
 OR3x1_ASAP7_75t_R _21085_ (.A(_00092_),
    .B(_08389_),
    .C(_08401_),
    .Y(_08458_));
 XOR2x2_ASAP7_75t_R _21086_ (.A(_00091_),
    .B(_08458_),
    .Y(_08459_));
 AND2x2_ASAP7_75t_R _21087_ (.A(_08877_),
    .B(_08459_),
    .Y(_04987_));
 OR4x1_ASAP7_75t_R _21088_ (.A(_00091_),
    .B(_00092_),
    .C(_08389_),
    .D(_08394_),
    .Y(_08460_));
 NAND2x1_ASAP7_75t_R _21089_ (.A(_00090_),
    .B(_08460_),
    .Y(_08461_));
 OA211x2_ASAP7_75t_R _21090_ (.A1(_08394_),
    .A2(_08395_),
    .B(_08461_),
    .C(_07260_),
    .Y(_04988_));
 OR3x1_ASAP7_75t_R _21091_ (.A(_00089_),
    .B(_08395_),
    .C(_08401_),
    .Y(_08462_));
 OAI21x1_ASAP7_75t_R _21092_ (.A1(_08395_),
    .A2(_08401_),
    .B(_00089_),
    .Y(_08463_));
 AND3x1_ASAP7_75t_R _21093_ (.A(_08999_),
    .B(_08462_),
    .C(_08463_),
    .Y(_04989_));
 AND2x2_ASAP7_75t_R _21094_ (.A(_08877_),
    .B(_00030_),
    .Y(_04990_));
 INVx2_ASAP7_75t_R _21095_ (.A(_02148_),
    .Y(_08464_));
 AND4x1_ASAP7_75t_R _21096_ (.A(\peo[18][36] ),
    .B(_00161_),
    .C(_00162_),
    .D(\peo[18][33] ),
    .Y(_08465_));
 AND3x1_ASAP7_75t_R _21097_ (.A(\peo[18][39] ),
    .B(\peo[18][32] ),
    .C(_08465_),
    .Y(_08466_));
 INVx1_ASAP7_75t_R _21098_ (.A(_02155_),
    .Y(_08467_));
 NAND2x1_ASAP7_75t_R _21099_ (.A(_00122_),
    .B(_00123_),
    .Y(_08468_));
 OR2x6_ASAP7_75t_R _21100_ (.A(_00121_),
    .B(_00124_),
    .Y(_08469_));
 OAI21x1_ASAP7_75t_R _21101_ (.A1(_08468_),
    .A2(_08469_),
    .B(\peo[19][39] ),
    .Y(_08470_));
 AND2x2_ASAP7_75t_R _21102_ (.A(_00122_),
    .B(_00123_),
    .Y(_08471_));
 AND5x2_ASAP7_75t_R _21103_ (.A(\peo[19][39] ),
    .B(\peo[19][36] ),
    .C(\peo[19][33] ),
    .D(_00125_),
    .E(_08471_),
    .Y(_08472_));
 AO21x1_ASAP7_75t_R _21104_ (.A1(_08467_),
    .A2(_08470_),
    .B(_08472_),
    .Y(_08473_));
 OA211x2_ASAP7_75t_R _21105_ (.A1(_00159_),
    .A2(_08465_),
    .B(_08472_),
    .C(_02155_),
    .Y(_08474_));
 AO21x2_ASAP7_75t_R _21106_ (.A1(_08466_),
    .A2(_08473_),
    .B(_08474_),
    .Y(_08475_));
 INVx2_ASAP7_75t_R _21107_ (.A(_02149_),
    .Y(_08476_));
 OR3x1_ASAP7_75t_R _21108_ (.A(_02148_),
    .B(_08476_),
    .C(_08467_),
    .Y(_08477_));
 AOI21x1_ASAP7_75t_R _21109_ (.A1(_08464_),
    .A2(_08475_),
    .B(_08477_),
    .Y(_08478_));
 NAND2x1_ASAP7_75t_R _21110_ (.A(_02159_),
    .B(_08478_),
    .Y(_08479_));
 OR2x2_ASAP7_75t_R _21111_ (.A(_08468_),
    .B(_08469_),
    .Y(_08480_));
 OR3x1_ASAP7_75t_R _21112_ (.A(_00120_),
    .B(\peo[19][32] ),
    .C(_08480_),
    .Y(_08481_));
 OR4x1_ASAP7_75t_R _21113_ (.A(_00160_),
    .B(\peo[18][35] ),
    .C(\peo[18][34] ),
    .D(_00163_),
    .Y(_08482_));
 AO32x1_ASAP7_75t_R _21114_ (.A1(\peo[18][39] ),
    .A2(_08482_),
    .A3(_08472_),
    .B1(_08480_),
    .B2(\peo[19][39] ),
    .Y(_08483_));
 OA31x2_ASAP7_75t_R _21115_ (.A1(_00125_),
    .A2(_08468_),
    .A3(_08469_),
    .B1(\peo[19][39] ),
    .Y(_08484_));
 AND2x2_ASAP7_75t_R _21116_ (.A(_02148_),
    .B(_00030_),
    .Y(_08485_));
 OA21x2_ASAP7_75t_R _21117_ (.A1(_08468_),
    .A2(_08469_),
    .B(\peo[19][39] ),
    .Y(_08486_));
 AO32x1_ASAP7_75t_R _21118_ (.A1(_08464_),
    .A2(_02155_),
    .A3(_08484_),
    .B1(_08485_),
    .B2(_08486_),
    .Y(_08487_));
 AND2x2_ASAP7_75t_R _21119_ (.A(\peo[18][39] ),
    .B(_08482_),
    .Y(_08488_));
 AO32x2_ASAP7_75t_R _21120_ (.A1(_08464_),
    .A2(_08476_),
    .A3(_08483_),
    .B1(_08487_),
    .B2(_08488_),
    .Y(_08489_));
 NOR2x1_ASAP7_75t_R _21121_ (.A(_08481_),
    .B(_08489_),
    .Y(_08490_));
 OR3x1_ASAP7_75t_R _21122_ (.A(\peo[18][0] ),
    .B(_08478_),
    .C(_08490_),
    .Y(_08491_));
 OR3x1_ASAP7_75t_R _21123_ (.A(\peo[19][0] ),
    .B(_08481_),
    .C(_08489_),
    .Y(_08492_));
 AND4x1_ASAP7_75t_R _21124_ (.A(_08585_),
    .B(_08479_),
    .C(_08491_),
    .D(_08492_),
    .Y(_04991_));
 NAND2x2_ASAP7_75t_R _21125_ (.A(_08528_),
    .B(_08478_),
    .Y(_08493_));
 NOR2x1_ASAP7_75t_R _21126_ (.A(_02158_),
    .B(_08493_),
    .Y(_04992_));
 NOR2x1_ASAP7_75t_R _21127_ (.A(_02157_),
    .B(_08493_),
    .Y(_04993_));
 NOR2x1_ASAP7_75t_R _21128_ (.A(_02156_),
    .B(_08493_),
    .Y(_04994_));
 NOR2x1_ASAP7_75t_R _21129_ (.A(_02147_),
    .B(_08493_),
    .Y(_04995_));
 NOR2x1_ASAP7_75t_R _21130_ (.A(_02146_),
    .B(_08493_),
    .Y(_04996_));
 OR3x1_ASAP7_75t_R _21131_ (.A(_02148_),
    .B(_08476_),
    .C(_02155_),
    .Y(_08494_));
 AO21x1_ASAP7_75t_R _21132_ (.A1(_08466_),
    .A2(_08470_),
    .B(_08494_),
    .Y(_08495_));
 NOR2x1_ASAP7_75t_R _21133_ (.A(_02159_),
    .B(_08495_),
    .Y(_08496_));
 AO21x1_ASAP7_75t_R _21134_ (.A1(\peo[18][0] ),
    .A2(_08495_),
    .B(_08496_),
    .Y(_08497_));
 NAND2x1_ASAP7_75t_R _21135_ (.A(_00127_),
    .B(_08489_),
    .Y(_08498_));
 OA211x2_ASAP7_75t_R _21136_ (.A1(_08489_),
    .A2(_08497_),
    .B(_08498_),
    .C(_08599_),
    .Y(_04997_));
 OR2x2_ASAP7_75t_R _21137_ (.A(_09220_),
    .B(_08495_),
    .Y(_08499_));
 BUFx3_ASAP7_75t_R _21138_ (.A(_08499_),
    .Y(_08500_));
 NOR2x1_ASAP7_75t_R _21139_ (.A(_02158_),
    .B(_08500_),
    .Y(_04998_));
 NOR2x1_ASAP7_75t_R _21140_ (.A(_02157_),
    .B(_08500_),
    .Y(_04999_));
 NOR2x1_ASAP7_75t_R _21141_ (.A(_02156_),
    .B(_08500_),
    .Y(_05000_));
 NOR2x1_ASAP7_75t_R _21142_ (.A(_02147_),
    .B(_08500_),
    .Y(_05001_));
 NOR2x1_ASAP7_75t_R _21143_ (.A(_02146_),
    .B(_08500_),
    .Y(_05002_));
 AO221x1_ASAP7_75t_R _21144_ (.A1(_08464_),
    .A2(_08476_),
    .B1(_08488_),
    .B2(_08487_),
    .C(_08470_),
    .Y(_08501_));
 BUFx6f_ASAP7_75t_R _21145_ (.A(_08501_),
    .Y(_08502_));
 OR2x2_ASAP7_75t_R _21146_ (.A(\peo[19][0] ),
    .B(_08502_),
    .Y(_08503_));
 NAND2x1_ASAP7_75t_R _21147_ (.A(_00166_),
    .B(_08502_),
    .Y(_08504_));
 OA21x2_ASAP7_75t_R _21148_ (.A1(_08476_),
    .A2(_08475_),
    .B(_08464_),
    .Y(_08505_));
 BUFx6f_ASAP7_75t_R _21149_ (.A(_08505_),
    .Y(_08506_));
 NOR2x1_ASAP7_75t_R _21150_ (.A(_10826_),
    .B(_08506_),
    .Y(_08507_));
 NOR2x1_ASAP7_75t_R _21151_ (.A(_06206_),
    .B(_02159_),
    .Y(_08508_));
 AO32x1_ASAP7_75t_R _21152_ (.A1(_08503_),
    .A2(_08504_),
    .A3(_08507_),
    .B1(_08508_),
    .B2(_08506_),
    .Y(_05003_));
 NAND2x2_ASAP7_75t_R _21153_ (.A(_09029_),
    .B(_08505_),
    .Y(_08509_));
 NOR2x1_ASAP7_75t_R _21154_ (.A(_02158_),
    .B(_08509_),
    .Y(_05004_));
 NOR2x1_ASAP7_75t_R _21155_ (.A(_02157_),
    .B(_08509_),
    .Y(_05005_));
 NOR2x1_ASAP7_75t_R _21156_ (.A(_02156_),
    .B(_08509_),
    .Y(_05006_));
 NOR2x1_ASAP7_75t_R _21157_ (.A(_00125_),
    .B(_08502_),
    .Y(_08510_));
 AO21x1_ASAP7_75t_R _21158_ (.A1(\peo[18][32] ),
    .A2(_08502_),
    .B(_08510_),
    .Y(_08511_));
 AND3x1_ASAP7_75t_R _21159_ (.A(_08599_),
    .B(_08467_),
    .C(_08506_),
    .Y(_08512_));
 AO21x1_ASAP7_75t_R _21160_ (.A1(_08507_),
    .A2(_08511_),
    .B(_08512_),
    .Y(_05007_));
 NOR2x1_ASAP7_75t_R _21161_ (.A(_00120_),
    .B(_08489_),
    .Y(_08513_));
 AOI22x1_ASAP7_75t_R _21162_ (.A1(_00163_),
    .A2(_08502_),
    .B1(_08513_),
    .B2(_00124_),
    .Y(_08514_));
 NAND2x1_ASAP7_75t_R _21163_ (.A(_02154_),
    .B(_08506_),
    .Y(_08515_));
 OA211x2_ASAP7_75t_R _21164_ (.A1(_08506_),
    .A2(_08514_),
    .B(_08515_),
    .C(_08599_),
    .Y(_05008_));
 OR2x2_ASAP7_75t_R _21165_ (.A(\peo[19][34] ),
    .B(_08502_),
    .Y(_08516_));
 NAND2x1_ASAP7_75t_R _21166_ (.A(_00162_),
    .B(_08502_),
    .Y(_08517_));
 NOR2x1_ASAP7_75t_R _21167_ (.A(_06206_),
    .B(_02153_),
    .Y(_08518_));
 AO32x1_ASAP7_75t_R _21168_ (.A1(_08507_),
    .A2(_08516_),
    .A3(_08517_),
    .B1(_08518_),
    .B2(_08506_),
    .Y(_05009_));
 OR2x2_ASAP7_75t_R _21169_ (.A(\peo[19][35] ),
    .B(_08502_),
    .Y(_08519_));
 NAND2x1_ASAP7_75t_R _21170_ (.A(_00161_),
    .B(_08502_),
    .Y(_08520_));
 NOR2x1_ASAP7_75t_R _21171_ (.A(_10047_),
    .B(_02152_),
    .Y(_08521_));
 AO32x1_ASAP7_75t_R _21172_ (.A1(_08507_),
    .A2(_08519_),
    .A3(_08520_),
    .B1(_08521_),
    .B2(_08506_),
    .Y(_05010_));
 AOI22x1_ASAP7_75t_R _21173_ (.A1(_00160_),
    .A2(_08502_),
    .B1(_08513_),
    .B2(_00121_),
    .Y(_08522_));
 NAND2x1_ASAP7_75t_R _21174_ (.A(_02151_),
    .B(_08506_),
    .Y(_08523_));
 OA211x2_ASAP7_75t_R _21175_ (.A1(_08506_),
    .A2(_08522_),
    .B(_08523_),
    .C(_08599_),
    .Y(_05011_));
 NOR2x1_ASAP7_75t_R _21176_ (.A(_02150_),
    .B(_08509_),
    .Y(_05012_));
 AND4x1_ASAP7_75t_R _21177_ (.A(_08585_),
    .B(_08464_),
    .C(_02149_),
    .D(_08475_),
    .Y(_05013_));
 AO21x1_ASAP7_75t_R _21178_ (.A1(\peo[18][39] ),
    .A2(_08482_),
    .B(_08486_),
    .Y(_08524_));
 OA21x2_ASAP7_75t_R _21179_ (.A1(_08506_),
    .A2(_08524_),
    .B(_08529_),
    .Y(_05014_));
 NOR2x1_ASAP7_75t_R _21180_ (.A(_02147_),
    .B(_08509_),
    .Y(_05015_));
 NOR2x1_ASAP7_75t_R _21181_ (.A(_02146_),
    .B(_08509_),
    .Y(_05016_));
 HAxp5_ASAP7_75t_R _21182_ (.A(\xs[8].cli1.r[0] ),
    .B(\xs[8].cli1.r[1] ),
    .CON(_02611_),
    .SN(_02612_));
 HAxp5_ASAP7_75t_R _21183_ (.A(\xs[13].cli1.r[0] ),
    .B(\xs[13].cli1.r[1] ),
    .CON(_02613_),
    .SN(_02614_));
 HAxp5_ASAP7_75t_R _21184_ (.A(\xs[1].cli0.r[0] ),
    .B(\xs[1].cli0.r[1] ),
    .CON(_02615_),
    .SN(_02616_));
 HAxp5_ASAP7_75t_R _21185_ (.A(\xs[15].cli1.r[0] ),
    .B(\xs[15].cli1.r[1] ),
    .CON(_02617_),
    .SN(_02618_));
 HAxp5_ASAP7_75t_R _21186_ (.A(\xs[5].cli1.r[0] ),
    .B(\xs[5].cli1.r[1] ),
    .CON(_02619_),
    .SN(_02620_));
 HAxp5_ASAP7_75t_R _21187_ (.A(\xs[6].cli0.r[0] ),
    .B(\xs[6].cli0.r[1] ),
    .CON(_02621_),
    .SN(_02622_));
 HAxp5_ASAP7_75t_R _21188_ (.A(\xs[0].cli1.r[0] ),
    .B(\xs[0].cli1.r[1] ),
    .CON(_02623_),
    .SN(_02624_));
 HAxp5_ASAP7_75t_R _21189_ (.A(\xs[12].cli1.r[0] ),
    .B(\xs[12].cli1.r[1] ),
    .CON(_02625_),
    .SN(_02626_));
 HAxp5_ASAP7_75t_R _21190_ (.A(\xs[10].cli0.r[0] ),
    .B(\xs[10].cli0.r[1] ),
    .CON(_02627_),
    .SN(_02628_));
 HAxp5_ASAP7_75t_R _21191_ (.A(\xs[15].cli0.r[0] ),
    .B(\xs[15].cli0.r[1] ),
    .CON(_02629_),
    .SN(_02630_));
 HAxp5_ASAP7_75t_R _21192_ (.A(\xs[0].cli0.r[0] ),
    .B(\xs[0].cli0.r[1] ),
    .CON(_02631_),
    .SN(_02632_));
 HAxp5_ASAP7_75t_R _21193_ (.A(\xs[14].cli1.r[0] ),
    .B(\xs[14].cli1.r[1] ),
    .CON(_02633_),
    .SN(_02634_));
 HAxp5_ASAP7_75t_R _21194_ (.A(\xs[10].cli1.r[0] ),
    .B(\xs[10].cli1.r[1] ),
    .CON(_02635_),
    .SN(_02636_));
 HAxp5_ASAP7_75t_R _21195_ (.A(\xs[11].cli0.r[0] ),
    .B(\xs[11].cli0.r[1] ),
    .CON(_02637_),
    .SN(_02638_));
 HAxp5_ASAP7_75t_R _21196_ (.A(\xs[6].cli1.r[0] ),
    .B(\xs[6].cli1.r[1] ),
    .CON(_02639_),
    .SN(_02640_));
 HAxp5_ASAP7_75t_R _21197_ (.A(\xs[4].cli1.r[0] ),
    .B(\xs[4].cli1.r[1] ),
    .CON(_02641_),
    .SN(_02642_));
 HAxp5_ASAP7_75t_R _21198_ (.A(\xs[11].cli1.r[0] ),
    .B(\xs[11].cli1.r[1] ),
    .CON(_02643_),
    .SN(_02644_));
 HAxp5_ASAP7_75t_R _21199_ (.A(\xs[13].cli0.r[0] ),
    .B(\xs[13].cli0.r[1] ),
    .CON(_02645_),
    .SN(_02646_));
 HAxp5_ASAP7_75t_R _21200_ (.A(\xs[9].cli0.r[0] ),
    .B(\xs[9].cli0.r[1] ),
    .CON(_02647_),
    .SN(_02648_));
 HAxp5_ASAP7_75t_R _21201_ (.A(\xs[5].cli0.r[0] ),
    .B(\xs[5].cli0.r[1] ),
    .CON(_02649_),
    .SN(_02650_));
 HAxp5_ASAP7_75t_R _21202_ (.A(\xs[7].cli0.r[0] ),
    .B(\xs[7].cli0.r[1] ),
    .CON(_02651_),
    .SN(_02652_));
 HAxp5_ASAP7_75t_R _21203_ (.A(\xs[9].cli1.r[0] ),
    .B(\xs[9].cli1.r[1] ),
    .CON(_02653_),
    .SN(_02654_));
 HAxp5_ASAP7_75t_R _21204_ (.A(\xs[12].cli0.r[0] ),
    .B(\xs[12].cli0.r[1] ),
    .CON(_02655_),
    .SN(_02656_));
 HAxp5_ASAP7_75t_R _21205_ (.A(\xs[3].cli0.r[0] ),
    .B(\xs[3].cli0.r[1] ),
    .CON(_02657_),
    .SN(_02658_));
 HAxp5_ASAP7_75t_R _21206_ (.A(\xs[1].cli1.r[0] ),
    .B(\xs[1].cli1.r[1] ),
    .CON(_02659_),
    .SN(_02660_));
 HAxp5_ASAP7_75t_R _21207_ (.A(\xs[4].cli0.r[0] ),
    .B(\xs[4].cli0.r[1] ),
    .CON(_02661_),
    .SN(_02662_));
 HAxp5_ASAP7_75t_R _21208_ (.A(\xs[14].cli0.r[0] ),
    .B(\xs[14].cli0.r[1] ),
    .CON(_02663_),
    .SN(_02664_));
 HAxp5_ASAP7_75t_R _21209_ (.A(\xs[7].cli1.r[0] ),
    .B(\xs[7].cli1.r[1] ),
    .CON(_02665_),
    .SN(_02666_));
 HAxp5_ASAP7_75t_R _21210_ (.A(\xs[3].cli1.r[0] ),
    .B(\xs[3].cli1.r[1] ),
    .CON(_02667_),
    .SN(_02668_));
 HAxp5_ASAP7_75t_R _21211_ (.A(\xs[2].cli0.r[0] ),
    .B(\xs[2].cli0.r[1] ),
    .CON(_02669_),
    .SN(_02670_));
 HAxp5_ASAP7_75t_R _21212_ (.A(\xs[8].cli0.r[0] ),
    .B(\xs[8].cli0.r[1] ),
    .CON(_02671_),
    .SN(_02672_));
 HAxp5_ASAP7_75t_R _21213_ (.A(\xs[2].cli1.r[0] ),
    .B(\xs[2].cli1.r[1] ),
    .CON(_02673_),
    .SN(_02674_));
 BUFx24_ASAP7_75t_R clkbuf_leaf_0_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_0_clk));
 BUFx2_ASAP7_75t_R _21215_ (.A(net326),
    .Y(done_all));
 BUFx2_ASAP7_75t_R _21216_ (.A(net327),
    .Y(out[1]));
 BUFx2_ASAP7_75t_R _21217_ (.A(net328),
    .Y(out[2]));
 BUFx2_ASAP7_75t_R _21218_ (.A(net329),
    .Y(out[3]));
 BUFx2_ASAP7_75t_R _21219_ (.A(net330),
    .Y(out[4]));
 BUFx2_ASAP7_75t_R _21220_ (.A(net331),
    .Y(out[5]));
 BUFx2_ASAP7_75t_R _21221_ (.A(net332),
    .Y(out[6]));
 BUFx2_ASAP7_75t_R _21222_ (.A(net333),
    .Y(out[7]));
 BUFx2_ASAP7_75t_R _21223_ (.A(net334),
    .Y(out[8]));
 BUFx2_ASAP7_75t_R _21224_ (.A(net335),
    .Y(out[9]));
 BUFx2_ASAP7_75t_R _21225_ (.A(net336),
    .Y(out[10]));
 BUFx2_ASAP7_75t_R _21226_ (.A(net337),
    .Y(out[11]));
 BUFx2_ASAP7_75t_R _21227_ (.A(net338),
    .Y(out[12]));
 BUFx2_ASAP7_75t_R _21228_ (.A(net339),
    .Y(out[13]));
 BUFx2_ASAP7_75t_R _21229_ (.A(net340),
    .Y(out[14]));
 BUFx2_ASAP7_75t_R _21230_ (.A(net341),
    .Y(out[15]));
 BUFx2_ASAP7_75t_R _21231_ (.A(net342),
    .Y(out[16]));
 BUFx2_ASAP7_75t_R _21232_ (.A(net343),
    .Y(out[17]));
 BUFx2_ASAP7_75t_R _21233_ (.A(net344),
    .Y(out[18]));
 BUFx2_ASAP7_75t_R _21234_ (.A(net345),
    .Y(out[19]));
 BUFx2_ASAP7_75t_R _21235_ (.A(net346),
    .Y(out[20]));
 BUFx2_ASAP7_75t_R _21236_ (.A(net347),
    .Y(out[21]));
 BUFx2_ASAP7_75t_R _21237_ (.A(net348),
    .Y(out[22]));
 BUFx2_ASAP7_75t_R _21238_ (.A(net349),
    .Y(out[23]));
 BUFx2_ASAP7_75t_R _21239_ (.A(net350),
    .Y(out[24]));
 BUFx2_ASAP7_75t_R _21240_ (.A(net351),
    .Y(out[25]));
 BUFx2_ASAP7_75t_R _21241_ (.A(net352),
    .Y(out[26]));
 BUFx2_ASAP7_75t_R _21242_ (.A(net353),
    .Y(out[27]));
 BUFx2_ASAP7_75t_R _21243_ (.A(net354),
    .Y(out[28]));
 BUFx2_ASAP7_75t_R _21244_ (.A(net355),
    .Y(out[29]));
 BUFx2_ASAP7_75t_R _21245_ (.A(net356),
    .Y(out[30]));
 BUFx2_ASAP7_75t_R _21246_ (.A(net357),
    .Y(out[31]));
 BUFx2_ASAP7_75t_R _21247_ (.A(net358),
    .Y(out[37]));
 BUFx2_ASAP7_75t_R _21248_ (.A(net359),
    .Y(out[38]));
 BUFx2_ASAP7_75t_R _21249_ (.A(net360),
    .Y(out[41]));
 BUFx2_ASAP7_75t_R _21250_ (.A(net361),
    .Y(out[42]));
 BUFx2_ASAP7_75t_R _21251_ (.A(net362),
    .Y(out[43]));
 BUFx2_ASAP7_75t_R _21252_ (.A(net363),
    .Y(out[44]));
 BUFx2_ASAP7_75t_R _21253_ (.A(net364),
    .Y(out[45]));
 BUFx2_ASAP7_75t_R _21254_ (.A(net365),
    .Y(out[46]));
 BUFx2_ASAP7_75t_R _21255_ (.A(net366),
    .Y(out[47]));
 BUFx2_ASAP7_75t_R _21256_ (.A(net367),
    .Y(out[48]));
 BUFx2_ASAP7_75t_R _21257_ (.A(net368),
    .Y(out[49]));
 BUFx2_ASAP7_75t_R _21258_ (.A(net369),
    .Y(out[51]));
 BUFx2_ASAP7_75t_R _21259_ (.A(net370),
    .Y(out[52]));
 BUFx2_ASAP7_75t_R _21260_ (.A(net371),
    .Y(out[53]));
 BUFx2_ASAP7_75t_R _21261_ (.A(net372),
    .Y(out[54]));
 BUFx2_ASAP7_75t_R _21262_ (.A(net373),
    .Y(out[55]));
 BUFx2_ASAP7_75t_R _21263_ (.A(net374),
    .Y(out[56]));
 BUFx2_ASAP7_75t_R _21264_ (.A(net375),
    .Y(out[57]));
 BUFx2_ASAP7_75t_R _21265_ (.A(net376),
    .Y(out[58]));
 BUFx2_ASAP7_75t_R _21266_ (.A(net377),
    .Y(out[59]));
 BUFx2_ASAP7_75t_R _21267_ (.A(net378),
    .Y(out[60]));
 BUFx2_ASAP7_75t_R _21268_ (.A(net379),
    .Y(out[61]));
 BUFx2_ASAP7_75t_R _21269_ (.A(net380),
    .Y(out[62]));
 BUFx2_ASAP7_75t_R _21270_ (.A(net381),
    .Y(out[63]));
 BUFx2_ASAP7_75t_R _21271_ (.A(net382),
    .Y(out[64]));
 BUFx2_ASAP7_75t_R _21272_ (.A(net383),
    .Y(out[65]));
 BUFx2_ASAP7_75t_R _21273_ (.A(net384),
    .Y(out[66]));
 BUFx2_ASAP7_75t_R _21274_ (.A(net385),
    .Y(out[67]));
 BUFx2_ASAP7_75t_R _21275_ (.A(net386),
    .Y(out[68]));
 BUFx2_ASAP7_75t_R _21276_ (.A(net387),
    .Y(out[69]));
 BUFx2_ASAP7_75t_R _21277_ (.A(net388),
    .Y(out[70]));
 BUFx2_ASAP7_75t_R _21278_ (.A(net389),
    .Y(out[71]));
 BUFx2_ASAP7_75t_R _21279_ (.A(net390),
    .Y(out[77]));
 BUFx2_ASAP7_75t_R _21280_ (.A(net391),
    .Y(out[78]));
 BUFx2_ASAP7_75t_R _21281_ (.A(net392),
    .Y(out[81]));
 BUFx2_ASAP7_75t_R _21282_ (.A(net393),
    .Y(out[82]));
 BUFx2_ASAP7_75t_R _21283_ (.A(net394),
    .Y(out[83]));
 BUFx2_ASAP7_75t_R _21284_ (.A(net395),
    .Y(out[84]));
 BUFx2_ASAP7_75t_R _21285_ (.A(net396),
    .Y(out[85]));
 BUFx2_ASAP7_75t_R _21286_ (.A(net397),
    .Y(out[86]));
 BUFx2_ASAP7_75t_R _21287_ (.A(net398),
    .Y(out[87]));
 BUFx2_ASAP7_75t_R _21288_ (.A(net399),
    .Y(out[88]));
 BUFx2_ASAP7_75t_R _21289_ (.A(net400),
    .Y(out[89]));
 BUFx2_ASAP7_75t_R _21290_ (.A(net401),
    .Y(out[90]));
 BUFx2_ASAP7_75t_R _21291_ (.A(net402),
    .Y(out[92]));
 BUFx2_ASAP7_75t_R _21292_ (.A(net403),
    .Y(out[93]));
 BUFx2_ASAP7_75t_R _21293_ (.A(net404),
    .Y(out[94]));
 BUFx2_ASAP7_75t_R _21294_ (.A(net405),
    .Y(out[95]));
 BUFx2_ASAP7_75t_R _21295_ (.A(net406),
    .Y(out[96]));
 BUFx2_ASAP7_75t_R _21296_ (.A(net407),
    .Y(out[97]));
 BUFx2_ASAP7_75t_R _21297_ (.A(net408),
    .Y(out[98]));
 BUFx2_ASAP7_75t_R _21298_ (.A(net409),
    .Y(out[99]));
 BUFx2_ASAP7_75t_R _21299_ (.A(net410),
    .Y(out[100]));
 BUFx2_ASAP7_75t_R _21300_ (.A(net411),
    .Y(out[101]));
 BUFx2_ASAP7_75t_R _21301_ (.A(net412),
    .Y(out[102]));
 BUFx2_ASAP7_75t_R _21302_ (.A(net413),
    .Y(out[103]));
 BUFx2_ASAP7_75t_R _21303_ (.A(net414),
    .Y(out[104]));
 BUFx2_ASAP7_75t_R _21304_ (.A(net415),
    .Y(out[105]));
 BUFx2_ASAP7_75t_R _21305_ (.A(net416),
    .Y(out[106]));
 BUFx2_ASAP7_75t_R _21306_ (.A(net417),
    .Y(out[107]));
 BUFx2_ASAP7_75t_R _21307_ (.A(net418),
    .Y(out[108]));
 BUFx2_ASAP7_75t_R _21308_ (.A(net419),
    .Y(out[109]));
 BUFx2_ASAP7_75t_R _21309_ (.A(net420),
    .Y(out[110]));
 BUFx2_ASAP7_75t_R _21310_ (.A(net421),
    .Y(out[111]));
 BUFx2_ASAP7_75t_R _21311_ (.A(net422),
    .Y(out[117]));
 BUFx2_ASAP7_75t_R _21312_ (.A(net423),
    .Y(out[118]));
 BUFx2_ASAP7_75t_R _21313_ (.A(net424),
    .Y(out[121]));
 BUFx2_ASAP7_75t_R _21314_ (.A(net425),
    .Y(out[122]));
 BUFx2_ASAP7_75t_R _21315_ (.A(net426),
    .Y(out[123]));
 BUFx2_ASAP7_75t_R _21316_ (.A(net427),
    .Y(out[124]));
 BUFx2_ASAP7_75t_R _21317_ (.A(net428),
    .Y(out[125]));
 BUFx2_ASAP7_75t_R _21318_ (.A(net429),
    .Y(out[126]));
 BUFx2_ASAP7_75t_R _21319_ (.A(net430),
    .Y(out[127]));
 BUFx2_ASAP7_75t_R _21320_ (.A(net431),
    .Y(out[128]));
 BUFx2_ASAP7_75t_R _21321_ (.A(net432),
    .Y(out[129]));
 BUFx3_ASAP7_75t_R _21322_ (.A(net106),
    .Y(net105));
 BUFx2_ASAP7_75t_R _21323_ (.A(net433),
    .Y(out[132]));
 BUFx2_ASAP7_75t_R _21324_ (.A(net434),
    .Y(out[133]));
 BUFx2_ASAP7_75t_R _21325_ (.A(net435),
    .Y(out[134]));
 BUFx2_ASAP7_75t_R _21326_ (.A(net436),
    .Y(out[135]));
 BUFx2_ASAP7_75t_R _21327_ (.A(net437),
    .Y(out[136]));
 BUFx2_ASAP7_75t_R _21328_ (.A(net438),
    .Y(out[137]));
 BUFx2_ASAP7_75t_R _21329_ (.A(net439),
    .Y(out[138]));
 BUFx2_ASAP7_75t_R _21330_ (.A(net440),
    .Y(out[139]));
 BUFx2_ASAP7_75t_R _21331_ (.A(net441),
    .Y(out[140]));
 BUFx2_ASAP7_75t_R _21332_ (.A(net442),
    .Y(out[141]));
 BUFx2_ASAP7_75t_R _21333_ (.A(net443),
    .Y(out[142]));
 BUFx2_ASAP7_75t_R _21334_ (.A(net444),
    .Y(out[143]));
 BUFx2_ASAP7_75t_R _21335_ (.A(net445),
    .Y(out[144]));
 BUFx2_ASAP7_75t_R _21336_ (.A(net446),
    .Y(out[145]));
 BUFx2_ASAP7_75t_R _21337_ (.A(net447),
    .Y(out[146]));
 BUFx2_ASAP7_75t_R _21338_ (.A(net448),
    .Y(out[147]));
 BUFx2_ASAP7_75t_R _21339_ (.A(net449),
    .Y(out[148]));
 BUFx2_ASAP7_75t_R _21340_ (.A(net450),
    .Y(out[149]));
 BUFx2_ASAP7_75t_R _21341_ (.A(net451),
    .Y(out[150]));
 BUFx2_ASAP7_75t_R _21342_ (.A(net452),
    .Y(out[151]));
 BUFx2_ASAP7_75t_R _21343_ (.A(net453),
    .Y(out[157]));
 BUFx2_ASAP7_75t_R _21344_ (.A(net454),
    .Y(out[158]));
 BUFx2_ASAP7_75t_R _21345_ (.A(net455),
    .Y(out[161]));
 BUFx2_ASAP7_75t_R _21346_ (.A(net456),
    .Y(out[162]));
 BUFx2_ASAP7_75t_R _21347_ (.A(net457),
    .Y(out[163]));
 BUFx2_ASAP7_75t_R _21348_ (.A(net458),
    .Y(out[164]));
 BUFx2_ASAP7_75t_R _21349_ (.A(net459),
    .Y(out[165]));
 BUFx2_ASAP7_75t_R _21350_ (.A(net460),
    .Y(out[166]));
 BUFx2_ASAP7_75t_R _21351_ (.A(net461),
    .Y(out[167]));
 BUFx2_ASAP7_75t_R _21352_ (.A(net462),
    .Y(out[168]));
 BUFx2_ASAP7_75t_R _21353_ (.A(net463),
    .Y(out[169]));
 BUFx2_ASAP7_75t_R _21354_ (.A(net464),
    .Y(out[170]));
 BUFx2_ASAP7_75t_R _21355_ (.A(net465),
    .Y(out[171]));
 BUFx2_ASAP7_75t_R _21356_ (.A(net466),
    .Y(out[173]));
 BUFx2_ASAP7_75t_R _21357_ (.A(net467),
    .Y(out[174]));
 BUFx2_ASAP7_75t_R _21358_ (.A(net468),
    .Y(out[175]));
 BUFx2_ASAP7_75t_R _21359_ (.A(net469),
    .Y(out[176]));
 BUFx2_ASAP7_75t_R _21360_ (.A(net470),
    .Y(out[177]));
 BUFx2_ASAP7_75t_R _21361_ (.A(net471),
    .Y(out[178]));
 BUFx2_ASAP7_75t_R _21362_ (.A(net472),
    .Y(out[179]));
 BUFx2_ASAP7_75t_R _21363_ (.A(net473),
    .Y(out[180]));
 BUFx2_ASAP7_75t_R _21364_ (.A(net474),
    .Y(out[181]));
 BUFx2_ASAP7_75t_R _21365_ (.A(net475),
    .Y(out[182]));
 BUFx2_ASAP7_75t_R _21366_ (.A(net476),
    .Y(out[183]));
 BUFx2_ASAP7_75t_R _21367_ (.A(net477),
    .Y(out[184]));
 BUFx2_ASAP7_75t_R _21368_ (.A(net478),
    .Y(out[185]));
 BUFx2_ASAP7_75t_R _21369_ (.A(net479),
    .Y(out[186]));
 BUFx2_ASAP7_75t_R _21370_ (.A(net480),
    .Y(out[187]));
 BUFx2_ASAP7_75t_R _21371_ (.A(net481),
    .Y(out[188]));
 BUFx2_ASAP7_75t_R _21372_ (.A(net482),
    .Y(out[189]));
 BUFx2_ASAP7_75t_R _21373_ (.A(net483),
    .Y(out[190]));
 BUFx2_ASAP7_75t_R _21374_ (.A(net484),
    .Y(out[191]));
 BUFx2_ASAP7_75t_R _21375_ (.A(net485),
    .Y(out[197]));
 BUFx2_ASAP7_75t_R _21376_ (.A(net486),
    .Y(out[198]));
 BUFx2_ASAP7_75t_R _21377_ (.A(net487),
    .Y(out[201]));
 BUFx2_ASAP7_75t_R _21378_ (.A(net488),
    .Y(out[202]));
 BUFx2_ASAP7_75t_R _21379_ (.A(net489),
    .Y(out[203]));
 BUFx2_ASAP7_75t_R _21380_ (.A(net490),
    .Y(out[204]));
 BUFx2_ASAP7_75t_R _21381_ (.A(net491),
    .Y(out[205]));
 BUFx2_ASAP7_75t_R _21382_ (.A(net492),
    .Y(out[206]));
 BUFx2_ASAP7_75t_R _21383_ (.A(net493),
    .Y(out[207]));
 BUFx2_ASAP7_75t_R _21384_ (.A(net494),
    .Y(out[208]));
 BUFx2_ASAP7_75t_R _21385_ (.A(net495),
    .Y(out[209]));
 BUFx3_ASAP7_75t_R _21386_ (.A(net123),
    .Y(net122));
 BUFx2_ASAP7_75t_R _21387_ (.A(net496),
    .Y(out[211]));
 BUFx2_ASAP7_75t_R _21388_ (.A(net497),
    .Y(out[213]));
 BUFx2_ASAP7_75t_R _21389_ (.A(net498),
    .Y(out[214]));
 BUFx2_ASAP7_75t_R _21390_ (.A(net499),
    .Y(out[215]));
 BUFx2_ASAP7_75t_R _21391_ (.A(net500),
    .Y(out[216]));
 BUFx2_ASAP7_75t_R _21392_ (.A(net501),
    .Y(out[217]));
 BUFx2_ASAP7_75t_R _21393_ (.A(net502),
    .Y(out[218]));
 BUFx2_ASAP7_75t_R _21394_ (.A(net503),
    .Y(out[219]));
 BUFx2_ASAP7_75t_R _21395_ (.A(net504),
    .Y(out[220]));
 BUFx2_ASAP7_75t_R _21396_ (.A(net505),
    .Y(out[221]));
 BUFx2_ASAP7_75t_R _21397_ (.A(net506),
    .Y(out[222]));
 BUFx2_ASAP7_75t_R _21398_ (.A(net507),
    .Y(out[223]));
 BUFx2_ASAP7_75t_R _21399_ (.A(net508),
    .Y(out[224]));
 BUFx2_ASAP7_75t_R _21400_ (.A(net509),
    .Y(out[225]));
 BUFx2_ASAP7_75t_R _21401_ (.A(net510),
    .Y(out[226]));
 BUFx2_ASAP7_75t_R _21402_ (.A(net511),
    .Y(out[227]));
 BUFx2_ASAP7_75t_R _21403_ (.A(net512),
    .Y(out[228]));
 BUFx2_ASAP7_75t_R _21404_ (.A(net513),
    .Y(out[229]));
 BUFx2_ASAP7_75t_R _21405_ (.A(net514),
    .Y(out[230]));
 BUFx2_ASAP7_75t_R _21406_ (.A(net515),
    .Y(out[231]));
 BUFx2_ASAP7_75t_R _21407_ (.A(net516),
    .Y(out[237]));
 BUFx2_ASAP7_75t_R _21408_ (.A(net517),
    .Y(out[238]));
 BUFx2_ASAP7_75t_R _21409_ (.A(net518),
    .Y(out[241]));
 BUFx2_ASAP7_75t_R _21410_ (.A(net519),
    .Y(out[242]));
 BUFx2_ASAP7_75t_R _21411_ (.A(net520),
    .Y(out[243]));
 BUFx2_ASAP7_75t_R _21412_ (.A(net521),
    .Y(out[244]));
 BUFx2_ASAP7_75t_R _21413_ (.A(net522),
    .Y(out[245]));
 BUFx2_ASAP7_75t_R _21414_ (.A(net523),
    .Y(out[246]));
 BUFx2_ASAP7_75t_R _21415_ (.A(net524),
    .Y(out[247]));
 BUFx2_ASAP7_75t_R _21416_ (.A(net525),
    .Y(out[248]));
 BUFx2_ASAP7_75t_R _21417_ (.A(net526),
    .Y(out[249]));
 BUFx2_ASAP7_75t_R _21418_ (.A(net527),
    .Y(out[250]));
 BUFx3_ASAP7_75t_R _21419_ (.A(net132),
    .Y(net131));
 BUFx2_ASAP7_75t_R _21420_ (.A(net528),
    .Y(out[253]));
 BUFx2_ASAP7_75t_R _21421_ (.A(net529),
    .Y(out[254]));
 BUFx2_ASAP7_75t_R _21422_ (.A(net530),
    .Y(out[255]));
 BUFx2_ASAP7_75t_R _21423_ (.A(net531),
    .Y(out[256]));
 BUFx2_ASAP7_75t_R _21424_ (.A(net532),
    .Y(out[257]));
 BUFx2_ASAP7_75t_R _21425_ (.A(net533),
    .Y(out[258]));
 BUFx2_ASAP7_75t_R _21426_ (.A(net534),
    .Y(out[259]));
 BUFx2_ASAP7_75t_R _21427_ (.A(net535),
    .Y(out[260]));
 BUFx2_ASAP7_75t_R _21428_ (.A(net536),
    .Y(out[261]));
 BUFx2_ASAP7_75t_R _21429_ (.A(net537),
    .Y(out[262]));
 BUFx2_ASAP7_75t_R _21430_ (.A(net538),
    .Y(out[263]));
 BUFx2_ASAP7_75t_R _21431_ (.A(net539),
    .Y(out[264]));
 BUFx2_ASAP7_75t_R _21432_ (.A(net540),
    .Y(out[265]));
 BUFx2_ASAP7_75t_R _21433_ (.A(net541),
    .Y(out[266]));
 BUFx2_ASAP7_75t_R _21434_ (.A(net542),
    .Y(out[267]));
 BUFx2_ASAP7_75t_R _21435_ (.A(net543),
    .Y(out[268]));
 BUFx2_ASAP7_75t_R _21436_ (.A(net544),
    .Y(out[269]));
 BUFx2_ASAP7_75t_R _21437_ (.A(net545),
    .Y(out[270]));
 BUFx2_ASAP7_75t_R _21438_ (.A(net546),
    .Y(out[271]));
 BUFx2_ASAP7_75t_R _21439_ (.A(net547),
    .Y(out[277]));
 BUFx2_ASAP7_75t_R _21440_ (.A(net548),
    .Y(out[278]));
 BUFx2_ASAP7_75t_R _21441_ (.A(net549),
    .Y(out[281]));
 BUFx2_ASAP7_75t_R _21442_ (.A(net550),
    .Y(out[282]));
 BUFx2_ASAP7_75t_R _21443_ (.A(net551),
    .Y(out[283]));
 BUFx2_ASAP7_75t_R _21444_ (.A(net552),
    .Y(out[284]));
 BUFx2_ASAP7_75t_R _21445_ (.A(net553),
    .Y(out[285]));
 BUFx2_ASAP7_75t_R _21446_ (.A(net554),
    .Y(out[286]));
 BUFx2_ASAP7_75t_R _21447_ (.A(net555),
    .Y(out[287]));
 BUFx2_ASAP7_75t_R _21448_ (.A(net556),
    .Y(out[288]));
 BUFx2_ASAP7_75t_R _21449_ (.A(net557),
    .Y(out[289]));
 BUFx3_ASAP7_75t_R _21450_ (.A(net142),
    .Y(net140));
 BUFx3_ASAP7_75t_R _21451_ (.A(net142),
    .Y(net141));
 BUFx2_ASAP7_75t_R _21452_ (.A(net558),
    .Y(out[293]));
 BUFx2_ASAP7_75t_R _21453_ (.A(net559),
    .Y(out[294]));
 BUFx2_ASAP7_75t_R _21454_ (.A(net560),
    .Y(out[295]));
 BUFx2_ASAP7_75t_R _21455_ (.A(net561),
    .Y(out[296]));
 BUFx2_ASAP7_75t_R _21456_ (.A(net562),
    .Y(out[297]));
 BUFx2_ASAP7_75t_R _21457_ (.A(net563),
    .Y(out[298]));
 BUFx2_ASAP7_75t_R _21458_ (.A(net564),
    .Y(out[299]));
 BUFx2_ASAP7_75t_R _21459_ (.A(net565),
    .Y(out[300]));
 BUFx2_ASAP7_75t_R _21460_ (.A(net566),
    .Y(out[301]));
 BUFx2_ASAP7_75t_R _21461_ (.A(net567),
    .Y(out[302]));
 BUFx2_ASAP7_75t_R _21462_ (.A(net568),
    .Y(out[303]));
 BUFx2_ASAP7_75t_R _21463_ (.A(net569),
    .Y(out[304]));
 BUFx2_ASAP7_75t_R _21464_ (.A(net570),
    .Y(out[305]));
 BUFx2_ASAP7_75t_R _21465_ (.A(net571),
    .Y(out[306]));
 BUFx2_ASAP7_75t_R _21466_ (.A(net572),
    .Y(out[307]));
 BUFx2_ASAP7_75t_R _21467_ (.A(net573),
    .Y(out[308]));
 BUFx2_ASAP7_75t_R _21468_ (.A(net574),
    .Y(out[309]));
 BUFx2_ASAP7_75t_R _21469_ (.A(net575),
    .Y(out[310]));
 BUFx2_ASAP7_75t_R _21470_ (.A(net576),
    .Y(out[311]));
 BUFx2_ASAP7_75t_R _21471_ (.A(net577),
    .Y(out[317]));
 BUFx2_ASAP7_75t_R _21472_ (.A(net578),
    .Y(out[318]));
 BUFx2_ASAP7_75t_R _21473_ (.A(net579),
    .Y(out[321]));
 BUFx2_ASAP7_75t_R _21474_ (.A(net580),
    .Y(out[322]));
 BUFx2_ASAP7_75t_R _21475_ (.A(net581),
    .Y(out[323]));
 BUFx2_ASAP7_75t_R _21476_ (.A(net582),
    .Y(out[324]));
 BUFx2_ASAP7_75t_R _21477_ (.A(net583),
    .Y(out[325]));
 BUFx2_ASAP7_75t_R _21478_ (.A(net584),
    .Y(out[326]));
 BUFx2_ASAP7_75t_R _21479_ (.A(net585),
    .Y(out[327]));
 BUFx2_ASAP7_75t_R _21480_ (.A(net586),
    .Y(out[328]));
 BUFx2_ASAP7_75t_R _21481_ (.A(net587),
    .Y(out[329]));
 BUFx2_ASAP7_75t_R _21482_ (.A(net588),
    .Y(out[330]));
 BUFx2_ASAP7_75t_R _21483_ (.A(net589),
    .Y(out[331]));
 BUFx2_ASAP7_75t_R _21484_ (.A(net590),
    .Y(out[332]));
 BUFx2_ASAP7_75t_R _21485_ (.A(net591),
    .Y(out[334]));
 BUFx2_ASAP7_75t_R _21486_ (.A(net592),
    .Y(out[335]));
 BUFx2_ASAP7_75t_R _21487_ (.A(net593),
    .Y(out[336]));
 BUFx2_ASAP7_75t_R _21488_ (.A(net594),
    .Y(out[337]));
 BUFx2_ASAP7_75t_R _21489_ (.A(net595),
    .Y(out[338]));
 BUFx2_ASAP7_75t_R _21490_ (.A(net596),
    .Y(out[339]));
 BUFx2_ASAP7_75t_R _21491_ (.A(net597),
    .Y(out[340]));
 BUFx2_ASAP7_75t_R _21492_ (.A(net598),
    .Y(out[341]));
 BUFx2_ASAP7_75t_R _21493_ (.A(net599),
    .Y(out[342]));
 BUFx2_ASAP7_75t_R _21494_ (.A(net600),
    .Y(out[343]));
 BUFx2_ASAP7_75t_R _21495_ (.A(net601),
    .Y(out[344]));
 BUFx2_ASAP7_75t_R _21496_ (.A(net602),
    .Y(out[345]));
 BUFx2_ASAP7_75t_R _21497_ (.A(net603),
    .Y(out[346]));
 BUFx2_ASAP7_75t_R _21498_ (.A(net604),
    .Y(out[347]));
 BUFx2_ASAP7_75t_R _21499_ (.A(net605),
    .Y(out[348]));
 BUFx2_ASAP7_75t_R _21500_ (.A(net606),
    .Y(out[349]));
 BUFx2_ASAP7_75t_R _21501_ (.A(net607),
    .Y(out[350]));
 BUFx2_ASAP7_75t_R _21502_ (.A(net608),
    .Y(out[351]));
 BUFx2_ASAP7_75t_R _21503_ (.A(net609),
    .Y(out[357]));
 BUFx2_ASAP7_75t_R _21504_ (.A(net610),
    .Y(out[358]));
 BUFx2_ASAP7_75t_R _21505_ (.A(net611),
    .Y(out[361]));
 BUFx2_ASAP7_75t_R _21506_ (.A(net612),
    .Y(out[362]));
 BUFx2_ASAP7_75t_R _21507_ (.A(net613),
    .Y(out[363]));
 BUFx2_ASAP7_75t_R _21508_ (.A(net614),
    .Y(out[364]));
 BUFx2_ASAP7_75t_R _21509_ (.A(net615),
    .Y(out[365]));
 BUFx2_ASAP7_75t_R _21510_ (.A(net616),
    .Y(out[366]));
 BUFx2_ASAP7_75t_R _21511_ (.A(net617),
    .Y(out[367]));
 BUFx2_ASAP7_75t_R _21512_ (.A(net618),
    .Y(out[368]));
 BUFx2_ASAP7_75t_R _21513_ (.A(net619),
    .Y(out[369]));
 BUFx3_ASAP7_75t_R _21514_ (.A(net164),
    .Y(net163));
 BUFx2_ASAP7_75t_R _21515_ (.A(net620),
    .Y(out[371]));
 BUFx2_ASAP7_75t_R _21516_ (.A(net621),
    .Y(out[372]));
 BUFx2_ASAP7_75t_R _21517_ (.A(net622),
    .Y(out[374]));
 BUFx2_ASAP7_75t_R _21518_ (.A(net623),
    .Y(out[375]));
 BUFx2_ASAP7_75t_R _21519_ (.A(net624),
    .Y(out[376]));
 BUFx2_ASAP7_75t_R _21520_ (.A(net625),
    .Y(out[377]));
 BUFx2_ASAP7_75t_R _21521_ (.A(net626),
    .Y(out[378]));
 BUFx2_ASAP7_75t_R _21522_ (.A(net627),
    .Y(out[379]));
 BUFx2_ASAP7_75t_R _21523_ (.A(net628),
    .Y(out[380]));
 BUFx2_ASAP7_75t_R _21524_ (.A(net629),
    .Y(out[381]));
 BUFx2_ASAP7_75t_R _21525_ (.A(net630),
    .Y(out[382]));
 BUFx2_ASAP7_75t_R _21526_ (.A(net631),
    .Y(out[383]));
 BUFx2_ASAP7_75t_R _21527_ (.A(net632),
    .Y(out[384]));
 BUFx2_ASAP7_75t_R _21528_ (.A(net633),
    .Y(out[385]));
 BUFx2_ASAP7_75t_R _21529_ (.A(net634),
    .Y(out[386]));
 BUFx2_ASAP7_75t_R _21530_ (.A(net635),
    .Y(out[387]));
 BUFx2_ASAP7_75t_R _21531_ (.A(net636),
    .Y(out[388]));
 BUFx2_ASAP7_75t_R _21532_ (.A(net637),
    .Y(out[389]));
 BUFx2_ASAP7_75t_R _21533_ (.A(net638),
    .Y(out[390]));
 BUFx2_ASAP7_75t_R _21534_ (.A(net639),
    .Y(out[391]));
 BUFx2_ASAP7_75t_R _21535_ (.A(net640),
    .Y(out[397]));
 BUFx2_ASAP7_75t_R _21536_ (.A(net641),
    .Y(out[398]));
 BUFx2_ASAP7_75t_R _21537_ (.A(net642),
    .Y(out[401]));
 BUFx2_ASAP7_75t_R _21538_ (.A(net643),
    .Y(out[402]));
 BUFx2_ASAP7_75t_R _21539_ (.A(net644),
    .Y(out[403]));
 BUFx2_ASAP7_75t_R _21540_ (.A(net645),
    .Y(out[404]));
 BUFx2_ASAP7_75t_R _21541_ (.A(net646),
    .Y(out[405]));
 BUFx2_ASAP7_75t_R _21542_ (.A(net647),
    .Y(out[406]));
 BUFx2_ASAP7_75t_R _21543_ (.A(net648),
    .Y(out[407]));
 BUFx2_ASAP7_75t_R _21544_ (.A(net649),
    .Y(out[408]));
 BUFx2_ASAP7_75t_R _21545_ (.A(net650),
    .Y(out[409]));
 BUFx2_ASAP7_75t_R _21546_ (.A(net651),
    .Y(out[410]));
 BUFx3_ASAP7_75t_R _21547_ (.A(net175),
    .Y(net174));
 BUFx2_ASAP7_75t_R _21548_ (.A(net652),
    .Y(out[412]));
 BUFx2_ASAP7_75t_R _21549_ (.A(net653),
    .Y(out[414]));
 BUFx2_ASAP7_75t_R _21550_ (.A(net654),
    .Y(out[415]));
 BUFx2_ASAP7_75t_R _21551_ (.A(net655),
    .Y(out[416]));
 BUFx2_ASAP7_75t_R _21552_ (.A(net656),
    .Y(out[417]));
 BUFx2_ASAP7_75t_R _21553_ (.A(net657),
    .Y(out[418]));
 BUFx2_ASAP7_75t_R _21554_ (.A(net658),
    .Y(out[419]));
 BUFx2_ASAP7_75t_R _21555_ (.A(net659),
    .Y(out[420]));
 BUFx2_ASAP7_75t_R _21556_ (.A(net660),
    .Y(out[421]));
 BUFx2_ASAP7_75t_R _21557_ (.A(net661),
    .Y(out[422]));
 BUFx2_ASAP7_75t_R _21558_ (.A(net662),
    .Y(out[423]));
 BUFx2_ASAP7_75t_R _21559_ (.A(net663),
    .Y(out[424]));
 BUFx2_ASAP7_75t_R _21560_ (.A(net664),
    .Y(out[425]));
 BUFx2_ASAP7_75t_R _21561_ (.A(net665),
    .Y(out[426]));
 BUFx2_ASAP7_75t_R _21562_ (.A(net666),
    .Y(out[427]));
 BUFx2_ASAP7_75t_R _21563_ (.A(net667),
    .Y(out[428]));
 BUFx2_ASAP7_75t_R _21564_ (.A(net668),
    .Y(out[429]));
 BUFx2_ASAP7_75t_R _21565_ (.A(net669),
    .Y(out[430]));
 BUFx2_ASAP7_75t_R _21566_ (.A(net670),
    .Y(out[431]));
 BUFx2_ASAP7_75t_R _21567_ (.A(net671),
    .Y(out[437]));
 BUFx2_ASAP7_75t_R _21568_ (.A(net672),
    .Y(out[438]));
 BUFx2_ASAP7_75t_R _21569_ (.A(net673),
    .Y(out[441]));
 BUFx2_ASAP7_75t_R _21570_ (.A(net674),
    .Y(out[442]));
 BUFx2_ASAP7_75t_R _21571_ (.A(net675),
    .Y(out[443]));
 BUFx2_ASAP7_75t_R _21572_ (.A(net676),
    .Y(out[444]));
 BUFx2_ASAP7_75t_R _21573_ (.A(net677),
    .Y(out[445]));
 BUFx2_ASAP7_75t_R _21574_ (.A(net678),
    .Y(out[446]));
 BUFx2_ASAP7_75t_R _21575_ (.A(net679),
    .Y(out[447]));
 BUFx2_ASAP7_75t_R _21576_ (.A(net680),
    .Y(out[448]));
 BUFx2_ASAP7_75t_R _21577_ (.A(net681),
    .Y(out[449]));
 BUFx3_ASAP7_75t_R _21578_ (.A(net185),
    .Y(net183));
 BUFx3_ASAP7_75t_R _21579_ (.A(net185),
    .Y(net184));
 BUFx2_ASAP7_75t_R _21580_ (.A(net682),
    .Y(out[452]));
 BUFx2_ASAP7_75t_R _21581_ (.A(net683),
    .Y(out[454]));
 BUFx2_ASAP7_75t_R _21582_ (.A(net684),
    .Y(out[455]));
 BUFx2_ASAP7_75t_R _21583_ (.A(net685),
    .Y(out[456]));
 BUFx2_ASAP7_75t_R _21584_ (.A(net686),
    .Y(out[457]));
 BUFx2_ASAP7_75t_R _21585_ (.A(net687),
    .Y(out[458]));
 BUFx2_ASAP7_75t_R _21586_ (.A(net688),
    .Y(out[459]));
 BUFx2_ASAP7_75t_R _21587_ (.A(net689),
    .Y(out[460]));
 BUFx2_ASAP7_75t_R _21588_ (.A(net690),
    .Y(out[461]));
 BUFx2_ASAP7_75t_R _21589_ (.A(net691),
    .Y(out[462]));
 BUFx2_ASAP7_75t_R _21590_ (.A(net692),
    .Y(out[463]));
 BUFx2_ASAP7_75t_R _21591_ (.A(net693),
    .Y(out[464]));
 BUFx2_ASAP7_75t_R _21592_ (.A(net694),
    .Y(out[465]));
 BUFx2_ASAP7_75t_R _21593_ (.A(net695),
    .Y(out[466]));
 BUFx2_ASAP7_75t_R _21594_ (.A(net696),
    .Y(out[467]));
 BUFx2_ASAP7_75t_R _21595_ (.A(net697),
    .Y(out[468]));
 BUFx2_ASAP7_75t_R _21596_ (.A(net698),
    .Y(out[469]));
 BUFx2_ASAP7_75t_R _21597_ (.A(net699),
    .Y(out[470]));
 BUFx2_ASAP7_75t_R _21598_ (.A(net700),
    .Y(out[471]));
 BUFx2_ASAP7_75t_R _21599_ (.A(net701),
    .Y(out[477]));
 BUFx2_ASAP7_75t_R _21600_ (.A(net702),
    .Y(out[478]));
 BUFx2_ASAP7_75t_R _21601_ (.A(net703),
    .Y(out[481]));
 BUFx2_ASAP7_75t_R _21602_ (.A(net704),
    .Y(out[482]));
 BUFx2_ASAP7_75t_R _21603_ (.A(net705),
    .Y(out[483]));
 BUFx2_ASAP7_75t_R _21604_ (.A(net706),
    .Y(out[484]));
 BUFx2_ASAP7_75t_R _21605_ (.A(net707),
    .Y(out[485]));
 BUFx2_ASAP7_75t_R _21606_ (.A(net708),
    .Y(out[486]));
 BUFx2_ASAP7_75t_R _21607_ (.A(net709),
    .Y(out[487]));
 BUFx2_ASAP7_75t_R _21608_ (.A(net710),
    .Y(out[488]));
 BUFx2_ASAP7_75t_R _21609_ (.A(net711),
    .Y(out[489]));
 BUFx2_ASAP7_75t_R _21610_ (.A(net712),
    .Y(out[490]));
 BUFx2_ASAP7_75t_R _21611_ (.A(net713),
    .Y(out[491]));
 BUFx3_ASAP7_75t_R _21612_ (.A(net194),
    .Y(net193));
 BUFx2_ASAP7_75t_R _21613_ (.A(net714),
    .Y(out[494]));
 BUFx2_ASAP7_75t_R _21614_ (.A(net715),
    .Y(out[495]));
 BUFx2_ASAP7_75t_R _21615_ (.A(net716),
    .Y(out[496]));
 BUFx2_ASAP7_75t_R _21616_ (.A(net717),
    .Y(out[497]));
 BUFx2_ASAP7_75t_R _21617_ (.A(net718),
    .Y(out[498]));
 BUFx2_ASAP7_75t_R _21618_ (.A(net719),
    .Y(out[499]));
 BUFx2_ASAP7_75t_R _21619_ (.A(net720),
    .Y(out[500]));
 BUFx2_ASAP7_75t_R _21620_ (.A(net721),
    .Y(out[501]));
 BUFx2_ASAP7_75t_R _21621_ (.A(net722),
    .Y(out[502]));
 BUFx2_ASAP7_75t_R _21622_ (.A(net723),
    .Y(out[503]));
 BUFx2_ASAP7_75t_R _21623_ (.A(net724),
    .Y(out[504]));
 BUFx2_ASAP7_75t_R _21624_ (.A(net725),
    .Y(out[505]));
 BUFx2_ASAP7_75t_R _21625_ (.A(net726),
    .Y(out[506]));
 BUFx2_ASAP7_75t_R _21626_ (.A(net727),
    .Y(out[507]));
 BUFx2_ASAP7_75t_R _21627_ (.A(net728),
    .Y(out[508]));
 BUFx2_ASAP7_75t_R _21628_ (.A(net729),
    .Y(out[509]));
 BUFx2_ASAP7_75t_R _21629_ (.A(net730),
    .Y(out[510]));
 BUFx2_ASAP7_75t_R _21630_ (.A(net731),
    .Y(out[511]));
 BUFx2_ASAP7_75t_R _21631_ (.A(net732),
    .Y(out[517]));
 BUFx2_ASAP7_75t_R _21632_ (.A(net733),
    .Y(out[518]));
 BUFx2_ASAP7_75t_R _21633_ (.A(net734),
    .Y(out[521]));
 BUFx2_ASAP7_75t_R _21634_ (.A(net735),
    .Y(out[522]));
 BUFx2_ASAP7_75t_R _21635_ (.A(net736),
    .Y(out[523]));
 BUFx2_ASAP7_75t_R _21636_ (.A(net737),
    .Y(out[524]));
 BUFx2_ASAP7_75t_R _21637_ (.A(net738),
    .Y(out[525]));
 BUFx2_ASAP7_75t_R _21638_ (.A(net739),
    .Y(out[526]));
 BUFx2_ASAP7_75t_R _21639_ (.A(net740),
    .Y(out[527]));
 BUFx2_ASAP7_75t_R _21640_ (.A(net741),
    .Y(out[528]));
 BUFx2_ASAP7_75t_R _21641_ (.A(net742),
    .Y(out[529]));
 BUFx3_ASAP7_75t_R _21642_ (.A(net205),
    .Y(net203));
 BUFx2_ASAP7_75t_R _21643_ (.A(net743),
    .Y(out[531]));
 BUFx3_ASAP7_75t_R _21644_ (.A(net205),
    .Y(net204));
 BUFx2_ASAP7_75t_R _21645_ (.A(net744),
    .Y(out[534]));
 BUFx2_ASAP7_75t_R _21646_ (.A(net745),
    .Y(out[535]));
 BUFx2_ASAP7_75t_R _21647_ (.A(net746),
    .Y(out[536]));
 BUFx2_ASAP7_75t_R _21648_ (.A(net747),
    .Y(out[537]));
 BUFx2_ASAP7_75t_R _21649_ (.A(net748),
    .Y(out[538]));
 BUFx2_ASAP7_75t_R _21650_ (.A(net749),
    .Y(out[539]));
 BUFx2_ASAP7_75t_R _21651_ (.A(net750),
    .Y(out[540]));
 BUFx2_ASAP7_75t_R _21652_ (.A(net751),
    .Y(out[541]));
 BUFx2_ASAP7_75t_R _21653_ (.A(net752),
    .Y(out[542]));
 BUFx2_ASAP7_75t_R _21654_ (.A(net753),
    .Y(out[543]));
 BUFx2_ASAP7_75t_R _21655_ (.A(net754),
    .Y(out[544]));
 BUFx2_ASAP7_75t_R _21656_ (.A(net755),
    .Y(out[545]));
 BUFx2_ASAP7_75t_R _21657_ (.A(net756),
    .Y(out[546]));
 BUFx2_ASAP7_75t_R _21658_ (.A(net757),
    .Y(out[547]));
 BUFx2_ASAP7_75t_R _21659_ (.A(net758),
    .Y(out[548]));
 BUFx2_ASAP7_75t_R _21660_ (.A(net759),
    .Y(out[549]));
 BUFx2_ASAP7_75t_R _21661_ (.A(net760),
    .Y(out[550]));
 BUFx2_ASAP7_75t_R _21662_ (.A(net761),
    .Y(out[551]));
 BUFx2_ASAP7_75t_R _21663_ (.A(net762),
    .Y(out[557]));
 BUFx2_ASAP7_75t_R _21664_ (.A(net763),
    .Y(out[558]));
 BUFx2_ASAP7_75t_R _21665_ (.A(net764),
    .Y(out[561]));
 BUFx2_ASAP7_75t_R _21666_ (.A(net765),
    .Y(out[562]));
 BUFx2_ASAP7_75t_R _21667_ (.A(net766),
    .Y(out[563]));
 BUFx2_ASAP7_75t_R _21668_ (.A(net767),
    .Y(out[564]));
 BUFx2_ASAP7_75t_R _21669_ (.A(net768),
    .Y(out[565]));
 BUFx2_ASAP7_75t_R _21670_ (.A(net769),
    .Y(out[566]));
 BUFx2_ASAP7_75t_R _21671_ (.A(net770),
    .Y(out[567]));
 BUFx2_ASAP7_75t_R _21672_ (.A(net771),
    .Y(out[568]));
 BUFx2_ASAP7_75t_R _21673_ (.A(net772),
    .Y(out[569]));
 BUFx2_ASAP7_75t_R _21674_ (.A(net773),
    .Y(out[570]));
 BUFx3_ASAP7_75t_R _21675_ (.A(net215),
    .Y(net213));
 BUFx3_ASAP7_75t_R _21676_ (.A(net215),
    .Y(net214));
 BUFx2_ASAP7_75t_R _21677_ (.A(net774),
    .Y(out[574]));
 BUFx2_ASAP7_75t_R _21678_ (.A(net775),
    .Y(out[575]));
 BUFx2_ASAP7_75t_R _21679_ (.A(net776),
    .Y(out[576]));
 BUFx2_ASAP7_75t_R _21680_ (.A(net777),
    .Y(out[577]));
 BUFx2_ASAP7_75t_R _21681_ (.A(net778),
    .Y(out[578]));
 BUFx2_ASAP7_75t_R _21682_ (.A(net779),
    .Y(out[579]));
 BUFx2_ASAP7_75t_R _21683_ (.A(net780),
    .Y(out[580]));
 BUFx2_ASAP7_75t_R _21684_ (.A(net781),
    .Y(out[581]));
 BUFx2_ASAP7_75t_R _21685_ (.A(net782),
    .Y(out[582]));
 BUFx2_ASAP7_75t_R _21686_ (.A(net783),
    .Y(out[583]));
 BUFx2_ASAP7_75t_R _21687_ (.A(net784),
    .Y(out[584]));
 BUFx2_ASAP7_75t_R _21688_ (.A(net785),
    .Y(out[585]));
 BUFx2_ASAP7_75t_R _21689_ (.A(net786),
    .Y(out[586]));
 BUFx2_ASAP7_75t_R _21690_ (.A(net787),
    .Y(out[587]));
 BUFx2_ASAP7_75t_R _21691_ (.A(net788),
    .Y(out[588]));
 BUFx2_ASAP7_75t_R _21692_ (.A(net789),
    .Y(out[589]));
 BUFx2_ASAP7_75t_R _21693_ (.A(net790),
    .Y(out[590]));
 BUFx2_ASAP7_75t_R _21694_ (.A(net791),
    .Y(out[591]));
 BUFx2_ASAP7_75t_R _21695_ (.A(net792),
    .Y(out[597]));
 BUFx2_ASAP7_75t_R _21696_ (.A(net793),
    .Y(out[598]));
 BUFx2_ASAP7_75t_R _21697_ (.A(net794),
    .Y(out[601]));
 BUFx2_ASAP7_75t_R _21698_ (.A(net795),
    .Y(out[602]));
 BUFx2_ASAP7_75t_R _21699_ (.A(net796),
    .Y(out[603]));
 BUFx2_ASAP7_75t_R _21700_ (.A(net797),
    .Y(out[604]));
 BUFx2_ASAP7_75t_R _21701_ (.A(net798),
    .Y(out[605]));
 BUFx2_ASAP7_75t_R _21702_ (.A(net799),
    .Y(out[606]));
 BUFx2_ASAP7_75t_R _21703_ (.A(net800),
    .Y(out[607]));
 BUFx2_ASAP7_75t_R _21704_ (.A(net801),
    .Y(out[608]));
 BUFx2_ASAP7_75t_R _21705_ (.A(net802),
    .Y(out[609]));
 BUFx3_ASAP7_75t_R _21706_ (.A(net226),
    .Y(net223));
 BUFx3_ASAP7_75t_R _21707_ (.A(net226),
    .Y(net224));
 BUFx3_ASAP7_75t_R _21708_ (.A(net226),
    .Y(net225));
 BUFx2_ASAP7_75t_R _21709_ (.A(net803),
    .Y(out[614]));
 BUFx2_ASAP7_75t_R _21710_ (.A(net804),
    .Y(out[615]));
 BUFx2_ASAP7_75t_R _21711_ (.A(net805),
    .Y(out[616]));
 BUFx2_ASAP7_75t_R _21712_ (.A(net806),
    .Y(out[617]));
 BUFx2_ASAP7_75t_R _21713_ (.A(net807),
    .Y(out[618]));
 BUFx2_ASAP7_75t_R _21714_ (.A(net808),
    .Y(out[619]));
 BUFx2_ASAP7_75t_R _21715_ (.A(net809),
    .Y(out[620]));
 BUFx2_ASAP7_75t_R _21716_ (.A(net810),
    .Y(out[621]));
 BUFx2_ASAP7_75t_R _21717_ (.A(net811),
    .Y(out[622]));
 BUFx2_ASAP7_75t_R _21718_ (.A(net812),
    .Y(out[623]));
 BUFx2_ASAP7_75t_R _21719_ (.A(net813),
    .Y(out[624]));
 BUFx2_ASAP7_75t_R _21720_ (.A(net814),
    .Y(out[625]));
 BUFx2_ASAP7_75t_R _21721_ (.A(net815),
    .Y(out[626]));
 BUFx2_ASAP7_75t_R _21722_ (.A(net816),
    .Y(out[627]));
 BUFx2_ASAP7_75t_R _21723_ (.A(net817),
    .Y(out[628]));
 BUFx2_ASAP7_75t_R _21724_ (.A(net818),
    .Y(out[629]));
 BUFx2_ASAP7_75t_R _21725_ (.A(net819),
    .Y(out[630]));
 BUFx2_ASAP7_75t_R _21726_ (.A(net820),
    .Y(out[631]));
 BUFx2_ASAP7_75t_R _21727_ (.A(net821),
    .Y(out[637]));
 BUFx2_ASAP7_75t_R _21728_ (.A(net822),
    .Y(out[638]));
 BUFx2_ASAP7_75t_R _21729_ (.A(net823),
    .Y(out[641]));
 BUFx2_ASAP7_75t_R _21730_ (.A(net824),
    .Y(out[642]));
 BUFx2_ASAP7_75t_R _21731_ (.A(net825),
    .Y(out[643]));
 BUFx2_ASAP7_75t_R _21732_ (.A(net826),
    .Y(out[644]));
 BUFx2_ASAP7_75t_R _21733_ (.A(net827),
    .Y(out[645]));
 BUFx2_ASAP7_75t_R _21734_ (.A(net828),
    .Y(out[646]));
 BUFx2_ASAP7_75t_R _21735_ (.A(net829),
    .Y(out[647]));
 BUFx2_ASAP7_75t_R _21736_ (.A(net830),
    .Y(out[648]));
 BUFx2_ASAP7_75t_R _21737_ (.A(net831),
    .Y(out[649]));
 BUFx2_ASAP7_75t_R _21738_ (.A(net832),
    .Y(out[650]));
 BUFx2_ASAP7_75t_R _21739_ (.A(net833),
    .Y(out[651]));
 BUFx2_ASAP7_75t_R _21740_ (.A(net834),
    .Y(out[652]));
 BUFx2_ASAP7_75t_R _21741_ (.A(net835),
    .Y(out[653]));
 BUFx2_ASAP7_75t_R _21742_ (.A(net836),
    .Y(out[655]));
 BUFx2_ASAP7_75t_R _21743_ (.A(net837),
    .Y(out[656]));
 BUFx2_ASAP7_75t_R _21744_ (.A(net838),
    .Y(out[657]));
 BUFx2_ASAP7_75t_R _21745_ (.A(net839),
    .Y(out[658]));
 BUFx2_ASAP7_75t_R _21746_ (.A(net840),
    .Y(out[659]));
 BUFx2_ASAP7_75t_R _21747_ (.A(net841),
    .Y(out[660]));
 BUFx2_ASAP7_75t_R _21748_ (.A(net842),
    .Y(out[661]));
 BUFx2_ASAP7_75t_R _21749_ (.A(net843),
    .Y(out[662]));
 BUFx2_ASAP7_75t_R _21750_ (.A(net844),
    .Y(out[663]));
 BUFx2_ASAP7_75t_R _21751_ (.A(net845),
    .Y(out[664]));
 BUFx2_ASAP7_75t_R _21752_ (.A(net846),
    .Y(out[665]));
 BUFx2_ASAP7_75t_R _21753_ (.A(net847),
    .Y(out[666]));
 BUFx2_ASAP7_75t_R _21754_ (.A(net848),
    .Y(out[667]));
 BUFx2_ASAP7_75t_R _21755_ (.A(net849),
    .Y(out[668]));
 BUFx2_ASAP7_75t_R _21756_ (.A(net850),
    .Y(out[669]));
 BUFx2_ASAP7_75t_R _21757_ (.A(net851),
    .Y(out[670]));
 BUFx2_ASAP7_75t_R _21758_ (.A(net852),
    .Y(out[671]));
 BUFx2_ASAP7_75t_R _21759_ (.A(net853),
    .Y(out[677]));
 BUFx2_ASAP7_75t_R _21760_ (.A(net854),
    .Y(out[678]));
 BUFx2_ASAP7_75t_R _21761_ (.A(net855),
    .Y(out[681]));
 BUFx2_ASAP7_75t_R _21762_ (.A(net856),
    .Y(out[682]));
 BUFx2_ASAP7_75t_R _21763_ (.A(net857),
    .Y(out[683]));
 BUFx2_ASAP7_75t_R _21764_ (.A(net858),
    .Y(out[684]));
 BUFx2_ASAP7_75t_R _21765_ (.A(net859),
    .Y(out[685]));
 BUFx2_ASAP7_75t_R _21766_ (.A(net860),
    .Y(out[686]));
 BUFx2_ASAP7_75t_R _21767_ (.A(net861),
    .Y(out[687]));
 BUFx2_ASAP7_75t_R _21768_ (.A(net862),
    .Y(out[688]));
 BUFx2_ASAP7_75t_R _21769_ (.A(net863),
    .Y(out[689]));
 BUFx3_ASAP7_75t_R _21770_ (.A(net243),
    .Y(net242));
 BUFx2_ASAP7_75t_R _21771_ (.A(net864),
    .Y(out[691]));
 BUFx2_ASAP7_75t_R _21772_ (.A(net865),
    .Y(out[692]));
 BUFx2_ASAP7_75t_R _21773_ (.A(net866),
    .Y(out[693]));
 BUFx2_ASAP7_75t_R _21774_ (.A(net867),
    .Y(out[695]));
 BUFx2_ASAP7_75t_R _21775_ (.A(net868),
    .Y(out[696]));
 BUFx2_ASAP7_75t_R _21776_ (.A(net869),
    .Y(out[697]));
 BUFx2_ASAP7_75t_R _21777_ (.A(net870),
    .Y(out[698]));
 BUFx2_ASAP7_75t_R _21778_ (.A(net871),
    .Y(out[699]));
 BUFx2_ASAP7_75t_R _21779_ (.A(net872),
    .Y(out[700]));
 BUFx2_ASAP7_75t_R _21780_ (.A(net873),
    .Y(out[701]));
 BUFx2_ASAP7_75t_R _21781_ (.A(net874),
    .Y(out[702]));
 BUFx2_ASAP7_75t_R _21782_ (.A(net875),
    .Y(out[703]));
 BUFx2_ASAP7_75t_R _21783_ (.A(net876),
    .Y(out[704]));
 BUFx2_ASAP7_75t_R _21784_ (.A(net877),
    .Y(out[705]));
 BUFx2_ASAP7_75t_R _21785_ (.A(net878),
    .Y(out[706]));
 BUFx2_ASAP7_75t_R _21786_ (.A(net879),
    .Y(out[707]));
 BUFx2_ASAP7_75t_R _21787_ (.A(net880),
    .Y(out[708]));
 BUFx2_ASAP7_75t_R _21788_ (.A(net881),
    .Y(out[709]));
 BUFx2_ASAP7_75t_R _21789_ (.A(net882),
    .Y(out[710]));
 BUFx2_ASAP7_75t_R _21790_ (.A(net883),
    .Y(out[711]));
 BUFx2_ASAP7_75t_R _21791_ (.A(net884),
    .Y(out[717]));
 BUFx2_ASAP7_75t_R _21792_ (.A(net885),
    .Y(out[718]));
 BUFx2_ASAP7_75t_R _21793_ (.A(net886),
    .Y(out[721]));
 BUFx2_ASAP7_75t_R _21794_ (.A(net887),
    .Y(out[722]));
 BUFx2_ASAP7_75t_R _21795_ (.A(net888),
    .Y(out[723]));
 BUFx2_ASAP7_75t_R _21796_ (.A(net889),
    .Y(out[724]));
 BUFx2_ASAP7_75t_R _21797_ (.A(net890),
    .Y(out[725]));
 BUFx2_ASAP7_75t_R _21798_ (.A(net891),
    .Y(out[726]));
 BUFx2_ASAP7_75t_R _21799_ (.A(net892),
    .Y(out[727]));
 BUFx2_ASAP7_75t_R _21800_ (.A(net893),
    .Y(out[728]));
 BUFx2_ASAP7_75t_R _21801_ (.A(net894),
    .Y(out[729]));
 BUFx2_ASAP7_75t_R _21802_ (.A(net895),
    .Y(out[730]));
 BUFx3_ASAP7_75t_R _21803_ (.A(net253),
    .Y(net252));
 BUFx2_ASAP7_75t_R _21804_ (.A(net896),
    .Y(out[732]));
 BUFx2_ASAP7_75t_R _21805_ (.A(net897),
    .Y(out[733]));
 BUFx2_ASAP7_75t_R _21806_ (.A(net898),
    .Y(out[735]));
 BUFx2_ASAP7_75t_R _21807_ (.A(net899),
    .Y(out[736]));
 BUFx2_ASAP7_75t_R _21808_ (.A(net900),
    .Y(out[737]));
 BUFx2_ASAP7_75t_R _21809_ (.A(net901),
    .Y(out[738]));
 BUFx2_ASAP7_75t_R _21810_ (.A(net902),
    .Y(out[739]));
 BUFx2_ASAP7_75t_R _21811_ (.A(net903),
    .Y(out[740]));
 BUFx2_ASAP7_75t_R _21812_ (.A(net904),
    .Y(out[741]));
 BUFx2_ASAP7_75t_R _21813_ (.A(net905),
    .Y(out[742]));
 BUFx2_ASAP7_75t_R _21814_ (.A(net906),
    .Y(out[743]));
 BUFx2_ASAP7_75t_R _21815_ (.A(net907),
    .Y(out[744]));
 BUFx2_ASAP7_75t_R _21816_ (.A(net908),
    .Y(out[745]));
 BUFx2_ASAP7_75t_R _21817_ (.A(net909),
    .Y(out[746]));
 BUFx2_ASAP7_75t_R _21818_ (.A(net910),
    .Y(out[747]));
 BUFx2_ASAP7_75t_R _21819_ (.A(net911),
    .Y(out[748]));
 BUFx2_ASAP7_75t_R _21820_ (.A(net912),
    .Y(out[749]));
 BUFx2_ASAP7_75t_R _21821_ (.A(net913),
    .Y(out[750]));
 BUFx2_ASAP7_75t_R _21822_ (.A(net914),
    .Y(out[751]));
 BUFx2_ASAP7_75t_R _21823_ (.A(net915),
    .Y(out[757]));
 BUFx2_ASAP7_75t_R _21824_ (.A(net916),
    .Y(out[758]));
 BUFx2_ASAP7_75t_R _21825_ (.A(net917),
    .Y(out[761]));
 BUFx2_ASAP7_75t_R _21826_ (.A(net918),
    .Y(out[762]));
 BUFx2_ASAP7_75t_R _21827_ (.A(net919),
    .Y(out[763]));
 BUFx2_ASAP7_75t_R _21828_ (.A(net920),
    .Y(out[764]));
 BUFx2_ASAP7_75t_R _21829_ (.A(net921),
    .Y(out[765]));
 BUFx2_ASAP7_75t_R _21830_ (.A(net922),
    .Y(out[766]));
 BUFx2_ASAP7_75t_R _21831_ (.A(net923),
    .Y(out[767]));
 BUFx2_ASAP7_75t_R _21832_ (.A(net924),
    .Y(out[768]));
 BUFx2_ASAP7_75t_R _21833_ (.A(net925),
    .Y(out[769]));
 BUFx3_ASAP7_75t_R _21834_ (.A(net267),
    .Y(net265));
 BUFx3_ASAP7_75t_R _21835_ (.A(net267),
    .Y(net266));
 BUFx2_ASAP7_75t_R _21836_ (.A(net926),
    .Y(out[772]));
 BUFx2_ASAP7_75t_R _21837_ (.A(net927),
    .Y(out[773]));
 BUFx2_ASAP7_75t_R _21838_ (.A(net928),
    .Y(out[775]));
 BUFx2_ASAP7_75t_R _21839_ (.A(net929),
    .Y(out[776]));
 BUFx2_ASAP7_75t_R _21840_ (.A(net930),
    .Y(out[777]));
 BUFx2_ASAP7_75t_R _21841_ (.A(net931),
    .Y(out[778]));
 BUFx2_ASAP7_75t_R _21842_ (.A(net932),
    .Y(out[779]));
 BUFx2_ASAP7_75t_R _21843_ (.A(net933),
    .Y(out[780]));
 BUFx2_ASAP7_75t_R _21844_ (.A(net934),
    .Y(out[781]));
 BUFx2_ASAP7_75t_R _21845_ (.A(net935),
    .Y(out[782]));
 BUFx2_ASAP7_75t_R _21846_ (.A(net936),
    .Y(out[783]));
 BUFx2_ASAP7_75t_R _21847_ (.A(net937),
    .Y(out[784]));
 BUFx2_ASAP7_75t_R _21848_ (.A(net938),
    .Y(out[785]));
 BUFx2_ASAP7_75t_R _21849_ (.A(net939),
    .Y(out[786]));
 BUFx2_ASAP7_75t_R _21850_ (.A(net940),
    .Y(out[787]));
 BUFx2_ASAP7_75t_R _21851_ (.A(net941),
    .Y(out[788]));
 BUFx2_ASAP7_75t_R _21852_ (.A(net942),
    .Y(out[789]));
 BUFx2_ASAP7_75t_R _21853_ (.A(net943),
    .Y(out[790]));
 BUFx2_ASAP7_75t_R _21854_ (.A(net944),
    .Y(out[791]));
 BUFx2_ASAP7_75t_R _21855_ (.A(net945),
    .Y(out[797]));
 BUFx2_ASAP7_75t_R _21856_ (.A(net946),
    .Y(out[798]));
 BUFx2_ASAP7_75t_R _21857_ (.A(net947),
    .Y(out[801]));
 BUFx2_ASAP7_75t_R _21858_ (.A(net948),
    .Y(out[802]));
 BUFx2_ASAP7_75t_R _21859_ (.A(net949),
    .Y(out[803]));
 BUFx2_ASAP7_75t_R _21860_ (.A(net950),
    .Y(out[804]));
 BUFx2_ASAP7_75t_R _21861_ (.A(net951),
    .Y(out[805]));
 BUFx2_ASAP7_75t_R _21862_ (.A(net952),
    .Y(out[806]));
 BUFx2_ASAP7_75t_R _21863_ (.A(net953),
    .Y(out[807]));
 BUFx2_ASAP7_75t_R _21864_ (.A(net954),
    .Y(out[808]));
 BUFx2_ASAP7_75t_R _21865_ (.A(net955),
    .Y(out[809]));
 BUFx2_ASAP7_75t_R _21866_ (.A(net956),
    .Y(out[810]));
 BUFx2_ASAP7_75t_R _21867_ (.A(net957),
    .Y(out[811]));
 BUFx3_ASAP7_75t_R _21868_ (.A(net278),
    .Y(net277));
 BUFx2_ASAP7_75t_R _21869_ (.A(net958),
    .Y(out[813]));
 BUFx2_ASAP7_75t_R _21870_ (.A(net959),
    .Y(out[815]));
 BUFx2_ASAP7_75t_R _21871_ (.A(net960),
    .Y(out[816]));
 BUFx2_ASAP7_75t_R _21872_ (.A(net961),
    .Y(out[817]));
 BUFx2_ASAP7_75t_R _21873_ (.A(net962),
    .Y(out[818]));
 BUFx2_ASAP7_75t_R _21874_ (.A(net963),
    .Y(out[819]));
 BUFx2_ASAP7_75t_R _21875_ (.A(net964),
    .Y(out[820]));
 BUFx2_ASAP7_75t_R _21876_ (.A(net965),
    .Y(out[821]));
 BUFx2_ASAP7_75t_R _21877_ (.A(net966),
    .Y(out[822]));
 BUFx2_ASAP7_75t_R _21878_ (.A(net967),
    .Y(out[823]));
 BUFx2_ASAP7_75t_R _21879_ (.A(net968),
    .Y(out[824]));
 BUFx2_ASAP7_75t_R _21880_ (.A(net969),
    .Y(out[825]));
 BUFx2_ASAP7_75t_R _21881_ (.A(net970),
    .Y(out[826]));
 BUFx2_ASAP7_75t_R _21882_ (.A(net971),
    .Y(out[827]));
 BUFx2_ASAP7_75t_R _21883_ (.A(net972),
    .Y(out[828]));
 BUFx2_ASAP7_75t_R _21884_ (.A(net973),
    .Y(out[829]));
 BUFx2_ASAP7_75t_R _21885_ (.A(net974),
    .Y(out[830]));
 BUFx2_ASAP7_75t_R _21886_ (.A(net975),
    .Y(out[831]));
 BUFx2_ASAP7_75t_R _21887_ (.A(net976),
    .Y(out[837]));
 BUFx2_ASAP7_75t_R _21888_ (.A(net977),
    .Y(out[838]));
 BUFx2_ASAP7_75t_R _21889_ (.A(net978),
    .Y(out[841]));
 BUFx2_ASAP7_75t_R _21890_ (.A(net979),
    .Y(out[842]));
 BUFx2_ASAP7_75t_R _21891_ (.A(net980),
    .Y(out[843]));
 BUFx2_ASAP7_75t_R _21892_ (.A(net981),
    .Y(out[844]));
 BUFx2_ASAP7_75t_R _21893_ (.A(net982),
    .Y(out[845]));
 BUFx2_ASAP7_75t_R _21894_ (.A(net983),
    .Y(out[846]));
 BUFx2_ASAP7_75t_R _21895_ (.A(net984),
    .Y(out[847]));
 BUFx2_ASAP7_75t_R _21896_ (.A(net985),
    .Y(out[848]));
 BUFx2_ASAP7_75t_R _21897_ (.A(net986),
    .Y(out[849]));
 BUFx3_ASAP7_75t_R _21898_ (.A(net288),
    .Y(net286));
 BUFx2_ASAP7_75t_R _21899_ (.A(net987),
    .Y(out[851]));
 BUFx3_ASAP7_75t_R _21900_ (.A(net288),
    .Y(net287));
 BUFx2_ASAP7_75t_R _21901_ (.A(net988),
    .Y(out[853]));
 BUFx2_ASAP7_75t_R _21902_ (.A(net989),
    .Y(out[855]));
 BUFx2_ASAP7_75t_R _21903_ (.A(net990),
    .Y(out[856]));
 BUFx2_ASAP7_75t_R _21904_ (.A(net991),
    .Y(out[857]));
 BUFx2_ASAP7_75t_R _21905_ (.A(net992),
    .Y(out[858]));
 BUFx2_ASAP7_75t_R _21906_ (.A(net993),
    .Y(out[859]));
 BUFx2_ASAP7_75t_R _21907_ (.A(net994),
    .Y(out[860]));
 BUFx2_ASAP7_75t_R _21908_ (.A(net995),
    .Y(out[861]));
 BUFx2_ASAP7_75t_R _21909_ (.A(net996),
    .Y(out[862]));
 BUFx2_ASAP7_75t_R _21910_ (.A(net997),
    .Y(out[863]));
 BUFx2_ASAP7_75t_R _21911_ (.A(net998),
    .Y(out[864]));
 BUFx2_ASAP7_75t_R _21912_ (.A(net999),
    .Y(out[865]));
 BUFx2_ASAP7_75t_R _21913_ (.A(net1000),
    .Y(out[866]));
 BUFx2_ASAP7_75t_R _21914_ (.A(net1001),
    .Y(out[867]));
 BUFx2_ASAP7_75t_R _21915_ (.A(net1002),
    .Y(out[868]));
 BUFx2_ASAP7_75t_R _21916_ (.A(net1003),
    .Y(out[869]));
 BUFx2_ASAP7_75t_R _21917_ (.A(net1004),
    .Y(out[870]));
 BUFx2_ASAP7_75t_R _21918_ (.A(net1005),
    .Y(out[871]));
 BUFx2_ASAP7_75t_R _21919_ (.A(net1006),
    .Y(out[877]));
 BUFx2_ASAP7_75t_R _21920_ (.A(net1007),
    .Y(out[878]));
 BUFx2_ASAP7_75t_R _21921_ (.A(net1008),
    .Y(out[881]));
 BUFx2_ASAP7_75t_R _21922_ (.A(net1009),
    .Y(out[882]));
 BUFx2_ASAP7_75t_R _21923_ (.A(net1010),
    .Y(out[883]));
 BUFx2_ASAP7_75t_R _21924_ (.A(net1011),
    .Y(out[884]));
 BUFx2_ASAP7_75t_R _21925_ (.A(net1012),
    .Y(out[885]));
 BUFx2_ASAP7_75t_R _21926_ (.A(net1013),
    .Y(out[886]));
 BUFx2_ASAP7_75t_R _21927_ (.A(net1014),
    .Y(out[887]));
 BUFx2_ASAP7_75t_R _21928_ (.A(net1015),
    .Y(out[888]));
 BUFx2_ASAP7_75t_R _21929_ (.A(net1016),
    .Y(out[889]));
 BUFx2_ASAP7_75t_R _21930_ (.A(net1017),
    .Y(out[890]));
 BUFx3_ASAP7_75t_R _21931_ (.A(net298),
    .Y(net296));
 BUFx3_ASAP7_75t_R _21932_ (.A(net298),
    .Y(net297));
 BUFx2_ASAP7_75t_R _21933_ (.A(net1018),
    .Y(out[893]));
 BUFx2_ASAP7_75t_R _21934_ (.A(net1019),
    .Y(out[895]));
 BUFx2_ASAP7_75t_R _21935_ (.A(net1020),
    .Y(out[896]));
 BUFx2_ASAP7_75t_R _21936_ (.A(net1021),
    .Y(out[897]));
 BUFx2_ASAP7_75t_R _21937_ (.A(net1022),
    .Y(out[898]));
 BUFx2_ASAP7_75t_R _21938_ (.A(net1023),
    .Y(out[899]));
 BUFx2_ASAP7_75t_R _21939_ (.A(net1024),
    .Y(out[900]));
 BUFx2_ASAP7_75t_R _21940_ (.A(net1025),
    .Y(out[901]));
 BUFx2_ASAP7_75t_R _21941_ (.A(net1026),
    .Y(out[902]));
 BUFx2_ASAP7_75t_R _21942_ (.A(net1027),
    .Y(out[903]));
 BUFx2_ASAP7_75t_R _21943_ (.A(net1028),
    .Y(out[904]));
 BUFx2_ASAP7_75t_R _21944_ (.A(net1029),
    .Y(out[905]));
 BUFx2_ASAP7_75t_R _21945_ (.A(net1030),
    .Y(out[906]));
 BUFx2_ASAP7_75t_R _21946_ (.A(net1031),
    .Y(out[907]));
 BUFx2_ASAP7_75t_R _21947_ (.A(net1032),
    .Y(out[908]));
 BUFx2_ASAP7_75t_R _21948_ (.A(net1033),
    .Y(out[909]));
 BUFx2_ASAP7_75t_R _21949_ (.A(net1034),
    .Y(out[910]));
 BUFx2_ASAP7_75t_R _21950_ (.A(net1035),
    .Y(out[911]));
 BUFx2_ASAP7_75t_R _21951_ (.A(net1036),
    .Y(out[917]));
 BUFx2_ASAP7_75t_R _21952_ (.A(net1037),
    .Y(out[918]));
 BUFx2_ASAP7_75t_R _21953_ (.A(net1038),
    .Y(out[921]));
 BUFx2_ASAP7_75t_R _21954_ (.A(net1039),
    .Y(out[922]));
 BUFx2_ASAP7_75t_R _21955_ (.A(net1040),
    .Y(out[923]));
 BUFx2_ASAP7_75t_R _21956_ (.A(net1041),
    .Y(out[924]));
 BUFx2_ASAP7_75t_R _21957_ (.A(net1042),
    .Y(out[925]));
 BUFx2_ASAP7_75t_R _21958_ (.A(net1043),
    .Y(out[926]));
 BUFx2_ASAP7_75t_R _21959_ (.A(net1044),
    .Y(out[927]));
 BUFx2_ASAP7_75t_R _21960_ (.A(net1045),
    .Y(out[928]));
 BUFx2_ASAP7_75t_R _21961_ (.A(net1046),
    .Y(out[929]));
 BUFx3_ASAP7_75t_R _21962_ (.A(net310),
    .Y(net307));
 BUFx3_ASAP7_75t_R _21963_ (.A(net310),
    .Y(net308));
 BUFx3_ASAP7_75t_R _21964_ (.A(net310),
    .Y(net309));
 BUFx2_ASAP7_75t_R _21965_ (.A(net1047),
    .Y(out[933]));
 BUFx2_ASAP7_75t_R _21966_ (.A(net1048),
    .Y(out[935]));
 BUFx2_ASAP7_75t_R _21967_ (.A(net1049),
    .Y(out[936]));
 BUFx2_ASAP7_75t_R _21968_ (.A(net1050),
    .Y(out[937]));
 BUFx2_ASAP7_75t_R _21969_ (.A(net1051),
    .Y(out[938]));
 BUFx2_ASAP7_75t_R _21970_ (.A(net1052),
    .Y(out[939]));
 BUFx2_ASAP7_75t_R _21971_ (.A(net1053),
    .Y(out[940]));
 BUFx2_ASAP7_75t_R _21972_ (.A(net1054),
    .Y(out[941]));
 BUFx2_ASAP7_75t_R _21973_ (.A(net1055),
    .Y(out[942]));
 BUFx2_ASAP7_75t_R _21974_ (.A(net1056),
    .Y(out[943]));
 BUFx2_ASAP7_75t_R _21975_ (.A(net1057),
    .Y(out[944]));
 BUFx2_ASAP7_75t_R _21976_ (.A(net1058),
    .Y(out[945]));
 BUFx2_ASAP7_75t_R _21977_ (.A(net1059),
    .Y(out[946]));
 BUFx2_ASAP7_75t_R _21978_ (.A(net1060),
    .Y(out[947]));
 BUFx2_ASAP7_75t_R _21979_ (.A(net1061),
    .Y(out[948]));
 BUFx2_ASAP7_75t_R _21980_ (.A(net1062),
    .Y(out[949]));
 BUFx2_ASAP7_75t_R _21981_ (.A(net1063),
    .Y(out[950]));
 BUFx2_ASAP7_75t_R _21982_ (.A(net1064),
    .Y(out[951]));
 BUFx2_ASAP7_75t_R _21983_ (.A(net1065),
    .Y(out[957]));
 BUFx2_ASAP7_75t_R _21984_ (.A(net1066),
    .Y(out[958]));
 BUFx2_ASAP7_75t_R _21985_ (.A(net1067),
    .Y(out[961]));
 BUFx2_ASAP7_75t_R _21986_ (.A(net1068),
    .Y(out[962]));
 BUFx2_ASAP7_75t_R _21987_ (.A(net1069),
    .Y(out[963]));
 BUFx2_ASAP7_75t_R _21988_ (.A(net1070),
    .Y(out[964]));
 BUFx2_ASAP7_75t_R _21989_ (.A(net1071),
    .Y(out[965]));
 BUFx2_ASAP7_75t_R _21990_ (.A(net1072),
    .Y(out[966]));
 BUFx2_ASAP7_75t_R _21991_ (.A(net1073),
    .Y(out[967]));
 BUFx2_ASAP7_75t_R _21992_ (.A(net1074),
    .Y(out[968]));
 BUFx2_ASAP7_75t_R _21993_ (.A(net1075),
    .Y(out[969]));
 BUFx2_ASAP7_75t_R _21994_ (.A(net1076),
    .Y(out[970]));
 BUFx2_ASAP7_75t_R _21995_ (.A(net1077),
    .Y(out[971]));
 BUFx2_ASAP7_75t_R _21996_ (.A(net1078),
    .Y(out[972]));
 BUFx3_ASAP7_75t_R _21997_ (.A(net319),
    .Y(net318));
 BUFx2_ASAP7_75t_R _21998_ (.A(net1079),
    .Y(out[975]));
 BUFx2_ASAP7_75t_R _21999_ (.A(net1080),
    .Y(out[976]));
 BUFx2_ASAP7_75t_R _22000_ (.A(net1081),
    .Y(out[977]));
 BUFx2_ASAP7_75t_R _22001_ (.A(net1082),
    .Y(out[978]));
 BUFx2_ASAP7_75t_R _22002_ (.A(net1083),
    .Y(out[979]));
 BUFx2_ASAP7_75t_R _22003_ (.A(net1084),
    .Y(out[980]));
 BUFx2_ASAP7_75t_R _22004_ (.A(net1085),
    .Y(out[981]));
 BUFx2_ASAP7_75t_R _22005_ (.A(net1086),
    .Y(out[982]));
 BUFx2_ASAP7_75t_R _22006_ (.A(net1087),
    .Y(out[983]));
 BUFx2_ASAP7_75t_R _22007_ (.A(net1088),
    .Y(out[984]));
 BUFx2_ASAP7_75t_R _22008_ (.A(net1089),
    .Y(out[985]));
 BUFx2_ASAP7_75t_R _22009_ (.A(net1090),
    .Y(out[986]));
 BUFx2_ASAP7_75t_R _22010_ (.A(net1091),
    .Y(out[987]));
 BUFx2_ASAP7_75t_R _22011_ (.A(net1092),
    .Y(out[988]));
 BUFx2_ASAP7_75t_R _22012_ (.A(net1093),
    .Y(out[989]));
 BUFx2_ASAP7_75t_R _22013_ (.A(net1094),
    .Y(out[990]));
 BUFx2_ASAP7_75t_R _22014_ (.A(net1095),
    .Y(out[991]));
 BUFx2_ASAP7_75t_R _22015_ (.A(net1096),
    .Y(out[997]));
 BUFx2_ASAP7_75t_R _22016_ (.A(net1097),
    .Y(out[998]));
 BUFx2_ASAP7_75t_R _22017_ (.A(net1098),
    .Y(out[1001]));
 BUFx2_ASAP7_75t_R _22018_ (.A(net1099),
    .Y(out[1002]));
 BUFx2_ASAP7_75t_R _22019_ (.A(net1100),
    .Y(out[1003]));
 BUFx2_ASAP7_75t_R _22020_ (.A(net1101),
    .Y(out[1004]));
 BUFx2_ASAP7_75t_R _22021_ (.A(net1102),
    .Y(out[1005]));
 BUFx2_ASAP7_75t_R _22022_ (.A(net1103),
    .Y(out[1006]));
 BUFx2_ASAP7_75t_R _22023_ (.A(net1104),
    .Y(out[1007]));
 BUFx2_ASAP7_75t_R _22024_ (.A(net1105),
    .Y(out[1008]));
 BUFx2_ASAP7_75t_R _22025_ (.A(net1106),
    .Y(out[1009]));
 BUFx3_ASAP7_75t_R _22026_ (.A(net26),
    .Y(net24));
 BUFx2_ASAP7_75t_R _22027_ (.A(net1107),
    .Y(out[1011]));
 BUFx2_ASAP7_75t_R _22028_ (.A(net1108),
    .Y(out[1012]));
 BUFx3_ASAP7_75t_R _22029_ (.A(net26),
    .Y(net25));
 BUFx2_ASAP7_75t_R _22030_ (.A(net1109),
    .Y(out[1015]));
 BUFx2_ASAP7_75t_R _22031_ (.A(net1110),
    .Y(out[1016]));
 BUFx2_ASAP7_75t_R _22032_ (.A(net1111),
    .Y(out[1017]));
 BUFx2_ASAP7_75t_R _22033_ (.A(net1112),
    .Y(out[1018]));
 BUFx2_ASAP7_75t_R _22034_ (.A(net1113),
    .Y(out[1019]));
 BUFx2_ASAP7_75t_R _22035_ (.A(net1114),
    .Y(out[1020]));
 BUFx2_ASAP7_75t_R _22036_ (.A(net1115),
    .Y(out[1021]));
 BUFx2_ASAP7_75t_R _22037_ (.A(net1116),
    .Y(out[1022]));
 BUFx2_ASAP7_75t_R _22038_ (.A(net1117),
    .Y(out[1023]));
 BUFx2_ASAP7_75t_R _22039_ (.A(net1118),
    .Y(out[1024]));
 BUFx2_ASAP7_75t_R _22040_ (.A(net1119),
    .Y(out[1025]));
 BUFx2_ASAP7_75t_R _22041_ (.A(net1120),
    .Y(out[1026]));
 BUFx2_ASAP7_75t_R _22042_ (.A(net1121),
    .Y(out[1027]));
 BUFx2_ASAP7_75t_R _22043_ (.A(net1122),
    .Y(out[1028]));
 BUFx2_ASAP7_75t_R _22044_ (.A(net1123),
    .Y(out[1029]));
 BUFx2_ASAP7_75t_R _22045_ (.A(net1124),
    .Y(out[1030]));
 BUFx2_ASAP7_75t_R _22046_ (.A(net1125),
    .Y(out[1031]));
 BUFx2_ASAP7_75t_R _22047_ (.A(net1126),
    .Y(out[1037]));
 BUFx2_ASAP7_75t_R _22048_ (.A(net1127),
    .Y(out[1038]));
 BUFx2_ASAP7_75t_R _22049_ (.A(net1128),
    .Y(out[1041]));
 BUFx2_ASAP7_75t_R _22050_ (.A(net1129),
    .Y(out[1042]));
 BUFx2_ASAP7_75t_R _22051_ (.A(net1130),
    .Y(out[1043]));
 BUFx2_ASAP7_75t_R _22052_ (.A(net1131),
    .Y(out[1044]));
 BUFx2_ASAP7_75t_R _22053_ (.A(net1132),
    .Y(out[1045]));
 BUFx2_ASAP7_75t_R _22054_ (.A(net1133),
    .Y(out[1046]));
 BUFx2_ASAP7_75t_R _22055_ (.A(net1134),
    .Y(out[1047]));
 BUFx2_ASAP7_75t_R _22056_ (.A(net1135),
    .Y(out[1048]));
 BUFx2_ASAP7_75t_R _22057_ (.A(net1136),
    .Y(out[1049]));
 BUFx2_ASAP7_75t_R _22058_ (.A(net1137),
    .Y(out[1050]));
 BUFx3_ASAP7_75t_R _22059_ (.A(net36),
    .Y(net34));
 BUFx2_ASAP7_75t_R _22060_ (.A(net1138),
    .Y(out[1052]));
 BUFx3_ASAP7_75t_R _22061_ (.A(net36),
    .Y(net35));
 BUFx2_ASAP7_75t_R _22062_ (.A(net1139),
    .Y(out[1055]));
 BUFx2_ASAP7_75t_R _22063_ (.A(net1140),
    .Y(out[1056]));
 BUFx2_ASAP7_75t_R _22064_ (.A(net1141),
    .Y(out[1057]));
 BUFx2_ASAP7_75t_R _22065_ (.A(net1142),
    .Y(out[1058]));
 BUFx2_ASAP7_75t_R _22066_ (.A(net1143),
    .Y(out[1059]));
 BUFx2_ASAP7_75t_R _22067_ (.A(net1144),
    .Y(out[1060]));
 BUFx2_ASAP7_75t_R _22068_ (.A(net1145),
    .Y(out[1061]));
 BUFx2_ASAP7_75t_R _22069_ (.A(net1146),
    .Y(out[1062]));
 BUFx2_ASAP7_75t_R _22070_ (.A(net1147),
    .Y(out[1063]));
 BUFx2_ASAP7_75t_R _22071_ (.A(net1148),
    .Y(out[1064]));
 BUFx2_ASAP7_75t_R _22072_ (.A(net1149),
    .Y(out[1065]));
 BUFx2_ASAP7_75t_R _22073_ (.A(net1150),
    .Y(out[1066]));
 BUFx2_ASAP7_75t_R _22074_ (.A(net1151),
    .Y(out[1067]));
 BUFx2_ASAP7_75t_R _22075_ (.A(net1152),
    .Y(out[1068]));
 BUFx2_ASAP7_75t_R _22076_ (.A(net1153),
    .Y(out[1069]));
 BUFx2_ASAP7_75t_R _22077_ (.A(net1154),
    .Y(out[1070]));
 BUFx2_ASAP7_75t_R _22078_ (.A(net1155),
    .Y(out[1071]));
 BUFx2_ASAP7_75t_R _22079_ (.A(net1156),
    .Y(out[1077]));
 BUFx2_ASAP7_75t_R _22080_ (.A(net1157),
    .Y(out[1078]));
 BUFx2_ASAP7_75t_R _22081_ (.A(net1158),
    .Y(out[1081]));
 BUFx2_ASAP7_75t_R _22082_ (.A(net1159),
    .Y(out[1082]));
 BUFx2_ASAP7_75t_R _22083_ (.A(net1160),
    .Y(out[1083]));
 BUFx2_ASAP7_75t_R _22084_ (.A(net1161),
    .Y(out[1084]));
 BUFx2_ASAP7_75t_R _22085_ (.A(net1162),
    .Y(out[1085]));
 BUFx2_ASAP7_75t_R _22086_ (.A(net1163),
    .Y(out[1086]));
 BUFx2_ASAP7_75t_R _22087_ (.A(net1164),
    .Y(out[1087]));
 BUFx2_ASAP7_75t_R _22088_ (.A(net1165),
    .Y(out[1088]));
 BUFx2_ASAP7_75t_R _22089_ (.A(net1166),
    .Y(out[1089]));
 BUFx3_ASAP7_75t_R _22090_ (.A(net47),
    .Y(net44));
 BUFx3_ASAP7_75t_R _22091_ (.A(net47),
    .Y(net45));
 BUFx2_ASAP7_75t_R _22092_ (.A(net1167),
    .Y(out[1092]));
 BUFx3_ASAP7_75t_R _22093_ (.A(net47),
    .Y(net46));
 BUFx2_ASAP7_75t_R _22094_ (.A(net1168),
    .Y(out[1095]));
 BUFx2_ASAP7_75t_R _22095_ (.A(net1169),
    .Y(out[1096]));
 BUFx2_ASAP7_75t_R _22096_ (.A(net1170),
    .Y(out[1097]));
 BUFx2_ASAP7_75t_R _22097_ (.A(net1171),
    .Y(out[1098]));
 BUFx2_ASAP7_75t_R _22098_ (.A(net1172),
    .Y(out[1099]));
 BUFx2_ASAP7_75t_R _22099_ (.A(net1173),
    .Y(out[1100]));
 BUFx2_ASAP7_75t_R _22100_ (.A(net1174),
    .Y(out[1101]));
 BUFx2_ASAP7_75t_R _22101_ (.A(net1175),
    .Y(out[1102]));
 BUFx2_ASAP7_75t_R _22102_ (.A(net1176),
    .Y(out[1103]));
 BUFx2_ASAP7_75t_R _22103_ (.A(net1177),
    .Y(out[1104]));
 BUFx2_ASAP7_75t_R _22104_ (.A(net1178),
    .Y(out[1105]));
 BUFx2_ASAP7_75t_R _22105_ (.A(net1179),
    .Y(out[1106]));
 BUFx2_ASAP7_75t_R _22106_ (.A(net1180),
    .Y(out[1107]));
 BUFx2_ASAP7_75t_R _22107_ (.A(net1181),
    .Y(out[1108]));
 BUFx2_ASAP7_75t_R _22108_ (.A(net1182),
    .Y(out[1109]));
 BUFx2_ASAP7_75t_R _22109_ (.A(net1183),
    .Y(out[1110]));
 BUFx2_ASAP7_75t_R _22110_ (.A(net1184),
    .Y(out[1111]));
 BUFx2_ASAP7_75t_R _22111_ (.A(net1185),
    .Y(out[1117]));
 BUFx2_ASAP7_75t_R _22112_ (.A(net1186),
    .Y(out[1118]));
 BUFx2_ASAP7_75t_R _22113_ (.A(net1187),
    .Y(out[1121]));
 BUFx2_ASAP7_75t_R _22114_ (.A(net1188),
    .Y(out[1122]));
 BUFx2_ASAP7_75t_R _22115_ (.A(net1189),
    .Y(out[1123]));
 BUFx2_ASAP7_75t_R _22116_ (.A(net1190),
    .Y(out[1124]));
 BUFx2_ASAP7_75t_R _22117_ (.A(net1191),
    .Y(out[1125]));
 BUFx2_ASAP7_75t_R _22118_ (.A(net1192),
    .Y(out[1126]));
 BUFx2_ASAP7_75t_R _22119_ (.A(net1193),
    .Y(out[1127]));
 BUFx2_ASAP7_75t_R _22120_ (.A(net1194),
    .Y(out[1128]));
 BUFx2_ASAP7_75t_R _22121_ (.A(net1195),
    .Y(out[1129]));
 BUFx2_ASAP7_75t_R _22122_ (.A(net1196),
    .Y(out[1130]));
 BUFx2_ASAP7_75t_R _22123_ (.A(net1197),
    .Y(out[1131]));
 BUFx3_ASAP7_75t_R _22124_ (.A(net58),
    .Y(net56));
 BUFx3_ASAP7_75t_R _22125_ (.A(net58),
    .Y(net57));
 BUFx2_ASAP7_75t_R _22126_ (.A(net1198),
    .Y(out[1135]));
 BUFx2_ASAP7_75t_R _22127_ (.A(net1199),
    .Y(out[1136]));
 BUFx2_ASAP7_75t_R _22128_ (.A(net1200),
    .Y(out[1137]));
 BUFx2_ASAP7_75t_R _22129_ (.A(net1201),
    .Y(out[1138]));
 BUFx2_ASAP7_75t_R _22130_ (.A(net1202),
    .Y(out[1139]));
 BUFx2_ASAP7_75t_R _22131_ (.A(net1203),
    .Y(out[1140]));
 BUFx2_ASAP7_75t_R _22132_ (.A(net1204),
    .Y(out[1141]));
 BUFx2_ASAP7_75t_R _22133_ (.A(net1205),
    .Y(out[1142]));
 BUFx2_ASAP7_75t_R _22134_ (.A(net1206),
    .Y(out[1143]));
 BUFx2_ASAP7_75t_R _22135_ (.A(net1207),
    .Y(out[1144]));
 BUFx2_ASAP7_75t_R _22136_ (.A(net1208),
    .Y(out[1145]));
 BUFx2_ASAP7_75t_R _22137_ (.A(net1209),
    .Y(out[1146]));
 BUFx2_ASAP7_75t_R _22138_ (.A(net1210),
    .Y(out[1147]));
 BUFx2_ASAP7_75t_R _22139_ (.A(net1211),
    .Y(out[1148]));
 BUFx2_ASAP7_75t_R _22140_ (.A(net1212),
    .Y(out[1149]));
 BUFx2_ASAP7_75t_R _22141_ (.A(net1213),
    .Y(out[1150]));
 BUFx2_ASAP7_75t_R _22142_ (.A(net1214),
    .Y(out[1151]));
 BUFx2_ASAP7_75t_R _22143_ (.A(net1215),
    .Y(out[1157]));
 BUFx2_ASAP7_75t_R _22144_ (.A(net1216),
    .Y(out[1158]));
 BUFx2_ASAP7_75t_R _22145_ (.A(net1217),
    .Y(out[1161]));
 BUFx2_ASAP7_75t_R _22146_ (.A(net1218),
    .Y(out[1162]));
 BUFx2_ASAP7_75t_R _22147_ (.A(net1219),
    .Y(out[1163]));
 BUFx2_ASAP7_75t_R _22148_ (.A(net1220),
    .Y(out[1164]));
 BUFx2_ASAP7_75t_R _22149_ (.A(net1221),
    .Y(out[1165]));
 BUFx2_ASAP7_75t_R _22150_ (.A(net1222),
    .Y(out[1166]));
 BUFx2_ASAP7_75t_R _22151_ (.A(net1223),
    .Y(out[1167]));
 BUFx2_ASAP7_75t_R _22152_ (.A(net1224),
    .Y(out[1168]));
 BUFx2_ASAP7_75t_R _22153_ (.A(net1225),
    .Y(out[1169]));
 BUFx3_ASAP7_75t_R _22154_ (.A(net73),
    .Y(net70));
 BUFx2_ASAP7_75t_R _22155_ (.A(net1226),
    .Y(out[1171]));
 BUFx3_ASAP7_75t_R _22156_ (.A(net73),
    .Y(net71));
 BUFx3_ASAP7_75t_R _22157_ (.A(net73),
    .Y(net72));
 BUFx2_ASAP7_75t_R _22158_ (.A(net1227),
    .Y(out[1175]));
 BUFx2_ASAP7_75t_R _22159_ (.A(net1228),
    .Y(out[1176]));
 BUFx2_ASAP7_75t_R _22160_ (.A(net1229),
    .Y(out[1177]));
 BUFx2_ASAP7_75t_R _22161_ (.A(net1230),
    .Y(out[1178]));
 BUFx2_ASAP7_75t_R _22162_ (.A(net1231),
    .Y(out[1179]));
 BUFx2_ASAP7_75t_R _22163_ (.A(net1232),
    .Y(out[1180]));
 BUFx2_ASAP7_75t_R _22164_ (.A(net1233),
    .Y(out[1181]));
 BUFx2_ASAP7_75t_R _22165_ (.A(net1234),
    .Y(out[1182]));
 BUFx2_ASAP7_75t_R _22166_ (.A(net1235),
    .Y(out[1183]));
 BUFx2_ASAP7_75t_R _22167_ (.A(net1236),
    .Y(out[1184]));
 BUFx2_ASAP7_75t_R _22168_ (.A(net1237),
    .Y(out[1185]));
 BUFx2_ASAP7_75t_R _22169_ (.A(net1238),
    .Y(out[1186]));
 BUFx2_ASAP7_75t_R _22170_ (.A(net1239),
    .Y(out[1187]));
 BUFx2_ASAP7_75t_R _22171_ (.A(net1240),
    .Y(out[1188]));
 BUFx2_ASAP7_75t_R _22172_ (.A(net1241),
    .Y(out[1189]));
 BUFx2_ASAP7_75t_R _22173_ (.A(net1242),
    .Y(out[1190]));
 BUFx2_ASAP7_75t_R _22174_ (.A(net1243),
    .Y(out[1191]));
 BUFx2_ASAP7_75t_R _22175_ (.A(net1244),
    .Y(out[1197]));
 BUFx2_ASAP7_75t_R _22176_ (.A(net1245),
    .Y(out[1198]));
 BUFx2_ASAP7_75t_R _22177_ (.A(net1246),
    .Y(out[1201]));
 BUFx2_ASAP7_75t_R _22178_ (.A(net1247),
    .Y(out[1202]));
 BUFx2_ASAP7_75t_R _22179_ (.A(net1248),
    .Y(out[1203]));
 BUFx2_ASAP7_75t_R _22180_ (.A(net1249),
    .Y(out[1204]));
 BUFx2_ASAP7_75t_R _22181_ (.A(net1250),
    .Y(out[1205]));
 BUFx2_ASAP7_75t_R _22182_ (.A(net1251),
    .Y(out[1206]));
 BUFx2_ASAP7_75t_R _22183_ (.A(net1252),
    .Y(out[1207]));
 BUFx2_ASAP7_75t_R _22184_ (.A(net1253),
    .Y(out[1208]));
 BUFx2_ASAP7_75t_R _22185_ (.A(net1254),
    .Y(out[1209]));
 BUFx2_ASAP7_75t_R _22186_ (.A(net1255),
    .Y(out[1210]));
 BUFx3_ASAP7_75t_R _22187_ (.A(net86),
    .Y(net83));
 BUFx3_ASAP7_75t_R _22188_ (.A(net86),
    .Y(net84));
 BUFx3_ASAP7_75t_R _22189_ (.A(net86),
    .Y(net85));
 BUFx2_ASAP7_75t_R _22190_ (.A(net1256),
    .Y(out[1215]));
 BUFx2_ASAP7_75t_R _22191_ (.A(net1257),
    .Y(out[1216]));
 BUFx2_ASAP7_75t_R _22192_ (.A(net1258),
    .Y(out[1217]));
 BUFx2_ASAP7_75t_R _22193_ (.A(net1259),
    .Y(out[1218]));
 BUFx2_ASAP7_75t_R _22194_ (.A(net1260),
    .Y(out[1219]));
 BUFx2_ASAP7_75t_R _22195_ (.A(net1261),
    .Y(out[1220]));
 BUFx2_ASAP7_75t_R _22196_ (.A(net1262),
    .Y(out[1221]));
 BUFx2_ASAP7_75t_R _22197_ (.A(net1263),
    .Y(out[1222]));
 BUFx2_ASAP7_75t_R _22198_ (.A(net1264),
    .Y(out[1223]));
 BUFx2_ASAP7_75t_R _22199_ (.A(net1265),
    .Y(out[1224]));
 BUFx2_ASAP7_75t_R _22200_ (.A(net1266),
    .Y(out[1225]));
 BUFx2_ASAP7_75t_R _22201_ (.A(net1267),
    .Y(out[1226]));
 BUFx2_ASAP7_75t_R _22202_ (.A(net1268),
    .Y(out[1227]));
 BUFx2_ASAP7_75t_R _22203_ (.A(net1269),
    .Y(out[1228]));
 BUFx2_ASAP7_75t_R _22204_ (.A(net1270),
    .Y(out[1229]));
 BUFx2_ASAP7_75t_R _22205_ (.A(net1271),
    .Y(out[1230]));
 BUFx2_ASAP7_75t_R _22206_ (.A(net1272),
    .Y(out[1231]));
 BUFx2_ASAP7_75t_R _22207_ (.A(net1273),
    .Y(out[1237]));
 BUFx2_ASAP7_75t_R _22208_ (.A(net1274),
    .Y(out[1238]));
 BUFx2_ASAP7_75t_R _22209_ (.A(net1275),
    .Y(out[1241]));
 BUFx2_ASAP7_75t_R _22210_ (.A(net1276),
    .Y(out[1242]));
 BUFx2_ASAP7_75t_R _22211_ (.A(net1277),
    .Y(out[1243]));
 BUFx2_ASAP7_75t_R _22212_ (.A(net1278),
    .Y(out[1244]));
 BUFx2_ASAP7_75t_R _22213_ (.A(net1279),
    .Y(out[1245]));
 BUFx2_ASAP7_75t_R _22214_ (.A(net1280),
    .Y(out[1246]));
 BUFx2_ASAP7_75t_R _22215_ (.A(net1281),
    .Y(out[1247]));
 BUFx2_ASAP7_75t_R _22216_ (.A(net1282),
    .Y(out[1248]));
 BUFx2_ASAP7_75t_R _22217_ (.A(net1283),
    .Y(out[1249]));
 BUFx3_ASAP7_75t_R _22218_ (.A(net98),
    .Y(net94));
 BUFx3_ASAP7_75t_R _22219_ (.A(net98),
    .Y(net95));
 BUFx3_ASAP7_75t_R _22220_ (.A(net98),
    .Y(net96));
 BUFx3_ASAP7_75t_R _22221_ (.A(net98),
    .Y(net97));
 BUFx2_ASAP7_75t_R _22222_ (.A(net1284),
    .Y(out[1255]));
 BUFx2_ASAP7_75t_R _22223_ (.A(net1285),
    .Y(out[1256]));
 BUFx2_ASAP7_75t_R _22224_ (.A(net1286),
    .Y(out[1257]));
 BUFx2_ASAP7_75t_R _22225_ (.A(net1287),
    .Y(out[1258]));
 BUFx2_ASAP7_75t_R _22226_ (.A(net1288),
    .Y(out[1259]));
 BUFx2_ASAP7_75t_R _22227_ (.A(net1289),
    .Y(out[1260]));
 BUFx2_ASAP7_75t_R _22228_ (.A(net1290),
    .Y(out[1261]));
 BUFx2_ASAP7_75t_R _22229_ (.A(net1291),
    .Y(out[1262]));
 BUFx2_ASAP7_75t_R _22230_ (.A(net1292),
    .Y(out[1263]));
 BUFx2_ASAP7_75t_R _22231_ (.A(net1293),
    .Y(out[1264]));
 BUFx2_ASAP7_75t_R _22232_ (.A(net1294),
    .Y(out[1265]));
 BUFx2_ASAP7_75t_R _22233_ (.A(net1295),
    .Y(out[1266]));
 BUFx2_ASAP7_75t_R _22234_ (.A(net1296),
    .Y(out[1267]));
 BUFx2_ASAP7_75t_R _22235_ (.A(net1297),
    .Y(out[1268]));
 BUFx2_ASAP7_75t_R _22236_ (.A(net1298),
    .Y(out[1269]));
 BUFx2_ASAP7_75t_R _22237_ (.A(net1299),
    .Y(out[1270]));
 BUFx2_ASAP7_75t_R _22238_ (.A(net1300),
    .Y(out[1271]));
 BUFx2_ASAP7_75t_R _22239_ (.A(net1301),
    .Y(out[1277]));
 BUFx2_ASAP7_75t_R _22240_ (.A(net1302),
    .Y(out[1278]));
 DFFHQNx1_ASAP7_75t_R \in_r[0]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(net7),
    .QN(_02343_));
 DFFHQNx1_ASAP7_75t_R \in_r[1]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(net8),
    .QN(_02344_));
 DFFHQNx3_ASAP7_75t_R \in_r[2]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(net9),
    .QN(_02345_));
 DFFHQNx3_ASAP7_75t_R \in_r[31]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(net10),
    .QN(_02346_));
 DFFHQNx3_ASAP7_75t_R \in_r[32]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(net11),
    .QN(_02347_));
 DFFHQNx1_ASAP7_75t_R \in_r[33]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(net12),
    .QN(_02348_));
 DFFHQNx1_ASAP7_75t_R \in_r[34]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(net13),
    .QN(_02349_));
 DFFHQNx1_ASAP7_75t_R \in_r[35]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(net14),
    .QN(_02350_));
 DFFHQNx1_ASAP7_75t_R \in_r[36]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(net15),
    .QN(_02351_));
 DFFHQNx1_ASAP7_75t_R \in_r[37]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(net16),
    .QN(_02352_));
 DFFHQNx3_ASAP7_75t_R \in_r[38]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(net17),
    .QN(_02353_));
 DFFHQNx3_ASAP7_75t_R \in_r[39]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(net18),
    .QN(_02354_));
 DFFHQNx1_ASAP7_75t_R \in_r[3]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(net19),
    .QN(_02355_));
 DFFHQNx3_ASAP7_75t_R \in_r[4]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(net20),
    .QN(_02342_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_02675_),
    .QN(_00000_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_02676_),
    .QN(_02341_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_02677_),
    .QN(_02340_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_02678_),
    .QN(_02339_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_02679_),
    .QN(_02338_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_02680_),
    .QN(_02337_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_02681_),
    .QN(_02336_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_02682_),
    .QN(_02335_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_02683_),
    .QN(_02334_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_02684_),
    .QN(_02333_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02685_),
    .QN(_02332_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_02686_),
    .QN(_02331_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_02687_),
    .QN(_02330_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_02688_),
    .QN(_02329_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_02689_),
    .QN(_02328_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_02690_),
    .QN(_02327_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_02691_),
    .QN(_02326_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02692_),
    .QN(_02325_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_02693_),
    .QN(_02324_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_02694_),
    .QN(_02323_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_02695_),
    .QN(_02322_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02696_),
    .QN(_02321_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_02697_),
    .QN(_02320_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_02698_),
    .QN(_02319_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02699_),
    .QN(_02318_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_02700_),
    .QN(_02317_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_02701_),
    .QN(_02316_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_02702_),
    .QN(_02315_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02703_),
    .QN(_02314_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02704_),
    .QN(_02313_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02705_),
    .QN(_02312_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02706_),
    .QN(_02311_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02707_),
    .QN(_02310_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02708_),
    .QN(_02309_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02709_),
    .QN(_02308_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02710_),
    .QN(_02307_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02711_),
    .QN(_02306_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02712_),
    .QN(_02305_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02713_),
    .QN(_02304_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02714_),
    .QN(_02303_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02715_),
    .QN(_02302_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02716_),
    .QN(_02301_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[0].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02717_),
    .QN(_02300_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_02718_),
    .QN(_00001_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_02719_),
    .QN(_02299_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_02720_),
    .QN(_02298_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_02721_),
    .QN(_02297_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_02722_),
    .QN(_02296_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_02723_),
    .QN(_02295_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02724_),
    .QN(_02294_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02725_),
    .QN(_02293_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_02726_),
    .QN(_02292_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_02727_),
    .QN(_02291_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_02728_),
    .QN(_02290_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02729_),
    .QN(_02289_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02730_),
    .QN(_02288_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_02731_),
    .QN(_02287_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_02732_),
    .QN(_02286_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_02733_),
    .QN(_02285_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_02734_),
    .QN(_02284_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_02735_),
    .QN(_02283_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_02736_),
    .QN(_02282_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_02737_),
    .QN(_02281_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_02738_),
    .QN(_02280_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_02739_),
    .QN(_02279_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_02740_),
    .QN(_02278_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_02741_),
    .QN(_02277_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_02742_),
    .QN(_02276_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_02743_),
    .QN(_02275_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_02744_),
    .QN(_02274_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_02745_),
    .QN(_02273_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_02746_),
    .QN(_02272_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_02747_),
    .QN(_02271_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_02748_),
    .QN(_02270_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_02749_),
    .QN(_02269_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_02750_),
    .QN(_02268_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_02751_),
    .QN(_02267_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_02752_),
    .QN(_02266_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_02753_),
    .QN(_02265_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_02754_),
    .QN(_02264_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_02755_),
    .QN(_02263_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_02756_),
    .QN(_02262_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_02757_),
    .QN(_02261_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_02758_),
    .QN(_02260_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_02759_),
    .QN(_02259_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[1].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_02760_),
    .QN(_02258_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_02761_),
    .QN(_00002_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_02762_),
    .QN(_02257_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_02763_),
    .QN(_02256_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_02764_),
    .QN(_02255_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_02765_),
    .QN(_02254_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_02766_),
    .QN(_02253_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02767_),
    .QN(_02252_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02768_),
    .QN(_02251_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_02769_),
    .QN(_02250_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02770_),
    .QN(_02249_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02771_),
    .QN(_02248_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02772_),
    .QN(_02247_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_02773_),
    .QN(_02246_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02774_),
    .QN(_02245_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_02775_),
    .QN(_02244_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_02776_),
    .QN(_02243_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_02777_),
    .QN(_02242_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_02778_),
    .QN(_02241_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_02779_),
    .QN(_02240_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_02780_),
    .QN(_02239_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_02781_),
    .QN(_02238_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_02782_),
    .QN(_02237_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_02783_),
    .QN(_02236_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_02784_),
    .QN(_02235_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02785_),
    .QN(_02234_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_02786_),
    .QN(_02233_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_02787_),
    .QN(_02232_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_02788_),
    .QN(_02231_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_02789_),
    .QN(_02230_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02790_),
    .QN(_02229_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02791_),
    .QN(_02228_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02792_),
    .QN(_02227_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02793_),
    .QN(_02226_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02794_),
    .QN(_02225_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02795_),
    .QN(_02224_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02796_),
    .QN(_02223_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02797_),
    .QN(_02222_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02798_),
    .QN(_02221_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02799_),
    .QN(_02220_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02800_),
    .QN(_02219_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02801_),
    .QN(_02218_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02802_),
    .QN(_02217_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[2].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_02803_),
    .QN(_02216_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02804_),
    .QN(_00003_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_02805_),
    .QN(_02215_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02806_),
    .QN(_02214_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02807_),
    .QN(_02213_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_02808_),
    .QN(_02212_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_02809_),
    .QN(_02211_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02810_),
    .QN(_02210_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_02811_),
    .QN(_02209_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_02812_),
    .QN(_02208_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02813_),
    .QN(_02207_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02814_),
    .QN(_02206_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_02815_),
    .QN(_02205_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02816_),
    .QN(_02204_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02817_),
    .QN(_02203_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02818_),
    .QN(_02202_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02819_),
    .QN(_02201_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02820_),
    .QN(_02200_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02821_),
    .QN(_02199_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02822_),
    .QN(_02198_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02823_),
    .QN(_02197_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_02824_),
    .QN(_02196_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02825_),
    .QN(_02195_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02826_),
    .QN(_02194_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02827_),
    .QN(_02193_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_02828_),
    .QN(_02192_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_02829_),
    .QN(_02191_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_02830_),
    .QN(_02190_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02831_),
    .QN(_02189_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02832_),
    .QN(_02188_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02833_),
    .QN(_02187_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02834_),
    .QN(_02186_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02835_),
    .QN(_02185_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02836_),
    .QN(_02184_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02837_),
    .QN(_02183_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02838_),
    .QN(_02182_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_02839_),
    .QN(_02181_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_02840_),
    .QN(_02180_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02841_),
    .QN(_02179_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02842_),
    .QN(_02178_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02843_),
    .QN(_02177_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02844_),
    .QN(_02176_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02845_),
    .QN(_02175_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[3].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_02846_),
    .QN(_02174_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02847_),
    .QN(_00004_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02848_),
    .QN(_02173_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_02849_),
    .QN(_02172_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_02850_),
    .QN(_02171_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02851_),
    .QN(_02170_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02852_),
    .QN(_02169_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_02853_),
    .QN(_02168_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02854_),
    .QN(_02167_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_02855_),
    .QN(_02166_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02856_),
    .QN(_02165_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02857_),
    .QN(_02164_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02858_),
    .QN(_02163_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02859_),
    .QN(_02162_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_02860_),
    .QN(_02161_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_02861_),
    .QN(_02160_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02862_),
    .QN(_02159_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02863_),
    .QN(_02158_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02864_),
    .QN(_02157_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02865_),
    .QN(_02156_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02866_),
    .QN(_02155_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02867_),
    .QN(_02154_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02868_),
    .QN(_02153_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02869_),
    .QN(_02152_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02870_),
    .QN(_02151_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02871_),
    .QN(_02150_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02872_),
    .QN(_02149_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02873_),
    .QN(_02148_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02874_),
    .QN(_02147_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_02875_),
    .QN(_02146_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02876_),
    .QN(_02145_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02877_),
    .QN(_02144_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02878_),
    .QN(_02143_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02879_),
    .QN(_02142_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02880_),
    .QN(_02141_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02881_),
    .QN(_02140_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02882_),
    .QN(_02139_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02883_),
    .QN(_02138_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02884_),
    .QN(_02137_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02885_),
    .QN(_02136_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02886_),
    .QN(_02135_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02887_),
    .QN(_02134_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02888_),
    .QN(_02133_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[4].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02889_),
    .QN(_02132_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_02890_),
    .QN(_00005_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02891_),
    .QN(_02131_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02892_),
    .QN(_02130_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02893_),
    .QN(_02129_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02894_),
    .QN(_02128_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02895_),
    .QN(_02127_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02896_),
    .QN(_02126_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02897_),
    .QN(_02125_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02898_),
    .QN(_02124_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02899_),
    .QN(_02123_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02900_),
    .QN(_02122_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02901_),
    .QN(_02121_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02902_),
    .QN(_02120_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02903_),
    .QN(_02119_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02904_),
    .QN(_02118_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02905_),
    .QN(_02117_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_02906_),
    .QN(_02116_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02907_),
    .QN(_02115_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_02908_),
    .QN(_02114_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02909_),
    .QN(_02113_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02910_),
    .QN(_02112_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02911_),
    .QN(_02111_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02912_),
    .QN(_02110_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02913_),
    .QN(_02109_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_02914_),
    .QN(_02108_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_02915_),
    .QN(_02107_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_02916_),
    .QN(_02106_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_02917_),
    .QN(_02105_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_02918_),
    .QN(_02104_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02919_),
    .QN(_02103_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02920_),
    .QN(_02102_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02921_),
    .QN(_02101_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02922_),
    .QN(_02100_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_02923_),
    .QN(_02099_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02924_),
    .QN(_02098_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02925_),
    .QN(_02097_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02926_),
    .QN(_02096_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02927_),
    .QN(_02095_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02928_),
    .QN(_02094_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02929_),
    .QN(_02093_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02930_),
    .QN(_02092_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02931_),
    .QN(_02091_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[5].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02932_),
    .QN(_02090_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02933_),
    .QN(_00006_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02934_),
    .QN(_02089_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02935_),
    .QN(_02088_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02936_),
    .QN(_02087_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02937_),
    .QN(_02086_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02938_),
    .QN(_02085_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02939_),
    .QN(_02084_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02940_),
    .QN(_02083_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02941_),
    .QN(_02082_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02942_),
    .QN(_02081_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02943_),
    .QN(_02080_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02944_),
    .QN(_02079_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_02945_),
    .QN(_02078_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02946_),
    .QN(_02077_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02947_),
    .QN(_02076_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02948_),
    .QN(_02075_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_02949_),
    .QN(_02074_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_02950_),
    .QN(_02073_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_02951_),
    .QN(_02072_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02952_),
    .QN(_02071_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02953_),
    .QN(_02070_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02954_),
    .QN(_02069_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02955_),
    .QN(_02068_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02956_),
    .QN(_02067_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02957_),
    .QN(_02066_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02958_),
    .QN(_02065_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02959_),
    .QN(_02064_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_02960_),
    .QN(_02063_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_02961_),
    .QN(_02062_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02962_),
    .QN(_02061_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02963_),
    .QN(_02060_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02964_),
    .QN(_02059_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02965_),
    .QN(_02058_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02966_),
    .QN(_02057_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02967_),
    .QN(_02056_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02968_),
    .QN(_02055_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02969_),
    .QN(_02054_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02970_),
    .QN(_02053_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02971_),
    .QN(_02052_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02972_),
    .QN(_02051_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_02973_),
    .QN(_02050_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_02974_),
    .QN(_02049_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[6].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_02975_),
    .QN(_02048_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02976_),
    .QN(_00007_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_02977_),
    .QN(_02047_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02978_),
    .QN(_02046_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02979_),
    .QN(_02045_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02980_),
    .QN(_02044_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02981_),
    .QN(_02043_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_02982_),
    .QN(_02042_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_02983_),
    .QN(_02041_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02984_),
    .QN(_02040_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02985_),
    .QN(_02039_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02986_),
    .QN(_02038_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_02987_),
    .QN(_02037_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02988_),
    .QN(_02036_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02989_),
    .QN(_02035_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02990_),
    .QN(_02034_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_02991_),
    .QN(_02033_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_02992_),
    .QN(_02032_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_02993_),
    .QN(_02031_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_02994_),
    .QN(_02030_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_02995_),
    .QN(_02029_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_02996_),
    .QN(_02028_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_02997_),
    .QN(_02027_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02998_),
    .QN(_02026_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_02999_),
    .QN(_02025_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03000_),
    .QN(_02024_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03001_),
    .QN(_02023_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03002_),
    .QN(_02022_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03003_),
    .QN(_02021_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03004_),
    .QN(_02020_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03005_),
    .QN(_02019_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03006_),
    .QN(_02018_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03007_),
    .QN(_02017_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03008_),
    .QN(_02016_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03009_),
    .QN(_02015_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03010_),
    .QN(_02014_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03011_),
    .QN(_02013_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03012_),
    .QN(_02012_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03013_),
    .QN(_02011_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03014_),
    .QN(_02010_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03015_),
    .QN(_02009_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03016_),
    .QN(_02008_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03017_),
    .QN(_02007_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[1].ms[7].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03018_),
    .QN(_02006_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03019_),
    .QN(_00008_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03020_),
    .QN(_02005_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03021_),
    .QN(_02004_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03022_),
    .QN(_02003_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03023_),
    .QN(_02002_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03024_),
    .QN(_02001_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03025_),
    .QN(_02000_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03026_),
    .QN(_01999_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03027_),
    .QN(_01998_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03028_),
    .QN(_01997_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03029_),
    .QN(_01996_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03030_),
    .QN(_01995_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03031_),
    .QN(_01994_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03032_),
    .QN(_01993_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03033_),
    .QN(_01992_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_03034_),
    .QN(_01991_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03035_),
    .QN(_01990_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_03036_),
    .QN(_01989_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03037_),
    .QN(_01988_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03038_),
    .QN(_01987_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03039_),
    .QN(_01986_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03040_),
    .QN(_01985_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03041_),
    .QN(_01984_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03042_),
    .QN(_01983_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03043_),
    .QN(_01982_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03044_),
    .QN(_01981_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03045_),
    .QN(_01980_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03046_),
    .QN(_01979_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03047_),
    .QN(_01978_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03048_),
    .QN(_01977_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03049_),
    .QN(_01976_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03050_),
    .QN(_01975_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03051_),
    .QN(_01974_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03052_),
    .QN(_01973_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03053_),
    .QN(_01972_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03054_),
    .QN(_01971_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03055_),
    .QN(_01970_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03056_),
    .QN(_01969_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03057_),
    .QN(_01968_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03058_),
    .QN(_01967_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03059_),
    .QN(_01966_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03060_),
    .QN(_01965_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[0].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03061_),
    .QN(_01964_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03062_),
    .QN(_00009_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03063_),
    .QN(_01963_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03064_),
    .QN(_01962_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03065_),
    .QN(_01961_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03066_),
    .QN(_01960_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03067_),
    .QN(_01959_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03068_),
    .QN(_01958_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03069_),
    .QN(_01957_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03070_),
    .QN(_01956_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03071_),
    .QN(_01955_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03072_),
    .QN(_01954_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03073_),
    .QN(_01953_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03074_),
    .QN(_01952_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03075_),
    .QN(_01951_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03076_),
    .QN(_01950_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03077_),
    .QN(_01949_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03078_),
    .QN(_01948_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03079_),
    .QN(_01947_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03080_),
    .QN(_01946_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03081_),
    .QN(_01945_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03082_),
    .QN(_01944_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03083_),
    .QN(_01943_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03084_),
    .QN(_01942_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03085_),
    .QN(_01941_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03086_),
    .QN(_01940_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03087_),
    .QN(_01939_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03088_),
    .QN(_01938_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03089_),
    .QN(_01937_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03090_),
    .QN(_01936_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03091_),
    .QN(_01935_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03092_),
    .QN(_01934_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03093_),
    .QN(_01933_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03094_),
    .QN(_01932_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03095_),
    .QN(_01931_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03096_),
    .QN(_01930_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03097_),
    .QN(_01929_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03098_),
    .QN(_01928_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03099_),
    .QN(_01927_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03100_),
    .QN(_01926_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03101_),
    .QN(_01925_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03102_),
    .QN(_01924_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03103_),
    .QN(_01923_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[1].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03104_),
    .QN(_01922_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03105_),
    .QN(_00010_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03106_),
    .QN(_01921_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03107_),
    .QN(_01920_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03108_),
    .QN(_01919_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03109_),
    .QN(_01918_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03110_),
    .QN(_01917_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03111_),
    .QN(_01916_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03112_),
    .QN(_01915_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03113_),
    .QN(_01914_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03114_),
    .QN(_01913_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03115_),
    .QN(_01912_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03116_),
    .QN(_01911_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03117_),
    .QN(_01910_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03118_),
    .QN(_01909_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03119_),
    .QN(_01908_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03120_),
    .QN(_01907_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03121_),
    .QN(_01906_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03122_),
    .QN(_01905_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03123_),
    .QN(_01904_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03124_),
    .QN(_01903_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03125_),
    .QN(_01902_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03126_),
    .QN(_01901_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03127_),
    .QN(_01900_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03128_),
    .QN(_01899_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03129_),
    .QN(_01898_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03130_),
    .QN(_01897_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03131_),
    .QN(_01896_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03132_),
    .QN(_01895_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03133_),
    .QN(_01894_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03134_),
    .QN(_01893_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03135_),
    .QN(_01892_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03136_),
    .QN(_01891_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03137_),
    .QN(_01890_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03138_),
    .QN(_01889_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03139_),
    .QN(_01888_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03140_),
    .QN(_01887_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03141_),
    .QN(_01886_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03142_),
    .QN(_01885_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03143_),
    .QN(_01884_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03144_),
    .QN(_01883_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03145_),
    .QN(_01882_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03146_),
    .QN(_01881_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[2].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03147_),
    .QN(_01880_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03148_),
    .QN(_00011_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03149_),
    .QN(_01879_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03150_),
    .QN(_01878_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03151_),
    .QN(_01877_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03152_),
    .QN(_01876_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03153_),
    .QN(_01875_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03154_),
    .QN(_01874_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03155_),
    .QN(_01873_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03156_),
    .QN(_01872_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03157_),
    .QN(_01871_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03158_),
    .QN(_01870_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03159_),
    .QN(_01869_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03160_),
    .QN(_01868_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03161_),
    .QN(_01867_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03162_),
    .QN(_01866_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03163_),
    .QN(_01865_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03164_),
    .QN(_01864_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03165_),
    .QN(_01863_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03166_),
    .QN(_01862_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03167_),
    .QN(_01861_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03168_),
    .QN(_01860_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03169_),
    .QN(_01859_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03170_),
    .QN(_01858_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_03171_),
    .QN(_01857_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03172_),
    .QN(_01856_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03173_),
    .QN(_01855_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03174_),
    .QN(_01854_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03175_),
    .QN(_01853_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03176_),
    .QN(_01852_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03177_),
    .QN(_01851_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03178_),
    .QN(_01850_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03179_),
    .QN(_01849_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03180_),
    .QN(_01848_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03181_),
    .QN(_01847_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03182_),
    .QN(_01846_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03183_),
    .QN(_01845_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03184_),
    .QN(_01844_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03185_),
    .QN(_01843_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03186_),
    .QN(_01842_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03187_),
    .QN(_01841_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03188_),
    .QN(_01840_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03189_),
    .QN(_01839_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[2].ms[3].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03190_),
    .QN(_01838_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_03191_),
    .QN(_00012_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03192_),
    .QN(_01837_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03193_),
    .QN(_01836_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03194_),
    .QN(_01835_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03195_),
    .QN(_01834_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03196_),
    .QN(_01833_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03197_),
    .QN(_01832_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03198_),
    .QN(_01831_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03199_),
    .QN(_01830_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03200_),
    .QN(_01829_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03201_),
    .QN(_01828_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03202_),
    .QN(_01827_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03203_),
    .QN(_01826_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03204_),
    .QN(_01825_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03205_),
    .QN(_01824_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03206_),
    .QN(_01823_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03207_),
    .QN(_01822_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03208_),
    .QN(_01821_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03209_),
    .QN(_01820_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03210_),
    .QN(_01819_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03211_),
    .QN(_01818_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03212_),
    .QN(_01817_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03213_),
    .QN(_01816_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03214_),
    .QN(_01815_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03215_),
    .QN(_01814_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03216_),
    .QN(_01813_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03217_),
    .QN(_01812_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03218_),
    .QN(_01811_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03219_),
    .QN(_01810_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03220_),
    .QN(_01809_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03221_),
    .QN(_01808_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03222_),
    .QN(_01807_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03223_),
    .QN(_01806_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03224_),
    .QN(_01805_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03225_),
    .QN(_01804_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03226_),
    .QN(_01803_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03227_),
    .QN(_01802_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03228_),
    .QN(_01801_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03229_),
    .QN(_01800_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03230_),
    .QN(_01799_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03231_),
    .QN(_01798_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03232_),
    .QN(_01797_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[0].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03233_),
    .QN(_01796_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03234_),
    .QN(_00013_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03235_),
    .QN(_01795_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03236_),
    .QN(_01794_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03237_),
    .QN(_01793_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03238_),
    .QN(_01792_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03239_),
    .QN(_01791_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03240_),
    .QN(_01790_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03241_),
    .QN(_01789_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03242_),
    .QN(_01788_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03243_),
    .QN(_01787_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03244_),
    .QN(_01786_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03245_),
    .QN(_01785_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03246_),
    .QN(_01784_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03247_),
    .QN(_01783_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03248_),
    .QN(_01782_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03249_),
    .QN(_01781_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03250_),
    .QN(_01780_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03251_),
    .QN(_01779_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03252_),
    .QN(_01778_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03253_),
    .QN(_01777_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03254_),
    .QN(_01776_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03255_),
    .QN(_01775_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03256_),
    .QN(_01774_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03257_),
    .QN(_01773_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03258_),
    .QN(_01772_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03259_),
    .QN(_01771_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03260_),
    .QN(_01770_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03261_),
    .QN(_01769_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03262_),
    .QN(_01768_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03263_),
    .QN(_01767_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03264_),
    .QN(_01766_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03265_),
    .QN(_01765_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03266_),
    .QN(_01764_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03267_),
    .QN(_01763_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03268_),
    .QN(_01762_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03269_),
    .QN(_01761_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03270_),
    .QN(_01760_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03271_),
    .QN(_01759_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03272_),
    .QN(_01758_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03273_),
    .QN(_01757_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03274_),
    .QN(_01756_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03275_),
    .QN(_01755_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[3].ms[1].ns[0].t_level.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03276_),
    .QN(_01754_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03277_),
    .QN(_00014_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03278_),
    .QN(_01753_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03279_),
    .QN(_01752_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03280_),
    .QN(_01751_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03281_),
    .QN(_01750_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03282_),
    .QN(_01749_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03283_),
    .QN(_01748_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03284_),
    .QN(_01747_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03285_),
    .QN(_01746_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03286_),
    .QN(_01745_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03287_),
    .QN(_01744_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03288_),
    .QN(_01743_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03289_),
    .QN(_01742_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03290_),
    .QN(_01741_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03291_),
    .QN(_01740_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03292_),
    .QN(_01739_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03293_),
    .QN(_01738_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03294_),
    .QN(_01737_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03295_),
    .QN(_01736_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03296_),
    .QN(_01735_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03297_),
    .QN(_01734_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_03298_),
    .QN(_01733_));
 DFFHQNx1_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03299_),
    .QN(_01732_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03300_),
    .QN(_01731_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03301_),
    .QN(_01730_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03302_),
    .QN(_01729_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03303_),
    .QN(_01728_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03304_),
    .QN(_01727_));
 DFFHQNx3_ASAP7_75t_R \n2.ls[4].ms[0].ns[0].t_level.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03305_),
    .QN(_02356_));
 DFFHQNx1_ASAP7_75t_R \out_r[0]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(\peo[0][0] ),
    .QN(_02357_));
 DFFHQNx1_ASAP7_75t_R \out_r[1000]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(\peo[25][0] ),
    .QN(_02358_));
 DFFHQNx1_ASAP7_75t_R \out_r[1014]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\peo[25][10] ),
    .QN(_02359_));
 DFFHQNx1_ASAP7_75t_R \out_r[1032]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(\peo[25][32] ),
    .QN(_02360_));
 DFFHQNx1_ASAP7_75t_R \out_r[1033]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\xs[12].cli1.i[33] ),
    .QN(_02361_));
 DFFHQNx1_ASAP7_75t_R \out_r[1034]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\xs[12].cli1.i[34] ),
    .QN(_02362_));
 DFFHQNx1_ASAP7_75t_R \out_r[1035]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(\xs[12].cli1.i[35] ),
    .QN(_02363_));
 DFFHQNx1_ASAP7_75t_R \out_r[1036]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(\xs[12].cli1.i[36] ),
    .QN(_02364_));
 DFFHQNx1_ASAP7_75t_R \out_r[1039]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(\xs[12].cli1.i[39] ),
    .QN(_02365_));
 DFFHQNx1_ASAP7_75t_R \out_r[1040]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\peo[26][0] ),
    .QN(_02366_));
 DFFHQNx1_ASAP7_75t_R \out_r[1054]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\peo[26][11] ),
    .QN(_02367_));
 DFFHQNx1_ASAP7_75t_R \out_r[1072]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\peo[26][32] ),
    .QN(_02368_));
 DFFHQNx1_ASAP7_75t_R \out_r[1073]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\peo[26][33] ),
    .QN(_02369_));
 DFFHQNx1_ASAP7_75t_R \out_r[1074]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\peo[26][34] ),
    .QN(_02370_));
 DFFHQNx1_ASAP7_75t_R \out_r[1075]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(\peo[26][35] ),
    .QN(_02371_));
 DFFHQNx1_ASAP7_75t_R \out_r[1076]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\peo[26][36] ),
    .QN(_02372_));
 DFFHQNx1_ASAP7_75t_R \out_r[1079]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\peo[26][39] ),
    .QN(_02373_));
 DFFHQNx1_ASAP7_75t_R \out_r[1080]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\peo[27][0] ),
    .QN(_02374_));
 DFFHQNx1_ASAP7_75t_R \out_r[1094]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(\peo[27][10] ),
    .QN(_02375_));
 DFFHQNx1_ASAP7_75t_R \out_r[1112]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\peo[27][32] ),
    .QN(_02376_));
 DFFHQNx1_ASAP7_75t_R \out_r[1113]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\xs[13].cli1.i[33] ),
    .QN(_02377_));
 DFFHQNx1_ASAP7_75t_R \out_r[1114]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\xs[13].cli1.i[34] ),
    .QN(_02378_));
 DFFHQNx1_ASAP7_75t_R \out_r[1115]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\xs[13].cli1.i[35] ),
    .QN(_02379_));
 DFFHQNx1_ASAP7_75t_R \out_r[1116]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\xs[13].cli1.i[36] ),
    .QN(_02380_));
 DFFHQNx1_ASAP7_75t_R \out_r[1119]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\xs[13].cli1.i[39] ),
    .QN(_02381_));
 DFFHQNx1_ASAP7_75t_R \out_r[1120]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .D(\peo[28][0] ),
    .QN(_02382_));
 DFFHQNx1_ASAP7_75t_R \out_r[112]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(\peo[2][32] ),
    .QN(_02383_));
 DFFHQNx1_ASAP7_75t_R \out_r[1134]$_DFF_P_  (.CLK(clknet_leaf_47_clk),
    .D(\peo[28][12] ),
    .QN(_02384_));
 DFFHQNx1_ASAP7_75t_R \out_r[113]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(\peo[2][33] ),
    .QN(_02385_));
 DFFHQNx1_ASAP7_75t_R \out_r[114]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(\peo[2][34] ),
    .QN(_02386_));
 DFFHQNx1_ASAP7_75t_R \out_r[1152]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .D(\peo[28][32] ),
    .QN(_02387_));
 DFFHQNx1_ASAP7_75t_R \out_r[1153]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .D(\peo[28][33] ),
    .QN(_02388_));
 DFFHQNx1_ASAP7_75t_R \out_r[1154]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .D(\peo[28][34] ),
    .QN(_02389_));
 DFFHQNx1_ASAP7_75t_R \out_r[1155]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .D(\peo[28][35] ),
    .QN(_02390_));
 DFFHQNx1_ASAP7_75t_R \out_r[1156]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .D(\peo[28][36] ),
    .QN(_02391_));
 DFFHQNx1_ASAP7_75t_R \out_r[1159]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .D(\peo[28][39] ),
    .QN(_02392_));
 DFFHQNx1_ASAP7_75t_R \out_r[115]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(\peo[2][35] ),
    .QN(_02393_));
 DFFHQNx1_ASAP7_75t_R \out_r[1160]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .D(\peo[29][0] ),
    .QN(_02394_));
 DFFHQNx1_ASAP7_75t_R \out_r[116]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(\peo[2][36] ),
    .QN(_02395_));
 DFFHQNx1_ASAP7_75t_R \out_r[1174]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .D(\peo[29][10] ),
    .QN(_02396_));
 DFFHQNx1_ASAP7_75t_R \out_r[1192]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .D(\peo[29][32] ),
    .QN(_02397_));
 DFFHQNx1_ASAP7_75t_R \out_r[1193]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .D(\xs[14].cli1.i[33] ),
    .QN(_02398_));
 DFFHQNx1_ASAP7_75t_R \out_r[1194]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .D(\xs[14].cli1.i[34] ),
    .QN(_02399_));
 DFFHQNx1_ASAP7_75t_R \out_r[1195]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .D(\xs[14].cli1.i[35] ),
    .QN(_02400_));
 DFFHQNx1_ASAP7_75t_R \out_r[1196]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .D(\xs[14].cli1.i[36] ),
    .QN(_02401_));
 DFFHQNx1_ASAP7_75t_R \out_r[1199]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .D(\xs[14].cli1.i[39] ),
    .QN(_02402_));
 DFFHQNx1_ASAP7_75t_R \out_r[119]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(\peo[2][39] ),
    .QN(_02403_));
 DFFHQNx1_ASAP7_75t_R \out_r[1200]$_DFF_P_  (.CLK(clknet_leaf_42_clk),
    .D(\peo[30][0] ),
    .QN(_02404_));
 DFFHQNx1_ASAP7_75t_R \out_r[120]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(\peo[3][0] ),
    .QN(_02405_));
 DFFHQNx1_ASAP7_75t_R \out_r[1214]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .D(\peo[30][11] ),
    .QN(_02406_));
 DFFHQNx1_ASAP7_75t_R \out_r[1232]$_DFF_P_  (.CLK(clknet_leaf_42_clk),
    .D(\peo[30][32] ),
    .QN(_02407_));
 DFFHQNx1_ASAP7_75t_R \out_r[1233]$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .D(\peo[30][33] ),
    .QN(_02408_));
 DFFHQNx1_ASAP7_75t_R \out_r[1234]$_DFF_P_  (.CLK(clknet_leaf_42_clk),
    .D(\peo[30][34] ),
    .QN(_02409_));
 DFFHQNx1_ASAP7_75t_R \out_r[1235]$_DFF_P_  (.CLK(clknet_leaf_42_clk),
    .D(\peo[30][35] ),
    .QN(_02410_));
 DFFHQNx1_ASAP7_75t_R \out_r[1236]$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .D(\peo[30][36] ),
    .QN(_02411_));
 DFFHQNx1_ASAP7_75t_R \out_r[1239]$_DFF_P_  (.CLK(clknet_leaf_42_clk),
    .D(\peo[30][39] ),
    .QN(_02412_));
 DFFHQNx1_ASAP7_75t_R \out_r[1240]$_DFF_P_  (.CLK(clknet_leaf_42_clk),
    .D(\peo[31][0] ),
    .QN(_02413_));
 DFFHQNx1_ASAP7_75t_R \out_r[1254]$_DFF_P_  (.CLK(clknet_leaf_53_clk),
    .D(\peo[31][10] ),
    .QN(_02414_));
 DFFHQNx1_ASAP7_75t_R \out_r[1272]$_DFF_P_  (.CLK(clknet_leaf_42_clk),
    .D(\peo[31][32] ),
    .QN(_02415_));
 DFFHQNx1_ASAP7_75t_R \out_r[1273]$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .D(\xs[15].cli1.i[33] ),
    .QN(_02416_));
 DFFHQNx1_ASAP7_75t_R \out_r[1274]$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .D(\xs[15].cli1.i[34] ),
    .QN(_02417_));
 DFFHQNx1_ASAP7_75t_R \out_r[1275]$_DFF_P_  (.CLK(clknet_leaf_42_clk),
    .D(\xs[15].cli1.i[35] ),
    .QN(_02418_));
 DFFHQNx1_ASAP7_75t_R \out_r[1276]$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .D(\xs[15].cli1.i[36] ),
    .QN(_02419_));
 DFFHQNx1_ASAP7_75t_R \out_r[1279]$_DFF_P_  (.CLK(clknet_leaf_45_clk),
    .D(\xs[15].cli1.i[39] ),
    .QN(_02420_));
 DFFHQNx1_ASAP7_75t_R \out_r[131]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(\xs[1].cli1.i[10] ),
    .QN(_02421_));
 DFFHQNx1_ASAP7_75t_R \out_r[152]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\xs[1].cli1.i[32] ),
    .QN(_02422_));
 DFFHQNx1_ASAP7_75t_R \out_r[153]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(\xs[1].cli1.i[33] ),
    .QN(_02423_));
 DFFHQNx1_ASAP7_75t_R \out_r[154]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(\xs[1].cli1.i[34] ),
    .QN(_02424_));
 DFFHQNx1_ASAP7_75t_R \out_r[155]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(\xs[1].cli1.i[35] ),
    .QN(_02425_));
 DFFHQNx1_ASAP7_75t_R \out_r[156]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(\xs[1].cli1.i[36] ),
    .QN(_02426_));
 DFFHQNx1_ASAP7_75t_R \out_r[159]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(\xs[1].cli1.i[39] ),
    .QN(_02427_));
 DFFHQNx1_ASAP7_75t_R \out_r[160]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\peo[4][0] ),
    .QN(_02428_));
 DFFHQNx1_ASAP7_75t_R \out_r[172]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\peo[4][12] ),
    .QN(_02429_));
 DFFHQNx1_ASAP7_75t_R \out_r[192]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\peo[4][32] ),
    .QN(_02430_));
 DFFHQNx1_ASAP7_75t_R \out_r[193]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\peo[4][33] ),
    .QN(_02431_));
 DFFHQNx1_ASAP7_75t_R \out_r[194]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\peo[4][34] ),
    .QN(_02432_));
 DFFHQNx1_ASAP7_75t_R \out_r[195]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\peo[4][35] ),
    .QN(_02433_));
 DFFHQNx1_ASAP7_75t_R \out_r[196]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\peo[4][36] ),
    .QN(_02434_));
 DFFHQNx1_ASAP7_75t_R \out_r[199]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\peo[4][39] ),
    .QN(_02435_));
 DFFHQNx1_ASAP7_75t_R \out_r[200]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\peo[5][0] ),
    .QN(_02436_));
 DFFHQNx1_ASAP7_75t_R \out_r[212]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\peo[5][10] ),
    .QN(_02437_));
 DFFHQNx1_ASAP7_75t_R \out_r[232]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\xs[2].cli1.i[32] ),
    .QN(_02438_));
 DFFHQNx1_ASAP7_75t_R \out_r[233]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\xs[2].cli1.i[33] ),
    .QN(_02439_));
 DFFHQNx1_ASAP7_75t_R \out_r[234]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\xs[2].cli1.i[34] ),
    .QN(_02440_));
 DFFHQNx1_ASAP7_75t_R \out_r[235]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(\xs[2].cli1.i[35] ),
    .QN(_02441_));
 DFFHQNx1_ASAP7_75t_R \out_r[236]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\xs[2].cli1.i[36] ),
    .QN(_02442_));
 DFFHQNx1_ASAP7_75t_R \out_r[239]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\xs[2].cli1.i[39] ),
    .QN(_02443_));
 DFFHQNx1_ASAP7_75t_R \out_r[240]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(\peo[6][0] ),
    .QN(_02444_));
 DFFHQNx1_ASAP7_75t_R \out_r[252]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(\peo[6][11] ),
    .QN(_02445_));
 DFFHQNx1_ASAP7_75t_R \out_r[272]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(\peo[6][32] ),
    .QN(_02446_));
 DFFHQNx1_ASAP7_75t_R \out_r[273]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(\peo[6][33] ),
    .QN(_02447_));
 DFFHQNx1_ASAP7_75t_R \out_r[274]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(\peo[6][34] ),
    .QN(_02448_));
 DFFHQNx1_ASAP7_75t_R \out_r[275]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(\peo[6][35] ),
    .QN(_02449_));
 DFFHQNx1_ASAP7_75t_R \out_r[276]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(\peo[6][36] ),
    .QN(_02450_));
 DFFHQNx1_ASAP7_75t_R \out_r[279]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(\peo[6][39] ),
    .QN(_02451_));
 DFFHQNx1_ASAP7_75t_R \out_r[280]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(\peo[7][0] ),
    .QN(_02452_));
 DFFHQNx1_ASAP7_75t_R \out_r[292]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(\peo[7][10] ),
    .QN(_02453_));
 DFFHQNx1_ASAP7_75t_R \out_r[312]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(\xs[3].cli1.i[32] ),
    .QN(_02454_));
 DFFHQNx1_ASAP7_75t_R \out_r[313]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(\xs[3].cli1.i[33] ),
    .QN(_02455_));
 DFFHQNx1_ASAP7_75t_R \out_r[314]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(\xs[3].cli1.i[34] ),
    .QN(_02456_));
 DFFHQNx1_ASAP7_75t_R \out_r[315]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(\xs[3].cli1.i[35] ),
    .QN(_02457_));
 DFFHQNx1_ASAP7_75t_R \out_r[316]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(\xs[3].cli1.i[36] ),
    .QN(_02458_));
 DFFHQNx1_ASAP7_75t_R \out_r[319]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(\xs[3].cli1.i[39] ),
    .QN(_02459_));
 DFFHQNx1_ASAP7_75t_R \out_r[320]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .D(\peo[8][0] ),
    .QN(_02460_));
 DFFHQNx1_ASAP7_75t_R \out_r[32]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(\peo[0][32] ),
    .QN(_02461_));
 DFFHQNx1_ASAP7_75t_R \out_r[333]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .D(\peo[8][13] ),
    .QN(_02462_));
 DFFHQNx1_ASAP7_75t_R \out_r[33]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(\peo[0][33] ),
    .QN(_02463_));
 DFFHQNx1_ASAP7_75t_R \out_r[34]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(\peo[0][34] ),
    .QN(_02464_));
 DFFHQNx1_ASAP7_75t_R \out_r[352]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .D(\peo[8][32] ),
    .QN(_02465_));
 DFFHQNx1_ASAP7_75t_R \out_r[353]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .D(\peo[8][33] ),
    .QN(_02466_));
 DFFHQNx1_ASAP7_75t_R \out_r[354]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .D(\peo[8][34] ),
    .QN(_02467_));
 DFFHQNx1_ASAP7_75t_R \out_r[355]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .D(\peo[8][35] ),
    .QN(_02468_));
 DFFHQNx1_ASAP7_75t_R \out_r[356]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .D(\peo[8][36] ),
    .QN(_02469_));
 DFFHQNx1_ASAP7_75t_R \out_r[359]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .D(\peo[8][39] ),
    .QN(_02470_));
 DFFHQNx1_ASAP7_75t_R \out_r[35]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(\peo[0][35] ),
    .QN(_02471_));
 DFFHQNx1_ASAP7_75t_R \out_r[360]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .D(\peo[9][0] ),
    .QN(_02472_));
 DFFHQNx1_ASAP7_75t_R \out_r[36]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(\peo[0][36] ),
    .QN(_02473_));
 DFFHQNx1_ASAP7_75t_R \out_r[373]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .D(\peo[9][10] ),
    .QN(_02474_));
 DFFHQNx1_ASAP7_75t_R \out_r[392]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .D(\xs[4].cli1.i[32] ),
    .QN(_02475_));
 DFFHQNx1_ASAP7_75t_R \out_r[393]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .D(\xs[4].cli1.i[33] ),
    .QN(_02476_));
 DFFHQNx1_ASAP7_75t_R \out_r[394]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .D(\xs[4].cli1.i[34] ),
    .QN(_02477_));
 DFFHQNx1_ASAP7_75t_R \out_r[395]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .D(\xs[4].cli1.i[35] ),
    .QN(_02478_));
 DFFHQNx1_ASAP7_75t_R \out_r[396]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .D(\xs[4].cli1.i[36] ),
    .QN(_02479_));
 DFFHQNx1_ASAP7_75t_R \out_r[399]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .D(\xs[4].cli1.i[39] ),
    .QN(_02480_));
 DFFHQNx1_ASAP7_75t_R \out_r[39]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(\peo[0][39] ),
    .QN(_02481_));
 DFFHQNx1_ASAP7_75t_R \out_r[400]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .D(\peo[10][0] ),
    .QN(_02482_));
 DFFHQNx1_ASAP7_75t_R \out_r[40]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(\peo[1][0] ),
    .QN(_02483_));
 DFFHQNx1_ASAP7_75t_R \out_r[413]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .D(\peo[10][11] ),
    .QN(_02484_));
 DFFHQNx1_ASAP7_75t_R \out_r[432]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .D(\peo[10][32] ),
    .QN(_02485_));
 DFFHQNx1_ASAP7_75t_R \out_r[433]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .D(\peo[10][33] ),
    .QN(_02486_));
 DFFHQNx1_ASAP7_75t_R \out_r[434]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .D(\peo[10][34] ),
    .QN(_02487_));
 DFFHQNx1_ASAP7_75t_R \out_r[435]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .D(\peo[10][35] ),
    .QN(_02488_));
 DFFHQNx1_ASAP7_75t_R \out_r[436]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .D(\peo[10][36] ),
    .QN(_02489_));
 DFFHQNx1_ASAP7_75t_R \out_r[439]$_DFF_P_  (.CLK(clknet_leaf_43_clk),
    .D(\peo[10][39] ),
    .QN(_02490_));
 DFFHQNx1_ASAP7_75t_R \out_r[440]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .D(\peo[11][0] ),
    .QN(_02491_));
 DFFHQNx1_ASAP7_75t_R \out_r[453]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .D(\peo[11][10] ),
    .QN(_02492_));
 DFFHQNx1_ASAP7_75t_R \out_r[472]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .D(\xs[5].cli1.i[32] ),
    .QN(_02493_));
 DFFHQNx1_ASAP7_75t_R \out_r[473]$_DFF_P_  (.CLK(clknet_leaf_43_clk),
    .D(\xs[5].cli1.i[33] ),
    .QN(_02494_));
 DFFHQNx1_ASAP7_75t_R \out_r[474]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .D(\xs[5].cli1.i[34] ),
    .QN(_02495_));
 DFFHQNx1_ASAP7_75t_R \out_r[475]$_DFF_P_  (.CLK(clknet_leaf_43_clk),
    .D(\xs[5].cli1.i[35] ),
    .QN(_02496_));
 DFFHQNx1_ASAP7_75t_R \out_r[476]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .D(\xs[5].cli1.i[36] ),
    .QN(_02497_));
 DFFHQNx1_ASAP7_75t_R \out_r[479]$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .D(\xs[5].cli1.i[39] ),
    .QN(_02498_));
 DFFHQNx1_ASAP7_75t_R \out_r[480]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\peo[12][0] ),
    .QN(_02499_));
 DFFHQNx1_ASAP7_75t_R \out_r[493]$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .D(\peo[12][12] ),
    .QN(_02500_));
 DFFHQNx1_ASAP7_75t_R \out_r[50]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(\peo[1][10] ),
    .QN(_02501_));
 DFFHQNx1_ASAP7_75t_R \out_r[512]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\peo[12][32] ),
    .QN(_02502_));
 DFFHQNx1_ASAP7_75t_R \out_r[513]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\peo[12][33] ),
    .QN(_02503_));
 DFFHQNx1_ASAP7_75t_R \out_r[514]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .D(\peo[12][34] ),
    .QN(_02504_));
 DFFHQNx1_ASAP7_75t_R \out_r[515]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\peo[12][35] ),
    .QN(_02505_));
 DFFHQNx1_ASAP7_75t_R \out_r[516]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\peo[12][36] ),
    .QN(_02506_));
 DFFHQNx1_ASAP7_75t_R \out_r[519]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .D(\peo[12][39] ),
    .QN(_02507_));
 DFFHQNx1_ASAP7_75t_R \out_r[520]$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .D(\peo[13][0] ),
    .QN(_02508_));
 DFFHQNx1_ASAP7_75t_R \out_r[533]$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .D(\peo[13][10] ),
    .QN(_02509_));
 DFFHQNx1_ASAP7_75t_R \out_r[552]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .D(\xs[6].cli1.i[32] ),
    .QN(_02510_));
 DFFHQNx1_ASAP7_75t_R \out_r[553]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .D(\xs[6].cli1.i[33] ),
    .QN(_02511_));
 DFFHQNx1_ASAP7_75t_R \out_r[554]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .D(\xs[6].cli1.i[34] ),
    .QN(_02512_));
 DFFHQNx1_ASAP7_75t_R \out_r[555]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .D(\xs[6].cli1.i[35] ),
    .QN(_02513_));
 DFFHQNx1_ASAP7_75t_R \out_r[556]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .D(\xs[6].cli1.i[36] ),
    .QN(_02514_));
 DFFHQNx1_ASAP7_75t_R \out_r[559]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .D(\xs[6].cli1.i[39] ),
    .QN(_02515_));
 DFFHQNx1_ASAP7_75t_R \out_r[560]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\peo[14][0] ),
    .QN(_02516_));
 DFFHQNx1_ASAP7_75t_R \out_r[573]$_DFF_P_  (.CLK(clknet_leaf_37_clk),
    .D(\peo[14][11] ),
    .QN(_02517_));
 DFFHQNx1_ASAP7_75t_R \out_r[592]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\peo[14][32] ),
    .QN(_02518_));
 DFFHQNx1_ASAP7_75t_R \out_r[593]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\peo[14][33] ),
    .QN(_02519_));
 DFFHQNx1_ASAP7_75t_R \out_r[594]$_DFF_P_  (.CLK(clknet_leaf_37_clk),
    .D(\peo[14][34] ),
    .QN(_02520_));
 DFFHQNx1_ASAP7_75t_R \out_r[595]$_DFF_P_  (.CLK(clknet_leaf_37_clk),
    .D(\peo[14][35] ),
    .QN(_02521_));
 DFFHQNx1_ASAP7_75t_R \out_r[596]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\peo[14][36] ),
    .QN(_02522_));
 DFFHQNx1_ASAP7_75t_R \out_r[599]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\peo[14][39] ),
    .QN(_02523_));
 DFFHQNx1_ASAP7_75t_R \out_r[600]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\peo[15][0] ),
    .QN(_02524_));
 DFFHQNx1_ASAP7_75t_R \out_r[613]$_DFF_P_  (.CLK(clknet_leaf_36_clk),
    .D(\peo[15][10] ),
    .QN(_02525_));
 DFFHQNx1_ASAP7_75t_R \out_r[632]$_DFF_P_  (.CLK(clknet_leaf_36_clk),
    .D(\xs[7].cli1.i[32] ),
    .QN(_02526_));
 DFFHQNx1_ASAP7_75t_R \out_r[633]$_DFF_P_  (.CLK(clknet_leaf_36_clk),
    .D(\xs[7].cli1.i[33] ),
    .QN(_02527_));
 DFFHQNx1_ASAP7_75t_R \out_r[634]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .D(\xs[7].cli1.i[34] ),
    .QN(_02528_));
 DFFHQNx1_ASAP7_75t_R \out_r[635]$_DFF_P_  (.CLK(clknet_leaf_37_clk),
    .D(\xs[7].cli1.i[35] ),
    .QN(_02529_));
 DFFHQNx1_ASAP7_75t_R \out_r[636]$_DFF_P_  (.CLK(clknet_leaf_36_clk),
    .D(\xs[7].cli1.i[36] ),
    .QN(_02530_));
 DFFHQNx1_ASAP7_75t_R \out_r[639]$_DFF_P_  (.CLK(clknet_leaf_37_clk),
    .D(\xs[7].cli1.i[39] ),
    .QN(_02531_));
 DFFHQNx1_ASAP7_75t_R \out_r[640]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\peo[16][0] ),
    .QN(_02532_));
 DFFHQNx1_ASAP7_75t_R \out_r[654]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[16][14] ),
    .QN(_02533_));
 DFFHQNx1_ASAP7_75t_R \out_r[672]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\peo[16][32] ),
    .QN(_02534_));
 DFFHQNx1_ASAP7_75t_R \out_r[673]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\peo[16][33] ),
    .QN(_02535_));
 DFFHQNx1_ASAP7_75t_R \out_r[674]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\peo[16][34] ),
    .QN(_02536_));
 DFFHQNx1_ASAP7_75t_R \out_r[675]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\peo[16][35] ),
    .QN(_02537_));
 DFFHQNx1_ASAP7_75t_R \out_r[676]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\peo[16][36] ),
    .QN(_02538_));
 DFFHQNx1_ASAP7_75t_R \out_r[679]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\peo[16][39] ),
    .QN(_02539_));
 DFFHQNx1_ASAP7_75t_R \out_r[680]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(\peo[17][0] ),
    .QN(_02540_));
 DFFHQNx1_ASAP7_75t_R \out_r[694]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[17][10] ),
    .QN(_02541_));
 DFFHQNx1_ASAP7_75t_R \out_r[712]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\xs[8].cli1.i[32] ),
    .QN(_02542_));
 DFFHQNx1_ASAP7_75t_R \out_r[713]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\xs[8].cli1.i[33] ),
    .QN(_02543_));
 DFFHQNx1_ASAP7_75t_R \out_r[714]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\xs[8].cli1.i[34] ),
    .QN(_02544_));
 DFFHQNx1_ASAP7_75t_R \out_r[715]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\xs[8].cli1.i[35] ),
    .QN(_02545_));
 DFFHQNx1_ASAP7_75t_R \out_r[716]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\xs[8].cli1.i[36] ),
    .QN(_02546_));
 DFFHQNx1_ASAP7_75t_R \out_r[719]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\xs[8].cli1.i[39] ),
    .QN(_02547_));
 DFFHQNx1_ASAP7_75t_R \out_r[720]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[18][0] ),
    .QN(_02548_));
 DFFHQNx1_ASAP7_75t_R \out_r[72]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(\peo[1][32] ),
    .QN(_02549_));
 DFFHQNx1_ASAP7_75t_R \out_r[734]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(\peo[18][11] ),
    .QN(_02550_));
 DFFHQNx1_ASAP7_75t_R \out_r[73]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(\xs[0].cli1.i[33] ),
    .QN(_02551_));
 DFFHQNx1_ASAP7_75t_R \out_r[74]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(\xs[0].cli1.i[34] ),
    .QN(_02552_));
 DFFHQNx1_ASAP7_75t_R \out_r[752]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[18][32] ),
    .QN(_02553_));
 DFFHQNx1_ASAP7_75t_R \out_r[753]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[18][33] ),
    .QN(_02554_));
 DFFHQNx1_ASAP7_75t_R \out_r[754]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[18][34] ),
    .QN(_02555_));
 DFFHQNx1_ASAP7_75t_R \out_r[755]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[18][35] ),
    .QN(_02556_));
 DFFHQNx1_ASAP7_75t_R \out_r[756]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[18][36] ),
    .QN(_02557_));
 DFFHQNx1_ASAP7_75t_R \out_r[759]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[18][39] ),
    .QN(_02558_));
 DFFHQNx1_ASAP7_75t_R \out_r[75]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(\xs[0].cli1.i[35] ),
    .QN(_02559_));
 DFFHQNx1_ASAP7_75t_R \out_r[760]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[19][0] ),
    .QN(_02560_));
 DFFHQNx1_ASAP7_75t_R \out_r[76]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(\xs[0].cli1.i[36] ),
    .QN(_02561_));
 DFFHQNx1_ASAP7_75t_R \out_r[774]$_DFF_P_  (.CLK(clknet_leaf_37_clk),
    .D(\peo[19][10] ),
    .QN(_02562_));
 DFFHQNx1_ASAP7_75t_R \out_r[792]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[19][32] ),
    .QN(_02563_));
 DFFHQNx1_ASAP7_75t_R \out_r[793]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[19][33] ),
    .QN(_02564_));
 DFFHQNx1_ASAP7_75t_R \out_r[794]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[19][34] ),
    .QN(_02565_));
 DFFHQNx1_ASAP7_75t_R \out_r[795]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[19][35] ),
    .QN(_02566_));
 DFFHQNx1_ASAP7_75t_R \out_r[796]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[19][36] ),
    .QN(_02567_));
 DFFHQNx1_ASAP7_75t_R \out_r[799]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(\peo[19][39] ),
    .QN(_02568_));
 DFFHQNx1_ASAP7_75t_R \out_r[79]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(\xs[0].cli1.i[39] ),
    .QN(_02569_));
 DFFHQNx1_ASAP7_75t_R \out_r[800]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(\peo[20][0] ),
    .QN(_02570_));
 DFFHQNx1_ASAP7_75t_R \out_r[80]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(\peo[2][0] ),
    .QN(_02571_));
 DFFHQNx1_ASAP7_75t_R \out_r[814]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\peo[20][12] ),
    .QN(_02572_));
 DFFHQNx1_ASAP7_75t_R \out_r[832]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\peo[20][32] ),
    .QN(_02573_));
 DFFHQNx1_ASAP7_75t_R \out_r[833]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\peo[20][33] ),
    .QN(_02574_));
 DFFHQNx1_ASAP7_75t_R \out_r[834]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\peo[20][34] ),
    .QN(_02575_));
 DFFHQNx1_ASAP7_75t_R \out_r[835]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\peo[20][35] ),
    .QN(_02576_));
 DFFHQNx1_ASAP7_75t_R \out_r[836]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\peo[20][36] ),
    .QN(_02577_));
 DFFHQNx1_ASAP7_75t_R \out_r[839]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(\peo[20][39] ),
    .QN(_02578_));
 DFFHQNx1_ASAP7_75t_R \out_r[840]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(\peo[21][0] ),
    .QN(_02579_));
 DFFHQNx1_ASAP7_75t_R \out_r[854]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(\peo[21][10] ),
    .QN(_02580_));
 DFFHQNx1_ASAP7_75t_R \out_r[872]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\peo[21][32] ),
    .QN(_02581_));
 DFFHQNx1_ASAP7_75t_R \out_r[873]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\xs[10].cli1.i[33] ),
    .QN(_02582_));
 DFFHQNx1_ASAP7_75t_R \out_r[874]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(\xs[10].cli1.i[34] ),
    .QN(_02583_));
 DFFHQNx1_ASAP7_75t_R \out_r[875]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\xs[10].cli1.i[35] ),
    .QN(_02584_));
 DFFHQNx1_ASAP7_75t_R \out_r[876]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(\xs[10].cli1.i[36] ),
    .QN(_02585_));
 DFFHQNx1_ASAP7_75t_R \out_r[879]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(\xs[10].cli1.i[39] ),
    .QN(_02586_));
 DFFHQNx1_ASAP7_75t_R \out_r[880]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(\peo[22][0] ),
    .QN(_02587_));
 DFFHQNx1_ASAP7_75t_R \out_r[894]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(\peo[22][11] ),
    .QN(_02588_));
 DFFHQNx1_ASAP7_75t_R \out_r[912]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(\peo[22][32] ),
    .QN(_02589_));
 DFFHQNx1_ASAP7_75t_R \out_r[913]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(\peo[22][33] ),
    .QN(_02590_));
 DFFHQNx1_ASAP7_75t_R \out_r[914]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(\peo[22][34] ),
    .QN(_02591_));
 DFFHQNx1_ASAP7_75t_R \out_r[915]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(\peo[22][35] ),
    .QN(_02592_));
 DFFHQNx1_ASAP7_75t_R \out_r[916]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(\peo[22][36] ),
    .QN(_02593_));
 DFFHQNx1_ASAP7_75t_R \out_r[919]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(\peo[22][39] ),
    .QN(_02594_));
 DFFHQNx1_ASAP7_75t_R \out_r[91]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(\peo[2][11] ),
    .QN(_02595_));
 DFFHQNx1_ASAP7_75t_R \out_r[920]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(\peo[23][0] ),
    .QN(_02596_));
 DFFHQNx1_ASAP7_75t_R \out_r[934]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(\peo[23][10] ),
    .QN(_02597_));
 DFFHQNx1_ASAP7_75t_R \out_r[952]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(\peo[23][32] ),
    .QN(_02598_));
 DFFHQNx1_ASAP7_75t_R \out_r[953]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(\xs[11].cli1.i[33] ),
    .QN(_02599_));
 DFFHQNx1_ASAP7_75t_R \out_r[954]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(\xs[11].cli1.i[34] ),
    .QN(_02600_));
 DFFHQNx1_ASAP7_75t_R \out_r[955]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(\xs[11].cli1.i[35] ),
    .QN(_02601_));
 DFFHQNx1_ASAP7_75t_R \out_r[956]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(\xs[11].cli1.i[36] ),
    .QN(_02602_));
 DFFHQNx1_ASAP7_75t_R \out_r[959]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(\xs[11].cli1.i[39] ),
    .QN(_02603_));
 DFFHQNx1_ASAP7_75t_R \out_r[960]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(\peo[24][0] ),
    .QN(_02604_));
 DFFHQNx1_ASAP7_75t_R \out_r[974]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(\peo[24][13] ),
    .QN(_02605_));
 DFFHQNx1_ASAP7_75t_R \out_r[992]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(\peo[24][32] ),
    .QN(_02606_));
 DFFHQNx1_ASAP7_75t_R \out_r[993]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\peo[24][33] ),
    .QN(_02607_));
 DFFHQNx1_ASAP7_75t_R \out_r[994]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\peo[24][34] ),
    .QN(_02608_));
 DFFHQNx1_ASAP7_75t_R \out_r[995]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(\peo[24][35] ),
    .QN(_02609_));
 DFFHQNx1_ASAP7_75t_R \out_r[996]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(\peo[24][36] ),
    .QN(_02610_));
 DFFHQNx1_ASAP7_75t_R \out_r[999]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(\peo[24][39] ),
    .QN(_01726_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03306_),
    .QN(_01725_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03307_),
    .QN(_01724_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03308_),
    .QN(_01723_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03309_),
    .QN(_01722_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03310_),
    .QN(_01721_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03311_),
    .QN(_01720_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03312_),
    .QN(_01719_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03313_),
    .QN(_00031_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03314_),
    .QN(_01718_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03315_),
    .QN(_01717_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03316_),
    .QN(_01716_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03317_),
    .QN(_01715_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03318_),
    .QN(_01714_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03319_),
    .QN(_01713_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03320_),
    .QN(_01712_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03321_),
    .QN(_01711_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03322_),
    .QN(_01710_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03323_),
    .QN(_01709_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03324_),
    .QN(_01708_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03325_),
    .QN(_01707_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03326_),
    .QN(_01706_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03327_),
    .QN(_01705_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03328_),
    .QN(_01704_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03329_),
    .QN(_01703_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03330_),
    .QN(_01702_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03331_),
    .QN(_01701_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03332_),
    .QN(_01700_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03333_),
    .QN(_01699_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03334_),
    .QN(_01698_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03335_),
    .QN(_01697_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03336_),
    .QN(_01696_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03337_),
    .QN(_01695_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03338_),
    .QN(_01694_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03339_),
    .QN(_01693_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03340_),
    .QN(_01692_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03341_),
    .QN(_01691_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03342_),
    .QN(_01690_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03343_),
    .QN(_01689_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03344_),
    .QN(_01688_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03345_),
    .QN(_01687_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli1.i[10]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03346_),
    .QN(_01686_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03347_),
    .QN(_01685_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03348_),
    .QN(_01684_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03349_),
    .QN(_01683_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03350_),
    .QN(_01682_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03351_),
    .QN(_01681_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03352_),
    .QN(_01680_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_03353_),
    .QN(_00032_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03354_),
    .QN(_01679_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03355_),
    .QN(_01678_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03356_),
    .QN(_01677_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03357_),
    .QN(_01676_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03358_),
    .QN(_01675_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03359_),
    .QN(_01674_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03360_),
    .QN(_01673_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03361_),
    .QN(_01672_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03362_),
    .QN(_01671_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03363_),
    .QN(_01670_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_03364_),
    .QN(_01669_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03365_),
    .QN(_01668_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03366_),
    .QN(_01667_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03367_),
    .QN(_01666_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03368_),
    .QN(_01665_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03369_),
    .QN(_01664_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03370_),
    .QN(_01663_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03371_),
    .QN(_01662_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03372_),
    .QN(_01661_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03373_),
    .QN(_01660_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_03374_),
    .QN(_01659_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_03375_),
    .QN(_01658_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_03376_),
    .QN(_01657_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03377_),
    .QN(_01656_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_03378_),
    .QN(_01655_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_03379_),
    .QN(_01654_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_03380_),
    .QN(_01653_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_03381_),
    .QN(_01652_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03382_),
    .QN(_01651_));
 DFFHQNx3_ASAP7_75t_R \xs[0].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03383_),
    .QN(_01650_));
 DFFHQNx1_ASAP7_75t_R \xs[0].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_03384_),
    .QN(_01649_));
 DFFHQNx3_ASAP7_75t_R \xs[0].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_03385_),
    .QN(_00015_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03386_),
    .QN(_01648_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03387_),
    .QN(_01647_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03388_),
    .QN(_01646_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03389_),
    .QN(_01645_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03390_),
    .QN(_01644_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03391_),
    .QN(_01643_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03392_),
    .QN(_01642_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03393_),
    .QN(_01641_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03394_),
    .QN(_01640_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03395_),
    .QN(_01639_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03396_),
    .QN(_01638_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03397_),
    .QN(_01637_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_03398_),
    .QN(_01636_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_03399_),
    .QN(_01635_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_03400_),
    .QN(_01634_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_03401_),
    .QN(_01633_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03402_),
    .QN(_01632_));
 DFFHQNx3_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03403_),
    .QN(_01631_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03404_),
    .QN(_01630_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03405_),
    .QN(_01629_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03406_),
    .QN(_01628_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03407_),
    .QN(_01627_));
 DFFHQNx3_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03408_),
    .QN(_01626_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_03409_),
    .QN(_01625_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_03410_),
    .QN(_01624_));
 DFFHQNx1_ASAP7_75t_R \xs[0].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_03411_),
    .QN(_01623_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03412_),
    .QN(_01622_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli0.i[12]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03413_),
    .QN(_01621_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03414_),
    .QN(_01620_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03415_),
    .QN(_01619_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03416_),
    .QN(_01618_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03417_),
    .QN(_01617_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03418_),
    .QN(_01616_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03419_),
    .QN(_01615_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03420_),
    .QN(_00033_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03421_),
    .QN(_01614_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03422_),
    .QN(_01613_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03423_),
    .QN(_01612_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03424_),
    .QN(_01611_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03425_),
    .QN(_01610_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03426_),
    .QN(_01609_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03427_),
    .QN(_01608_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03428_),
    .QN(_01607_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03429_),
    .QN(_01606_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03430_),
    .QN(_01605_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03431_),
    .QN(_01604_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03432_),
    .QN(_01603_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03433_),
    .QN(_01602_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03434_),
    .QN(_01601_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03435_),
    .QN(_01600_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03436_),
    .QN(_01599_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03437_),
    .QN(_01598_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03438_),
    .QN(_01597_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03439_),
    .QN(_01596_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03440_),
    .QN(_01595_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03441_),
    .QN(_01594_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03442_),
    .QN(_01593_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03443_),
    .QN(_01592_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03444_),
    .QN(_01591_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03445_),
    .QN(_01590_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03446_),
    .QN(_01589_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03447_),
    .QN(_01588_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03448_),
    .QN(_01587_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03449_),
    .QN(_01586_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03450_),
    .QN(_01585_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03451_),
    .QN(_01584_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03452_),
    .QN(_01583_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli1.i[12]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03453_),
    .QN(_01582_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03454_),
    .QN(_01581_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03455_),
    .QN(_01580_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03456_),
    .QN(_01579_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03457_),
    .QN(_01578_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03458_),
    .QN(_01577_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03459_),
    .QN(_01576_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03460_),
    .QN(_00034_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03461_),
    .QN(_01575_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03462_),
    .QN(_01574_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03463_),
    .QN(_01573_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03464_),
    .QN(_01572_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03465_),
    .QN(_01571_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03466_),
    .QN(_01570_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03467_),
    .QN(_01569_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03468_),
    .QN(_01568_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03469_),
    .QN(_01567_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03470_),
    .QN(_01566_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03471_),
    .QN(_01565_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03472_),
    .QN(_01564_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03473_),
    .QN(_01563_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03474_),
    .QN(_01562_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03475_),
    .QN(_01561_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03476_),
    .QN(_01560_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03477_),
    .QN(_01559_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03478_),
    .QN(_01558_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03479_),
    .QN(_01557_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03480_),
    .QN(_01556_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03481_),
    .QN(_01555_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03482_),
    .QN(_01554_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03483_),
    .QN(_01553_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03484_),
    .QN(_01552_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03485_),
    .QN(_01551_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03486_),
    .QN(_01550_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03487_),
    .QN(_01549_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03488_),
    .QN(_01548_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03489_),
    .QN(_01547_));
 DFFHQNx3_ASAP7_75t_R \xs[10].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .D(_03490_),
    .QN(_01546_));
 DFFHQNx1_ASAP7_75t_R \xs[10].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03491_),
    .QN(_01545_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03492_),
    .QN(_00016_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03493_),
    .QN(_01544_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03494_),
    .QN(_01543_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03495_),
    .QN(_01542_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03496_),
    .QN(_01541_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03497_),
    .QN(_01540_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03498_),
    .QN(_01539_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03499_),
    .QN(_01538_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03500_),
    .QN(_01537_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03501_),
    .QN(_01536_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03502_),
    .QN(_01535_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03503_),
    .QN(_01534_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03504_),
    .QN(_01533_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03505_),
    .QN(_01532_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03506_),
    .QN(_01531_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03507_),
    .QN(_01530_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03508_),
    .QN(_01529_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03509_),
    .QN(_01528_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03510_),
    .QN(_01527_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03511_),
    .QN(_01526_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03512_),
    .QN(_01525_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03513_),
    .QN(_01524_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03514_),
    .QN(_01523_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03515_),
    .QN(_01522_));
 DFFHQNx1_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03516_),
    .QN(_01521_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03517_),
    .QN(_01520_));
 DFFHQNx3_ASAP7_75t_R \xs[10].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03518_),
    .QN(_01519_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03519_),
    .QN(_01518_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli0.i[12]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03520_),
    .QN(_01517_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03521_),
    .QN(_01516_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03522_),
    .QN(_01515_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03523_),
    .QN(_01514_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03524_),
    .QN(_01513_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03525_),
    .QN(_01512_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03526_),
    .QN(_01511_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03527_),
    .QN(_00035_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03528_),
    .QN(_01510_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03529_),
    .QN(_01509_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03530_),
    .QN(_01508_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03531_),
    .QN(_01507_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03532_),
    .QN(_01506_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03533_),
    .QN(_01505_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03534_),
    .QN(_01504_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03535_),
    .QN(_01503_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03536_),
    .QN(_01502_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03537_),
    .QN(_01501_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03538_),
    .QN(_01500_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03539_),
    .QN(_01499_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03540_),
    .QN(_01498_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03541_),
    .QN(_01497_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03542_),
    .QN(_01496_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03543_),
    .QN(_01495_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03544_),
    .QN(_01494_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03545_),
    .QN(_01493_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03546_),
    .QN(_01492_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03547_),
    .QN(_01491_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03548_),
    .QN(_01490_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03549_),
    .QN(_01489_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03550_),
    .QN(_01488_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03551_),
    .QN(_01487_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03552_),
    .QN(_01486_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03553_),
    .QN(_01485_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03554_),
    .QN(_01484_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03555_),
    .QN(_01483_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03556_),
    .QN(_01482_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03557_),
    .QN(_01481_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03558_),
    .QN(_01480_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03559_),
    .QN(_01479_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli1.i[12]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03560_),
    .QN(_01478_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03561_),
    .QN(_01477_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03562_),
    .QN(_01476_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03563_),
    .QN(_01475_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03564_),
    .QN(_01474_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03565_),
    .QN(_01473_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03566_),
    .QN(_01472_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03567_),
    .QN(_00036_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03568_),
    .QN(_01471_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03569_),
    .QN(_01470_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03570_),
    .QN(_01469_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03571_),
    .QN(_01468_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03572_),
    .QN(_01467_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03573_),
    .QN(_01466_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .D(_03574_),
    .QN(_01465_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03575_),
    .QN(_01464_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03576_),
    .QN(_01463_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03577_),
    .QN(_01462_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03578_),
    .QN(_01461_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03579_),
    .QN(_01460_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03580_),
    .QN(_01459_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03581_),
    .QN(_01458_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03582_),
    .QN(_01457_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03583_),
    .QN(_01456_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03584_),
    .QN(_01455_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03585_),
    .QN(_01454_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03586_),
    .QN(_01453_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03587_),
    .QN(_01452_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03588_),
    .QN(_01451_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03589_),
    .QN(_01450_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03590_),
    .QN(_01449_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03591_),
    .QN(_01448_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03592_),
    .QN(_01447_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03593_),
    .QN(_01446_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03594_),
    .QN(_01445_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03595_),
    .QN(_01444_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03596_),
    .QN(_01443_));
 DFFHQNx3_ASAP7_75t_R \xs[11].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03597_),
    .QN(_01442_));
 DFFHQNx1_ASAP7_75t_R \xs[11].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03598_),
    .QN(_01441_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03599_),
    .QN(_00017_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03600_),
    .QN(_01440_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03601_),
    .QN(_01439_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03602_),
    .QN(_01438_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03603_),
    .QN(_01437_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03604_),
    .QN(_01436_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03605_),
    .QN(_01435_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03606_),
    .QN(_01434_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03607_),
    .QN(_01433_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03608_),
    .QN(_01432_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03609_),
    .QN(_01431_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03610_),
    .QN(_01430_));
 DFFHQNx1_ASAP7_75t_R \xs[11].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03611_),
    .QN(_01429_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03612_),
    .QN(_01428_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03613_),
    .QN(_01427_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03614_),
    .QN(_01426_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03615_),
    .QN(_01425_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03616_),
    .QN(_01424_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03617_),
    .QN(_01423_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03618_),
    .QN(_01422_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03619_),
    .QN(_01421_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03620_),
    .QN(_01420_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03621_),
    .QN(_01419_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03622_),
    .QN(_01418_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03623_),
    .QN(_01417_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03624_),
    .QN(_01416_));
 DFFHQNx3_ASAP7_75t_R \xs[11].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03625_),
    .QN(_01415_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .D(_03626_),
    .QN(_01414_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli0.i[13]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03627_),
    .QN(_01413_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_03628_),
    .QN(_01412_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03629_),
    .QN(_01411_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03630_),
    .QN(_01410_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03631_),
    .QN(_01409_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03632_),
    .QN(_01408_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03633_),
    .QN(_01407_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03634_),
    .QN(_00037_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03635_),
    .QN(_01406_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03636_),
    .QN(_01405_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03637_),
    .QN(_01404_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03638_),
    .QN(_01403_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03639_),
    .QN(_01402_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03640_),
    .QN(_01401_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03641_),
    .QN(_01400_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03642_),
    .QN(_01399_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03643_),
    .QN(_01398_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03644_),
    .QN(_01397_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03645_),
    .QN(_01396_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03646_),
    .QN(_01395_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03647_),
    .QN(_01394_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03648_),
    .QN(_01393_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03649_),
    .QN(_01392_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03650_),
    .QN(_01391_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03651_),
    .QN(_01390_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03652_),
    .QN(_01389_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03653_),
    .QN(_01388_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03654_),
    .QN(_01387_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03655_),
    .QN(_01386_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03656_),
    .QN(_01385_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03657_),
    .QN(_01384_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03658_),
    .QN(_01383_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03659_),
    .QN(_01382_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03660_),
    .QN(_01381_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03661_),
    .QN(_01380_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03662_),
    .QN(_01379_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03663_),
    .QN(_01378_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03664_),
    .QN(_01377_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .D(_03665_),
    .QN(_01376_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03666_),
    .QN(_01375_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli1.i[13]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03667_),
    .QN(_01374_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03668_),
    .QN(_01373_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03669_),
    .QN(_01372_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03670_),
    .QN(_01371_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03671_),
    .QN(_01370_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03672_),
    .QN(_01369_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03673_),
    .QN(_01368_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03674_),
    .QN(_00038_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03675_),
    .QN(_01367_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03676_),
    .QN(_01366_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .D(_03677_),
    .QN(_01365_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03678_),
    .QN(_01364_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03679_),
    .QN(_01363_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03680_),
    .QN(_01362_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03681_),
    .QN(_01361_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03682_),
    .QN(_01360_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03683_),
    .QN(_01359_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03684_),
    .QN(_01358_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03685_),
    .QN(_01357_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03686_),
    .QN(_01356_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03687_),
    .QN(_01355_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03688_),
    .QN(_01354_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03689_),
    .QN(_01353_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03690_),
    .QN(_01352_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03691_),
    .QN(_01351_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03692_),
    .QN(_01350_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03693_),
    .QN(_01349_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03694_),
    .QN(_01348_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03695_),
    .QN(_01347_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03696_),
    .QN(_01346_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03697_),
    .QN(_01345_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03698_),
    .QN(_01344_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03699_),
    .QN(_01343_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03700_),
    .QN(_01342_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03701_),
    .QN(_01341_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03702_),
    .QN(_01340_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03703_),
    .QN(_01339_));
 DFFHQNx3_ASAP7_75t_R \xs[12].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03704_),
    .QN(_01338_));
 DFFHQNx1_ASAP7_75t_R \xs[12].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03705_),
    .QN(_01337_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03706_),
    .QN(_00018_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03707_),
    .QN(_01336_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03708_),
    .QN(_01335_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03709_),
    .QN(_01334_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03710_),
    .QN(_01333_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03711_),
    .QN(_01332_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03712_),
    .QN(_01331_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03713_),
    .QN(_01330_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03714_),
    .QN(_01329_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03715_),
    .QN(_01328_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03716_),
    .QN(_01327_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03717_),
    .QN(_01326_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03718_),
    .QN(_01325_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03719_),
    .QN(_01324_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03720_),
    .QN(_01323_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03721_),
    .QN(_01322_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .D(_03722_),
    .QN(_01321_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03723_),
    .QN(_01320_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03724_),
    .QN(_01319_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03725_),
    .QN(_01318_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03726_),
    .QN(_01317_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03727_),
    .QN(_01316_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03728_),
    .QN(_01315_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03729_),
    .QN(_01314_));
 DFFHQNx1_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .D(_03730_),
    .QN(_01313_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03731_),
    .QN(_01312_));
 DFFHQNx3_ASAP7_75t_R \xs[12].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_03732_),
    .QN(_01311_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03733_),
    .QN(_01310_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli0.i[13]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03734_),
    .QN(_01309_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_03735_),
    .QN(_01308_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03736_),
    .QN(_01307_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03737_),
    .QN(_01306_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03738_),
    .QN(_01305_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03739_),
    .QN(_01304_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_03740_),
    .QN(_01303_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03741_),
    .QN(_00039_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03742_),
    .QN(_01302_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03743_),
    .QN(_01301_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03744_),
    .QN(_01300_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03745_),
    .QN(_01299_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03746_),
    .QN(_01298_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03747_),
    .QN(_01297_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03748_),
    .QN(_01296_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03749_),
    .QN(_01295_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03750_),
    .QN(_01294_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03751_),
    .QN(_01293_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03752_),
    .QN(_01292_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03753_),
    .QN(_01291_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03754_),
    .QN(_01290_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03755_),
    .QN(_01289_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03756_),
    .QN(_01288_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03757_),
    .QN(_01287_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03758_),
    .QN(_01286_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03759_),
    .QN(_01285_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03760_),
    .QN(_01284_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03761_),
    .QN(_01283_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03762_),
    .QN(_01282_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03763_),
    .QN(_01281_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03764_),
    .QN(_01280_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03765_),
    .QN(_01279_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03766_),
    .QN(_01278_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03767_),
    .QN(_01277_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03768_),
    .QN(_01276_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03769_),
    .QN(_01275_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .D(_03770_),
    .QN(_01274_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03771_),
    .QN(_01273_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .D(_03772_),
    .QN(_01272_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03773_),
    .QN(_01271_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli1.i[13]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_03774_),
    .QN(_01270_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03775_),
    .QN(_01269_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03776_),
    .QN(_01268_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03777_),
    .QN(_01267_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03778_),
    .QN(_01266_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03779_),
    .QN(_01265_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03780_),
    .QN(_01264_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03781_),
    .QN(_00040_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03782_),
    .QN(_01263_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03783_),
    .QN(_01262_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03784_),
    .QN(_01261_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03785_),
    .QN(_01260_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03786_),
    .QN(_01259_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03787_),
    .QN(_01258_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03788_),
    .QN(_01257_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03789_),
    .QN(_01256_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03790_),
    .QN(_01255_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03791_),
    .QN(_01254_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .D(_03792_),
    .QN(_01253_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .D(_03793_),
    .QN(_01252_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03794_),
    .QN(_01251_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03795_),
    .QN(_01250_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03796_),
    .QN(_01249_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03797_),
    .QN(_01248_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03798_),
    .QN(_01247_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03799_),
    .QN(_01246_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03800_),
    .QN(_01245_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03801_),
    .QN(_01244_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03802_),
    .QN(_01243_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03803_),
    .QN(_01242_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03804_),
    .QN(_01241_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03805_),
    .QN(_01240_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03806_),
    .QN(_01239_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03807_),
    .QN(_01238_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03808_),
    .QN(_01237_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03809_),
    .QN(_01236_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03810_),
    .QN(_01235_));
 DFFHQNx3_ASAP7_75t_R \xs[13].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03811_),
    .QN(_01234_));
 DFFHQNx1_ASAP7_75t_R \xs[13].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .D(_03812_),
    .QN(_01233_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .D(_03813_),
    .QN(_00019_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_03814_),
    .QN(_01232_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03815_),
    .QN(_01231_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03816_),
    .QN(_01230_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03817_),
    .QN(_01229_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03818_),
    .QN(_01228_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03819_),
    .QN(_01227_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03820_),
    .QN(_01226_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03821_),
    .QN(_01225_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03822_),
    .QN(_01224_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03823_),
    .QN(_01223_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03824_),
    .QN(_01222_));
 DFFHQNx1_ASAP7_75t_R \xs[13].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03825_),
    .QN(_01221_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03826_),
    .QN(_01220_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03827_),
    .QN(_01219_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03828_),
    .QN(_01218_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_03829_),
    .QN(_01217_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03830_),
    .QN(_01216_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03831_),
    .QN(_01215_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03832_),
    .QN(_01214_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_03833_),
    .QN(_01213_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03834_),
    .QN(_01212_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03835_),
    .QN(_01211_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_03836_),
    .QN(_01210_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03837_),
    .QN(_01209_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03838_),
    .QN(_01208_));
 DFFHQNx3_ASAP7_75t_R \xs[13].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_03839_),
    .QN(_01207_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03840_),
    .QN(_01206_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli0.i[13]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03841_),
    .QN(_01205_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03842_),
    .QN(_01204_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03843_),
    .QN(_01203_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03844_),
    .QN(_01202_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03845_),
    .QN(_01201_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03846_),
    .QN(_01200_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03847_),
    .QN(_01199_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03848_),
    .QN(_00041_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03849_),
    .QN(_01198_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03850_),
    .QN(_01197_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03851_),
    .QN(_01196_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03852_),
    .QN(_01195_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03853_),
    .QN(_01194_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03854_),
    .QN(_01193_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03855_),
    .QN(_01192_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .D(_03856_),
    .QN(_01191_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03857_),
    .QN(_01190_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .D(_03858_),
    .QN(_01189_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03859_),
    .QN(_01188_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03860_),
    .QN(_01187_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03861_),
    .QN(_01186_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03862_),
    .QN(_01185_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03863_),
    .QN(_01184_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03864_),
    .QN(_01183_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03865_),
    .QN(_01182_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03866_),
    .QN(_01181_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03867_),
    .QN(_01180_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03868_),
    .QN(_01179_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03869_),
    .QN(_01178_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03870_),
    .QN(_01177_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03871_),
    .QN(_01176_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03872_),
    .QN(_01175_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03873_),
    .QN(_01174_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03874_),
    .QN(_01173_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03875_),
    .QN(_01172_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03876_),
    .QN(_01171_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03877_),
    .QN(_01170_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03878_),
    .QN(_01169_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03879_),
    .QN(_01168_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03880_),
    .QN(_01167_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli1.i[13]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_03881_),
    .QN(_01166_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03882_),
    .QN(_01165_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03883_),
    .QN(_01164_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03884_),
    .QN(_01163_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03885_),
    .QN(_01162_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03886_),
    .QN(_01161_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03887_),
    .QN(_01160_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03888_),
    .QN(_00042_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03889_),
    .QN(_01159_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03890_),
    .QN(_01158_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03891_),
    .QN(_01157_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_03892_),
    .QN(_01156_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_03893_),
    .QN(_01155_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03894_),
    .QN(_01154_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_03895_),
    .QN(_01153_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_03896_),
    .QN(_01152_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_03897_),
    .QN(_01151_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03898_),
    .QN(_01150_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03899_),
    .QN(_01149_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03900_),
    .QN(_01148_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_03901_),
    .QN(_01147_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_03902_),
    .QN(_01146_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_03903_),
    .QN(_01145_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03904_),
    .QN(_01144_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_03905_),
    .QN(_01143_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03906_),
    .QN(_01142_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03907_),
    .QN(_01141_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03908_),
    .QN(_01140_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_03909_),
    .QN(_01139_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03910_),
    .QN(_01138_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03911_),
    .QN(_01137_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03912_),
    .QN(_01136_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03913_),
    .QN(_01135_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_03914_),
    .QN(_01134_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03915_),
    .QN(_01133_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03916_),
    .QN(_01132_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03917_),
    .QN(_01131_));
 DFFHQNx3_ASAP7_75t_R \xs[14].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03918_),
    .QN(_01130_));
 DFFHQNx1_ASAP7_75t_R \xs[14].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03919_),
    .QN(_01129_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_03920_),
    .QN(_00020_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03921_),
    .QN(_01128_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03922_),
    .QN(_01127_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03923_),
    .QN(_01126_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03924_),
    .QN(_01125_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03925_),
    .QN(_01124_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03926_),
    .QN(_01123_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03927_),
    .QN(_01122_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03928_),
    .QN(_01121_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03929_),
    .QN(_01120_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03930_),
    .QN(_01119_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03931_),
    .QN(_01118_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03932_),
    .QN(_01117_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03933_),
    .QN(_01116_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03934_),
    .QN(_01115_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03935_),
    .QN(_01114_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03936_),
    .QN(_01113_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03937_),
    .QN(_01112_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03938_),
    .QN(_01111_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03939_),
    .QN(_01110_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_03940_),
    .QN(_01109_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03941_),
    .QN(_01108_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03942_),
    .QN(_01107_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03943_),
    .QN(_01106_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03944_),
    .QN(_01105_));
 DFFHQNx3_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03945_),
    .QN(_01104_));
 DFFHQNx1_ASAP7_75t_R \xs[14].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_03946_),
    .QN(_01103_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03947_),
    .QN(_01102_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli0.i[13]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_03948_),
    .QN(_01101_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_03949_),
    .QN(_01100_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_03950_),
    .QN(_01099_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_03951_),
    .QN(_01098_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_03952_),
    .QN(_01097_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_03953_),
    .QN(_01096_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_03954_),
    .QN(_01095_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03955_),
    .QN(_00043_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03956_),
    .QN(_01094_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03957_),
    .QN(_01093_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03958_),
    .QN(_01092_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03959_),
    .QN(_01091_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03960_),
    .QN(_01090_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03961_),
    .QN(_01089_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03962_),
    .QN(_01088_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03963_),
    .QN(_01087_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03964_),
    .QN(_01086_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03965_),
    .QN(_01085_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03966_),
    .QN(_01084_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03967_),
    .QN(_01083_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03968_),
    .QN(_01082_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03969_),
    .QN(_01081_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03970_),
    .QN(_01080_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03971_),
    .QN(_01079_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03972_),
    .QN(_01078_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03973_),
    .QN(_01077_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03974_),
    .QN(_01076_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03975_),
    .QN(_01075_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03976_),
    .QN(_01074_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03977_),
    .QN(_01073_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03978_),
    .QN(_01072_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03979_),
    .QN(_01071_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03980_),
    .QN(_01070_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03981_),
    .QN(_01069_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03982_),
    .QN(_01068_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03983_),
    .QN(_01067_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03984_),
    .QN(_01066_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03985_),
    .QN(_01065_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_03986_),
    .QN(_01064_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_03987_),
    .QN(_01063_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli1.i[13]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_03988_),
    .QN(_01062_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03989_),
    .QN(_01061_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_03990_),
    .QN(_01060_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_03991_),
    .QN(_01059_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_03992_),
    .QN(_01058_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_03993_),
    .QN(_01057_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_03994_),
    .QN(_01056_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03995_),
    .QN(_00044_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03996_),
    .QN(_01055_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03997_),
    .QN(_01054_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03998_),
    .QN(_01053_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_03999_),
    .QN(_01052_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04000_),
    .QN(_01051_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04001_),
    .QN(_01050_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04002_),
    .QN(_01049_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04003_),
    .QN(_01048_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04004_),
    .QN(_01047_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04005_),
    .QN(_01046_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04006_),
    .QN(_01045_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04007_),
    .QN(_01044_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04008_),
    .QN(_01043_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04009_),
    .QN(_01042_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04010_),
    .QN(_01041_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04011_),
    .QN(_01040_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04012_),
    .QN(_01039_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04013_),
    .QN(_01038_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04014_),
    .QN(_01037_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04015_),
    .QN(_01036_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04016_),
    .QN(_01035_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04017_),
    .QN(_01034_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04018_),
    .QN(_01033_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04019_),
    .QN(_01032_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04020_),
    .QN(_01031_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04021_),
    .QN(_01030_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04022_),
    .QN(_01029_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04023_),
    .QN(_01028_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04024_),
    .QN(_01027_));
 DFFHQNx3_ASAP7_75t_R \xs[15].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04025_),
    .QN(_01026_));
 DFFHQNx1_ASAP7_75t_R \xs[15].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04026_),
    .QN(_01025_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04027_),
    .QN(_00021_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04028_),
    .QN(_01024_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04029_),
    .QN(_01023_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04030_),
    .QN(_01022_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04031_),
    .QN(_01021_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04032_),
    .QN(_01020_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04033_),
    .QN(_01019_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04034_),
    .QN(_01018_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04035_),
    .QN(_01017_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04036_),
    .QN(_01016_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04037_),
    .QN(_01015_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04038_),
    .QN(_01014_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04039_),
    .QN(_01013_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04040_),
    .QN(_01012_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04041_),
    .QN(_01011_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04042_),
    .QN(_01010_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04043_),
    .QN(_01009_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04044_),
    .QN(_01008_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_04045_),
    .QN(_01007_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04046_),
    .QN(_01006_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_04047_),
    .QN(_01005_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_04048_),
    .QN(_01004_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_04049_),
    .QN(_01003_));
 DFFHQNx1_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04050_),
    .QN(_01002_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04051_),
    .QN(_01001_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04052_),
    .QN(_01000_));
 DFFHQNx3_ASAP7_75t_R \xs[15].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04053_),
    .QN(_00999_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04054_),
    .QN(_00998_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli0.i[11]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04055_),
    .QN(_00997_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04056_),
    .QN(_00996_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04057_),
    .QN(_00995_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04058_),
    .QN(_00994_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04059_),
    .QN(_00993_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04060_),
    .QN(_00992_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04061_),
    .QN(_00991_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04062_),
    .QN(_00045_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04063_),
    .QN(_00990_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04064_),
    .QN(_00989_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04065_),
    .QN(_00988_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04066_),
    .QN(_00987_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04067_),
    .QN(_00986_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04068_),
    .QN(_00985_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04069_),
    .QN(_00984_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04070_),
    .QN(_00983_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04071_),
    .QN(_00982_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04072_),
    .QN(_00981_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04073_),
    .QN(_00980_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04074_),
    .QN(_00979_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04075_),
    .QN(_00978_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04076_),
    .QN(_00977_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04077_),
    .QN(_00976_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04078_),
    .QN(_00975_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04079_),
    .QN(_00974_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04080_),
    .QN(_00973_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04081_),
    .QN(_00972_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04082_),
    .QN(_00971_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04083_),
    .QN(_00970_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04084_),
    .QN(_00969_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04085_),
    .QN(_00968_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04086_),
    .QN(_00967_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04087_),
    .QN(_00966_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04088_),
    .QN(_00965_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04089_),
    .QN(_00964_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04090_),
    .QN(_00963_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04091_),
    .QN(_00962_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04092_),
    .QN(_00961_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04093_),
    .QN(_00960_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04094_),
    .QN(_00959_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli1.i[10]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04095_),
    .QN(_00958_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04096_),
    .QN(_00957_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04097_),
    .QN(_00956_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04098_),
    .QN(_00955_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04099_),
    .QN(_00954_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04100_),
    .QN(_00953_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04101_),
    .QN(_00952_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04102_),
    .QN(_00046_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04103_),
    .QN(_00951_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04104_),
    .QN(_00950_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04105_),
    .QN(_00949_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04106_),
    .QN(_00948_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04107_),
    .QN(_00947_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04108_),
    .QN(_00946_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04109_),
    .QN(_00945_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04110_),
    .QN(_00944_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04111_),
    .QN(_00943_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04112_),
    .QN(_00942_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04113_),
    .QN(_00941_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04114_),
    .QN(_00940_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04115_),
    .QN(_00939_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04116_),
    .QN(_00938_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04117_),
    .QN(_00937_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04118_),
    .QN(_00936_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04119_),
    .QN(_00935_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04120_),
    .QN(_00934_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04121_),
    .QN(_00933_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04122_),
    .QN(_00932_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04123_),
    .QN(_00931_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04124_),
    .QN(_00930_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04125_),
    .QN(_00929_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04126_),
    .QN(_00928_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04127_),
    .QN(_00927_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04128_),
    .QN(_00926_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04129_),
    .QN(_00925_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04130_),
    .QN(_00924_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04131_),
    .QN(_00923_));
 DFFHQNx3_ASAP7_75t_R \xs[1].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04132_),
    .QN(_00922_));
 DFFHQNx1_ASAP7_75t_R \xs[1].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04133_),
    .QN(_00921_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04134_),
    .QN(_00022_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04135_),
    .QN(_00920_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04136_),
    .QN(_00919_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04137_),
    .QN(_00918_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04138_),
    .QN(_00917_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04139_),
    .QN(_00916_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04140_),
    .QN(_00915_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04141_),
    .QN(_00914_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04142_),
    .QN(_00913_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04143_),
    .QN(_00912_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04144_),
    .QN(_00911_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04145_),
    .QN(_00910_));
 DFFHQNx1_ASAP7_75t_R \xs[1].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .D(_04146_),
    .QN(_00909_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04147_),
    .QN(_00908_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04148_),
    .QN(_00907_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04149_),
    .QN(_00906_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04150_),
    .QN(_00905_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04151_),
    .QN(_00904_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04152_),
    .QN(_00903_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_04153_),
    .QN(_00902_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04154_),
    .QN(_00901_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .D(_04155_),
    .QN(_00900_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_04156_),
    .QN(_00899_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_04157_),
    .QN(_00898_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .D(_04158_),
    .QN(_00897_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04159_),
    .QN(_00896_));
 DFFHQNx3_ASAP7_75t_R \xs[1].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_04160_),
    .QN(_00895_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04161_),
    .QN(_00894_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli0.i[12]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04162_),
    .QN(_00893_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04163_),
    .QN(_00892_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04164_),
    .QN(_00891_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04165_),
    .QN(_00890_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04166_),
    .QN(_00889_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04167_),
    .QN(_00888_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04168_),
    .QN(_00887_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04169_),
    .QN(_00047_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04170_),
    .QN(_00886_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04171_),
    .QN(_00885_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04172_),
    .QN(_00884_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04173_),
    .QN(_00883_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04174_),
    .QN(_00882_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04175_),
    .QN(_00881_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04176_),
    .QN(_00880_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04177_),
    .QN(_00879_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04178_),
    .QN(_00878_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04179_),
    .QN(_00877_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04180_),
    .QN(_00876_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04181_),
    .QN(_00875_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04182_),
    .QN(_00874_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04183_),
    .QN(_00873_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04184_),
    .QN(_00872_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04185_),
    .QN(_00871_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04186_),
    .QN(_00870_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04187_),
    .QN(_00869_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04188_),
    .QN(_00868_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04189_),
    .QN(_00867_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04190_),
    .QN(_00866_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04191_),
    .QN(_00865_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04192_),
    .QN(_00864_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04193_),
    .QN(_00863_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04194_),
    .QN(_00862_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04195_),
    .QN(_00861_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04196_),
    .QN(_00860_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04197_),
    .QN(_00859_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04198_),
    .QN(_00858_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .D(_04199_),
    .QN(_00857_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04200_),
    .QN(_00856_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04201_),
    .QN(_00855_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli1.i[10]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04202_),
    .QN(_00854_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04203_),
    .QN(_00853_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04204_),
    .QN(_00852_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04205_),
    .QN(_00851_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04206_),
    .QN(_00850_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04207_),
    .QN(_00849_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04208_),
    .QN(_00848_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04209_),
    .QN(_00048_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04210_),
    .QN(_00847_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04211_),
    .QN(_00846_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04212_),
    .QN(_00845_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04213_),
    .QN(_00844_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04214_),
    .QN(_00843_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04215_),
    .QN(_00842_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04216_),
    .QN(_00841_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04217_),
    .QN(_00840_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04218_),
    .QN(_00839_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04219_),
    .QN(_00838_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04220_),
    .QN(_00837_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04221_),
    .QN(_00836_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04222_),
    .QN(_00835_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04223_),
    .QN(_00834_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04224_),
    .QN(_00833_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04225_),
    .QN(_00832_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04226_),
    .QN(_00831_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04227_),
    .QN(_00830_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04228_),
    .QN(_00829_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04229_),
    .QN(_00828_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04230_),
    .QN(_00827_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04231_),
    .QN(_00826_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04232_),
    .QN(_00825_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04233_),
    .QN(_00824_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04234_),
    .QN(_00823_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04235_),
    .QN(_00822_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04236_),
    .QN(_00821_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04237_),
    .QN(_00820_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04238_),
    .QN(_00819_));
 DFFHQNx3_ASAP7_75t_R \xs[2].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04239_),
    .QN(_00818_));
 DFFHQNx1_ASAP7_75t_R \xs[2].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04240_),
    .QN(_00817_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04241_),
    .QN(_00023_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04242_),
    .QN(_00816_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04243_),
    .QN(_00815_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04244_),
    .QN(_00814_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04245_),
    .QN(_00813_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04246_),
    .QN(_00812_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04247_),
    .QN(_00811_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04248_),
    .QN(_00810_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04249_),
    .QN(_00809_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04250_),
    .QN(_00808_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04251_),
    .QN(_00807_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04252_),
    .QN(_00806_));
 DFFHQNx1_ASAP7_75t_R \xs[2].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .D(_04253_),
    .QN(_00805_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04254_),
    .QN(_00804_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04255_),
    .QN(_00803_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04256_),
    .QN(_00802_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04257_),
    .QN(_00801_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .D(_04258_),
    .QN(_00800_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_04259_),
    .QN(_00799_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_04260_),
    .QN(_00798_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04261_),
    .QN(_00797_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_04262_),
    .QN(_00796_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04263_),
    .QN(_00795_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .D(_04264_),
    .QN(_00794_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04265_),
    .QN(_00793_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04266_),
    .QN(_00792_));
 DFFHQNx3_ASAP7_75t_R \xs[2].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04267_),
    .QN(_00791_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04268_),
    .QN(_00790_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli0.i[11]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04269_),
    .QN(_00789_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04270_),
    .QN(_00788_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04271_),
    .QN(_00787_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04272_),
    .QN(_00786_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04273_),
    .QN(_00785_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04274_),
    .QN(_00784_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04275_),
    .QN(_00783_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04276_),
    .QN(_00049_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04277_),
    .QN(_00782_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04278_),
    .QN(_00781_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04279_),
    .QN(_00780_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04280_),
    .QN(_00779_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04281_),
    .QN(_00778_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04282_),
    .QN(_00777_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04283_),
    .QN(_00776_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04284_),
    .QN(_00775_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04285_),
    .QN(_00774_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04286_),
    .QN(_00773_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04287_),
    .QN(_00772_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04288_),
    .QN(_00771_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04289_),
    .QN(_00770_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04290_),
    .QN(_00769_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04291_),
    .QN(_00768_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04292_),
    .QN(_00767_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04293_),
    .QN(_00766_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04294_),
    .QN(_00765_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04295_),
    .QN(_00764_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04296_),
    .QN(_00763_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04297_),
    .QN(_00762_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04298_),
    .QN(_00761_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04299_),
    .QN(_00760_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04300_),
    .QN(_00759_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04301_),
    .QN(_00758_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04302_),
    .QN(_00757_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04303_),
    .QN(_00756_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04304_),
    .QN(_00755_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04305_),
    .QN(_00754_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04306_),
    .QN(_00753_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04307_),
    .QN(_00752_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04308_),
    .QN(_00751_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli1.i[11]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04309_),
    .QN(_00750_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04310_),
    .QN(_00749_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04311_),
    .QN(_00748_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04312_),
    .QN(_00747_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04313_),
    .QN(_00746_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_04314_),
    .QN(_00745_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_04315_),
    .QN(_00744_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04316_),
    .QN(_00050_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04317_),
    .QN(_00743_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04318_),
    .QN(_00742_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04319_),
    .QN(_00741_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04320_),
    .QN(_00740_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04321_),
    .QN(_00739_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04322_),
    .QN(_00738_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04323_),
    .QN(_00737_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04324_),
    .QN(_00736_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04325_),
    .QN(_00735_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04326_),
    .QN(_00734_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04327_),
    .QN(_00733_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04328_),
    .QN(_00732_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04329_),
    .QN(_00731_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04330_),
    .QN(_00730_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04331_),
    .QN(_00729_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04332_),
    .QN(_00728_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04333_),
    .QN(_00727_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04334_),
    .QN(_00726_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04335_),
    .QN(_00725_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04336_),
    .QN(_00724_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04337_),
    .QN(_00723_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04338_),
    .QN(_00722_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04339_),
    .QN(_00721_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04340_),
    .QN(_00720_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04341_),
    .QN(_00719_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04342_),
    .QN(_00718_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04343_),
    .QN(_00717_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04344_),
    .QN(_00716_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04345_),
    .QN(_00715_));
 DFFHQNx3_ASAP7_75t_R \xs[3].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .D(_04346_),
    .QN(_00714_));
 DFFHQNx1_ASAP7_75t_R \xs[3].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04347_),
    .QN(_00713_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04348_),
    .QN(_00024_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04349_),
    .QN(_00712_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04350_),
    .QN(_00711_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04351_),
    .QN(_00710_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04352_),
    .QN(_00709_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04353_),
    .QN(_00708_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04354_),
    .QN(_00707_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04355_),
    .QN(_00706_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04356_),
    .QN(_00705_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04357_),
    .QN(_00704_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04358_),
    .QN(_00703_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04359_),
    .QN(_00702_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .D(_04360_),
    .QN(_00701_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04361_),
    .QN(_00700_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04362_),
    .QN(_00699_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04363_),
    .QN(_00698_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .D(_04364_),
    .QN(_00697_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04365_),
    .QN(_00696_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_04366_),
    .QN(_00695_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_04367_),
    .QN(_00694_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04368_),
    .QN(_00693_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04369_),
    .QN(_00692_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04370_),
    .QN(_00691_));
 DFFHQNx1_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_04371_),
    .QN(_00690_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .D(_04372_),
    .QN(_00689_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04373_),
    .QN(_00688_));
 DFFHQNx3_ASAP7_75t_R \xs[3].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .D(_04374_),
    .QN(_00687_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04375_),
    .QN(_00686_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli0.i[13]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04376_),
    .QN(_00685_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04377_),
    .QN(_00684_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04378_),
    .QN(_00683_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04379_),
    .QN(_00682_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04380_),
    .QN(_00681_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04381_),
    .QN(_00680_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04382_),
    .QN(_00679_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04383_),
    .QN(_00051_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04384_),
    .QN(_00678_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04385_),
    .QN(_00677_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04386_),
    .QN(_00676_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04387_),
    .QN(_00675_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04388_),
    .QN(_00674_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04389_),
    .QN(_00673_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04390_),
    .QN(_00672_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04391_),
    .QN(_00671_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04392_),
    .QN(_00670_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04393_),
    .QN(_00669_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04394_),
    .QN(_00668_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04395_),
    .QN(_00667_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04396_),
    .QN(_00666_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04397_),
    .QN(_00665_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04398_),
    .QN(_00664_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04399_),
    .QN(_00663_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04400_),
    .QN(_00662_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04401_),
    .QN(_00661_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04402_),
    .QN(_00660_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04403_),
    .QN(_00659_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04404_),
    .QN(_00658_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04405_),
    .QN(_00657_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04406_),
    .QN(_00656_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04407_),
    .QN(_00655_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04408_),
    .QN(_00654_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04409_),
    .QN(_00653_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04410_),
    .QN(_00652_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04411_),
    .QN(_00651_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04412_),
    .QN(_00650_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04413_),
    .QN(_00649_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04414_),
    .QN(_00648_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04415_),
    .QN(_00647_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli1.i[10]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04416_),
    .QN(_00646_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04417_),
    .QN(_00645_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04418_),
    .QN(_00644_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04419_),
    .QN(_00643_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04420_),
    .QN(_00642_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04421_),
    .QN(_00641_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04422_),
    .QN(_00640_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04423_),
    .QN(_00052_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04424_),
    .QN(_00639_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04425_),
    .QN(_00638_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04426_),
    .QN(_00637_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04427_),
    .QN(_00636_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04428_),
    .QN(_00635_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04429_),
    .QN(_00634_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04430_),
    .QN(_00633_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04431_),
    .QN(_00632_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04432_),
    .QN(_00631_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04433_),
    .QN(_00630_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04434_),
    .QN(_00629_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04435_),
    .QN(_00628_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04436_),
    .QN(_00627_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04437_),
    .QN(_00626_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04438_),
    .QN(_00625_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04439_),
    .QN(_00624_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04440_),
    .QN(_00623_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04441_),
    .QN(_00622_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04442_),
    .QN(_00621_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04443_),
    .QN(_00620_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04444_),
    .QN(_00619_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04445_),
    .QN(_00618_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04446_),
    .QN(_00617_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04447_),
    .QN(_00616_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04448_),
    .QN(_00615_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04449_),
    .QN(_00614_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04450_),
    .QN(_00613_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04451_),
    .QN(_00612_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04452_),
    .QN(_00611_));
 DFFHQNx3_ASAP7_75t_R \xs[4].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04453_),
    .QN(_00610_));
 DFFHQNx1_ASAP7_75t_R \xs[4].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04454_),
    .QN(_00609_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04455_),
    .QN(_00025_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04456_),
    .QN(_00608_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(_04457_),
    .QN(_00607_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04458_),
    .QN(_00606_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04459_),
    .QN(_00605_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04460_),
    .QN(_00604_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04461_),
    .QN(_00603_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04462_),
    .QN(_00602_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04463_),
    .QN(_00601_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04464_),
    .QN(_00600_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04465_),
    .QN(_00599_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04466_),
    .QN(_00598_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(_04467_),
    .QN(_00597_));
 DFFHQNx3_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04468_),
    .QN(_00596_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04469_),
    .QN(_00595_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04470_),
    .QN(_00594_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04471_),
    .QN(_00593_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04472_),
    .QN(_00592_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_04473_),
    .QN(_00591_));
 DFFHQNx3_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_04474_),
    .QN(_00590_));
 DFFHQNx3_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_04475_),
    .QN(_00589_));
 DFFHQNx3_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_04476_),
    .QN(_00588_));
 DFFHQNx3_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_04477_),
    .QN(_00587_));
 DFFHQNx3_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04478_),
    .QN(_00586_));
 DFFHQNx3_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_04479_),
    .QN(_00585_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_48_clk),
    .D(_04480_),
    .QN(_00584_));
 DFFHQNx1_ASAP7_75t_R \xs[4].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04481_),
    .QN(_00583_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04482_),
    .QN(_00582_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli0.i[11]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04483_),
    .QN(_00581_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04484_),
    .QN(_00580_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04485_),
    .QN(_00579_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04486_),
    .QN(_00578_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04487_),
    .QN(_00577_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04488_),
    .QN(_00576_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04489_),
    .QN(_00575_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04490_),
    .QN(_00053_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04491_),
    .QN(_00574_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04492_),
    .QN(_00573_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04493_),
    .QN(_00572_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04494_),
    .QN(_00571_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04495_),
    .QN(_00570_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04496_),
    .QN(_00569_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04497_),
    .QN(_00568_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04498_),
    .QN(_00567_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04499_),
    .QN(_00566_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04500_),
    .QN(_00565_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04501_),
    .QN(_00564_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04502_),
    .QN(_00563_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04503_),
    .QN(_00562_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04504_),
    .QN(_00561_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04505_),
    .QN(_00560_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04506_),
    .QN(_00559_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04507_),
    .QN(_00558_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04508_),
    .QN(_00557_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04509_),
    .QN(_00556_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04510_),
    .QN(_00555_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04511_),
    .QN(_00554_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04512_),
    .QN(_00553_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04513_),
    .QN(_00552_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04514_),
    .QN(_00551_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04515_),
    .QN(_00550_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04516_),
    .QN(_00549_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04517_),
    .QN(_00548_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04518_),
    .QN(_00547_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04519_),
    .QN(_00546_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04520_),
    .QN(_00545_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04521_),
    .QN(_00544_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04522_),
    .QN(_00543_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli1.i[11]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04523_),
    .QN(_00542_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04524_),
    .QN(_00541_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04525_),
    .QN(_00540_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04526_),
    .QN(_00539_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04527_),
    .QN(_00538_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04528_),
    .QN(_00537_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04529_),
    .QN(_00536_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04530_),
    .QN(_00054_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04531_),
    .QN(_00535_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04532_),
    .QN(_00534_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04533_),
    .QN(_00533_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04534_),
    .QN(_00532_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04535_),
    .QN(_00531_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04536_),
    .QN(_00530_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04537_),
    .QN(_00529_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04538_),
    .QN(_00528_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04539_),
    .QN(_00527_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04540_),
    .QN(_00526_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04541_),
    .QN(_00525_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04542_),
    .QN(_00524_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04543_),
    .QN(_00523_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04544_),
    .QN(_00522_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04545_),
    .QN(_00521_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04546_),
    .QN(_00520_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04547_),
    .QN(_00519_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04548_),
    .QN(_00518_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04549_),
    .QN(_00517_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04550_),
    .QN(_00516_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04551_),
    .QN(_00515_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04552_),
    .QN(_00514_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04553_),
    .QN(_00513_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04554_),
    .QN(_00512_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04555_),
    .QN(_00511_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04556_),
    .QN(_00510_));
 DFFHQNx1_ASAP7_75t_R \xs[5].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04557_),
    .QN(_00509_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04558_),
    .QN(_00508_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04559_),
    .QN(_00507_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04560_),
    .QN(_00506_));
 DFFHQNx3_ASAP7_75t_R \xs[5].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04561_),
    .QN(_00505_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04562_),
    .QN(_00026_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04563_),
    .QN(_00504_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04564_),
    .QN(_00503_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04565_),
    .QN(_00502_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04566_),
    .QN(_00501_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04567_),
    .QN(_00500_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04568_),
    .QN(_00499_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04569_),
    .QN(_00498_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .D(_04570_),
    .QN(_00497_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04571_),
    .QN(_00496_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04572_),
    .QN(_00495_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04573_),
    .QN(_00494_));
 DFFHQNx1_ASAP7_75t_R \xs[5].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04574_),
    .QN(_00493_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04575_),
    .QN(_00492_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04576_),
    .QN(_00491_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_49_clk),
    .D(_04577_),
    .QN(_00490_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04578_),
    .QN(_00489_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04579_),
    .QN(_00488_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04580_),
    .QN(_00487_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04581_),
    .QN(_00486_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04582_),
    .QN(_00485_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .D(_04583_),
    .QN(_00484_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_04584_),
    .QN(_00483_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_04585_),
    .QN(_00482_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .D(_04586_),
    .QN(_00481_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04587_),
    .QN(_00480_));
 DFFHQNx3_ASAP7_75t_R \xs[5].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_50_clk),
    .D(_04588_),
    .QN(_00479_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04589_),
    .QN(_00478_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli0.i[12]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04590_),
    .QN(_00477_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04591_),
    .QN(_00476_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04592_),
    .QN(_00475_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04593_),
    .QN(_00474_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04594_),
    .QN(_00473_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04595_),
    .QN(_00472_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04596_),
    .QN(_00471_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04597_),
    .QN(_00055_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04598_),
    .QN(_00470_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04599_),
    .QN(_00469_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04600_),
    .QN(_00468_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04601_),
    .QN(_00467_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04602_),
    .QN(_00466_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04603_),
    .QN(_00465_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04604_),
    .QN(_00464_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04605_),
    .QN(_00463_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04606_),
    .QN(_00462_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04607_),
    .QN(_00461_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04608_),
    .QN(_00460_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04609_),
    .QN(_00459_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04610_),
    .QN(_00458_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04611_),
    .QN(_00457_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04612_),
    .QN(_00456_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04613_),
    .QN(_00455_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04614_),
    .QN(_00454_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04615_),
    .QN(_00453_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04616_),
    .QN(_00452_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04617_),
    .QN(_00451_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04618_),
    .QN(_00450_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04619_),
    .QN(_00449_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04620_),
    .QN(_00448_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04621_),
    .QN(_00447_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04622_),
    .QN(_00446_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04623_),
    .QN(_00445_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04624_),
    .QN(_00444_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04625_),
    .QN(_00443_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .D(_04626_),
    .QN(_00442_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04627_),
    .QN(_00441_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04628_),
    .QN(_00440_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04629_),
    .QN(_00439_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli1.i[12]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04630_),
    .QN(_00438_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04631_),
    .QN(_00437_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04632_),
    .QN(_00436_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04633_),
    .QN(_00435_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04634_),
    .QN(_00434_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04635_),
    .QN(_00433_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04636_),
    .QN(_00432_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04637_),
    .QN(_00056_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04638_),
    .QN(_00431_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04639_),
    .QN(_00430_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04640_),
    .QN(_00429_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04641_),
    .QN(_00428_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04642_),
    .QN(_00427_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04643_),
    .QN(_00426_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04644_),
    .QN(_00425_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04645_),
    .QN(_00424_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04646_),
    .QN(_00423_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04647_),
    .QN(_00422_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04648_),
    .QN(_00421_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04649_),
    .QN(_00420_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04650_),
    .QN(_00419_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04651_),
    .QN(_00418_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04652_),
    .QN(_00417_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04653_),
    .QN(_00416_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04654_),
    .QN(_00415_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04655_),
    .QN(_00414_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04656_),
    .QN(_00413_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04657_),
    .QN(_00412_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04658_),
    .QN(_00411_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04659_),
    .QN(_00410_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04660_),
    .QN(_00409_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04661_),
    .QN(_00408_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04662_),
    .QN(_00407_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04663_),
    .QN(_00406_));
 DFFHQNx1_ASAP7_75t_R \xs[6].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04664_),
    .QN(_00405_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04665_),
    .QN(_00404_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04666_),
    .QN(_00403_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04667_),
    .QN(_00402_));
 DFFHQNx3_ASAP7_75t_R \xs[6].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04668_),
    .QN(_00401_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04669_),
    .QN(_00027_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04670_),
    .QN(_00400_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04671_),
    .QN(_00399_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04672_),
    .QN(_00398_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04673_),
    .QN(_00397_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04674_),
    .QN(_00396_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04675_),
    .QN(_00395_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04676_),
    .QN(_00394_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04677_),
    .QN(_00393_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04678_),
    .QN(_00392_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04679_),
    .QN(_00391_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04680_),
    .QN(_00390_));
 DFFHQNx1_ASAP7_75t_R \xs[6].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .D(_04681_),
    .QN(_00389_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04682_),
    .QN(_00388_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_04683_),
    .QN(_00387_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_04684_),
    .QN(_00386_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_04685_),
    .QN(_00385_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04686_),
    .QN(_00384_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04687_),
    .QN(_00383_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04688_),
    .QN(_00382_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04689_),
    .QN(_00381_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04690_),
    .QN(_00380_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_04691_),
    .QN(_00379_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04692_),
    .QN(_00378_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_45_clk),
    .D(_04693_),
    .QN(_00377_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_04694_),
    .QN(_00376_));
 DFFHQNx3_ASAP7_75t_R \xs[6].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_04695_),
    .QN(_00375_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04696_),
    .QN(_00374_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli0.i[12]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04697_),
    .QN(_00373_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04698_),
    .QN(_00372_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04699_),
    .QN(_00371_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04700_),
    .QN(_00370_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04701_),
    .QN(_00369_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04702_),
    .QN(_00368_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04703_),
    .QN(_00367_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04704_),
    .QN(_00057_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04705_),
    .QN(_00366_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04706_),
    .QN(_00365_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04707_),
    .QN(_00364_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04708_),
    .QN(_00363_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04709_),
    .QN(_00362_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04710_),
    .QN(_00361_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .D(_04711_),
    .QN(_00360_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04712_),
    .QN(_00359_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04713_),
    .QN(_00358_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04714_),
    .QN(_00357_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04715_),
    .QN(_00356_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04716_),
    .QN(_00355_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04717_),
    .QN(_00354_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04718_),
    .QN(_00353_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04719_),
    .QN(_00352_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04720_),
    .QN(_00351_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04721_),
    .QN(_00350_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04722_),
    .QN(_00349_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04723_),
    .QN(_00348_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04724_),
    .QN(_00347_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04725_),
    .QN(_00346_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04726_),
    .QN(_00345_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04727_),
    .QN(_00344_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04728_),
    .QN(_00343_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04729_),
    .QN(_00342_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04730_),
    .QN(_00341_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04731_),
    .QN(_00340_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04732_),
    .QN(_00339_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04733_),
    .QN(_00338_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04734_),
    .QN(_00337_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04735_),
    .QN(_00336_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04736_),
    .QN(_00335_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli1.i[12]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04737_),
    .QN(_00334_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04738_),
    .QN(_00333_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04739_),
    .QN(_00332_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04740_),
    .QN(_00331_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04741_),
    .QN(_00330_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04742_),
    .QN(_00329_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04743_),
    .QN(_00328_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04744_),
    .QN(_00058_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04745_),
    .QN(_00327_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04746_),
    .QN(_00326_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04747_),
    .QN(_00325_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04748_),
    .QN(_00324_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04749_),
    .QN(_00323_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04750_),
    .QN(_00322_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04751_),
    .QN(_00321_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .D(_04752_),
    .QN(_00320_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04753_),
    .QN(_00319_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04754_),
    .QN(_00318_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04755_),
    .QN(_00317_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .D(_04756_),
    .QN(_00316_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04757_),
    .QN(_00315_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04758_),
    .QN(_00314_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04759_),
    .QN(_00313_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04760_),
    .QN(_00312_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04761_),
    .QN(_00311_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04762_),
    .QN(_00310_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04763_),
    .QN(_00309_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04764_),
    .QN(_00308_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04765_),
    .QN(_00307_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04766_),
    .QN(_00306_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04767_),
    .QN(_00305_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04768_),
    .QN(_00304_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04769_),
    .QN(_00303_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04770_),
    .QN(_00302_));
 DFFHQNx1_ASAP7_75t_R \xs[7].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04771_),
    .QN(_00301_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04772_),
    .QN(_00300_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04773_),
    .QN(_00299_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04774_),
    .QN(_00298_));
 DFFHQNx3_ASAP7_75t_R \xs[7].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04775_),
    .QN(_00297_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04776_),
    .QN(_00028_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04777_),
    .QN(_00296_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04778_),
    .QN(_00295_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04779_),
    .QN(_00294_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04780_),
    .QN(_00293_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04781_),
    .QN(_00292_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04782_),
    .QN(_00291_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04783_),
    .QN(_00290_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04784_),
    .QN(_00289_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04785_),
    .QN(_00288_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04786_),
    .QN(_00287_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04787_),
    .QN(_00286_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04788_),
    .QN(_00285_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04789_),
    .QN(_00284_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04790_),
    .QN(_00283_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04791_),
    .QN(_00282_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04792_),
    .QN(_00281_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04793_),
    .QN(_00280_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04794_),
    .QN(_00279_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04795_),
    .QN(_00278_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04796_),
    .QN(_00277_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_04797_),
    .QN(_00276_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04798_),
    .QN(_00275_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04799_),
    .QN(_00274_));
 DFFHQNx1_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04800_),
    .QN(_00273_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04801_),
    .QN(_00272_));
 DFFHQNx3_ASAP7_75t_R \xs[7].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .D(_04802_),
    .QN(_00271_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04803_),
    .QN(_00270_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli0.i[14]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04804_),
    .QN(_00269_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04805_),
    .QN(_00268_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04806_),
    .QN(_00267_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04807_),
    .QN(_00266_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04808_),
    .QN(_00265_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04809_),
    .QN(_00264_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04810_),
    .QN(_00263_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04811_),
    .QN(_00059_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04812_),
    .QN(_00262_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04813_),
    .QN(_00261_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .D(_04814_),
    .QN(_00260_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04815_),
    .QN(_00259_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04816_),
    .QN(_00258_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04817_),
    .QN(_00257_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04818_),
    .QN(_00256_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04819_),
    .QN(_00255_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04820_),
    .QN(_00254_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04821_),
    .QN(_00253_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04822_),
    .QN(_00252_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04823_),
    .QN(_00251_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04824_),
    .QN(_00250_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04825_),
    .QN(_00249_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04826_),
    .QN(_00248_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04827_),
    .QN(_00247_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04828_),
    .QN(_00246_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04829_),
    .QN(_00245_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04830_),
    .QN(_00244_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04831_),
    .QN(_00243_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04832_),
    .QN(_00242_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04833_),
    .QN(_00241_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04834_),
    .QN(_00240_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04835_),
    .QN(_00239_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04836_),
    .QN(_00238_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04837_),
    .QN(_00237_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04838_),
    .QN(_00236_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04839_),
    .QN(_00235_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04840_),
    .QN(_00234_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04841_),
    .QN(_00233_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04842_),
    .QN(_00232_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04843_),
    .QN(_00231_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli1.i[10]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04844_),
    .QN(_00230_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04845_),
    .QN(_00229_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04846_),
    .QN(_00228_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04847_),
    .QN(_00227_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04848_),
    .QN(_00226_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04849_),
    .QN(_00225_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04850_),
    .QN(_00224_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04851_),
    .QN(_00060_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04852_),
    .QN(_00223_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04853_),
    .QN(_00222_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04854_),
    .QN(_00221_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04855_),
    .QN(_00220_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04856_),
    .QN(_00219_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04857_),
    .QN(_00218_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04858_),
    .QN(_00217_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04859_),
    .QN(_00216_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04860_),
    .QN(_00215_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04861_),
    .QN(_00214_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04862_),
    .QN(_00213_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04863_),
    .QN(_00212_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04864_),
    .QN(_00211_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04865_),
    .QN(_00210_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04866_),
    .QN(_00209_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04867_),
    .QN(_00208_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04868_),
    .QN(_00207_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04869_),
    .QN(_00206_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04870_),
    .QN(_00205_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04871_),
    .QN(_00204_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04872_),
    .QN(_00203_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04873_),
    .QN(_00202_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04874_),
    .QN(_00201_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04875_),
    .QN(_00200_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04876_),
    .QN(_00199_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04877_),
    .QN(_00198_));
 DFFHQNx1_ASAP7_75t_R \xs[8].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04878_),
    .QN(_00197_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04879_),
    .QN(_00196_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04880_),
    .QN(_00195_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04881_),
    .QN(_00194_));
 DFFHQNx3_ASAP7_75t_R \xs[8].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04882_),
    .QN(_00193_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04883_),
    .QN(_00029_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04884_),
    .QN(_00192_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_04885_),
    .QN(_00191_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_04886_),
    .QN(_00190_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04887_),
    .QN(_00189_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_04888_),
    .QN(_00188_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_04889_),
    .QN(_00187_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04890_),
    .QN(_00186_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04891_),
    .QN(_00185_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .D(_04892_),
    .QN(_00184_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04893_),
    .QN(_00183_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04894_),
    .QN(_00182_));
 DFFHQNx1_ASAP7_75t_R \xs[8].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04895_),
    .QN(_00181_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04896_),
    .QN(_00180_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04897_),
    .QN(_00179_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04898_),
    .QN(_00178_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04899_),
    .QN(_00177_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04900_),
    .QN(_00176_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04901_),
    .QN(_00175_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04902_),
    .QN(_00174_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04903_),
    .QN(_00173_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04904_),
    .QN(_00172_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04905_),
    .QN(_00171_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04906_),
    .QN(_00170_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04907_),
    .QN(_00169_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04908_),
    .QN(_00168_));
 DFFHQNx3_ASAP7_75t_R \xs[8].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .D(_04909_),
    .QN(_00167_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli0.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04910_),
    .QN(_00166_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli0.i[11]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04911_),
    .QN(_00165_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli0.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04912_),
    .QN(_00164_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04913_),
    .QN(_00163_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04914_),
    .QN(_00162_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04915_),
    .QN(_00161_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04916_),
    .QN(_00160_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli0.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04917_),
    .QN(_00159_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04918_),
    .QN(_00061_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04919_),
    .QN(_00158_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04920_),
    .QN(_00157_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04921_),
    .QN(_00156_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli0.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04922_),
    .QN(_00155_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04923_),
    .QN(_00154_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04924_),
    .QN(_00153_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04925_),
    .QN(_00152_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04926_),
    .QN(_00151_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04927_),
    .QN(_00150_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04928_),
    .QN(_00149_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli0.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04929_),
    .QN(_00148_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04930_),
    .QN(_00147_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04931_),
    .QN(_00146_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04932_),
    .QN(_00145_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04933_),
    .QN(_00144_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04934_),
    .QN(_00143_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04935_),
    .QN(_00142_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04936_),
    .QN(_00141_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04937_),
    .QN(_00140_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04938_),
    .QN(_00139_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04939_),
    .QN(_00138_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04940_),
    .QN(_00137_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04941_),
    .QN(_00136_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli0.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04942_),
    .QN(_00135_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04943_),
    .QN(_00134_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04944_),
    .QN(_00133_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04945_),
    .QN(_00132_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04946_),
    .QN(_00131_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04947_),
    .QN(_00130_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli0.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04948_),
    .QN(_00129_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli0.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_04949_),
    .QN(_00128_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli1.i[0]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04950_),
    .QN(_00127_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli1.i[11]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04951_),
    .QN(_00126_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.i[32]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04952_),
    .QN(_00125_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.i[33]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04953_),
    .QN(_00124_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.i[34]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04954_),
    .QN(_00123_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.i[35]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04955_),
    .QN(_00122_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.i[36]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04956_),
    .QN(_00121_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.i[39]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04957_),
    .QN(_00120_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04958_),
    .QN(_00062_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[10]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04959_),
    .QN(_00119_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli1.r[11]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04960_),
    .QN(_00118_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[12]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04961_),
    .QN(_00117_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[13]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04962_),
    .QN(_00116_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[14]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04963_),
    .QN(_00115_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[15]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04964_),
    .QN(_00114_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[16]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04965_),
    .QN(_00113_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[17]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04966_),
    .QN(_00112_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[18]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .D(_04967_),
    .QN(_00111_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[19]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04968_),
    .QN(_00110_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli1.r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04969_),
    .QN(_00109_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[20]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04970_),
    .QN(_00108_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[21]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04971_),
    .QN(_00107_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[22]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04972_),
    .QN(_00106_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli1.r[23]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04973_),
    .QN(_00105_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[24]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04974_),
    .QN(_00104_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[25]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04975_),
    .QN(_00103_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[26]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04976_),
    .QN(_00102_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[27]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04977_),
    .QN(_00101_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[28]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04978_),
    .QN(_00100_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[29]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04979_),
    .QN(_00099_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04980_),
    .QN(_00098_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[30]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04981_),
    .QN(_00097_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli1.r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04982_),
    .QN(_00096_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04983_),
    .QN(_00095_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04984_),
    .QN(_00094_));
 DFFHQNx1_ASAP7_75t_R \xs[9].cli1.r[5]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04985_),
    .QN(_00093_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[6]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04986_),
    .QN(_00092_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[7]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04987_),
    .QN(_00091_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[8]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .D(_04988_),
    .QN(_00090_));
 DFFHQNx3_ASAP7_75t_R \xs[9].cli1.r[9]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .D(_04989_),
    .QN(_00089_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.full.r.toggle$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_04990_),
    .QN(_00030_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.l_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04991_),
    .QN(_00088_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.l_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04992_),
    .QN(_00087_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.l_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04993_),
    .QN(_00086_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.l_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04994_),
    .QN(_00085_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.l_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04995_),
    .QN(_00084_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.l_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04996_),
    .QN(_00083_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.r_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_04997_),
    .QN(_00082_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.r_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04998_),
    .QN(_00081_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.r_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_04999_),
    .QN(_00080_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.r_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05000_),
    .QN(_00079_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.r_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05001_),
    .QN(_00078_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.r_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05002_),
    .QN(_00077_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[0]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05003_),
    .QN(_00076_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[1]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05004_),
    .QN(_00075_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[2]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05005_),
    .QN(_00074_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[31]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05006_),
    .QN(_00073_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[32]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05007_),
    .QN(_00072_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[33]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05008_),
    .QN(_00071_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[34]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05009_),
    .QN(_00070_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[35]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05010_),
    .QN(_00069_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[36]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05011_),
    .QN(_00068_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[37]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_05012_),
    .QN(_00067_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[38]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .D(_05013_),
    .QN(_00066_));
 DFFHQNx1_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[39]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_05014_),
    .QN(_00065_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[3]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05015_),
    .QN(_00064_));
 DFFHQNx3_ASAP7_75t_R \xs[9].t_level0.sb.u0_o_r[4]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_05016_),
    .QN(_00063_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_Right_227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_Right_228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_Right_229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_Right_230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_Right_231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_Right_232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_Right_233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_Right_234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_Right_235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_Right_236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_Right_237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_Right_238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_Right_239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_Right_240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_Right_241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_Right_242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_Right_243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Left_299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Left_300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Left_301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Left_302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Left_303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Left_304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Left_305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Left_306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Left_307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Left_308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Left_309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Left_310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Left_311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Left_312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Left_313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Left_314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Left_315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Left_316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Left_317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Left_318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Left_319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Left_320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Left_321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Left_322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Left_323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Left_324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Left_325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Left_326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Left_327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Left_328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Left_329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Left_330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Left_331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Left_332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Left_333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Left_334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Left_335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Left_336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Left_337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Left_338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Left_339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Left_340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Left_341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Left_342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Left_343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Left_344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Left_345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Left_346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Left_347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Left_348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Left_349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Left_350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Left_351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Left_352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Left_353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Left_354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Left_355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Left_356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Left_357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Left_358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Left_359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Left_360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Left_361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Left_362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Left_363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Left_364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Left_365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Left_366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Left_367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Left_368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Left_369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Left_370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Left_371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Left_372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Left_373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Left_374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Left_375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Left_376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Left_377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Left_378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Left_379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Left_380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Left_381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Left_382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Left_383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Left_384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Left_385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Left_386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Left_387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Left_388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Left_389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Left_390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Left_391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Left_392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Left_393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Left_394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Left_395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_Left_396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_Left_397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_Left_398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_Left_399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_Left_400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_Left_401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_Left_402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_Left_403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_Left_404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_Left_405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Left_406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Left_407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Left_408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Left_409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Left_410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Left_411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Left_412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Left_413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Left_414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Left_415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Left_416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Left_417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_Left_418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_Left_419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_Left_420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_Left_421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Left_422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_Left_423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_Left_424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_Left_425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_Left_426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_Left_427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_Left_428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_Left_429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_Left_430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_Left_431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_Left_432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_Left_433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_Left_434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_Left_435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_Left_436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_Left_437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_Left_438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_Left_439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_Left_440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_Left_441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_Left_442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_Left_443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_Left_444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_Left_445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_Left_446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_Left_447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_Left_448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_Left_449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_Left_450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_Left_451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_Left_452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_Left_453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_Left_454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_Left_455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_Left_456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_Left_457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_Left_458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_Left_459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_Left_460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_Left_461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_Left_462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_Left_463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_Left_464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_Left_465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_Left_466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_Left_467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_Left_468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_Left_469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_Left_470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_Left_471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_Left_472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_Left_473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_Left_474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_Left_475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_Left_476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_Left_477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_Left_478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_Left_479 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_Left_480 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_Left_481 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_Left_482 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_Left_483 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_Left_484 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_Left_485 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_Left_486 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_Left_487 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_488 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_489 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_490 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_491 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_492 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_493 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_494 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_495 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_496 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_497 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_498 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_499 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_500 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_501 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_502 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_14_503 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_15_504 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_16_505 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_17_506 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_18_507 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_19_508 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_20_509 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_21_510 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_22_511 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_23_512 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_24_513 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_25_514 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_26_515 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_27_516 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_28_517 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_29_518 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_30_519 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_31_520 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_32_521 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_33_522 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_34_523 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_35_524 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_36_525 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_37_526 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_38_527 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_39_528 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_40_529 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_41_530 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_42_531 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_43_532 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_44_533 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_45_534 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_46_535 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_47_536 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_48_537 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_49_538 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_50_539 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_51_540 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_52_541 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_53_542 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_54_543 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_55_544 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_56_545 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_57_546 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_58_547 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_59_548 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_60_549 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_61_550 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_62_551 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_63_552 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_64_553 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_65_554 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_66_555 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_67_556 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_68_557 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_69_558 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_70_559 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_71_560 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_72_561 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_73_562 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_74_563 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_75_564 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_76_565 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_77_566 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_78_567 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_79_568 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_80_569 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_81_570 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_571 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_83_572 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_84_573 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_85_574 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_86_575 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_87_576 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_88_577 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_89_578 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_90_579 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_91_580 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_92_581 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_93_582 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_94_583 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_95_584 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_96_585 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_97_586 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_98_587 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_99_588 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_100_589 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_101_590 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_102_591 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_103_592 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_104_593 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_105_594 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_106_595 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_107_596 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_108_597 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_109_598 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_110_599 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_111_600 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_112_601 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_113_602 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_114_603 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_115_604 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_116_605 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_117_606 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_118_607 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_119_608 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_120_609 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_121_610 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_122_611 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_123_612 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_124_613 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_125_614 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_126_615 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_127_616 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_128_617 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_129_618 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_130_619 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_131_620 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_132_621 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_133_622 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_134_623 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_135_624 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_136_625 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_137_626 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_138_627 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_139_628 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_140_629 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_141_630 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_142_631 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_143_632 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_144_633 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_145_634 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_146_635 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_147_636 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_148_637 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_149_638 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_150_639 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_151_640 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_152_641 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_153_642 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_154_643 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_155_644 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_156_645 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_157_646 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_158_647 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_159_648 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_160_649 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_161_650 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_162_651 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_163_652 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_164_653 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_165_654 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_166_655 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_167_656 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_168_657 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_169_658 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_170_659 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_171_660 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_172_661 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_173_662 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_174_663 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_175_664 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_176_665 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_177_666 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_667 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_668 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_669 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_670 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_671 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_672 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_673 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_674 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_675 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_676 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_677 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_678 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_190_679 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_191_680 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_192_681 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_193_682 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_194_683 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_195_684 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_196_685 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_197_686 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_198_687 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_199_688 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_200_689 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_201_690 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_202_691 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_203_692 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_204_693 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_205_694 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_206_695 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_207_696 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_208_697 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_209_698 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_210_699 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_211_700 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_212_701 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_213_702 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_214_703 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_215_704 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_216_705 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_217_706 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_218_707 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_219_708 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_220_709 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_221_710 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_222_711 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_223_712 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_224_713 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_225_714 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_226_715 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_227_716 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_228_717 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_229_718 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_230_719 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_231_720 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_232_721 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_233_722 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_234_723 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_235_724 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_236_725 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_237_726 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_238_727 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_239_728 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_240_729 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_241_730 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_242_731 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_243_732 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_243_733 ();
 BUFx6f_ASAP7_75t_R input1 (.A(cmd[0]),
    .Y(net1));
 BUFx6f_ASAP7_75t_R input2 (.A(cmd[1]),
    .Y(net2));
 BUFx6f_ASAP7_75t_R input3 (.A(cmd[2]),
    .Y(net3));
 BUFx6f_ASAP7_75t_R input4 (.A(cmd[3]),
    .Y(net4));
 BUFx6f_ASAP7_75t_R input5 (.A(cmd[4]),
    .Y(net5));
 BUFx6f_ASAP7_75t_R input6 (.A(cmd[5]),
    .Y(net6));
 BUFx3_ASAP7_75t_R input7 (.A(in[0]),
    .Y(net7));
 BUFx3_ASAP7_75t_R input8 (.A(in[1]),
    .Y(net8));
 BUFx3_ASAP7_75t_R input9 (.A(in[2]),
    .Y(net9));
 BUFx6f_ASAP7_75t_R input10 (.A(in[31]),
    .Y(net10));
 BUFx6f_ASAP7_75t_R input11 (.A(in[32]),
    .Y(net11));
 BUFx3_ASAP7_75t_R input12 (.A(in[33]),
    .Y(net12));
 BUFx3_ASAP7_75t_R input13 (.A(in[34]),
    .Y(net13));
 BUFx3_ASAP7_75t_R input14 (.A(in[35]),
    .Y(net14));
 BUFx3_ASAP7_75t_R input15 (.A(in[36]),
    .Y(net15));
 BUFx3_ASAP7_75t_R input16 (.A(in[37]),
    .Y(net16));
 BUFx3_ASAP7_75t_R input17 (.A(in[38]),
    .Y(net17));
 BUFx3_ASAP7_75t_R input18 (.A(in[39]),
    .Y(net18));
 BUFx3_ASAP7_75t_R input19 (.A(in[3]),
    .Y(net19));
 BUFx3_ASAP7_75t_R input20 (.A(in[4]),
    .Y(net20));
 BUFx6f_ASAP7_75t_R input21 (.A(rst),
    .Y(net21));
 BUFx3_ASAP7_75t_R output22 (.A(net22),
    .Y(out[0]));
 BUFx3_ASAP7_75t_R output23 (.A(net23),
    .Y(out[1000]));
 BUFx3_ASAP7_75t_R output24 (.A(net24),
    .Y(out[1010]));
 BUFx3_ASAP7_75t_R output25 (.A(net25),
    .Y(out[1013]));
 BUFx3_ASAP7_75t_R output26 (.A(net26),
    .Y(out[1014]));
 BUFx3_ASAP7_75t_R output27 (.A(net27),
    .Y(out[1032]));
 BUFx3_ASAP7_75t_R output28 (.A(net28),
    .Y(out[1033]));
 BUFx3_ASAP7_75t_R output29 (.A(net29),
    .Y(out[1034]));
 BUFx3_ASAP7_75t_R output30 (.A(net30),
    .Y(out[1035]));
 BUFx3_ASAP7_75t_R output31 (.A(net31),
    .Y(out[1036]));
 BUFx3_ASAP7_75t_R output32 (.A(net32),
    .Y(out[1039]));
 BUFx3_ASAP7_75t_R output33 (.A(net33),
    .Y(out[1040]));
 BUFx3_ASAP7_75t_R output34 (.A(net34),
    .Y(out[1051]));
 BUFx3_ASAP7_75t_R output35 (.A(net35),
    .Y(out[1053]));
 BUFx3_ASAP7_75t_R output36 (.A(net36),
    .Y(out[1054]));
 BUFx3_ASAP7_75t_R output37 (.A(net37),
    .Y(out[1072]));
 BUFx3_ASAP7_75t_R output38 (.A(net38),
    .Y(out[1073]));
 BUFx3_ASAP7_75t_R output39 (.A(net39),
    .Y(out[1074]));
 BUFx3_ASAP7_75t_R output40 (.A(net40),
    .Y(out[1075]));
 BUFx3_ASAP7_75t_R output41 (.A(net41),
    .Y(out[1076]));
 BUFx3_ASAP7_75t_R output42 (.A(net42),
    .Y(out[1079]));
 BUFx3_ASAP7_75t_R output43 (.A(net43),
    .Y(out[1080]));
 BUFx3_ASAP7_75t_R output44 (.A(net44),
    .Y(out[1090]));
 BUFx3_ASAP7_75t_R output45 (.A(net45),
    .Y(out[1091]));
 BUFx3_ASAP7_75t_R output46 (.A(net46),
    .Y(out[1093]));
 BUFx3_ASAP7_75t_R output47 (.A(net47),
    .Y(out[1094]));
 BUFx3_ASAP7_75t_R output48 (.A(net48),
    .Y(out[1112]));
 BUFx3_ASAP7_75t_R output49 (.A(net49),
    .Y(out[1113]));
 BUFx3_ASAP7_75t_R output50 (.A(net50),
    .Y(out[1114]));
 BUFx3_ASAP7_75t_R output51 (.A(net51),
    .Y(out[1115]));
 BUFx3_ASAP7_75t_R output52 (.A(net52),
    .Y(out[1116]));
 BUFx3_ASAP7_75t_R output53 (.A(net53),
    .Y(out[1119]));
 BUFx3_ASAP7_75t_R output54 (.A(net54),
    .Y(out[1120]));
 BUFx3_ASAP7_75t_R output55 (.A(net55),
    .Y(out[112]));
 BUFx3_ASAP7_75t_R output56 (.A(net56),
    .Y(out[1132]));
 BUFx3_ASAP7_75t_R output57 (.A(net57),
    .Y(out[1133]));
 BUFx3_ASAP7_75t_R output58 (.A(net58),
    .Y(out[1134]));
 BUFx3_ASAP7_75t_R output59 (.A(net59),
    .Y(out[113]));
 BUFx3_ASAP7_75t_R output60 (.A(net60),
    .Y(out[114]));
 BUFx3_ASAP7_75t_R output61 (.A(net61),
    .Y(out[1152]));
 BUFx3_ASAP7_75t_R output62 (.A(net62),
    .Y(out[1153]));
 BUFx3_ASAP7_75t_R output63 (.A(net63),
    .Y(out[1154]));
 BUFx3_ASAP7_75t_R output64 (.A(net64),
    .Y(out[1155]));
 BUFx3_ASAP7_75t_R output65 (.A(net65),
    .Y(out[1156]));
 BUFx3_ASAP7_75t_R output66 (.A(net66),
    .Y(out[1159]));
 BUFx3_ASAP7_75t_R output67 (.A(net67),
    .Y(out[115]));
 BUFx3_ASAP7_75t_R output68 (.A(net68),
    .Y(out[1160]));
 BUFx3_ASAP7_75t_R output69 (.A(net69),
    .Y(out[116]));
 BUFx3_ASAP7_75t_R output70 (.A(net70),
    .Y(out[1170]));
 BUFx3_ASAP7_75t_R output71 (.A(net71),
    .Y(out[1172]));
 BUFx3_ASAP7_75t_R output72 (.A(net72),
    .Y(out[1173]));
 BUFx3_ASAP7_75t_R output73 (.A(net73),
    .Y(out[1174]));
 BUFx3_ASAP7_75t_R output74 (.A(net74),
    .Y(out[1192]));
 BUFx3_ASAP7_75t_R output75 (.A(net75),
    .Y(out[1193]));
 BUFx3_ASAP7_75t_R output76 (.A(net76),
    .Y(out[1194]));
 BUFx3_ASAP7_75t_R output77 (.A(net77),
    .Y(out[1195]));
 BUFx3_ASAP7_75t_R output78 (.A(net78),
    .Y(out[1196]));
 BUFx3_ASAP7_75t_R output79 (.A(net79),
    .Y(out[1199]));
 BUFx3_ASAP7_75t_R output80 (.A(net80),
    .Y(out[119]));
 BUFx3_ASAP7_75t_R output81 (.A(net81),
    .Y(out[1200]));
 BUFx3_ASAP7_75t_R output82 (.A(net82),
    .Y(out[120]));
 BUFx3_ASAP7_75t_R output83 (.A(net83),
    .Y(out[1211]));
 BUFx3_ASAP7_75t_R output84 (.A(net84),
    .Y(out[1212]));
 BUFx3_ASAP7_75t_R output85 (.A(net85),
    .Y(out[1213]));
 BUFx3_ASAP7_75t_R output86 (.A(net86),
    .Y(out[1214]));
 BUFx3_ASAP7_75t_R output87 (.A(net87),
    .Y(out[1232]));
 BUFx3_ASAP7_75t_R output88 (.A(net88),
    .Y(out[1233]));
 BUFx3_ASAP7_75t_R output89 (.A(net89),
    .Y(out[1234]));
 BUFx3_ASAP7_75t_R output90 (.A(net90),
    .Y(out[1235]));
 BUFx3_ASAP7_75t_R output91 (.A(net91),
    .Y(out[1236]));
 BUFx3_ASAP7_75t_R output92 (.A(net92),
    .Y(out[1239]));
 BUFx3_ASAP7_75t_R output93 (.A(net93),
    .Y(out[1240]));
 BUFx3_ASAP7_75t_R output94 (.A(net94),
    .Y(out[1250]));
 BUFx3_ASAP7_75t_R output95 (.A(net95),
    .Y(out[1251]));
 BUFx3_ASAP7_75t_R output96 (.A(net96),
    .Y(out[1252]));
 BUFx3_ASAP7_75t_R output97 (.A(net97),
    .Y(out[1253]));
 BUFx3_ASAP7_75t_R output98 (.A(net98),
    .Y(out[1254]));
 BUFx3_ASAP7_75t_R output99 (.A(net99),
    .Y(out[1272]));
 BUFx3_ASAP7_75t_R output100 (.A(net100),
    .Y(out[1273]));
 BUFx3_ASAP7_75t_R output101 (.A(net101),
    .Y(out[1274]));
 BUFx3_ASAP7_75t_R output102 (.A(net102),
    .Y(out[1275]));
 BUFx3_ASAP7_75t_R output103 (.A(net103),
    .Y(out[1276]));
 BUFx3_ASAP7_75t_R output104 (.A(net104),
    .Y(out[1279]));
 BUFx3_ASAP7_75t_R output105 (.A(net105),
    .Y(out[130]));
 BUFx3_ASAP7_75t_R output106 (.A(net106),
    .Y(out[131]));
 BUFx3_ASAP7_75t_R output107 (.A(net107),
    .Y(out[152]));
 BUFx3_ASAP7_75t_R output108 (.A(net108),
    .Y(out[153]));
 BUFx3_ASAP7_75t_R output109 (.A(net109),
    .Y(out[154]));
 BUFx3_ASAP7_75t_R output110 (.A(net110),
    .Y(out[155]));
 BUFx3_ASAP7_75t_R output111 (.A(net111),
    .Y(out[156]));
 BUFx3_ASAP7_75t_R output112 (.A(net112),
    .Y(out[159]));
 BUFx3_ASAP7_75t_R output113 (.A(net113),
    .Y(out[160]));
 BUFx3_ASAP7_75t_R output114 (.A(net114),
    .Y(out[172]));
 BUFx3_ASAP7_75t_R output115 (.A(net115),
    .Y(out[192]));
 BUFx3_ASAP7_75t_R output116 (.A(net116),
    .Y(out[193]));
 BUFx3_ASAP7_75t_R output117 (.A(net117),
    .Y(out[194]));
 BUFx3_ASAP7_75t_R output118 (.A(net118),
    .Y(out[195]));
 BUFx3_ASAP7_75t_R output119 (.A(net119),
    .Y(out[196]));
 BUFx3_ASAP7_75t_R output120 (.A(net120),
    .Y(out[199]));
 BUFx3_ASAP7_75t_R output121 (.A(net121),
    .Y(out[200]));
 BUFx3_ASAP7_75t_R output122 (.A(net122),
    .Y(out[210]));
 BUFx3_ASAP7_75t_R output123 (.A(net123),
    .Y(out[212]));
 BUFx3_ASAP7_75t_R output124 (.A(net124),
    .Y(out[232]));
 BUFx3_ASAP7_75t_R output125 (.A(net125),
    .Y(out[233]));
 BUFx3_ASAP7_75t_R output126 (.A(net126),
    .Y(out[234]));
 BUFx3_ASAP7_75t_R output127 (.A(net127),
    .Y(out[235]));
 BUFx3_ASAP7_75t_R output128 (.A(net128),
    .Y(out[236]));
 BUFx3_ASAP7_75t_R output129 (.A(net129),
    .Y(out[239]));
 BUFx3_ASAP7_75t_R output130 (.A(net130),
    .Y(out[240]));
 BUFx3_ASAP7_75t_R output131 (.A(net131),
    .Y(out[251]));
 BUFx3_ASAP7_75t_R output132 (.A(net132),
    .Y(out[252]));
 BUFx3_ASAP7_75t_R output133 (.A(net133),
    .Y(out[272]));
 BUFx3_ASAP7_75t_R output134 (.A(net134),
    .Y(out[273]));
 BUFx3_ASAP7_75t_R output135 (.A(net135),
    .Y(out[274]));
 BUFx3_ASAP7_75t_R output136 (.A(net136),
    .Y(out[275]));
 BUFx3_ASAP7_75t_R output137 (.A(net137),
    .Y(out[276]));
 BUFx3_ASAP7_75t_R output138 (.A(net138),
    .Y(out[279]));
 BUFx3_ASAP7_75t_R output139 (.A(net139),
    .Y(out[280]));
 BUFx3_ASAP7_75t_R output140 (.A(net140),
    .Y(out[290]));
 BUFx3_ASAP7_75t_R output141 (.A(net141),
    .Y(out[291]));
 BUFx3_ASAP7_75t_R output142 (.A(net142),
    .Y(out[292]));
 BUFx3_ASAP7_75t_R output143 (.A(net143),
    .Y(out[312]));
 BUFx3_ASAP7_75t_R output144 (.A(net144),
    .Y(out[313]));
 BUFx3_ASAP7_75t_R output145 (.A(net145),
    .Y(out[314]));
 BUFx3_ASAP7_75t_R output146 (.A(net146),
    .Y(out[315]));
 BUFx3_ASAP7_75t_R output147 (.A(net147),
    .Y(out[316]));
 BUFx3_ASAP7_75t_R output148 (.A(net148),
    .Y(out[319]));
 BUFx3_ASAP7_75t_R output149 (.A(net149),
    .Y(out[320]));
 BUFx3_ASAP7_75t_R output150 (.A(net150),
    .Y(out[32]));
 BUFx3_ASAP7_75t_R output151 (.A(net151),
    .Y(out[333]));
 BUFx3_ASAP7_75t_R output152 (.A(net152),
    .Y(out[33]));
 BUFx3_ASAP7_75t_R output153 (.A(net153),
    .Y(out[34]));
 BUFx3_ASAP7_75t_R output154 (.A(net154),
    .Y(out[352]));
 BUFx3_ASAP7_75t_R output155 (.A(net155),
    .Y(out[353]));
 BUFx3_ASAP7_75t_R output156 (.A(net156),
    .Y(out[354]));
 BUFx3_ASAP7_75t_R output157 (.A(net157),
    .Y(out[355]));
 BUFx3_ASAP7_75t_R output158 (.A(net158),
    .Y(out[356]));
 BUFx3_ASAP7_75t_R output159 (.A(net159),
    .Y(out[359]));
 BUFx3_ASAP7_75t_R output160 (.A(net160),
    .Y(out[35]));
 BUFx3_ASAP7_75t_R output161 (.A(net161),
    .Y(out[360]));
 BUFx3_ASAP7_75t_R output162 (.A(net162),
    .Y(out[36]));
 BUFx3_ASAP7_75t_R output163 (.A(net163),
    .Y(out[370]));
 BUFx3_ASAP7_75t_R output164 (.A(net164),
    .Y(out[373]));
 BUFx3_ASAP7_75t_R output165 (.A(net165),
    .Y(out[392]));
 BUFx3_ASAP7_75t_R output166 (.A(net166),
    .Y(out[393]));
 BUFx3_ASAP7_75t_R output167 (.A(net167),
    .Y(out[394]));
 BUFx3_ASAP7_75t_R output168 (.A(net168),
    .Y(out[395]));
 BUFx3_ASAP7_75t_R output169 (.A(net169),
    .Y(out[396]));
 BUFx3_ASAP7_75t_R output170 (.A(net170),
    .Y(out[399]));
 BUFx3_ASAP7_75t_R output171 (.A(net171),
    .Y(out[39]));
 BUFx3_ASAP7_75t_R output172 (.A(net172),
    .Y(out[400]));
 BUFx3_ASAP7_75t_R output173 (.A(net173),
    .Y(out[40]));
 BUFx3_ASAP7_75t_R output174 (.A(net174),
    .Y(out[411]));
 BUFx3_ASAP7_75t_R output175 (.A(net175),
    .Y(out[413]));
 BUFx3_ASAP7_75t_R output176 (.A(net176),
    .Y(out[432]));
 BUFx3_ASAP7_75t_R output177 (.A(net177),
    .Y(out[433]));
 BUFx3_ASAP7_75t_R output178 (.A(net178),
    .Y(out[434]));
 BUFx3_ASAP7_75t_R output179 (.A(net179),
    .Y(out[435]));
 BUFx3_ASAP7_75t_R output180 (.A(net180),
    .Y(out[436]));
 BUFx3_ASAP7_75t_R output181 (.A(net181),
    .Y(out[439]));
 BUFx3_ASAP7_75t_R output182 (.A(net182),
    .Y(out[440]));
 BUFx3_ASAP7_75t_R output183 (.A(net183),
    .Y(out[450]));
 BUFx3_ASAP7_75t_R output184 (.A(net184),
    .Y(out[451]));
 BUFx3_ASAP7_75t_R output185 (.A(net185),
    .Y(out[453]));
 BUFx3_ASAP7_75t_R output186 (.A(net186),
    .Y(out[472]));
 BUFx3_ASAP7_75t_R output187 (.A(net187),
    .Y(out[473]));
 BUFx3_ASAP7_75t_R output188 (.A(net188),
    .Y(out[474]));
 BUFx3_ASAP7_75t_R output189 (.A(net189),
    .Y(out[475]));
 BUFx3_ASAP7_75t_R output190 (.A(net190),
    .Y(out[476]));
 BUFx3_ASAP7_75t_R output191 (.A(net191),
    .Y(out[479]));
 BUFx3_ASAP7_75t_R output192 (.A(net192),
    .Y(out[480]));
 BUFx3_ASAP7_75t_R output193 (.A(net193),
    .Y(out[492]));
 BUFx3_ASAP7_75t_R output194 (.A(net194),
    .Y(out[493]));
 BUFx3_ASAP7_75t_R output195 (.A(net195),
    .Y(out[50]));
 BUFx3_ASAP7_75t_R output196 (.A(net196),
    .Y(out[512]));
 BUFx3_ASAP7_75t_R output197 (.A(net197),
    .Y(out[513]));
 BUFx3_ASAP7_75t_R output198 (.A(net198),
    .Y(out[514]));
 BUFx3_ASAP7_75t_R output199 (.A(net199),
    .Y(out[515]));
 BUFx3_ASAP7_75t_R output200 (.A(net200),
    .Y(out[516]));
 BUFx3_ASAP7_75t_R output201 (.A(net201),
    .Y(out[519]));
 BUFx3_ASAP7_75t_R output202 (.A(net202),
    .Y(out[520]));
 BUFx3_ASAP7_75t_R output203 (.A(net203),
    .Y(out[530]));
 BUFx3_ASAP7_75t_R output204 (.A(net204),
    .Y(out[532]));
 BUFx3_ASAP7_75t_R output205 (.A(net205),
    .Y(out[533]));
 BUFx3_ASAP7_75t_R output206 (.A(net206),
    .Y(out[552]));
 BUFx3_ASAP7_75t_R output207 (.A(net207),
    .Y(out[553]));
 BUFx3_ASAP7_75t_R output208 (.A(net208),
    .Y(out[554]));
 BUFx3_ASAP7_75t_R output209 (.A(net209),
    .Y(out[555]));
 BUFx3_ASAP7_75t_R output210 (.A(net210),
    .Y(out[556]));
 BUFx3_ASAP7_75t_R output211 (.A(net211),
    .Y(out[559]));
 BUFx3_ASAP7_75t_R output212 (.A(net212),
    .Y(out[560]));
 BUFx3_ASAP7_75t_R output213 (.A(net213),
    .Y(out[571]));
 BUFx3_ASAP7_75t_R output214 (.A(net214),
    .Y(out[572]));
 BUFx3_ASAP7_75t_R output215 (.A(net215),
    .Y(out[573]));
 BUFx3_ASAP7_75t_R output216 (.A(net216),
    .Y(out[592]));
 BUFx3_ASAP7_75t_R output217 (.A(net217),
    .Y(out[593]));
 BUFx3_ASAP7_75t_R output218 (.A(net218),
    .Y(out[594]));
 BUFx3_ASAP7_75t_R output219 (.A(net219),
    .Y(out[595]));
 BUFx3_ASAP7_75t_R output220 (.A(net220),
    .Y(out[596]));
 BUFx3_ASAP7_75t_R output221 (.A(net221),
    .Y(out[599]));
 BUFx3_ASAP7_75t_R output222 (.A(net222),
    .Y(out[600]));
 BUFx3_ASAP7_75t_R output223 (.A(net223),
    .Y(out[610]));
 BUFx3_ASAP7_75t_R output224 (.A(net224),
    .Y(out[611]));
 BUFx3_ASAP7_75t_R output225 (.A(net225),
    .Y(out[612]));
 BUFx3_ASAP7_75t_R output226 (.A(net226),
    .Y(out[613]));
 BUFx3_ASAP7_75t_R output227 (.A(net227),
    .Y(out[632]));
 BUFx3_ASAP7_75t_R output228 (.A(net228),
    .Y(out[633]));
 BUFx3_ASAP7_75t_R output229 (.A(net229),
    .Y(out[634]));
 BUFx3_ASAP7_75t_R output230 (.A(net230),
    .Y(out[635]));
 BUFx3_ASAP7_75t_R output231 (.A(net231),
    .Y(out[636]));
 BUFx3_ASAP7_75t_R output232 (.A(net232),
    .Y(out[639]));
 BUFx3_ASAP7_75t_R output233 (.A(net233),
    .Y(out[640]));
 BUFx3_ASAP7_75t_R output234 (.A(net234),
    .Y(out[654]));
 BUFx3_ASAP7_75t_R output235 (.A(net235),
    .Y(out[672]));
 BUFx3_ASAP7_75t_R output236 (.A(net236),
    .Y(out[673]));
 BUFx3_ASAP7_75t_R output237 (.A(net237),
    .Y(out[674]));
 BUFx3_ASAP7_75t_R output238 (.A(net238),
    .Y(out[675]));
 BUFx3_ASAP7_75t_R output239 (.A(net239),
    .Y(out[676]));
 BUFx3_ASAP7_75t_R output240 (.A(net240),
    .Y(out[679]));
 BUFx3_ASAP7_75t_R output241 (.A(net241),
    .Y(out[680]));
 BUFx3_ASAP7_75t_R output242 (.A(net242),
    .Y(out[690]));
 BUFx3_ASAP7_75t_R output243 (.A(net243),
    .Y(out[694]));
 BUFx3_ASAP7_75t_R output244 (.A(net244),
    .Y(out[712]));
 BUFx3_ASAP7_75t_R output245 (.A(net245),
    .Y(out[713]));
 BUFx3_ASAP7_75t_R output246 (.A(net246),
    .Y(out[714]));
 BUFx3_ASAP7_75t_R output247 (.A(net247),
    .Y(out[715]));
 BUFx3_ASAP7_75t_R output248 (.A(net248),
    .Y(out[716]));
 BUFx3_ASAP7_75t_R output249 (.A(net249),
    .Y(out[719]));
 BUFx3_ASAP7_75t_R output250 (.A(net250),
    .Y(out[720]));
 BUFx3_ASAP7_75t_R output251 (.A(net251),
    .Y(out[72]));
 BUFx3_ASAP7_75t_R output252 (.A(net252),
    .Y(out[731]));
 BUFx3_ASAP7_75t_R output253 (.A(net253),
    .Y(out[734]));
 BUFx3_ASAP7_75t_R output254 (.A(net254),
    .Y(out[73]));
 BUFx3_ASAP7_75t_R output255 (.A(net255),
    .Y(out[74]));
 BUFx3_ASAP7_75t_R output256 (.A(net256),
    .Y(out[752]));
 BUFx3_ASAP7_75t_R output257 (.A(net257),
    .Y(out[753]));
 BUFx3_ASAP7_75t_R output258 (.A(net258),
    .Y(out[754]));
 BUFx3_ASAP7_75t_R output259 (.A(net259),
    .Y(out[755]));
 BUFx3_ASAP7_75t_R output260 (.A(net260),
    .Y(out[756]));
 BUFx3_ASAP7_75t_R output261 (.A(net261),
    .Y(out[759]));
 BUFx3_ASAP7_75t_R output262 (.A(net262),
    .Y(out[75]));
 BUFx3_ASAP7_75t_R output263 (.A(net263),
    .Y(out[760]));
 BUFx3_ASAP7_75t_R output264 (.A(net264),
    .Y(out[76]));
 BUFx3_ASAP7_75t_R output265 (.A(net265),
    .Y(out[770]));
 BUFx3_ASAP7_75t_R output266 (.A(net266),
    .Y(out[771]));
 BUFx3_ASAP7_75t_R output267 (.A(net267),
    .Y(out[774]));
 BUFx3_ASAP7_75t_R output268 (.A(net268),
    .Y(out[792]));
 BUFx3_ASAP7_75t_R output269 (.A(net269),
    .Y(out[793]));
 BUFx3_ASAP7_75t_R output270 (.A(net270),
    .Y(out[794]));
 BUFx3_ASAP7_75t_R output271 (.A(net271),
    .Y(out[795]));
 BUFx3_ASAP7_75t_R output272 (.A(net272),
    .Y(out[796]));
 BUFx3_ASAP7_75t_R output273 (.A(net273),
    .Y(out[799]));
 BUFx3_ASAP7_75t_R output274 (.A(net274),
    .Y(out[79]));
 BUFx3_ASAP7_75t_R output275 (.A(net275),
    .Y(out[800]));
 BUFx3_ASAP7_75t_R output276 (.A(net276),
    .Y(out[80]));
 BUFx3_ASAP7_75t_R output277 (.A(net277),
    .Y(out[812]));
 BUFx3_ASAP7_75t_R output278 (.A(net278),
    .Y(out[814]));
 BUFx3_ASAP7_75t_R output279 (.A(net279),
    .Y(out[832]));
 BUFx3_ASAP7_75t_R output280 (.A(net280),
    .Y(out[833]));
 BUFx3_ASAP7_75t_R output281 (.A(net281),
    .Y(out[834]));
 BUFx3_ASAP7_75t_R output282 (.A(net282),
    .Y(out[835]));
 BUFx3_ASAP7_75t_R output283 (.A(net283),
    .Y(out[836]));
 BUFx3_ASAP7_75t_R output284 (.A(net284),
    .Y(out[839]));
 BUFx3_ASAP7_75t_R output285 (.A(net285),
    .Y(out[840]));
 BUFx3_ASAP7_75t_R output286 (.A(net286),
    .Y(out[850]));
 BUFx3_ASAP7_75t_R output287 (.A(net287),
    .Y(out[852]));
 BUFx3_ASAP7_75t_R output288 (.A(net288),
    .Y(out[854]));
 BUFx3_ASAP7_75t_R output289 (.A(net289),
    .Y(out[872]));
 BUFx3_ASAP7_75t_R output290 (.A(net290),
    .Y(out[873]));
 BUFx3_ASAP7_75t_R output291 (.A(net291),
    .Y(out[874]));
 BUFx3_ASAP7_75t_R output292 (.A(net292),
    .Y(out[875]));
 BUFx3_ASAP7_75t_R output293 (.A(net293),
    .Y(out[876]));
 BUFx3_ASAP7_75t_R output294 (.A(net294),
    .Y(out[879]));
 BUFx3_ASAP7_75t_R output295 (.A(net295),
    .Y(out[880]));
 BUFx3_ASAP7_75t_R output296 (.A(net296),
    .Y(out[891]));
 BUFx3_ASAP7_75t_R output297 (.A(net297),
    .Y(out[892]));
 BUFx3_ASAP7_75t_R output298 (.A(net298),
    .Y(out[894]));
 BUFx3_ASAP7_75t_R output299 (.A(net299),
    .Y(out[912]));
 BUFx3_ASAP7_75t_R output300 (.A(net300),
    .Y(out[913]));
 BUFx3_ASAP7_75t_R output301 (.A(net301),
    .Y(out[914]));
 BUFx3_ASAP7_75t_R output302 (.A(net302),
    .Y(out[915]));
 BUFx3_ASAP7_75t_R output303 (.A(net303),
    .Y(out[916]));
 BUFx3_ASAP7_75t_R output304 (.A(net304),
    .Y(out[919]));
 BUFx3_ASAP7_75t_R output305 (.A(net305),
    .Y(out[91]));
 BUFx3_ASAP7_75t_R output306 (.A(net306),
    .Y(out[920]));
 BUFx3_ASAP7_75t_R output307 (.A(net307),
    .Y(out[930]));
 BUFx3_ASAP7_75t_R output308 (.A(net308),
    .Y(out[931]));
 BUFx3_ASAP7_75t_R output309 (.A(net309),
    .Y(out[932]));
 BUFx3_ASAP7_75t_R output310 (.A(net310),
    .Y(out[934]));
 BUFx3_ASAP7_75t_R output311 (.A(net311),
    .Y(out[952]));
 BUFx3_ASAP7_75t_R output312 (.A(net312),
    .Y(out[953]));
 BUFx3_ASAP7_75t_R output313 (.A(net313),
    .Y(out[954]));
 BUFx3_ASAP7_75t_R output314 (.A(net314),
    .Y(out[955]));
 BUFx3_ASAP7_75t_R output315 (.A(net315),
    .Y(out[956]));
 BUFx3_ASAP7_75t_R output316 (.A(net316),
    .Y(out[959]));
 BUFx3_ASAP7_75t_R output317 (.A(net317),
    .Y(out[960]));
 BUFx3_ASAP7_75t_R output318 (.A(net318),
    .Y(out[973]));
 BUFx3_ASAP7_75t_R output319 (.A(net319),
    .Y(out[974]));
 BUFx3_ASAP7_75t_R output320 (.A(net320),
    .Y(out[992]));
 BUFx3_ASAP7_75t_R output321 (.A(net321),
    .Y(out[993]));
 BUFx3_ASAP7_75t_R output322 (.A(net322),
    .Y(out[994]));
 BUFx3_ASAP7_75t_R output323 (.A(net323),
    .Y(out[995]));
 BUFx3_ASAP7_75t_R output324 (.A(net324),
    .Y(out[996]));
 BUFx3_ASAP7_75t_R output325 (.A(net325),
    .Y(out[999]));
 TIELOx1_ASAP7_75t_R _21215__326 (.L(net326));
 TIELOx1_ASAP7_75t_R _21216__327 (.L(net327));
 TIELOx1_ASAP7_75t_R _21217__328 (.L(net328));
 TIELOx1_ASAP7_75t_R _21218__329 (.L(net329));
 TIELOx1_ASAP7_75t_R _21219__330 (.L(net330));
 TIELOx1_ASAP7_75t_R _21220__331 (.L(net331));
 TIELOx1_ASAP7_75t_R _21221__332 (.L(net332));
 TIELOx1_ASAP7_75t_R _21222__333 (.L(net333));
 TIELOx1_ASAP7_75t_R _21223__334 (.L(net334));
 TIELOx1_ASAP7_75t_R _21224__335 (.L(net335));
 TIELOx1_ASAP7_75t_R _21225__336 (.L(net336));
 TIELOx1_ASAP7_75t_R _21226__337 (.L(net337));
 TIELOx1_ASAP7_75t_R _21227__338 (.L(net338));
 TIELOx1_ASAP7_75t_R _21228__339 (.L(net339));
 TIELOx1_ASAP7_75t_R _21229__340 (.L(net340));
 TIELOx1_ASAP7_75t_R _21230__341 (.L(net341));
 TIELOx1_ASAP7_75t_R _21231__342 (.L(net342));
 TIELOx1_ASAP7_75t_R _21232__343 (.L(net343));
 TIELOx1_ASAP7_75t_R _21233__344 (.L(net344));
 TIELOx1_ASAP7_75t_R _21234__345 (.L(net345));
 TIELOx1_ASAP7_75t_R _21235__346 (.L(net346));
 TIELOx1_ASAP7_75t_R _21236__347 (.L(net347));
 TIELOx1_ASAP7_75t_R _21237__348 (.L(net348));
 TIELOx1_ASAP7_75t_R _21238__349 (.L(net349));
 TIELOx1_ASAP7_75t_R _21239__350 (.L(net350));
 TIELOx1_ASAP7_75t_R _21240__351 (.L(net351));
 TIELOx1_ASAP7_75t_R _21241__352 (.L(net352));
 TIELOx1_ASAP7_75t_R _21242__353 (.L(net353));
 TIELOx1_ASAP7_75t_R _21243__354 (.L(net354));
 TIELOx1_ASAP7_75t_R _21244__355 (.L(net355));
 TIELOx1_ASAP7_75t_R _21245__356 (.L(net356));
 TIELOx1_ASAP7_75t_R _21246__357 (.L(net357));
 TIELOx1_ASAP7_75t_R _21247__358 (.L(net358));
 TIELOx1_ASAP7_75t_R _21248__359 (.L(net359));
 TIELOx1_ASAP7_75t_R _21249__360 (.L(net360));
 TIELOx1_ASAP7_75t_R _21250__361 (.L(net361));
 TIELOx1_ASAP7_75t_R _21251__362 (.L(net362));
 TIELOx1_ASAP7_75t_R _21252__363 (.L(net363));
 TIELOx1_ASAP7_75t_R _21253__364 (.L(net364));
 TIELOx1_ASAP7_75t_R _21254__365 (.L(net365));
 TIELOx1_ASAP7_75t_R _21255__366 (.L(net366));
 TIELOx1_ASAP7_75t_R _21256__367 (.L(net367));
 TIELOx1_ASAP7_75t_R _21257__368 (.L(net368));
 TIELOx1_ASAP7_75t_R _21258__369 (.L(net369));
 TIELOx1_ASAP7_75t_R _21259__370 (.L(net370));
 TIELOx1_ASAP7_75t_R _21260__371 (.L(net371));
 TIELOx1_ASAP7_75t_R _21261__372 (.L(net372));
 TIELOx1_ASAP7_75t_R _21262__373 (.L(net373));
 TIELOx1_ASAP7_75t_R _21263__374 (.L(net374));
 TIELOx1_ASAP7_75t_R _21264__375 (.L(net375));
 TIELOx1_ASAP7_75t_R _21265__376 (.L(net376));
 TIELOx1_ASAP7_75t_R _21266__377 (.L(net377));
 TIELOx1_ASAP7_75t_R _21267__378 (.L(net378));
 TIELOx1_ASAP7_75t_R _21268__379 (.L(net379));
 TIELOx1_ASAP7_75t_R _21269__380 (.L(net380));
 TIELOx1_ASAP7_75t_R _21270__381 (.L(net381));
 TIELOx1_ASAP7_75t_R _21271__382 (.L(net382));
 TIELOx1_ASAP7_75t_R _21272__383 (.L(net383));
 TIELOx1_ASAP7_75t_R _21273__384 (.L(net384));
 TIELOx1_ASAP7_75t_R _21274__385 (.L(net385));
 TIELOx1_ASAP7_75t_R _21275__386 (.L(net386));
 TIELOx1_ASAP7_75t_R _21276__387 (.L(net387));
 TIELOx1_ASAP7_75t_R _21277__388 (.L(net388));
 TIELOx1_ASAP7_75t_R _21278__389 (.L(net389));
 TIELOx1_ASAP7_75t_R _21279__390 (.L(net390));
 TIELOx1_ASAP7_75t_R _21280__391 (.L(net391));
 TIELOx1_ASAP7_75t_R _21281__392 (.L(net392));
 TIELOx1_ASAP7_75t_R _21282__393 (.L(net393));
 TIELOx1_ASAP7_75t_R _21283__394 (.L(net394));
 TIELOx1_ASAP7_75t_R _21284__395 (.L(net395));
 TIELOx1_ASAP7_75t_R _21285__396 (.L(net396));
 TIELOx1_ASAP7_75t_R _21286__397 (.L(net397));
 TIELOx1_ASAP7_75t_R _21287__398 (.L(net398));
 TIELOx1_ASAP7_75t_R _21288__399 (.L(net399));
 TIELOx1_ASAP7_75t_R _21289__400 (.L(net400));
 TIELOx1_ASAP7_75t_R _21290__401 (.L(net401));
 TIELOx1_ASAP7_75t_R _21291__402 (.L(net402));
 TIELOx1_ASAP7_75t_R _21292__403 (.L(net403));
 TIELOx1_ASAP7_75t_R _21293__404 (.L(net404));
 TIELOx1_ASAP7_75t_R _21294__405 (.L(net405));
 TIELOx1_ASAP7_75t_R _21295__406 (.L(net406));
 TIELOx1_ASAP7_75t_R _21296__407 (.L(net407));
 TIELOx1_ASAP7_75t_R _21297__408 (.L(net408));
 TIELOx1_ASAP7_75t_R _21298__409 (.L(net409));
 TIELOx1_ASAP7_75t_R _21299__410 (.L(net410));
 TIELOx1_ASAP7_75t_R _21300__411 (.L(net411));
 TIELOx1_ASAP7_75t_R _21301__412 (.L(net412));
 TIELOx1_ASAP7_75t_R _21302__413 (.L(net413));
 TIELOx1_ASAP7_75t_R _21303__414 (.L(net414));
 TIELOx1_ASAP7_75t_R _21304__415 (.L(net415));
 TIELOx1_ASAP7_75t_R _21305__416 (.L(net416));
 TIELOx1_ASAP7_75t_R _21306__417 (.L(net417));
 TIELOx1_ASAP7_75t_R _21307__418 (.L(net418));
 TIELOx1_ASAP7_75t_R _21308__419 (.L(net419));
 TIELOx1_ASAP7_75t_R _21309__420 (.L(net420));
 TIELOx1_ASAP7_75t_R _21310__421 (.L(net421));
 TIELOx1_ASAP7_75t_R _21311__422 (.L(net422));
 TIELOx1_ASAP7_75t_R _21312__423 (.L(net423));
 TIELOx1_ASAP7_75t_R _21313__424 (.L(net424));
 TIELOx1_ASAP7_75t_R _21314__425 (.L(net425));
 TIELOx1_ASAP7_75t_R _21315__426 (.L(net426));
 TIELOx1_ASAP7_75t_R _21316__427 (.L(net427));
 TIELOx1_ASAP7_75t_R _21317__428 (.L(net428));
 TIELOx1_ASAP7_75t_R _21318__429 (.L(net429));
 TIELOx1_ASAP7_75t_R _21319__430 (.L(net430));
 TIELOx1_ASAP7_75t_R _21320__431 (.L(net431));
 TIELOx1_ASAP7_75t_R _21321__432 (.L(net432));
 TIELOx1_ASAP7_75t_R _21323__433 (.L(net433));
 TIELOx1_ASAP7_75t_R _21324__434 (.L(net434));
 TIELOx1_ASAP7_75t_R _21325__435 (.L(net435));
 TIELOx1_ASAP7_75t_R _21326__436 (.L(net436));
 TIELOx1_ASAP7_75t_R _21327__437 (.L(net437));
 TIELOx1_ASAP7_75t_R _21328__438 (.L(net438));
 TIELOx1_ASAP7_75t_R _21329__439 (.L(net439));
 TIELOx1_ASAP7_75t_R _21330__440 (.L(net440));
 TIELOx1_ASAP7_75t_R _21331__441 (.L(net441));
 TIELOx1_ASAP7_75t_R _21332__442 (.L(net442));
 TIELOx1_ASAP7_75t_R _21333__443 (.L(net443));
 TIELOx1_ASAP7_75t_R _21334__444 (.L(net444));
 TIELOx1_ASAP7_75t_R _21335__445 (.L(net445));
 TIELOx1_ASAP7_75t_R _21336__446 (.L(net446));
 TIELOx1_ASAP7_75t_R _21337__447 (.L(net447));
 TIELOx1_ASAP7_75t_R _21338__448 (.L(net448));
 TIELOx1_ASAP7_75t_R _21339__449 (.L(net449));
 TIELOx1_ASAP7_75t_R _21340__450 (.L(net450));
 TIELOx1_ASAP7_75t_R _21341__451 (.L(net451));
 TIELOx1_ASAP7_75t_R _21342__452 (.L(net452));
 TIELOx1_ASAP7_75t_R _21343__453 (.L(net453));
 TIELOx1_ASAP7_75t_R _21344__454 (.L(net454));
 TIELOx1_ASAP7_75t_R _21345__455 (.L(net455));
 TIELOx1_ASAP7_75t_R _21346__456 (.L(net456));
 TIELOx1_ASAP7_75t_R _21347__457 (.L(net457));
 TIELOx1_ASAP7_75t_R _21348__458 (.L(net458));
 TIELOx1_ASAP7_75t_R _21349__459 (.L(net459));
 TIELOx1_ASAP7_75t_R _21350__460 (.L(net460));
 TIELOx1_ASAP7_75t_R _21351__461 (.L(net461));
 TIELOx1_ASAP7_75t_R _21352__462 (.L(net462));
 TIELOx1_ASAP7_75t_R _21353__463 (.L(net463));
 TIELOx1_ASAP7_75t_R _21354__464 (.L(net464));
 TIELOx1_ASAP7_75t_R _21355__465 (.L(net465));
 TIELOx1_ASAP7_75t_R _21356__466 (.L(net466));
 TIELOx1_ASAP7_75t_R _21357__467 (.L(net467));
 TIELOx1_ASAP7_75t_R _21358__468 (.L(net468));
 TIELOx1_ASAP7_75t_R _21359__469 (.L(net469));
 TIELOx1_ASAP7_75t_R _21360__470 (.L(net470));
 TIELOx1_ASAP7_75t_R _21361__471 (.L(net471));
 TIELOx1_ASAP7_75t_R _21362__472 (.L(net472));
 TIELOx1_ASAP7_75t_R _21363__473 (.L(net473));
 TIELOx1_ASAP7_75t_R _21364__474 (.L(net474));
 TIELOx1_ASAP7_75t_R _21365__475 (.L(net475));
 TIELOx1_ASAP7_75t_R _21366__476 (.L(net476));
 TIELOx1_ASAP7_75t_R _21367__477 (.L(net477));
 TIELOx1_ASAP7_75t_R _21368__478 (.L(net478));
 TIELOx1_ASAP7_75t_R _21369__479 (.L(net479));
 TIELOx1_ASAP7_75t_R _21370__480 (.L(net480));
 TIELOx1_ASAP7_75t_R _21371__481 (.L(net481));
 TIELOx1_ASAP7_75t_R _21372__482 (.L(net482));
 TIELOx1_ASAP7_75t_R _21373__483 (.L(net483));
 TIELOx1_ASAP7_75t_R _21374__484 (.L(net484));
 TIELOx1_ASAP7_75t_R _21375__485 (.L(net485));
 TIELOx1_ASAP7_75t_R _21376__486 (.L(net486));
 TIELOx1_ASAP7_75t_R _21377__487 (.L(net487));
 TIELOx1_ASAP7_75t_R _21378__488 (.L(net488));
 TIELOx1_ASAP7_75t_R _21379__489 (.L(net489));
 TIELOx1_ASAP7_75t_R _21380__490 (.L(net490));
 TIELOx1_ASAP7_75t_R _21381__491 (.L(net491));
 TIELOx1_ASAP7_75t_R _21382__492 (.L(net492));
 TIELOx1_ASAP7_75t_R _21383__493 (.L(net493));
 TIELOx1_ASAP7_75t_R _21384__494 (.L(net494));
 TIELOx1_ASAP7_75t_R _21385__495 (.L(net495));
 TIELOx1_ASAP7_75t_R _21387__496 (.L(net496));
 TIELOx1_ASAP7_75t_R _21388__497 (.L(net497));
 TIELOx1_ASAP7_75t_R _21389__498 (.L(net498));
 TIELOx1_ASAP7_75t_R _21390__499 (.L(net499));
 TIELOx1_ASAP7_75t_R _21391__500 (.L(net500));
 TIELOx1_ASAP7_75t_R _21392__501 (.L(net501));
 TIELOx1_ASAP7_75t_R _21393__502 (.L(net502));
 TIELOx1_ASAP7_75t_R _21394__503 (.L(net503));
 TIELOx1_ASAP7_75t_R _21395__504 (.L(net504));
 TIELOx1_ASAP7_75t_R _21396__505 (.L(net505));
 TIELOx1_ASAP7_75t_R _21397__506 (.L(net506));
 TIELOx1_ASAP7_75t_R _21398__507 (.L(net507));
 TIELOx1_ASAP7_75t_R _21399__508 (.L(net508));
 TIELOx1_ASAP7_75t_R _21400__509 (.L(net509));
 TIELOx1_ASAP7_75t_R _21401__510 (.L(net510));
 TIELOx1_ASAP7_75t_R _21402__511 (.L(net511));
 TIELOx1_ASAP7_75t_R _21403__512 (.L(net512));
 TIELOx1_ASAP7_75t_R _21404__513 (.L(net513));
 TIELOx1_ASAP7_75t_R _21405__514 (.L(net514));
 TIELOx1_ASAP7_75t_R _21406__515 (.L(net515));
 TIELOx1_ASAP7_75t_R _21407__516 (.L(net516));
 TIELOx1_ASAP7_75t_R _21408__517 (.L(net517));
 TIELOx1_ASAP7_75t_R _21409__518 (.L(net518));
 TIELOx1_ASAP7_75t_R _21410__519 (.L(net519));
 TIELOx1_ASAP7_75t_R _21411__520 (.L(net520));
 TIELOx1_ASAP7_75t_R _21412__521 (.L(net521));
 TIELOx1_ASAP7_75t_R _21413__522 (.L(net522));
 TIELOx1_ASAP7_75t_R _21414__523 (.L(net523));
 TIELOx1_ASAP7_75t_R _21415__524 (.L(net524));
 TIELOx1_ASAP7_75t_R _21416__525 (.L(net525));
 TIELOx1_ASAP7_75t_R _21417__526 (.L(net526));
 TIELOx1_ASAP7_75t_R _21418__527 (.L(net527));
 TIELOx1_ASAP7_75t_R _21420__528 (.L(net528));
 TIELOx1_ASAP7_75t_R _21421__529 (.L(net529));
 TIELOx1_ASAP7_75t_R _21422__530 (.L(net530));
 TIELOx1_ASAP7_75t_R _21423__531 (.L(net531));
 TIELOx1_ASAP7_75t_R _21424__532 (.L(net532));
 TIELOx1_ASAP7_75t_R _21425__533 (.L(net533));
 TIELOx1_ASAP7_75t_R _21426__534 (.L(net534));
 TIELOx1_ASAP7_75t_R _21427__535 (.L(net535));
 TIELOx1_ASAP7_75t_R _21428__536 (.L(net536));
 TIELOx1_ASAP7_75t_R _21429__537 (.L(net537));
 TIELOx1_ASAP7_75t_R _21430__538 (.L(net538));
 TIELOx1_ASAP7_75t_R _21431__539 (.L(net539));
 TIELOx1_ASAP7_75t_R _21432__540 (.L(net540));
 TIELOx1_ASAP7_75t_R _21433__541 (.L(net541));
 TIELOx1_ASAP7_75t_R _21434__542 (.L(net542));
 TIELOx1_ASAP7_75t_R _21435__543 (.L(net543));
 TIELOx1_ASAP7_75t_R _21436__544 (.L(net544));
 TIELOx1_ASAP7_75t_R _21437__545 (.L(net545));
 TIELOx1_ASAP7_75t_R _21438__546 (.L(net546));
 TIELOx1_ASAP7_75t_R _21439__547 (.L(net547));
 TIELOx1_ASAP7_75t_R _21440__548 (.L(net548));
 TIELOx1_ASAP7_75t_R _21441__549 (.L(net549));
 TIELOx1_ASAP7_75t_R _21442__550 (.L(net550));
 TIELOx1_ASAP7_75t_R _21443__551 (.L(net551));
 TIELOx1_ASAP7_75t_R _21444__552 (.L(net552));
 TIELOx1_ASAP7_75t_R _21445__553 (.L(net553));
 TIELOx1_ASAP7_75t_R _21446__554 (.L(net554));
 TIELOx1_ASAP7_75t_R _21447__555 (.L(net555));
 TIELOx1_ASAP7_75t_R _21448__556 (.L(net556));
 TIELOx1_ASAP7_75t_R _21449__557 (.L(net557));
 TIELOx1_ASAP7_75t_R _21452__558 (.L(net558));
 TIELOx1_ASAP7_75t_R _21453__559 (.L(net559));
 TIELOx1_ASAP7_75t_R _21454__560 (.L(net560));
 TIELOx1_ASAP7_75t_R _21455__561 (.L(net561));
 TIELOx1_ASAP7_75t_R _21456__562 (.L(net562));
 TIELOx1_ASAP7_75t_R _21457__563 (.L(net563));
 TIELOx1_ASAP7_75t_R _21458__564 (.L(net564));
 TIELOx1_ASAP7_75t_R _21459__565 (.L(net565));
 TIELOx1_ASAP7_75t_R _21460__566 (.L(net566));
 TIELOx1_ASAP7_75t_R _21461__567 (.L(net567));
 TIELOx1_ASAP7_75t_R _21462__568 (.L(net568));
 TIELOx1_ASAP7_75t_R _21463__569 (.L(net569));
 TIELOx1_ASAP7_75t_R _21464__570 (.L(net570));
 TIELOx1_ASAP7_75t_R _21465__571 (.L(net571));
 TIELOx1_ASAP7_75t_R _21466__572 (.L(net572));
 TIELOx1_ASAP7_75t_R _21467__573 (.L(net573));
 TIELOx1_ASAP7_75t_R _21468__574 (.L(net574));
 TIELOx1_ASAP7_75t_R _21469__575 (.L(net575));
 TIELOx1_ASAP7_75t_R _21470__576 (.L(net576));
 TIELOx1_ASAP7_75t_R _21471__577 (.L(net577));
 TIELOx1_ASAP7_75t_R _21472__578 (.L(net578));
 TIELOx1_ASAP7_75t_R _21473__579 (.L(net579));
 TIELOx1_ASAP7_75t_R _21474__580 (.L(net580));
 TIELOx1_ASAP7_75t_R _21475__581 (.L(net581));
 TIELOx1_ASAP7_75t_R _21476__582 (.L(net582));
 TIELOx1_ASAP7_75t_R _21477__583 (.L(net583));
 TIELOx1_ASAP7_75t_R _21478__584 (.L(net584));
 TIELOx1_ASAP7_75t_R _21479__585 (.L(net585));
 TIELOx1_ASAP7_75t_R _21480__586 (.L(net586));
 TIELOx1_ASAP7_75t_R _21481__587 (.L(net587));
 TIELOx1_ASAP7_75t_R _21482__588 (.L(net588));
 TIELOx1_ASAP7_75t_R _21483__589 (.L(net589));
 TIELOx1_ASAP7_75t_R _21484__590 (.L(net590));
 TIELOx1_ASAP7_75t_R _21485__591 (.L(net591));
 TIELOx1_ASAP7_75t_R _21486__592 (.L(net592));
 TIELOx1_ASAP7_75t_R _21487__593 (.L(net593));
 TIELOx1_ASAP7_75t_R _21488__594 (.L(net594));
 TIELOx1_ASAP7_75t_R _21489__595 (.L(net595));
 TIELOx1_ASAP7_75t_R _21490__596 (.L(net596));
 TIELOx1_ASAP7_75t_R _21491__597 (.L(net597));
 TIELOx1_ASAP7_75t_R _21492__598 (.L(net598));
 TIELOx1_ASAP7_75t_R _21493__599 (.L(net599));
 TIELOx1_ASAP7_75t_R _21494__600 (.L(net600));
 TIELOx1_ASAP7_75t_R _21495__601 (.L(net601));
 TIELOx1_ASAP7_75t_R _21496__602 (.L(net602));
 TIELOx1_ASAP7_75t_R _21497__603 (.L(net603));
 TIELOx1_ASAP7_75t_R _21498__604 (.L(net604));
 TIELOx1_ASAP7_75t_R _21499__605 (.L(net605));
 TIELOx1_ASAP7_75t_R _21500__606 (.L(net606));
 TIELOx1_ASAP7_75t_R _21501__607 (.L(net607));
 TIELOx1_ASAP7_75t_R _21502__608 (.L(net608));
 TIELOx1_ASAP7_75t_R _21503__609 (.L(net609));
 TIELOx1_ASAP7_75t_R _21504__610 (.L(net610));
 TIELOx1_ASAP7_75t_R _21505__611 (.L(net611));
 TIELOx1_ASAP7_75t_R _21506__612 (.L(net612));
 TIELOx1_ASAP7_75t_R _21507__613 (.L(net613));
 TIELOx1_ASAP7_75t_R _21508__614 (.L(net614));
 TIELOx1_ASAP7_75t_R _21509__615 (.L(net615));
 TIELOx1_ASAP7_75t_R _21510__616 (.L(net616));
 TIELOx1_ASAP7_75t_R _21511__617 (.L(net617));
 TIELOx1_ASAP7_75t_R _21512__618 (.L(net618));
 TIELOx1_ASAP7_75t_R _21513__619 (.L(net619));
 TIELOx1_ASAP7_75t_R _21515__620 (.L(net620));
 TIELOx1_ASAP7_75t_R _21516__621 (.L(net621));
 TIELOx1_ASAP7_75t_R _21517__622 (.L(net622));
 TIELOx1_ASAP7_75t_R _21518__623 (.L(net623));
 TIELOx1_ASAP7_75t_R _21519__624 (.L(net624));
 TIELOx1_ASAP7_75t_R _21520__625 (.L(net625));
 TIELOx1_ASAP7_75t_R _21521__626 (.L(net626));
 TIELOx1_ASAP7_75t_R _21522__627 (.L(net627));
 TIELOx1_ASAP7_75t_R _21523__628 (.L(net628));
 TIELOx1_ASAP7_75t_R _21524__629 (.L(net629));
 TIELOx1_ASAP7_75t_R _21525__630 (.L(net630));
 TIELOx1_ASAP7_75t_R _21526__631 (.L(net631));
 TIELOx1_ASAP7_75t_R _21527__632 (.L(net632));
 TIELOx1_ASAP7_75t_R _21528__633 (.L(net633));
 TIELOx1_ASAP7_75t_R _21529__634 (.L(net634));
 TIELOx1_ASAP7_75t_R _21530__635 (.L(net635));
 TIELOx1_ASAP7_75t_R _21531__636 (.L(net636));
 TIELOx1_ASAP7_75t_R _21532__637 (.L(net637));
 TIELOx1_ASAP7_75t_R _21533__638 (.L(net638));
 TIELOx1_ASAP7_75t_R _21534__639 (.L(net639));
 TIELOx1_ASAP7_75t_R _21535__640 (.L(net640));
 TIELOx1_ASAP7_75t_R _21536__641 (.L(net641));
 TIELOx1_ASAP7_75t_R _21537__642 (.L(net642));
 TIELOx1_ASAP7_75t_R _21538__643 (.L(net643));
 TIELOx1_ASAP7_75t_R _21539__644 (.L(net644));
 TIELOx1_ASAP7_75t_R _21540__645 (.L(net645));
 TIELOx1_ASAP7_75t_R _21541__646 (.L(net646));
 TIELOx1_ASAP7_75t_R _21542__647 (.L(net647));
 TIELOx1_ASAP7_75t_R _21543__648 (.L(net648));
 TIELOx1_ASAP7_75t_R _21544__649 (.L(net649));
 TIELOx1_ASAP7_75t_R _21545__650 (.L(net650));
 TIELOx1_ASAP7_75t_R _21546__651 (.L(net651));
 TIELOx1_ASAP7_75t_R _21548__652 (.L(net652));
 TIELOx1_ASAP7_75t_R _21549__653 (.L(net653));
 TIELOx1_ASAP7_75t_R _21550__654 (.L(net654));
 TIELOx1_ASAP7_75t_R _21551__655 (.L(net655));
 TIELOx1_ASAP7_75t_R _21552__656 (.L(net656));
 TIELOx1_ASAP7_75t_R _21553__657 (.L(net657));
 TIELOx1_ASAP7_75t_R _21554__658 (.L(net658));
 TIELOx1_ASAP7_75t_R _21555__659 (.L(net659));
 TIELOx1_ASAP7_75t_R _21556__660 (.L(net660));
 TIELOx1_ASAP7_75t_R _21557__661 (.L(net661));
 TIELOx1_ASAP7_75t_R _21558__662 (.L(net662));
 TIELOx1_ASAP7_75t_R _21559__663 (.L(net663));
 TIELOx1_ASAP7_75t_R _21560__664 (.L(net664));
 TIELOx1_ASAP7_75t_R _21561__665 (.L(net665));
 TIELOx1_ASAP7_75t_R _21562__666 (.L(net666));
 TIELOx1_ASAP7_75t_R _21563__667 (.L(net667));
 TIELOx1_ASAP7_75t_R _21564__668 (.L(net668));
 TIELOx1_ASAP7_75t_R _21565__669 (.L(net669));
 TIELOx1_ASAP7_75t_R _21566__670 (.L(net670));
 TIELOx1_ASAP7_75t_R _21567__671 (.L(net671));
 TIELOx1_ASAP7_75t_R _21568__672 (.L(net672));
 TIELOx1_ASAP7_75t_R _21569__673 (.L(net673));
 TIELOx1_ASAP7_75t_R _21570__674 (.L(net674));
 TIELOx1_ASAP7_75t_R _21571__675 (.L(net675));
 TIELOx1_ASAP7_75t_R _21572__676 (.L(net676));
 TIELOx1_ASAP7_75t_R _21573__677 (.L(net677));
 TIELOx1_ASAP7_75t_R _21574__678 (.L(net678));
 TIELOx1_ASAP7_75t_R _21575__679 (.L(net679));
 TIELOx1_ASAP7_75t_R _21576__680 (.L(net680));
 TIELOx1_ASAP7_75t_R _21577__681 (.L(net681));
 TIELOx1_ASAP7_75t_R _21580__682 (.L(net682));
 TIELOx1_ASAP7_75t_R _21581__683 (.L(net683));
 TIELOx1_ASAP7_75t_R _21582__684 (.L(net684));
 TIELOx1_ASAP7_75t_R _21583__685 (.L(net685));
 TIELOx1_ASAP7_75t_R _21584__686 (.L(net686));
 TIELOx1_ASAP7_75t_R _21585__687 (.L(net687));
 TIELOx1_ASAP7_75t_R _21586__688 (.L(net688));
 TIELOx1_ASAP7_75t_R _21587__689 (.L(net689));
 TIELOx1_ASAP7_75t_R _21588__690 (.L(net690));
 TIELOx1_ASAP7_75t_R _21589__691 (.L(net691));
 TIELOx1_ASAP7_75t_R _21590__692 (.L(net692));
 TIELOx1_ASAP7_75t_R _21591__693 (.L(net693));
 TIELOx1_ASAP7_75t_R _21592__694 (.L(net694));
 TIELOx1_ASAP7_75t_R _21593__695 (.L(net695));
 TIELOx1_ASAP7_75t_R _21594__696 (.L(net696));
 TIELOx1_ASAP7_75t_R _21595__697 (.L(net697));
 TIELOx1_ASAP7_75t_R _21596__698 (.L(net698));
 TIELOx1_ASAP7_75t_R _21597__699 (.L(net699));
 TIELOx1_ASAP7_75t_R _21598__700 (.L(net700));
 TIELOx1_ASAP7_75t_R _21599__701 (.L(net701));
 TIELOx1_ASAP7_75t_R _21600__702 (.L(net702));
 TIELOx1_ASAP7_75t_R _21601__703 (.L(net703));
 TIELOx1_ASAP7_75t_R _21602__704 (.L(net704));
 TIELOx1_ASAP7_75t_R _21603__705 (.L(net705));
 TIELOx1_ASAP7_75t_R _21604__706 (.L(net706));
 TIELOx1_ASAP7_75t_R _21605__707 (.L(net707));
 TIELOx1_ASAP7_75t_R _21606__708 (.L(net708));
 TIELOx1_ASAP7_75t_R _21607__709 (.L(net709));
 TIELOx1_ASAP7_75t_R _21608__710 (.L(net710));
 TIELOx1_ASAP7_75t_R _21609__711 (.L(net711));
 TIELOx1_ASAP7_75t_R _21610__712 (.L(net712));
 TIELOx1_ASAP7_75t_R _21611__713 (.L(net713));
 TIELOx1_ASAP7_75t_R _21613__714 (.L(net714));
 TIELOx1_ASAP7_75t_R _21614__715 (.L(net715));
 TIELOx1_ASAP7_75t_R _21615__716 (.L(net716));
 TIELOx1_ASAP7_75t_R _21616__717 (.L(net717));
 TIELOx1_ASAP7_75t_R _21617__718 (.L(net718));
 TIELOx1_ASAP7_75t_R _21618__719 (.L(net719));
 TIELOx1_ASAP7_75t_R _21619__720 (.L(net720));
 TIELOx1_ASAP7_75t_R _21620__721 (.L(net721));
 TIELOx1_ASAP7_75t_R _21621__722 (.L(net722));
 TIELOx1_ASAP7_75t_R _21622__723 (.L(net723));
 TIELOx1_ASAP7_75t_R _21623__724 (.L(net724));
 TIELOx1_ASAP7_75t_R _21624__725 (.L(net725));
 TIELOx1_ASAP7_75t_R _21625__726 (.L(net726));
 TIELOx1_ASAP7_75t_R _21626__727 (.L(net727));
 TIELOx1_ASAP7_75t_R _21627__728 (.L(net728));
 TIELOx1_ASAP7_75t_R _21628__729 (.L(net729));
 TIELOx1_ASAP7_75t_R _21629__730 (.L(net730));
 TIELOx1_ASAP7_75t_R _21630__731 (.L(net731));
 TIELOx1_ASAP7_75t_R _21631__732 (.L(net732));
 TIELOx1_ASAP7_75t_R _21632__733 (.L(net733));
 TIELOx1_ASAP7_75t_R _21633__734 (.L(net734));
 TIELOx1_ASAP7_75t_R _21634__735 (.L(net735));
 TIELOx1_ASAP7_75t_R _21635__736 (.L(net736));
 TIELOx1_ASAP7_75t_R _21636__737 (.L(net737));
 TIELOx1_ASAP7_75t_R _21637__738 (.L(net738));
 TIELOx1_ASAP7_75t_R _21638__739 (.L(net739));
 TIELOx1_ASAP7_75t_R _21639__740 (.L(net740));
 TIELOx1_ASAP7_75t_R _21640__741 (.L(net741));
 TIELOx1_ASAP7_75t_R _21641__742 (.L(net742));
 TIELOx1_ASAP7_75t_R _21643__743 (.L(net743));
 TIELOx1_ASAP7_75t_R _21645__744 (.L(net744));
 TIELOx1_ASAP7_75t_R _21646__745 (.L(net745));
 TIELOx1_ASAP7_75t_R _21647__746 (.L(net746));
 TIELOx1_ASAP7_75t_R _21648__747 (.L(net747));
 TIELOx1_ASAP7_75t_R _21649__748 (.L(net748));
 TIELOx1_ASAP7_75t_R _21650__749 (.L(net749));
 TIELOx1_ASAP7_75t_R _21651__750 (.L(net750));
 TIELOx1_ASAP7_75t_R _21652__751 (.L(net751));
 TIELOx1_ASAP7_75t_R _21653__752 (.L(net752));
 TIELOx1_ASAP7_75t_R _21654__753 (.L(net753));
 TIELOx1_ASAP7_75t_R _21655__754 (.L(net754));
 TIELOx1_ASAP7_75t_R _21656__755 (.L(net755));
 TIELOx1_ASAP7_75t_R _21657__756 (.L(net756));
 TIELOx1_ASAP7_75t_R _21658__757 (.L(net757));
 TIELOx1_ASAP7_75t_R _21659__758 (.L(net758));
 TIELOx1_ASAP7_75t_R _21660__759 (.L(net759));
 TIELOx1_ASAP7_75t_R _21661__760 (.L(net760));
 TIELOx1_ASAP7_75t_R _21662__761 (.L(net761));
 TIELOx1_ASAP7_75t_R _21663__762 (.L(net762));
 TIELOx1_ASAP7_75t_R _21664__763 (.L(net763));
 TIELOx1_ASAP7_75t_R _21665__764 (.L(net764));
 TIELOx1_ASAP7_75t_R _21666__765 (.L(net765));
 TIELOx1_ASAP7_75t_R _21667__766 (.L(net766));
 TIELOx1_ASAP7_75t_R _21668__767 (.L(net767));
 TIELOx1_ASAP7_75t_R _21669__768 (.L(net768));
 TIELOx1_ASAP7_75t_R _21670__769 (.L(net769));
 TIELOx1_ASAP7_75t_R _21671__770 (.L(net770));
 TIELOx1_ASAP7_75t_R _21672__771 (.L(net771));
 TIELOx1_ASAP7_75t_R _21673__772 (.L(net772));
 TIELOx1_ASAP7_75t_R _21674__773 (.L(net773));
 TIELOx1_ASAP7_75t_R _21677__774 (.L(net774));
 TIELOx1_ASAP7_75t_R _21678__775 (.L(net775));
 TIELOx1_ASAP7_75t_R _21679__776 (.L(net776));
 TIELOx1_ASAP7_75t_R _21680__777 (.L(net777));
 TIELOx1_ASAP7_75t_R _21681__778 (.L(net778));
 TIELOx1_ASAP7_75t_R _21682__779 (.L(net779));
 TIELOx1_ASAP7_75t_R _21683__780 (.L(net780));
 TIELOx1_ASAP7_75t_R _21684__781 (.L(net781));
 TIELOx1_ASAP7_75t_R _21685__782 (.L(net782));
 TIELOx1_ASAP7_75t_R _21686__783 (.L(net783));
 TIELOx1_ASAP7_75t_R _21687__784 (.L(net784));
 TIELOx1_ASAP7_75t_R _21688__785 (.L(net785));
 TIELOx1_ASAP7_75t_R _21689__786 (.L(net786));
 TIELOx1_ASAP7_75t_R _21690__787 (.L(net787));
 TIELOx1_ASAP7_75t_R _21691__788 (.L(net788));
 TIELOx1_ASAP7_75t_R _21692__789 (.L(net789));
 TIELOx1_ASAP7_75t_R _21693__790 (.L(net790));
 TIELOx1_ASAP7_75t_R _21694__791 (.L(net791));
 TIELOx1_ASAP7_75t_R _21695__792 (.L(net792));
 TIELOx1_ASAP7_75t_R _21696__793 (.L(net793));
 TIELOx1_ASAP7_75t_R _21697__794 (.L(net794));
 TIELOx1_ASAP7_75t_R _21698__795 (.L(net795));
 TIELOx1_ASAP7_75t_R _21699__796 (.L(net796));
 TIELOx1_ASAP7_75t_R _21700__797 (.L(net797));
 TIELOx1_ASAP7_75t_R _21701__798 (.L(net798));
 TIELOx1_ASAP7_75t_R _21702__799 (.L(net799));
 TIELOx1_ASAP7_75t_R _21703__800 (.L(net800));
 TIELOx1_ASAP7_75t_R _21704__801 (.L(net801));
 TIELOx1_ASAP7_75t_R _21705__802 (.L(net802));
 TIELOx1_ASAP7_75t_R _21709__803 (.L(net803));
 TIELOx1_ASAP7_75t_R _21710__804 (.L(net804));
 TIELOx1_ASAP7_75t_R _21711__805 (.L(net805));
 TIELOx1_ASAP7_75t_R _21712__806 (.L(net806));
 TIELOx1_ASAP7_75t_R _21713__807 (.L(net807));
 TIELOx1_ASAP7_75t_R _21714__808 (.L(net808));
 TIELOx1_ASAP7_75t_R _21715__809 (.L(net809));
 TIELOx1_ASAP7_75t_R _21716__810 (.L(net810));
 TIELOx1_ASAP7_75t_R _21717__811 (.L(net811));
 TIELOx1_ASAP7_75t_R _21718__812 (.L(net812));
 TIELOx1_ASAP7_75t_R _21719__813 (.L(net813));
 TIELOx1_ASAP7_75t_R _21720__814 (.L(net814));
 TIELOx1_ASAP7_75t_R _21721__815 (.L(net815));
 TIELOx1_ASAP7_75t_R _21722__816 (.L(net816));
 TIELOx1_ASAP7_75t_R _21723__817 (.L(net817));
 TIELOx1_ASAP7_75t_R _21724__818 (.L(net818));
 TIELOx1_ASAP7_75t_R _21725__819 (.L(net819));
 TIELOx1_ASAP7_75t_R _21726__820 (.L(net820));
 TIELOx1_ASAP7_75t_R _21727__821 (.L(net821));
 TIELOx1_ASAP7_75t_R _21728__822 (.L(net822));
 TIELOx1_ASAP7_75t_R _21729__823 (.L(net823));
 TIELOx1_ASAP7_75t_R _21730__824 (.L(net824));
 TIELOx1_ASAP7_75t_R _21731__825 (.L(net825));
 TIELOx1_ASAP7_75t_R _21732__826 (.L(net826));
 TIELOx1_ASAP7_75t_R _21733__827 (.L(net827));
 TIELOx1_ASAP7_75t_R _21734__828 (.L(net828));
 TIELOx1_ASAP7_75t_R _21735__829 (.L(net829));
 TIELOx1_ASAP7_75t_R _21736__830 (.L(net830));
 TIELOx1_ASAP7_75t_R _21737__831 (.L(net831));
 TIELOx1_ASAP7_75t_R _21738__832 (.L(net832));
 TIELOx1_ASAP7_75t_R _21739__833 (.L(net833));
 TIELOx1_ASAP7_75t_R _21740__834 (.L(net834));
 TIELOx1_ASAP7_75t_R _21741__835 (.L(net835));
 TIELOx1_ASAP7_75t_R _21742__836 (.L(net836));
 TIELOx1_ASAP7_75t_R _21743__837 (.L(net837));
 TIELOx1_ASAP7_75t_R _21744__838 (.L(net838));
 TIELOx1_ASAP7_75t_R _21745__839 (.L(net839));
 TIELOx1_ASAP7_75t_R _21746__840 (.L(net840));
 TIELOx1_ASAP7_75t_R _21747__841 (.L(net841));
 TIELOx1_ASAP7_75t_R _21748__842 (.L(net842));
 TIELOx1_ASAP7_75t_R _21749__843 (.L(net843));
 TIELOx1_ASAP7_75t_R _21750__844 (.L(net844));
 TIELOx1_ASAP7_75t_R _21751__845 (.L(net845));
 TIELOx1_ASAP7_75t_R _21752__846 (.L(net846));
 TIELOx1_ASAP7_75t_R _21753__847 (.L(net847));
 TIELOx1_ASAP7_75t_R _21754__848 (.L(net848));
 TIELOx1_ASAP7_75t_R _21755__849 (.L(net849));
 TIELOx1_ASAP7_75t_R _21756__850 (.L(net850));
 TIELOx1_ASAP7_75t_R _21757__851 (.L(net851));
 TIELOx1_ASAP7_75t_R _21758__852 (.L(net852));
 TIELOx1_ASAP7_75t_R _21759__853 (.L(net853));
 TIELOx1_ASAP7_75t_R _21760__854 (.L(net854));
 TIELOx1_ASAP7_75t_R _21761__855 (.L(net855));
 TIELOx1_ASAP7_75t_R _21762__856 (.L(net856));
 TIELOx1_ASAP7_75t_R _21763__857 (.L(net857));
 TIELOx1_ASAP7_75t_R _21764__858 (.L(net858));
 TIELOx1_ASAP7_75t_R _21765__859 (.L(net859));
 TIELOx1_ASAP7_75t_R _21766__860 (.L(net860));
 TIELOx1_ASAP7_75t_R _21767__861 (.L(net861));
 TIELOx1_ASAP7_75t_R _21768__862 (.L(net862));
 TIELOx1_ASAP7_75t_R _21769__863 (.L(net863));
 TIELOx1_ASAP7_75t_R _21771__864 (.L(net864));
 TIELOx1_ASAP7_75t_R _21772__865 (.L(net865));
 TIELOx1_ASAP7_75t_R _21773__866 (.L(net866));
 TIELOx1_ASAP7_75t_R _21774__867 (.L(net867));
 TIELOx1_ASAP7_75t_R _21775__868 (.L(net868));
 TIELOx1_ASAP7_75t_R _21776__869 (.L(net869));
 TIELOx1_ASAP7_75t_R _21777__870 (.L(net870));
 TIELOx1_ASAP7_75t_R _21778__871 (.L(net871));
 TIELOx1_ASAP7_75t_R _21779__872 (.L(net872));
 TIELOx1_ASAP7_75t_R _21780__873 (.L(net873));
 TIELOx1_ASAP7_75t_R _21781__874 (.L(net874));
 TIELOx1_ASAP7_75t_R _21782__875 (.L(net875));
 TIELOx1_ASAP7_75t_R _21783__876 (.L(net876));
 TIELOx1_ASAP7_75t_R _21784__877 (.L(net877));
 TIELOx1_ASAP7_75t_R _21785__878 (.L(net878));
 TIELOx1_ASAP7_75t_R _21786__879 (.L(net879));
 TIELOx1_ASAP7_75t_R _21787__880 (.L(net880));
 TIELOx1_ASAP7_75t_R _21788__881 (.L(net881));
 TIELOx1_ASAP7_75t_R _21789__882 (.L(net882));
 TIELOx1_ASAP7_75t_R _21790__883 (.L(net883));
 TIELOx1_ASAP7_75t_R _21791__884 (.L(net884));
 TIELOx1_ASAP7_75t_R _21792__885 (.L(net885));
 TIELOx1_ASAP7_75t_R _21793__886 (.L(net886));
 TIELOx1_ASAP7_75t_R _21794__887 (.L(net887));
 TIELOx1_ASAP7_75t_R _21795__888 (.L(net888));
 TIELOx1_ASAP7_75t_R _21796__889 (.L(net889));
 TIELOx1_ASAP7_75t_R _21797__890 (.L(net890));
 TIELOx1_ASAP7_75t_R _21798__891 (.L(net891));
 TIELOx1_ASAP7_75t_R _21799__892 (.L(net892));
 TIELOx1_ASAP7_75t_R _21800__893 (.L(net893));
 TIELOx1_ASAP7_75t_R _21801__894 (.L(net894));
 TIELOx1_ASAP7_75t_R _21802__895 (.L(net895));
 TIELOx1_ASAP7_75t_R _21804__896 (.L(net896));
 TIELOx1_ASAP7_75t_R _21805__897 (.L(net897));
 TIELOx1_ASAP7_75t_R _21806__898 (.L(net898));
 TIELOx1_ASAP7_75t_R _21807__899 (.L(net899));
 TIELOx1_ASAP7_75t_R _21808__900 (.L(net900));
 TIELOx1_ASAP7_75t_R _21809__901 (.L(net901));
 TIELOx1_ASAP7_75t_R _21810__902 (.L(net902));
 TIELOx1_ASAP7_75t_R _21811__903 (.L(net903));
 TIELOx1_ASAP7_75t_R _21812__904 (.L(net904));
 TIELOx1_ASAP7_75t_R _21813__905 (.L(net905));
 TIELOx1_ASAP7_75t_R _21814__906 (.L(net906));
 TIELOx1_ASAP7_75t_R _21815__907 (.L(net907));
 TIELOx1_ASAP7_75t_R _21816__908 (.L(net908));
 TIELOx1_ASAP7_75t_R _21817__909 (.L(net909));
 TIELOx1_ASAP7_75t_R _21818__910 (.L(net910));
 TIELOx1_ASAP7_75t_R _21819__911 (.L(net911));
 TIELOx1_ASAP7_75t_R _21820__912 (.L(net912));
 TIELOx1_ASAP7_75t_R _21821__913 (.L(net913));
 TIELOx1_ASAP7_75t_R _21822__914 (.L(net914));
 TIELOx1_ASAP7_75t_R _21823__915 (.L(net915));
 TIELOx1_ASAP7_75t_R _21824__916 (.L(net916));
 TIELOx1_ASAP7_75t_R _21825__917 (.L(net917));
 TIELOx1_ASAP7_75t_R _21826__918 (.L(net918));
 TIELOx1_ASAP7_75t_R _21827__919 (.L(net919));
 TIELOx1_ASAP7_75t_R _21828__920 (.L(net920));
 TIELOx1_ASAP7_75t_R _21829__921 (.L(net921));
 TIELOx1_ASAP7_75t_R _21830__922 (.L(net922));
 TIELOx1_ASAP7_75t_R _21831__923 (.L(net923));
 TIELOx1_ASAP7_75t_R _21832__924 (.L(net924));
 TIELOx1_ASAP7_75t_R _21833__925 (.L(net925));
 TIELOx1_ASAP7_75t_R _21836__926 (.L(net926));
 TIELOx1_ASAP7_75t_R _21837__927 (.L(net927));
 TIELOx1_ASAP7_75t_R _21838__928 (.L(net928));
 TIELOx1_ASAP7_75t_R _21839__929 (.L(net929));
 TIELOx1_ASAP7_75t_R _21840__930 (.L(net930));
 TIELOx1_ASAP7_75t_R _21841__931 (.L(net931));
 TIELOx1_ASAP7_75t_R _21842__932 (.L(net932));
 TIELOx1_ASAP7_75t_R _21843__933 (.L(net933));
 TIELOx1_ASAP7_75t_R _21844__934 (.L(net934));
 TIELOx1_ASAP7_75t_R _21845__935 (.L(net935));
 TIELOx1_ASAP7_75t_R _21846__936 (.L(net936));
 TIELOx1_ASAP7_75t_R _21847__937 (.L(net937));
 TIELOx1_ASAP7_75t_R _21848__938 (.L(net938));
 TIELOx1_ASAP7_75t_R _21849__939 (.L(net939));
 TIELOx1_ASAP7_75t_R _21850__940 (.L(net940));
 TIELOx1_ASAP7_75t_R _21851__941 (.L(net941));
 TIELOx1_ASAP7_75t_R _21852__942 (.L(net942));
 TIELOx1_ASAP7_75t_R _21853__943 (.L(net943));
 TIELOx1_ASAP7_75t_R _21854__944 (.L(net944));
 TIELOx1_ASAP7_75t_R _21855__945 (.L(net945));
 TIELOx1_ASAP7_75t_R _21856__946 (.L(net946));
 TIELOx1_ASAP7_75t_R _21857__947 (.L(net947));
 TIELOx1_ASAP7_75t_R _21858__948 (.L(net948));
 TIELOx1_ASAP7_75t_R _21859__949 (.L(net949));
 TIELOx1_ASAP7_75t_R _21860__950 (.L(net950));
 TIELOx1_ASAP7_75t_R _21861__951 (.L(net951));
 TIELOx1_ASAP7_75t_R _21862__952 (.L(net952));
 TIELOx1_ASAP7_75t_R _21863__953 (.L(net953));
 TIELOx1_ASAP7_75t_R _21864__954 (.L(net954));
 TIELOx1_ASAP7_75t_R _21865__955 (.L(net955));
 TIELOx1_ASAP7_75t_R _21866__956 (.L(net956));
 TIELOx1_ASAP7_75t_R _21867__957 (.L(net957));
 TIELOx1_ASAP7_75t_R _21869__958 (.L(net958));
 TIELOx1_ASAP7_75t_R _21870__959 (.L(net959));
 TIELOx1_ASAP7_75t_R _21871__960 (.L(net960));
 TIELOx1_ASAP7_75t_R _21872__961 (.L(net961));
 TIELOx1_ASAP7_75t_R _21873__962 (.L(net962));
 TIELOx1_ASAP7_75t_R _21874__963 (.L(net963));
 TIELOx1_ASAP7_75t_R _21875__964 (.L(net964));
 TIELOx1_ASAP7_75t_R _21876__965 (.L(net965));
 TIELOx1_ASAP7_75t_R _21877__966 (.L(net966));
 TIELOx1_ASAP7_75t_R _21878__967 (.L(net967));
 TIELOx1_ASAP7_75t_R _21879__968 (.L(net968));
 TIELOx1_ASAP7_75t_R _21880__969 (.L(net969));
 TIELOx1_ASAP7_75t_R _21881__970 (.L(net970));
 TIELOx1_ASAP7_75t_R _21882__971 (.L(net971));
 TIELOx1_ASAP7_75t_R _21883__972 (.L(net972));
 TIELOx1_ASAP7_75t_R _21884__973 (.L(net973));
 TIELOx1_ASAP7_75t_R _21885__974 (.L(net974));
 TIELOx1_ASAP7_75t_R _21886__975 (.L(net975));
 TIELOx1_ASAP7_75t_R _21887__976 (.L(net976));
 TIELOx1_ASAP7_75t_R _21888__977 (.L(net977));
 TIELOx1_ASAP7_75t_R _21889__978 (.L(net978));
 TIELOx1_ASAP7_75t_R _21890__979 (.L(net979));
 TIELOx1_ASAP7_75t_R _21891__980 (.L(net980));
 TIELOx1_ASAP7_75t_R _21892__981 (.L(net981));
 TIELOx1_ASAP7_75t_R _21893__982 (.L(net982));
 TIELOx1_ASAP7_75t_R _21894__983 (.L(net983));
 TIELOx1_ASAP7_75t_R _21895__984 (.L(net984));
 TIELOx1_ASAP7_75t_R _21896__985 (.L(net985));
 TIELOx1_ASAP7_75t_R _21897__986 (.L(net986));
 TIELOx1_ASAP7_75t_R _21899__987 (.L(net987));
 TIELOx1_ASAP7_75t_R _21901__988 (.L(net988));
 TIELOx1_ASAP7_75t_R _21902__989 (.L(net989));
 TIELOx1_ASAP7_75t_R _21903__990 (.L(net990));
 TIELOx1_ASAP7_75t_R _21904__991 (.L(net991));
 TIELOx1_ASAP7_75t_R _21905__992 (.L(net992));
 TIELOx1_ASAP7_75t_R _21906__993 (.L(net993));
 TIELOx1_ASAP7_75t_R _21907__994 (.L(net994));
 TIELOx1_ASAP7_75t_R _21908__995 (.L(net995));
 TIELOx1_ASAP7_75t_R _21909__996 (.L(net996));
 TIELOx1_ASAP7_75t_R _21910__997 (.L(net997));
 TIELOx1_ASAP7_75t_R _21911__998 (.L(net998));
 TIELOx1_ASAP7_75t_R _21912__999 (.L(net999));
 TIELOx1_ASAP7_75t_R _21913__1000 (.L(net1000));
 TIELOx1_ASAP7_75t_R _21914__1001 (.L(net1001));
 TIELOx1_ASAP7_75t_R _21915__1002 (.L(net1002));
 TIELOx1_ASAP7_75t_R _21916__1003 (.L(net1003));
 TIELOx1_ASAP7_75t_R _21917__1004 (.L(net1004));
 TIELOx1_ASAP7_75t_R _21918__1005 (.L(net1005));
 TIELOx1_ASAP7_75t_R _21919__1006 (.L(net1006));
 TIELOx1_ASAP7_75t_R _21920__1007 (.L(net1007));
 TIELOx1_ASAP7_75t_R _21921__1008 (.L(net1008));
 TIELOx1_ASAP7_75t_R _21922__1009 (.L(net1009));
 TIELOx1_ASAP7_75t_R _21923__1010 (.L(net1010));
 TIELOx1_ASAP7_75t_R _21924__1011 (.L(net1011));
 TIELOx1_ASAP7_75t_R _21925__1012 (.L(net1012));
 TIELOx1_ASAP7_75t_R _21926__1013 (.L(net1013));
 TIELOx1_ASAP7_75t_R _21927__1014 (.L(net1014));
 TIELOx1_ASAP7_75t_R _21928__1015 (.L(net1015));
 TIELOx1_ASAP7_75t_R _21929__1016 (.L(net1016));
 TIELOx1_ASAP7_75t_R _21930__1017 (.L(net1017));
 TIELOx1_ASAP7_75t_R _21933__1018 (.L(net1018));
 TIELOx1_ASAP7_75t_R _21934__1019 (.L(net1019));
 TIELOx1_ASAP7_75t_R _21935__1020 (.L(net1020));
 TIELOx1_ASAP7_75t_R _21936__1021 (.L(net1021));
 TIELOx1_ASAP7_75t_R _21937__1022 (.L(net1022));
 TIELOx1_ASAP7_75t_R _21938__1023 (.L(net1023));
 TIELOx1_ASAP7_75t_R _21939__1024 (.L(net1024));
 TIELOx1_ASAP7_75t_R _21940__1025 (.L(net1025));
 TIELOx1_ASAP7_75t_R _21941__1026 (.L(net1026));
 TIELOx1_ASAP7_75t_R _21942__1027 (.L(net1027));
 TIELOx1_ASAP7_75t_R _21943__1028 (.L(net1028));
 TIELOx1_ASAP7_75t_R _21944__1029 (.L(net1029));
 TIELOx1_ASAP7_75t_R _21945__1030 (.L(net1030));
 TIELOx1_ASAP7_75t_R _21946__1031 (.L(net1031));
 TIELOx1_ASAP7_75t_R _21947__1032 (.L(net1032));
 TIELOx1_ASAP7_75t_R _21948__1033 (.L(net1033));
 TIELOx1_ASAP7_75t_R _21949__1034 (.L(net1034));
 TIELOx1_ASAP7_75t_R _21950__1035 (.L(net1035));
 TIELOx1_ASAP7_75t_R _21951__1036 (.L(net1036));
 TIELOx1_ASAP7_75t_R _21952__1037 (.L(net1037));
 TIELOx1_ASAP7_75t_R _21953__1038 (.L(net1038));
 TIELOx1_ASAP7_75t_R _21954__1039 (.L(net1039));
 TIELOx1_ASAP7_75t_R _21955__1040 (.L(net1040));
 TIELOx1_ASAP7_75t_R _21956__1041 (.L(net1041));
 TIELOx1_ASAP7_75t_R _21957__1042 (.L(net1042));
 TIELOx1_ASAP7_75t_R _21958__1043 (.L(net1043));
 TIELOx1_ASAP7_75t_R _21959__1044 (.L(net1044));
 TIELOx1_ASAP7_75t_R _21960__1045 (.L(net1045));
 TIELOx1_ASAP7_75t_R _21961__1046 (.L(net1046));
 TIELOx1_ASAP7_75t_R _21965__1047 (.L(net1047));
 TIELOx1_ASAP7_75t_R _21966__1048 (.L(net1048));
 TIELOx1_ASAP7_75t_R _21967__1049 (.L(net1049));
 TIELOx1_ASAP7_75t_R _21968__1050 (.L(net1050));
 TIELOx1_ASAP7_75t_R _21969__1051 (.L(net1051));
 TIELOx1_ASAP7_75t_R _21970__1052 (.L(net1052));
 TIELOx1_ASAP7_75t_R _21971__1053 (.L(net1053));
 TIELOx1_ASAP7_75t_R _21972__1054 (.L(net1054));
 TIELOx1_ASAP7_75t_R _21973__1055 (.L(net1055));
 TIELOx1_ASAP7_75t_R _21974__1056 (.L(net1056));
 TIELOx1_ASAP7_75t_R _21975__1057 (.L(net1057));
 TIELOx1_ASAP7_75t_R _21976__1058 (.L(net1058));
 TIELOx1_ASAP7_75t_R _21977__1059 (.L(net1059));
 TIELOx1_ASAP7_75t_R _21978__1060 (.L(net1060));
 TIELOx1_ASAP7_75t_R _21979__1061 (.L(net1061));
 TIELOx1_ASAP7_75t_R _21980__1062 (.L(net1062));
 TIELOx1_ASAP7_75t_R _21981__1063 (.L(net1063));
 TIELOx1_ASAP7_75t_R _21982__1064 (.L(net1064));
 TIELOx1_ASAP7_75t_R _21983__1065 (.L(net1065));
 TIELOx1_ASAP7_75t_R _21984__1066 (.L(net1066));
 TIELOx1_ASAP7_75t_R _21985__1067 (.L(net1067));
 TIELOx1_ASAP7_75t_R _21986__1068 (.L(net1068));
 TIELOx1_ASAP7_75t_R _21987__1069 (.L(net1069));
 TIELOx1_ASAP7_75t_R _21988__1070 (.L(net1070));
 TIELOx1_ASAP7_75t_R _21989__1071 (.L(net1071));
 TIELOx1_ASAP7_75t_R _21990__1072 (.L(net1072));
 TIELOx1_ASAP7_75t_R _21991__1073 (.L(net1073));
 TIELOx1_ASAP7_75t_R _21992__1074 (.L(net1074));
 TIELOx1_ASAP7_75t_R _21993__1075 (.L(net1075));
 TIELOx1_ASAP7_75t_R _21994__1076 (.L(net1076));
 TIELOx1_ASAP7_75t_R _21995__1077 (.L(net1077));
 TIELOx1_ASAP7_75t_R _21996__1078 (.L(net1078));
 TIELOx1_ASAP7_75t_R _21998__1079 (.L(net1079));
 TIELOx1_ASAP7_75t_R _21999__1080 (.L(net1080));
 TIELOx1_ASAP7_75t_R _22000__1081 (.L(net1081));
 TIELOx1_ASAP7_75t_R _22001__1082 (.L(net1082));
 TIELOx1_ASAP7_75t_R _22002__1083 (.L(net1083));
 TIELOx1_ASAP7_75t_R _22003__1084 (.L(net1084));
 TIELOx1_ASAP7_75t_R _22004__1085 (.L(net1085));
 TIELOx1_ASAP7_75t_R _22005__1086 (.L(net1086));
 TIELOx1_ASAP7_75t_R _22006__1087 (.L(net1087));
 TIELOx1_ASAP7_75t_R _22007__1088 (.L(net1088));
 TIELOx1_ASAP7_75t_R _22008__1089 (.L(net1089));
 TIELOx1_ASAP7_75t_R _22009__1090 (.L(net1090));
 TIELOx1_ASAP7_75t_R _22010__1091 (.L(net1091));
 TIELOx1_ASAP7_75t_R _22011__1092 (.L(net1092));
 TIELOx1_ASAP7_75t_R _22012__1093 (.L(net1093));
 TIELOx1_ASAP7_75t_R _22013__1094 (.L(net1094));
 TIELOx1_ASAP7_75t_R _22014__1095 (.L(net1095));
 TIELOx1_ASAP7_75t_R _22015__1096 (.L(net1096));
 TIELOx1_ASAP7_75t_R _22016__1097 (.L(net1097));
 TIELOx1_ASAP7_75t_R _22017__1098 (.L(net1098));
 TIELOx1_ASAP7_75t_R _22018__1099 (.L(net1099));
 TIELOx1_ASAP7_75t_R _22019__1100 (.L(net1100));
 TIELOx1_ASAP7_75t_R _22020__1101 (.L(net1101));
 TIELOx1_ASAP7_75t_R _22021__1102 (.L(net1102));
 TIELOx1_ASAP7_75t_R _22022__1103 (.L(net1103));
 TIELOx1_ASAP7_75t_R _22023__1104 (.L(net1104));
 TIELOx1_ASAP7_75t_R _22024__1105 (.L(net1105));
 TIELOx1_ASAP7_75t_R _22025__1106 (.L(net1106));
 TIELOx1_ASAP7_75t_R _22027__1107 (.L(net1107));
 TIELOx1_ASAP7_75t_R _22028__1108 (.L(net1108));
 TIELOx1_ASAP7_75t_R _22030__1109 (.L(net1109));
 TIELOx1_ASAP7_75t_R _22031__1110 (.L(net1110));
 TIELOx1_ASAP7_75t_R _22032__1111 (.L(net1111));
 TIELOx1_ASAP7_75t_R _22033__1112 (.L(net1112));
 TIELOx1_ASAP7_75t_R _22034__1113 (.L(net1113));
 TIELOx1_ASAP7_75t_R _22035__1114 (.L(net1114));
 TIELOx1_ASAP7_75t_R _22036__1115 (.L(net1115));
 TIELOx1_ASAP7_75t_R _22037__1116 (.L(net1116));
 TIELOx1_ASAP7_75t_R _22038__1117 (.L(net1117));
 TIELOx1_ASAP7_75t_R _22039__1118 (.L(net1118));
 TIELOx1_ASAP7_75t_R _22040__1119 (.L(net1119));
 TIELOx1_ASAP7_75t_R _22041__1120 (.L(net1120));
 TIELOx1_ASAP7_75t_R _22042__1121 (.L(net1121));
 TIELOx1_ASAP7_75t_R _22043__1122 (.L(net1122));
 TIELOx1_ASAP7_75t_R _22044__1123 (.L(net1123));
 TIELOx1_ASAP7_75t_R _22045__1124 (.L(net1124));
 TIELOx1_ASAP7_75t_R _22046__1125 (.L(net1125));
 TIELOx1_ASAP7_75t_R _22047__1126 (.L(net1126));
 TIELOx1_ASAP7_75t_R _22048__1127 (.L(net1127));
 TIELOx1_ASAP7_75t_R _22049__1128 (.L(net1128));
 TIELOx1_ASAP7_75t_R _22050__1129 (.L(net1129));
 TIELOx1_ASAP7_75t_R _22051__1130 (.L(net1130));
 TIELOx1_ASAP7_75t_R _22052__1131 (.L(net1131));
 TIELOx1_ASAP7_75t_R _22053__1132 (.L(net1132));
 TIELOx1_ASAP7_75t_R _22054__1133 (.L(net1133));
 TIELOx1_ASAP7_75t_R _22055__1134 (.L(net1134));
 TIELOx1_ASAP7_75t_R _22056__1135 (.L(net1135));
 TIELOx1_ASAP7_75t_R _22057__1136 (.L(net1136));
 TIELOx1_ASAP7_75t_R _22058__1137 (.L(net1137));
 TIELOx1_ASAP7_75t_R _22060__1138 (.L(net1138));
 TIELOx1_ASAP7_75t_R _22062__1139 (.L(net1139));
 TIELOx1_ASAP7_75t_R _22063__1140 (.L(net1140));
 TIELOx1_ASAP7_75t_R _22064__1141 (.L(net1141));
 TIELOx1_ASAP7_75t_R _22065__1142 (.L(net1142));
 TIELOx1_ASAP7_75t_R _22066__1143 (.L(net1143));
 TIELOx1_ASAP7_75t_R _22067__1144 (.L(net1144));
 TIELOx1_ASAP7_75t_R _22068__1145 (.L(net1145));
 TIELOx1_ASAP7_75t_R _22069__1146 (.L(net1146));
 TIELOx1_ASAP7_75t_R _22070__1147 (.L(net1147));
 TIELOx1_ASAP7_75t_R _22071__1148 (.L(net1148));
 TIELOx1_ASAP7_75t_R _22072__1149 (.L(net1149));
 TIELOx1_ASAP7_75t_R _22073__1150 (.L(net1150));
 TIELOx1_ASAP7_75t_R _22074__1151 (.L(net1151));
 TIELOx1_ASAP7_75t_R _22075__1152 (.L(net1152));
 TIELOx1_ASAP7_75t_R _22076__1153 (.L(net1153));
 TIELOx1_ASAP7_75t_R _22077__1154 (.L(net1154));
 TIELOx1_ASAP7_75t_R _22078__1155 (.L(net1155));
 TIELOx1_ASAP7_75t_R _22079__1156 (.L(net1156));
 TIELOx1_ASAP7_75t_R _22080__1157 (.L(net1157));
 TIELOx1_ASAP7_75t_R _22081__1158 (.L(net1158));
 TIELOx1_ASAP7_75t_R _22082__1159 (.L(net1159));
 TIELOx1_ASAP7_75t_R _22083__1160 (.L(net1160));
 TIELOx1_ASAP7_75t_R _22084__1161 (.L(net1161));
 TIELOx1_ASAP7_75t_R _22085__1162 (.L(net1162));
 TIELOx1_ASAP7_75t_R _22086__1163 (.L(net1163));
 TIELOx1_ASAP7_75t_R _22087__1164 (.L(net1164));
 TIELOx1_ASAP7_75t_R _22088__1165 (.L(net1165));
 TIELOx1_ASAP7_75t_R _22089__1166 (.L(net1166));
 TIELOx1_ASAP7_75t_R _22092__1167 (.L(net1167));
 TIELOx1_ASAP7_75t_R _22094__1168 (.L(net1168));
 TIELOx1_ASAP7_75t_R _22095__1169 (.L(net1169));
 TIELOx1_ASAP7_75t_R _22096__1170 (.L(net1170));
 TIELOx1_ASAP7_75t_R _22097__1171 (.L(net1171));
 TIELOx1_ASAP7_75t_R _22098__1172 (.L(net1172));
 TIELOx1_ASAP7_75t_R _22099__1173 (.L(net1173));
 TIELOx1_ASAP7_75t_R _22100__1174 (.L(net1174));
 TIELOx1_ASAP7_75t_R _22101__1175 (.L(net1175));
 TIELOx1_ASAP7_75t_R _22102__1176 (.L(net1176));
 TIELOx1_ASAP7_75t_R _22103__1177 (.L(net1177));
 TIELOx1_ASAP7_75t_R _22104__1178 (.L(net1178));
 TIELOx1_ASAP7_75t_R _22105__1179 (.L(net1179));
 TIELOx1_ASAP7_75t_R _22106__1180 (.L(net1180));
 TIELOx1_ASAP7_75t_R _22107__1181 (.L(net1181));
 TIELOx1_ASAP7_75t_R _22108__1182 (.L(net1182));
 TIELOx1_ASAP7_75t_R _22109__1183 (.L(net1183));
 TIELOx1_ASAP7_75t_R _22110__1184 (.L(net1184));
 TIELOx1_ASAP7_75t_R _22111__1185 (.L(net1185));
 TIELOx1_ASAP7_75t_R _22112__1186 (.L(net1186));
 TIELOx1_ASAP7_75t_R _22113__1187 (.L(net1187));
 TIELOx1_ASAP7_75t_R _22114__1188 (.L(net1188));
 TIELOx1_ASAP7_75t_R _22115__1189 (.L(net1189));
 TIELOx1_ASAP7_75t_R _22116__1190 (.L(net1190));
 TIELOx1_ASAP7_75t_R _22117__1191 (.L(net1191));
 TIELOx1_ASAP7_75t_R _22118__1192 (.L(net1192));
 TIELOx1_ASAP7_75t_R _22119__1193 (.L(net1193));
 TIELOx1_ASAP7_75t_R _22120__1194 (.L(net1194));
 TIELOx1_ASAP7_75t_R _22121__1195 (.L(net1195));
 TIELOx1_ASAP7_75t_R _22122__1196 (.L(net1196));
 TIELOx1_ASAP7_75t_R _22123__1197 (.L(net1197));
 TIELOx1_ASAP7_75t_R _22126__1198 (.L(net1198));
 TIELOx1_ASAP7_75t_R _22127__1199 (.L(net1199));
 TIELOx1_ASAP7_75t_R _22128__1200 (.L(net1200));
 TIELOx1_ASAP7_75t_R _22129__1201 (.L(net1201));
 TIELOx1_ASAP7_75t_R _22130__1202 (.L(net1202));
 TIELOx1_ASAP7_75t_R _22131__1203 (.L(net1203));
 TIELOx1_ASAP7_75t_R _22132__1204 (.L(net1204));
 TIELOx1_ASAP7_75t_R _22133__1205 (.L(net1205));
 TIELOx1_ASAP7_75t_R _22134__1206 (.L(net1206));
 TIELOx1_ASAP7_75t_R _22135__1207 (.L(net1207));
 TIELOx1_ASAP7_75t_R _22136__1208 (.L(net1208));
 TIELOx1_ASAP7_75t_R _22137__1209 (.L(net1209));
 TIELOx1_ASAP7_75t_R _22138__1210 (.L(net1210));
 TIELOx1_ASAP7_75t_R _22139__1211 (.L(net1211));
 TIELOx1_ASAP7_75t_R _22140__1212 (.L(net1212));
 TIELOx1_ASAP7_75t_R _22141__1213 (.L(net1213));
 TIELOx1_ASAP7_75t_R _22142__1214 (.L(net1214));
 TIELOx1_ASAP7_75t_R _22143__1215 (.L(net1215));
 TIELOx1_ASAP7_75t_R _22144__1216 (.L(net1216));
 TIELOx1_ASAP7_75t_R _22145__1217 (.L(net1217));
 TIELOx1_ASAP7_75t_R _22146__1218 (.L(net1218));
 TIELOx1_ASAP7_75t_R _22147__1219 (.L(net1219));
 TIELOx1_ASAP7_75t_R _22148__1220 (.L(net1220));
 TIELOx1_ASAP7_75t_R _22149__1221 (.L(net1221));
 TIELOx1_ASAP7_75t_R _22150__1222 (.L(net1222));
 TIELOx1_ASAP7_75t_R _22151__1223 (.L(net1223));
 TIELOx1_ASAP7_75t_R _22152__1224 (.L(net1224));
 TIELOx1_ASAP7_75t_R _22153__1225 (.L(net1225));
 TIELOx1_ASAP7_75t_R _22155__1226 (.L(net1226));
 TIELOx1_ASAP7_75t_R _22158__1227 (.L(net1227));
 TIELOx1_ASAP7_75t_R _22159__1228 (.L(net1228));
 TIELOx1_ASAP7_75t_R _22160__1229 (.L(net1229));
 TIELOx1_ASAP7_75t_R _22161__1230 (.L(net1230));
 TIELOx1_ASAP7_75t_R _22162__1231 (.L(net1231));
 TIELOx1_ASAP7_75t_R _22163__1232 (.L(net1232));
 TIELOx1_ASAP7_75t_R _22164__1233 (.L(net1233));
 TIELOx1_ASAP7_75t_R _22165__1234 (.L(net1234));
 TIELOx1_ASAP7_75t_R _22166__1235 (.L(net1235));
 TIELOx1_ASAP7_75t_R _22167__1236 (.L(net1236));
 TIELOx1_ASAP7_75t_R _22168__1237 (.L(net1237));
 TIELOx1_ASAP7_75t_R _22169__1238 (.L(net1238));
 TIELOx1_ASAP7_75t_R _22170__1239 (.L(net1239));
 TIELOx1_ASAP7_75t_R _22171__1240 (.L(net1240));
 TIELOx1_ASAP7_75t_R _22172__1241 (.L(net1241));
 TIELOx1_ASAP7_75t_R _22173__1242 (.L(net1242));
 TIELOx1_ASAP7_75t_R _22174__1243 (.L(net1243));
 TIELOx1_ASAP7_75t_R _22175__1244 (.L(net1244));
 TIELOx1_ASAP7_75t_R _22176__1245 (.L(net1245));
 TIELOx1_ASAP7_75t_R _22177__1246 (.L(net1246));
 TIELOx1_ASAP7_75t_R _22178__1247 (.L(net1247));
 TIELOx1_ASAP7_75t_R _22179__1248 (.L(net1248));
 TIELOx1_ASAP7_75t_R _22180__1249 (.L(net1249));
 TIELOx1_ASAP7_75t_R _22181__1250 (.L(net1250));
 TIELOx1_ASAP7_75t_R _22182__1251 (.L(net1251));
 TIELOx1_ASAP7_75t_R _22183__1252 (.L(net1252));
 TIELOx1_ASAP7_75t_R _22184__1253 (.L(net1253));
 TIELOx1_ASAP7_75t_R _22185__1254 (.L(net1254));
 TIELOx1_ASAP7_75t_R _22186__1255 (.L(net1255));
 TIELOx1_ASAP7_75t_R _22190__1256 (.L(net1256));
 TIELOx1_ASAP7_75t_R _22191__1257 (.L(net1257));
 TIELOx1_ASAP7_75t_R _22192__1258 (.L(net1258));
 TIELOx1_ASAP7_75t_R _22193__1259 (.L(net1259));
 TIELOx1_ASAP7_75t_R _22194__1260 (.L(net1260));
 TIELOx1_ASAP7_75t_R _22195__1261 (.L(net1261));
 TIELOx1_ASAP7_75t_R _22196__1262 (.L(net1262));
 TIELOx1_ASAP7_75t_R _22197__1263 (.L(net1263));
 TIELOx1_ASAP7_75t_R _22198__1264 (.L(net1264));
 TIELOx1_ASAP7_75t_R _22199__1265 (.L(net1265));
 TIELOx1_ASAP7_75t_R _22200__1266 (.L(net1266));
 TIELOx1_ASAP7_75t_R _22201__1267 (.L(net1267));
 TIELOx1_ASAP7_75t_R _22202__1268 (.L(net1268));
 TIELOx1_ASAP7_75t_R _22203__1269 (.L(net1269));
 TIELOx1_ASAP7_75t_R _22204__1270 (.L(net1270));
 TIELOx1_ASAP7_75t_R _22205__1271 (.L(net1271));
 TIELOx1_ASAP7_75t_R _22206__1272 (.L(net1272));
 TIELOx1_ASAP7_75t_R _22207__1273 (.L(net1273));
 TIELOx1_ASAP7_75t_R _22208__1274 (.L(net1274));
 TIELOx1_ASAP7_75t_R _22209__1275 (.L(net1275));
 TIELOx1_ASAP7_75t_R _22210__1276 (.L(net1276));
 TIELOx1_ASAP7_75t_R _22211__1277 (.L(net1277));
 TIELOx1_ASAP7_75t_R _22212__1278 (.L(net1278));
 TIELOx1_ASAP7_75t_R _22213__1279 (.L(net1279));
 TIELOx1_ASAP7_75t_R _22214__1280 (.L(net1280));
 TIELOx1_ASAP7_75t_R _22215__1281 (.L(net1281));
 TIELOx1_ASAP7_75t_R _22216__1282 (.L(net1282));
 TIELOx1_ASAP7_75t_R _22217__1283 (.L(net1283));
 TIELOx1_ASAP7_75t_R _22222__1284 (.L(net1284));
 TIELOx1_ASAP7_75t_R _22223__1285 (.L(net1285));
 TIELOx1_ASAP7_75t_R _22224__1286 (.L(net1286));
 TIELOx1_ASAP7_75t_R _22225__1287 (.L(net1287));
 TIELOx1_ASAP7_75t_R _22226__1288 (.L(net1288));
 TIELOx1_ASAP7_75t_R _22227__1289 (.L(net1289));
 TIELOx1_ASAP7_75t_R _22228__1290 (.L(net1290));
 TIELOx1_ASAP7_75t_R _22229__1291 (.L(net1291));
 TIELOx1_ASAP7_75t_R _22230__1292 (.L(net1292));
 TIELOx1_ASAP7_75t_R _22231__1293 (.L(net1293));
 TIELOx1_ASAP7_75t_R _22232__1294 (.L(net1294));
 TIELOx1_ASAP7_75t_R _22233__1295 (.L(net1295));
 TIELOx1_ASAP7_75t_R _22234__1296 (.L(net1296));
 TIELOx1_ASAP7_75t_R _22235__1297 (.L(net1297));
 TIELOx1_ASAP7_75t_R _22236__1298 (.L(net1298));
 TIELOx1_ASAP7_75t_R _22237__1299 (.L(net1299));
 TIELOx1_ASAP7_75t_R _22238__1300 (.L(net1300));
 TIELOx1_ASAP7_75t_R _22239__1301 (.L(net1301));
 TIELOx1_ASAP7_75t_R _22240__1302 (.L(net1302));
 BUFx24_ASAP7_75t_R clkbuf_leaf_1_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_1_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_2_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_2_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_3_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_3_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_4_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_4_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_5_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_5_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_6_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_6_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_7_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_7_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_8_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_8_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_9_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_9_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_10_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_10_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_11_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_11_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_12_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_12_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_13_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_13_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_14_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_14_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_15_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_15_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_16_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_16_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_17_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_17_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_18_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_18_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_19_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_19_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_20_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_20_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_21_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_21_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_22_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_22_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_23_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_23_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_24_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_24_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_25_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_25_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_26_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_26_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_27_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_27_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_28_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_28_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_29_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_29_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_30_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_30_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_31_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_31_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_32_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_32_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_33_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_33_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_34_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_34_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_35_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_35_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_36_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_36_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_37_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_37_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_38_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_38_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_39_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_39_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_40_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_40_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_41_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_41_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_42_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_42_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_43_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_43_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_44_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_44_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_45_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_45_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_46_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_46_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_47_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_47_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_48_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_48_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_49_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_49_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_50_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_50_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_51_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_51_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_52_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_52_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_53_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_53_clk));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_0_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_1_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_2_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_3_0_clk));
 BUFx24_ASAP7_75t_R clkload0 (.A(clknet_2_0_0_clk));
 BUFx24_ASAP7_75t_R clkload1 (.A(clknet_2_2_0_clk));
 INVxp33_ASAP7_75t_R clkload2 (.A(clknet_leaf_0_clk));
 INVxp33_ASAP7_75t_R clkload3 (.A(clknet_leaf_1_clk));
 INVxp33_ASAP7_75t_R clkload4 (.A(clknet_leaf_3_clk));
 INVxp33_ASAP7_75t_R clkload5 (.A(clknet_leaf_4_clk));
 INVxp33_ASAP7_75t_R clkload6 (.A(clknet_leaf_5_clk));
 INVxp33_ASAP7_75t_R clkload7 (.A(clknet_leaf_47_clk));
 INVxp33_ASAP7_75t_R clkload8 (.A(clknet_leaf_48_clk));
 INVxp33_ASAP7_75t_R clkload9 (.A(clknet_leaf_49_clk));
 INVxp33_ASAP7_75t_R clkload10 (.A(clknet_leaf_50_clk));
 INVxp33_ASAP7_75t_R clkload11 (.A(clknet_leaf_51_clk));
 INVxp33_ASAP7_75t_R clkload12 (.A(clknet_leaf_52_clk));
 INVx3_ASAP7_75t_R clkload13 (.A(clknet_leaf_53_clk));
 INVxp33_ASAP7_75t_R clkload14 (.A(clknet_leaf_33_clk));
 INVxp33_ASAP7_75t_R clkload15 (.A(clknet_leaf_35_clk));
 INVxp33_ASAP7_75t_R clkload16 (.A(clknet_leaf_37_clk));
 INVxp33_ASAP7_75t_R clkload17 (.A(clknet_leaf_38_clk));
 INVxp33_ASAP7_75t_R clkload18 (.A(clknet_leaf_39_clk));
 CKINVDCx20_ASAP7_75t_R clkload19 (.A(clknet_leaf_40_clk));
 INVxp33_ASAP7_75t_R clkload20 (.A(clknet_leaf_41_clk));
 INVxp33_ASAP7_75t_R clkload21 (.A(clknet_leaf_42_clk));
 INVxp33_ASAP7_75t_R clkload22 (.A(clknet_leaf_43_clk));
 INVxp33_ASAP7_75t_R clkload23 (.A(clknet_leaf_44_clk));
 INVxp33_ASAP7_75t_R clkload24 (.A(clknet_leaf_45_clk));
 INVxp33_ASAP7_75t_R clkload25 (.A(clknet_leaf_46_clk));
 INVxp33_ASAP7_75t_R clkload26 (.A(clknet_leaf_6_clk));
 INVxp33_ASAP7_75t_R clkload27 (.A(clknet_leaf_7_clk));
 INVxp33_ASAP7_75t_R clkload28 (.A(clknet_leaf_8_clk));
 INVxp33_ASAP7_75t_R clkload29 (.A(clknet_leaf_9_clk));
 CKINVDCx12_ASAP7_75t_R clkload30 (.A(clknet_leaf_11_clk));
 INVxp33_ASAP7_75t_R clkload31 (.A(clknet_leaf_12_clk));
 INVxp33_ASAP7_75t_R clkload32 (.A(clknet_leaf_14_clk));
 INVxp33_ASAP7_75t_R clkload33 (.A(clknet_leaf_15_clk));
 INVxp33_ASAP7_75t_R clkload34 (.A(clknet_leaf_16_clk));
 INVxp33_ASAP7_75t_R clkload35 (.A(clknet_leaf_17_clk));
 INVxp33_ASAP7_75t_R clkload36 (.A(clknet_leaf_18_clk));
 INVxp33_ASAP7_75t_R clkload37 (.A(clknet_leaf_20_clk));
 INVxp33_ASAP7_75t_R clkload38 (.A(clknet_leaf_21_clk));
 INVxp33_ASAP7_75t_R clkload39 (.A(clknet_leaf_22_clk));
 INVxp33_ASAP7_75t_R clkload40 (.A(clknet_leaf_23_clk));
 INVxp33_ASAP7_75t_R clkload41 (.A(clknet_leaf_24_clk));
 CKINVDCx20_ASAP7_75t_R clkload42 (.A(clknet_leaf_25_clk));
 INVxp33_ASAP7_75t_R clkload43 (.A(clknet_leaf_26_clk));
 INVxp33_ASAP7_75t_R clkload44 (.A(clknet_leaf_28_clk));
 INVxp33_ASAP7_75t_R clkload45 (.A(clknet_leaf_29_clk));
 INVxp33_ASAP7_75t_R clkload46 (.A(clknet_leaf_32_clk));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_337 ();
 DECAPx10_ASAP7_75t_R FILLER_0_344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_388 ();
 DECAPx2_ASAP7_75t_R FILLER_0_410 ();
 FILLER_ASAP7_75t_R FILLER_0_416 ();
 DECAPx4_ASAP7_75t_R FILLER_0_424 ();
 FILLER_ASAP7_75t_R FILLER_0_440 ();
 FILLER_ASAP7_75t_R FILLER_0_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_483 ();
 FILLER_ASAP7_75t_R FILLER_0_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_539 ();
 DECAPx2_ASAP7_75t_R FILLER_0_546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_586 ();
 DECAPx2_ASAP7_75t_R FILLER_0_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_617 ();
 FILLER_ASAP7_75t_R FILLER_0_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_646 ();
 FILLER_ASAP7_75t_R FILLER_0_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_662 ();
 FILLER_ASAP7_75t_R FILLER_0_669 ();
 FILLER_ASAP7_75t_R FILLER_0_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_696 ();
 FILLER_ASAP7_75t_R FILLER_0_707 ();
 FILLER_ASAP7_75t_R FILLER_0_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_724 ();
 FILLER_ASAP7_75t_R FILLER_0_759 ();
 FILLER_ASAP7_75t_R FILLER_0_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_791 ();
 FILLER_ASAP7_75t_R FILLER_0_795 ();
 FILLER_ASAP7_75t_R FILLER_0_808 ();
 FILLER_ASAP7_75t_R FILLER_0_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_841 ();
 FILLER_ASAP7_75t_R FILLER_0_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_865 ();
 FILLER_ASAP7_75t_R FILLER_0_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_876 ();
 FILLER_ASAP7_75t_R FILLER_0_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_888 ();
 FILLER_ASAP7_75t_R FILLER_0_902 ();
 FILLER_ASAP7_75t_R FILLER_0_914 ();
 FILLER_ASAP7_75t_R FILLER_0_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_928 ();
 FILLER_ASAP7_75t_R FILLER_0_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_967 ();
 FILLER_ASAP7_75t_R FILLER_0_1018 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_1135 ();
 FILLER_ASAP7_75t_R FILLER_0_1153 ();
 FILLER_ASAP7_75t_R FILLER_0_1168 ();
 FILLER_ASAP7_75t_R FILLER_0_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1188 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1215 ();
 FILLER_ASAP7_75t_R FILLER_0_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_1_112 ();
 DECAPx10_ASAP7_75t_R FILLER_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_1_156 ();
 DECAPx10_ASAP7_75t_R FILLER_1_178 ();
 DECAPx10_ASAP7_75t_R FILLER_1_200 ();
 DECAPx10_ASAP7_75t_R FILLER_1_222 ();
 DECAPx10_ASAP7_75t_R FILLER_1_244 ();
 DECAPx10_ASAP7_75t_R FILLER_1_266 ();
 DECAPx10_ASAP7_75t_R FILLER_1_288 ();
 DECAPx1_ASAP7_75t_R FILLER_1_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_314 ();
 FILLER_ASAP7_75t_R FILLER_1_333 ();
 DECAPx10_ASAP7_75t_R FILLER_1_341 ();
 DECAPx10_ASAP7_75t_R FILLER_1_363 ();
 DECAPx10_ASAP7_75t_R FILLER_1_385 ();
 DECAPx10_ASAP7_75t_R FILLER_1_407 ();
 DECAPx10_ASAP7_75t_R FILLER_1_429 ();
 DECAPx6_ASAP7_75t_R FILLER_1_457 ();
 DECAPx2_ASAP7_75t_R FILLER_1_471 ();
 FILLER_ASAP7_75t_R FILLER_1_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_507 ();
 DECAPx10_ASAP7_75t_R FILLER_1_520 ();
 DECAPx4_ASAP7_75t_R FILLER_1_542 ();
 FILLER_ASAP7_75t_R FILLER_1_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_554 ();
 DECAPx10_ASAP7_75t_R FILLER_1_561 ();
 DECAPx10_ASAP7_75t_R FILLER_1_583 ();
 DECAPx4_ASAP7_75t_R FILLER_1_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_615 ();
 DECAPx1_ASAP7_75t_R FILLER_1_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_640 ();
 DECAPx1_ASAP7_75t_R FILLER_1_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_673 ();
 DECAPx1_ASAP7_75t_R FILLER_1_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_684 ();
 FILLER_ASAP7_75t_R FILLER_1_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_718 ();
 DECAPx1_ASAP7_75t_R FILLER_1_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_728 ();
 FILLER_ASAP7_75t_R FILLER_1_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_734 ();
 FILLER_ASAP7_75t_R FILLER_1_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_758 ();
 FILLER_ASAP7_75t_R FILLER_1_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_847 ();
 DECAPx1_ASAP7_75t_R FILLER_1_880 ();
 FILLER_ASAP7_75t_R FILLER_1_895 ();
 FILLER_ASAP7_75t_R FILLER_1_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_930 ();
 FILLER_ASAP7_75t_R FILLER_1_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_947 ();
 FILLER_ASAP7_75t_R FILLER_1_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_968 ();
 FILLER_ASAP7_75t_R FILLER_1_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1008 ();
 FILLER_ASAP7_75t_R FILLER_1_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1042 ();
 FILLER_ASAP7_75t_R FILLER_1_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_1_1080 ();
 FILLER_ASAP7_75t_R FILLER_1_1094 ();
 FILLER_ASAP7_75t_R FILLER_1_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_1_1129 ();
 FILLER_ASAP7_75t_R FILLER_1_1138 ();
 FILLER_ASAP7_75t_R FILLER_1_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_1_1151 ();
 FILLER_ASAP7_75t_R FILLER_1_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_1_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_1_1185 ();
 FILLER_ASAP7_75t_R FILLER_1_1192 ();
 DECAPx6_ASAP7_75t_R FILLER_1_1199 ();
 FILLER_ASAP7_75t_R FILLER_1_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_2_112 ();
 DECAPx10_ASAP7_75t_R FILLER_2_134 ();
 DECAPx10_ASAP7_75t_R FILLER_2_156 ();
 DECAPx10_ASAP7_75t_R FILLER_2_178 ();
 DECAPx10_ASAP7_75t_R FILLER_2_200 ();
 DECAPx10_ASAP7_75t_R FILLER_2_222 ();
 DECAPx10_ASAP7_75t_R FILLER_2_244 ();
 DECAPx10_ASAP7_75t_R FILLER_2_266 ();
 DECAPx10_ASAP7_75t_R FILLER_2_288 ();
 DECAPx6_ASAP7_75t_R FILLER_2_310 ();
 DECAPx10_ASAP7_75t_R FILLER_2_330 ();
 DECAPx10_ASAP7_75t_R FILLER_2_352 ();
 DECAPx10_ASAP7_75t_R FILLER_2_374 ();
 DECAPx10_ASAP7_75t_R FILLER_2_396 ();
 DECAPx10_ASAP7_75t_R FILLER_2_418 ();
 DECAPx10_ASAP7_75t_R FILLER_2_440 ();
 DECAPx2_ASAP7_75t_R FILLER_2_464 ();
 FILLER_ASAP7_75t_R FILLER_2_470 ();
 DECAPx10_ASAP7_75t_R FILLER_2_489 ();
 DECAPx10_ASAP7_75t_R FILLER_2_511 ();
 DECAPx10_ASAP7_75t_R FILLER_2_533 ();
 DECAPx10_ASAP7_75t_R FILLER_2_555 ();
 DECAPx10_ASAP7_75t_R FILLER_2_577 ();
 DECAPx10_ASAP7_75t_R FILLER_2_599 ();
 DECAPx4_ASAP7_75t_R FILLER_2_621 ();
 FILLER_ASAP7_75t_R FILLER_2_631 ();
 DECAPx6_ASAP7_75t_R FILLER_2_636 ();
 FILLER_ASAP7_75t_R FILLER_2_653 ();
 DECAPx1_ASAP7_75t_R FILLER_2_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_667 ();
 DECAPx10_ASAP7_75t_R FILLER_2_673 ();
 DECAPx4_ASAP7_75t_R FILLER_2_695 ();
 FILLER_ASAP7_75t_R FILLER_2_705 ();
 DECAPx4_ASAP7_75t_R FILLER_2_724 ();
 FILLER_ASAP7_75t_R FILLER_2_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_736 ();
 FILLER_ASAP7_75t_R FILLER_2_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_774 ();
 FILLER_ASAP7_75t_R FILLER_2_789 ();
 FILLER_ASAP7_75t_R FILLER_2_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_811 ();
 DECAPx1_ASAP7_75t_R FILLER_2_815 ();
 FILLER_ASAP7_75t_R FILLER_2_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_839 ();
 DECAPx1_ASAP7_75t_R FILLER_2_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_850 ();
 DECAPx1_ASAP7_75t_R FILLER_2_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_868 ();
 DECAPx2_ASAP7_75t_R FILLER_2_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_883 ();
 DECAPx2_ASAP7_75t_R FILLER_2_889 ();
 FILLER_ASAP7_75t_R FILLER_2_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_897 ();
 FILLER_ASAP7_75t_R FILLER_2_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_922 ();
 FILLER_ASAP7_75t_R FILLER_2_931 ();
 FILLER_ASAP7_75t_R FILLER_2_941 ();
 FILLER_ASAP7_75t_R FILLER_2_946 ();
 FILLER_ASAP7_75t_R FILLER_2_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_957 ();
 DECAPx2_ASAP7_75t_R FILLER_2_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_972 ();
 DECAPx2_ASAP7_75t_R FILLER_2_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_995 ();
 DECAPx6_ASAP7_75t_R FILLER_2_999 ();
 FILLER_ASAP7_75t_R FILLER_2_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1031 ();
 FILLER_ASAP7_75t_R FILLER_2_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1050 ();
 FILLER_ASAP7_75t_R FILLER_2_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_2_1080 ();
 FILLER_ASAP7_75t_R FILLER_2_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1097 ();
 DECAPx1_ASAP7_75t_R FILLER_2_1103 ();
 FILLER_ASAP7_75t_R FILLER_2_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1125 ();
 DECAPx1_ASAP7_75t_R FILLER_2_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_2_1155 ();
 FILLER_ASAP7_75t_R FILLER_2_1166 ();
 FILLER_ASAP7_75t_R FILLER_2_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1205 ();
 FILLER_ASAP7_75t_R FILLER_2_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_3_112 ();
 DECAPx10_ASAP7_75t_R FILLER_3_134 ();
 DECAPx10_ASAP7_75t_R FILLER_3_156 ();
 DECAPx10_ASAP7_75t_R FILLER_3_178 ();
 DECAPx10_ASAP7_75t_R FILLER_3_200 ();
 DECAPx10_ASAP7_75t_R FILLER_3_222 ();
 DECAPx10_ASAP7_75t_R FILLER_3_244 ();
 DECAPx10_ASAP7_75t_R FILLER_3_266 ();
 DECAPx10_ASAP7_75t_R FILLER_3_288 ();
 DECAPx10_ASAP7_75t_R FILLER_3_310 ();
 DECAPx10_ASAP7_75t_R FILLER_3_332 ();
 DECAPx10_ASAP7_75t_R FILLER_3_354 ();
 DECAPx10_ASAP7_75t_R FILLER_3_376 ();
 DECAPx10_ASAP7_75t_R FILLER_3_398 ();
 DECAPx10_ASAP7_75t_R FILLER_3_420 ();
 DECAPx6_ASAP7_75t_R FILLER_3_442 ();
 DECAPx1_ASAP7_75t_R FILLER_3_456 ();
 DECAPx10_ASAP7_75t_R FILLER_3_480 ();
 DECAPx10_ASAP7_75t_R FILLER_3_502 ();
 DECAPx10_ASAP7_75t_R FILLER_3_524 ();
 DECAPx10_ASAP7_75t_R FILLER_3_546 ();
 DECAPx1_ASAP7_75t_R FILLER_3_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_572 ();
 DECAPx10_ASAP7_75t_R FILLER_3_584 ();
 DECAPx10_ASAP7_75t_R FILLER_3_606 ();
 DECAPx6_ASAP7_75t_R FILLER_3_628 ();
 DECAPx2_ASAP7_75t_R FILLER_3_642 ();
 DECAPx6_ASAP7_75t_R FILLER_3_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_667 ();
 DECAPx10_ASAP7_75t_R FILLER_3_686 ();
 FILLER_ASAP7_75t_R FILLER_3_708 ();
 FILLER_ASAP7_75t_R FILLER_3_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_717 ();
 DECAPx10_ASAP7_75t_R FILLER_3_721 ();
 DECAPx6_ASAP7_75t_R FILLER_3_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_757 ();
 DECAPx2_ASAP7_75t_R FILLER_3_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_767 ();
 FILLER_ASAP7_75t_R FILLER_3_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_819 ();
 FILLER_ASAP7_75t_R FILLER_3_823 ();
 FILLER_ASAP7_75t_R FILLER_3_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_835 ();
 DECAPx1_ASAP7_75t_R FILLER_3_846 ();
 DECAPx6_ASAP7_75t_R FILLER_3_853 ();
 DECAPx2_ASAP7_75t_R FILLER_3_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_882 ();
 DECAPx6_ASAP7_75t_R FILLER_3_888 ();
 FILLER_ASAP7_75t_R FILLER_3_902 ();
 DECAPx6_ASAP7_75t_R FILLER_3_907 ();
 FILLER_ASAP7_75t_R FILLER_3_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_923 ();
 DECAPx6_ASAP7_75t_R FILLER_3_926 ();
 DECAPx2_ASAP7_75t_R FILLER_3_940 ();
 FILLER_ASAP7_75t_R FILLER_3_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_951 ();
 DECAPx10_ASAP7_75t_R FILLER_3_957 ();
 DECAPx10_ASAP7_75t_R FILLER_3_979 ();
 DECAPx1_ASAP7_75t_R FILLER_3_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1019 ();
 FILLER_ASAP7_75t_R FILLER_3_1028 ();
 DECAPx2_ASAP7_75t_R FILLER_3_1035 ();
 DECAPx4_ASAP7_75t_R FILLER_3_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_3_1060 ();
 FILLER_ASAP7_75t_R FILLER_3_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_3_1081 ();
 FILLER_ASAP7_75t_R FILLER_3_1087 ();
 FILLER_ASAP7_75t_R FILLER_3_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_3_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_3_1115 ();
 FILLER_ASAP7_75t_R FILLER_3_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1129 ();
 FILLER_ASAP7_75t_R FILLER_3_1133 ();
 FILLER_ASAP7_75t_R FILLER_3_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_3_1161 ();
 FILLER_ASAP7_75t_R FILLER_3_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_3_1192 ();
 FILLER_ASAP7_75t_R FILLER_3_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1200 ();
 DECAPx6_ASAP7_75t_R FILLER_3_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_4_112 ();
 DECAPx10_ASAP7_75t_R FILLER_4_134 ();
 DECAPx10_ASAP7_75t_R FILLER_4_156 ();
 DECAPx10_ASAP7_75t_R FILLER_4_178 ();
 DECAPx10_ASAP7_75t_R FILLER_4_200 ();
 DECAPx10_ASAP7_75t_R FILLER_4_222 ();
 DECAPx10_ASAP7_75t_R FILLER_4_244 ();
 DECAPx10_ASAP7_75t_R FILLER_4_266 ();
 DECAPx10_ASAP7_75t_R FILLER_4_288 ();
 DECAPx10_ASAP7_75t_R FILLER_4_310 ();
 DECAPx10_ASAP7_75t_R FILLER_4_332 ();
 DECAPx10_ASAP7_75t_R FILLER_4_354 ();
 DECAPx10_ASAP7_75t_R FILLER_4_376 ();
 DECAPx10_ASAP7_75t_R FILLER_4_398 ();
 DECAPx10_ASAP7_75t_R FILLER_4_420 ();
 DECAPx6_ASAP7_75t_R FILLER_4_442 ();
 DECAPx2_ASAP7_75t_R FILLER_4_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_477 ();
 DECAPx10_ASAP7_75t_R FILLER_4_528 ();
 DECAPx4_ASAP7_75t_R FILLER_4_550 ();
 FILLER_ASAP7_75t_R FILLER_4_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_596 ();
 DECAPx10_ASAP7_75t_R FILLER_4_619 ();
 DECAPx4_ASAP7_75t_R FILLER_4_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_654 ();
 FILLER_ASAP7_75t_R FILLER_4_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_662 ();
 DECAPx4_ASAP7_75t_R FILLER_4_669 ();
 DECAPx6_ASAP7_75t_R FILLER_4_682 ();
 DECAPx1_ASAP7_75t_R FILLER_4_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_700 ();
 DECAPx2_ASAP7_75t_R FILLER_4_704 ();
 DECAPx10_ASAP7_75t_R FILLER_4_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_740 ();
 DECAPx2_ASAP7_75t_R FILLER_4_749 ();
 FILLER_ASAP7_75t_R FILLER_4_755 ();
 DECAPx10_ASAP7_75t_R FILLER_4_762 ();
 DECAPx6_ASAP7_75t_R FILLER_4_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_798 ();
 FILLER_ASAP7_75t_R FILLER_4_804 ();
 DECAPx4_ASAP7_75t_R FILLER_4_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_827 ();
 DECAPx10_ASAP7_75t_R FILLER_4_831 ();
 DECAPx4_ASAP7_75t_R FILLER_4_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_863 ();
 DECAPx6_ASAP7_75t_R FILLER_4_869 ();
 DECAPx6_ASAP7_75t_R FILLER_4_886 ();
 FILLER_ASAP7_75t_R FILLER_4_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_902 ();
 DECAPx10_ASAP7_75t_R FILLER_4_908 ();
 DECAPx10_ASAP7_75t_R FILLER_4_930 ();
 DECAPx10_ASAP7_75t_R FILLER_4_952 ();
 DECAPx6_ASAP7_75t_R FILLER_4_974 ();
 FILLER_ASAP7_75t_R FILLER_4_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_990 ();
 DECAPx2_ASAP7_75t_R FILLER_4_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_4_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_4_1031 ();
 FILLER_ASAP7_75t_R FILLER_4_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1076 ();
 DECAPx6_ASAP7_75t_R FILLER_4_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_4_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_4_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_4_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1152 ();
 DECAPx1_ASAP7_75t_R FILLER_4_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1162 ();
 DECAPx1_ASAP7_75t_R FILLER_4_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1202 ();
 DECAPx6_ASAP7_75t_R FILLER_4_1208 ();
 FILLER_ASAP7_75t_R FILLER_4_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_5_68 ();
 DECAPx10_ASAP7_75t_R FILLER_5_90 ();
 DECAPx10_ASAP7_75t_R FILLER_5_112 ();
 DECAPx10_ASAP7_75t_R FILLER_5_134 ();
 DECAPx10_ASAP7_75t_R FILLER_5_156 ();
 DECAPx10_ASAP7_75t_R FILLER_5_178 ();
 DECAPx10_ASAP7_75t_R FILLER_5_200 ();
 DECAPx10_ASAP7_75t_R FILLER_5_222 ();
 DECAPx10_ASAP7_75t_R FILLER_5_244 ();
 DECAPx10_ASAP7_75t_R FILLER_5_266 ();
 DECAPx10_ASAP7_75t_R FILLER_5_288 ();
 DECAPx10_ASAP7_75t_R FILLER_5_310 ();
 DECAPx10_ASAP7_75t_R FILLER_5_332 ();
 DECAPx10_ASAP7_75t_R FILLER_5_354 ();
 DECAPx10_ASAP7_75t_R FILLER_5_376 ();
 DECAPx10_ASAP7_75t_R FILLER_5_398 ();
 DECAPx10_ASAP7_75t_R FILLER_5_420 ();
 DECAPx1_ASAP7_75t_R FILLER_5_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_452 ();
 FILLER_ASAP7_75t_R FILLER_5_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_472 ();
 DECAPx6_ASAP7_75t_R FILLER_5_516 ();
 DECAPx2_ASAP7_75t_R FILLER_5_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_536 ();
 DECAPx10_ASAP7_75t_R FILLER_5_557 ();
 DECAPx1_ASAP7_75t_R FILLER_5_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_583 ();
 DECAPx6_ASAP7_75t_R FILLER_5_595 ();
 FILLER_ASAP7_75t_R FILLER_5_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_611 ();
 DECAPx6_ASAP7_75t_R FILLER_5_632 ();
 DECAPx2_ASAP7_75t_R FILLER_5_646 ();
 DECAPx6_ASAP7_75t_R FILLER_5_655 ();
 DECAPx1_ASAP7_75t_R FILLER_5_669 ();
 FILLER_ASAP7_75t_R FILLER_5_694 ();
 FILLER_ASAP7_75t_R FILLER_5_709 ();
 FILLER_ASAP7_75t_R FILLER_5_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_716 ();
 DECAPx4_ASAP7_75t_R FILLER_5_722 ();
 DECAPx2_ASAP7_75t_R FILLER_5_737 ();
 FILLER_ASAP7_75t_R FILLER_5_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_745 ();
 FILLER_ASAP7_75t_R FILLER_5_749 ();
 DECAPx1_ASAP7_75t_R FILLER_5_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_766 ();
 DECAPx4_ASAP7_75t_R FILLER_5_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_782 ();
 DECAPx2_ASAP7_75t_R FILLER_5_793 ();
 DECAPx10_ASAP7_75t_R FILLER_5_802 ();
 DECAPx6_ASAP7_75t_R FILLER_5_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_838 ();
 FILLER_ASAP7_75t_R FILLER_5_847 ();
 DECAPx2_ASAP7_75t_R FILLER_5_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_860 ();
 DECAPx10_ASAP7_75t_R FILLER_5_864 ();
 DECAPx6_ASAP7_75t_R FILLER_5_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_900 ();
 FILLER_ASAP7_75t_R FILLER_5_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_906 ();
 DECAPx1_ASAP7_75t_R FILLER_5_915 ();
 DECAPx10_ASAP7_75t_R FILLER_5_926 ();
 DECAPx10_ASAP7_75t_R FILLER_5_948 ();
 DECAPx4_ASAP7_75t_R FILLER_5_970 ();
 FILLER_ASAP7_75t_R FILLER_5_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_982 ();
 FILLER_ASAP7_75t_R FILLER_5_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_999 ();
 DECAPx6_ASAP7_75t_R FILLER_5_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_5_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_5_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_5_1035 ();
 FILLER_ASAP7_75t_R FILLER_5_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1043 ();
 DECAPx6_ASAP7_75t_R FILLER_5_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_5_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_5_1105 ();
 FILLER_ASAP7_75t_R FILLER_5_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_5_1119 ();
 FILLER_ASAP7_75t_R FILLER_5_1126 ();
 FILLER_ASAP7_75t_R FILLER_5_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_5_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1156 ();
 DECAPx6_ASAP7_75t_R FILLER_5_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_5_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_5_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1197 ();
 DECAPx4_ASAP7_75t_R FILLER_5_1201 ();
 FILLER_ASAP7_75t_R FILLER_5_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_6_68 ();
 DECAPx10_ASAP7_75t_R FILLER_6_90 ();
 DECAPx10_ASAP7_75t_R FILLER_6_112 ();
 DECAPx10_ASAP7_75t_R FILLER_6_134 ();
 DECAPx10_ASAP7_75t_R FILLER_6_156 ();
 DECAPx10_ASAP7_75t_R FILLER_6_178 ();
 DECAPx10_ASAP7_75t_R FILLER_6_200 ();
 DECAPx10_ASAP7_75t_R FILLER_6_222 ();
 DECAPx10_ASAP7_75t_R FILLER_6_244 ();
 DECAPx10_ASAP7_75t_R FILLER_6_266 ();
 DECAPx10_ASAP7_75t_R FILLER_6_288 ();
 DECAPx10_ASAP7_75t_R FILLER_6_310 ();
 DECAPx10_ASAP7_75t_R FILLER_6_332 ();
 DECAPx10_ASAP7_75t_R FILLER_6_354 ();
 DECAPx10_ASAP7_75t_R FILLER_6_376 ();
 DECAPx10_ASAP7_75t_R FILLER_6_398 ();
 DECAPx6_ASAP7_75t_R FILLER_6_420 ();
 DECAPx2_ASAP7_75t_R FILLER_6_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_486 ();
 DECAPx4_ASAP7_75t_R FILLER_6_495 ();
 FILLER_ASAP7_75t_R FILLER_6_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_507 ();
 DECAPx4_ASAP7_75t_R FILLER_6_530 ();
 FILLER_ASAP7_75t_R FILLER_6_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_542 ();
 DECAPx2_ASAP7_75t_R FILLER_6_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_555 ();
 DECAPx1_ASAP7_75t_R FILLER_6_591 ();
 DECAPx1_ASAP7_75t_R FILLER_6_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_624 ();
 DECAPx10_ASAP7_75t_R FILLER_6_631 ();
 FILLER_ASAP7_75t_R FILLER_6_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_655 ();
 FILLER_ASAP7_75t_R FILLER_6_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_663 ();
 DECAPx10_ASAP7_75t_R FILLER_6_667 ();
 DECAPx6_ASAP7_75t_R FILLER_6_689 ();
 DECAPx10_ASAP7_75t_R FILLER_6_706 ();
 DECAPx1_ASAP7_75t_R FILLER_6_728 ();
 DECAPx10_ASAP7_75t_R FILLER_6_735 ();
 DECAPx6_ASAP7_75t_R FILLER_6_757 ();
 DECAPx1_ASAP7_75t_R FILLER_6_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_775 ();
 DECAPx1_ASAP7_75t_R FILLER_6_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_783 ();
 DECAPx10_ASAP7_75t_R FILLER_6_787 ();
 DECAPx10_ASAP7_75t_R FILLER_6_809 ();
 DECAPx6_ASAP7_75t_R FILLER_6_831 ();
 FILLER_ASAP7_75t_R FILLER_6_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_847 ();
 DECAPx10_ASAP7_75t_R FILLER_6_851 ();
 DECAPx10_ASAP7_75t_R FILLER_6_873 ();
 FILLER_ASAP7_75t_R FILLER_6_895 ();
 DECAPx4_ASAP7_75t_R FILLER_6_902 ();
 FILLER_ASAP7_75t_R FILLER_6_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_914 ();
 DECAPx10_ASAP7_75t_R FILLER_6_926 ();
 DECAPx10_ASAP7_75t_R FILLER_6_948 ();
 DECAPx10_ASAP7_75t_R FILLER_6_970 ();
 DECAPx10_ASAP7_75t_R FILLER_6_992 ();
 DECAPx6_ASAP7_75t_R FILLER_6_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_6_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1046 ();
 DECAPx6_ASAP7_75t_R FILLER_6_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_6_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1079 ();
 FILLER_ASAP7_75t_R FILLER_6_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1103 ();
 DECAPx4_ASAP7_75t_R FILLER_6_1107 ();
 FILLER_ASAP7_75t_R FILLER_6_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1119 ();
 FILLER_ASAP7_75t_R FILLER_6_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_6_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_6_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_6_1170 ();
 FILLER_ASAP7_75t_R FILLER_6_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_6_1185 ();
 DECAPx6_ASAP7_75t_R FILLER_6_1195 ();
 DECAPx1_ASAP7_75t_R FILLER_6_1209 ();
 FILLER_ASAP7_75t_R FILLER_6_1216 ();
 FILLER_ASAP7_75t_R FILLER_6_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_7_90 ();
 DECAPx10_ASAP7_75t_R FILLER_7_112 ();
 DECAPx10_ASAP7_75t_R FILLER_7_134 ();
 DECAPx10_ASAP7_75t_R FILLER_7_156 ();
 DECAPx10_ASAP7_75t_R FILLER_7_178 ();
 DECAPx10_ASAP7_75t_R FILLER_7_200 ();
 DECAPx10_ASAP7_75t_R FILLER_7_222 ();
 DECAPx10_ASAP7_75t_R FILLER_7_244 ();
 DECAPx10_ASAP7_75t_R FILLER_7_266 ();
 DECAPx10_ASAP7_75t_R FILLER_7_288 ();
 DECAPx10_ASAP7_75t_R FILLER_7_310 ();
 DECAPx10_ASAP7_75t_R FILLER_7_332 ();
 DECAPx10_ASAP7_75t_R FILLER_7_354 ();
 DECAPx10_ASAP7_75t_R FILLER_7_376 ();
 DECAPx10_ASAP7_75t_R FILLER_7_398 ();
 DECAPx6_ASAP7_75t_R FILLER_7_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_434 ();
 DECAPx6_ASAP7_75t_R FILLER_7_446 ();
 DECAPx1_ASAP7_75t_R FILLER_7_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_464 ();
 DECAPx6_ASAP7_75t_R FILLER_7_471 ();
 FILLER_ASAP7_75t_R FILLER_7_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_487 ();
 FILLER_ASAP7_75t_R FILLER_7_495 ();
 DECAPx10_ASAP7_75t_R FILLER_7_514 ();
 FILLER_ASAP7_75t_R FILLER_7_536 ();
 DECAPx2_ASAP7_75t_R FILLER_7_549 ();
 DECAPx2_ASAP7_75t_R FILLER_7_565 ();
 FILLER_ASAP7_75t_R FILLER_7_571 ();
 DECAPx6_ASAP7_75t_R FILLER_7_579 ();
 FILLER_ASAP7_75t_R FILLER_7_593 ();
 DECAPx10_ASAP7_75t_R FILLER_7_617 ();
 DECAPx1_ASAP7_75t_R FILLER_7_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_643 ();
 DECAPx1_ASAP7_75t_R FILLER_7_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_657 ();
 FILLER_ASAP7_75t_R FILLER_7_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_681 ();
 DECAPx10_ASAP7_75t_R FILLER_7_690 ();
 DECAPx10_ASAP7_75t_R FILLER_7_712 ();
 DECAPx10_ASAP7_75t_R FILLER_7_734 ();
 DECAPx10_ASAP7_75t_R FILLER_7_756 ();
 DECAPx10_ASAP7_75t_R FILLER_7_778 ();
 DECAPx10_ASAP7_75t_R FILLER_7_800 ();
 DECAPx10_ASAP7_75t_R FILLER_7_822 ();
 DECAPx10_ASAP7_75t_R FILLER_7_844 ();
 DECAPx10_ASAP7_75t_R FILLER_7_866 ();
 FILLER_ASAP7_75t_R FILLER_7_888 ();
 DECAPx10_ASAP7_75t_R FILLER_7_893 ();
 DECAPx2_ASAP7_75t_R FILLER_7_915 ();
 FILLER_ASAP7_75t_R FILLER_7_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_923 ();
 DECAPx10_ASAP7_75t_R FILLER_7_926 ();
 DECAPx10_ASAP7_75t_R FILLER_7_948 ();
 DECAPx4_ASAP7_75t_R FILLER_7_970 ();
 FILLER_ASAP7_75t_R FILLER_7_980 ();
 DECAPx1_ASAP7_75t_R FILLER_7_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_991 ();
 DECAPx10_ASAP7_75t_R FILLER_7_997 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_7_1041 ();
 FILLER_ASAP7_75t_R FILLER_7_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_7_1052 ();
 DECAPx4_ASAP7_75t_R FILLER_7_1061 ();
 FILLER_ASAP7_75t_R FILLER_7_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_7_1078 ();
 FILLER_ASAP7_75t_R FILLER_7_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_7_1100 ();
 FILLER_ASAP7_75t_R FILLER_7_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_7_1136 ();
 FILLER_ASAP7_75t_R FILLER_7_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1167 ();
 DECAPx6_ASAP7_75t_R FILLER_7_1189 ();
 FILLER_ASAP7_75t_R FILLER_7_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_8_112 ();
 DECAPx10_ASAP7_75t_R FILLER_8_134 ();
 DECAPx10_ASAP7_75t_R FILLER_8_156 ();
 DECAPx10_ASAP7_75t_R FILLER_8_178 ();
 DECAPx10_ASAP7_75t_R FILLER_8_200 ();
 DECAPx10_ASAP7_75t_R FILLER_8_222 ();
 DECAPx10_ASAP7_75t_R FILLER_8_244 ();
 DECAPx10_ASAP7_75t_R FILLER_8_266 ();
 DECAPx10_ASAP7_75t_R FILLER_8_288 ();
 DECAPx10_ASAP7_75t_R FILLER_8_310 ();
 DECAPx10_ASAP7_75t_R FILLER_8_332 ();
 DECAPx10_ASAP7_75t_R FILLER_8_354 ();
 DECAPx10_ASAP7_75t_R FILLER_8_376 ();
 DECAPx4_ASAP7_75t_R FILLER_8_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_408 ();
 FILLER_ASAP7_75t_R FILLER_8_435 ();
 DECAPx6_ASAP7_75t_R FILLER_8_443 ();
 DECAPx1_ASAP7_75t_R FILLER_8_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_461 ();
 DECAPx6_ASAP7_75t_R FILLER_8_464 ();
 DECAPx2_ASAP7_75t_R FILLER_8_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_484 ();
 FILLER_ASAP7_75t_R FILLER_8_492 ();
 DECAPx6_ASAP7_75t_R FILLER_8_502 ();
 DECAPx2_ASAP7_75t_R FILLER_8_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_541 ();
 FILLER_ASAP7_75t_R FILLER_8_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_572 ();
 DECAPx1_ASAP7_75t_R FILLER_8_588 ();
 DECAPx1_ASAP7_75t_R FILLER_8_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_608 ();
 DECAPx10_ASAP7_75t_R FILLER_8_615 ();
 DECAPx2_ASAP7_75t_R FILLER_8_637 ();
 FILLER_ASAP7_75t_R FILLER_8_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_645 ();
 DECAPx6_ASAP7_75t_R FILLER_8_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_663 ();
 FILLER_ASAP7_75t_R FILLER_8_672 ();
 DECAPx10_ASAP7_75t_R FILLER_8_696 ();
 DECAPx10_ASAP7_75t_R FILLER_8_718 ();
 DECAPx10_ASAP7_75t_R FILLER_8_740 ();
 DECAPx10_ASAP7_75t_R FILLER_8_762 ();
 DECAPx6_ASAP7_75t_R FILLER_8_784 ();
 DECAPx10_ASAP7_75t_R FILLER_8_806 ();
 DECAPx1_ASAP7_75t_R FILLER_8_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_835 ();
 DECAPx10_ASAP7_75t_R FILLER_8_841 ();
 DECAPx10_ASAP7_75t_R FILLER_8_863 ();
 DECAPx10_ASAP7_75t_R FILLER_8_885 ();
 DECAPx10_ASAP7_75t_R FILLER_8_907 ();
 DECAPx10_ASAP7_75t_R FILLER_8_929 ();
 DECAPx10_ASAP7_75t_R FILLER_8_951 ();
 DECAPx2_ASAP7_75t_R FILLER_8_973 ();
 FILLER_ASAP7_75t_R FILLER_8_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_981 ();
 DECAPx2_ASAP7_75t_R FILLER_8_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_991 ();
 DECAPx4_ASAP7_75t_R FILLER_8_995 ();
 FILLER_ASAP7_75t_R FILLER_8_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1018 ();
 FILLER_ASAP7_75t_R FILLER_8_1040 ();
 FILLER_ASAP7_75t_R FILLER_8_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_8_1056 ();
 FILLER_ASAP7_75t_R FILLER_8_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1072 ();
 DECAPx6_ASAP7_75t_R FILLER_8_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_8_1090 ();
 FILLER_ASAP7_75t_R FILLER_8_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1106 ();
 DECAPx4_ASAP7_75t_R FILLER_8_1110 ();
 FILLER_ASAP7_75t_R FILLER_8_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_8_1130 ();
 FILLER_ASAP7_75t_R FILLER_8_1136 ();
 DECAPx1_ASAP7_75t_R FILLER_8_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1145 ();
 FILLER_ASAP7_75t_R FILLER_8_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1154 ();
 DECAPx1_ASAP7_75t_R FILLER_8_1158 ();
 DECAPx1_ASAP7_75t_R FILLER_8_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1175 ();
 DECAPx6_ASAP7_75t_R FILLER_8_1197 ();
 FILLER_ASAP7_75t_R FILLER_8_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_9_68 ();
 DECAPx10_ASAP7_75t_R FILLER_9_90 ();
 DECAPx10_ASAP7_75t_R FILLER_9_112 ();
 DECAPx10_ASAP7_75t_R FILLER_9_134 ();
 DECAPx10_ASAP7_75t_R FILLER_9_156 ();
 DECAPx10_ASAP7_75t_R FILLER_9_178 ();
 DECAPx10_ASAP7_75t_R FILLER_9_200 ();
 DECAPx10_ASAP7_75t_R FILLER_9_222 ();
 DECAPx10_ASAP7_75t_R FILLER_9_244 ();
 DECAPx10_ASAP7_75t_R FILLER_9_266 ();
 DECAPx10_ASAP7_75t_R FILLER_9_288 ();
 DECAPx10_ASAP7_75t_R FILLER_9_310 ();
 DECAPx10_ASAP7_75t_R FILLER_9_332 ();
 DECAPx10_ASAP7_75t_R FILLER_9_354 ();
 DECAPx10_ASAP7_75t_R FILLER_9_376 ();
 DECAPx4_ASAP7_75t_R FILLER_9_398 ();
 FILLER_ASAP7_75t_R FILLER_9_408 ();
 DECAPx4_ASAP7_75t_R FILLER_9_416 ();
 FILLER_ASAP7_75t_R FILLER_9_426 ();
 DECAPx1_ASAP7_75t_R FILLER_9_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_453 ();
 FILLER_ASAP7_75t_R FILLER_9_483 ();
 DECAPx10_ASAP7_75t_R FILLER_9_493 ();
 DECAPx1_ASAP7_75t_R FILLER_9_515 ();
 FILLER_ASAP7_75t_R FILLER_9_541 ();
 DECAPx6_ASAP7_75t_R FILLER_9_554 ();
 DECAPx2_ASAP7_75t_R FILLER_9_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_580 ();
 DECAPx6_ASAP7_75t_R FILLER_9_589 ();
 DECAPx2_ASAP7_75t_R FILLER_9_603 ();
 DECAPx6_ASAP7_75t_R FILLER_9_626 ();
 DECAPx10_ASAP7_75t_R FILLER_9_646 ();
 DECAPx2_ASAP7_75t_R FILLER_9_668 ();
 FILLER_ASAP7_75t_R FILLER_9_674 ();
 DECAPx10_ASAP7_75t_R FILLER_9_710 ();
 DECAPx10_ASAP7_75t_R FILLER_9_732 ();
 DECAPx10_ASAP7_75t_R FILLER_9_754 ();
 DECAPx10_ASAP7_75t_R FILLER_9_776 ();
 DECAPx10_ASAP7_75t_R FILLER_9_798 ();
 DECAPx6_ASAP7_75t_R FILLER_9_820 ();
 DECAPx1_ASAP7_75t_R FILLER_9_834 ();
 DECAPx10_ASAP7_75t_R FILLER_9_848 ();
 DECAPx10_ASAP7_75t_R FILLER_9_870 ();
 DECAPx10_ASAP7_75t_R FILLER_9_892 ();
 DECAPx4_ASAP7_75t_R FILLER_9_914 ();
 DECAPx10_ASAP7_75t_R FILLER_9_926 ();
 DECAPx10_ASAP7_75t_R FILLER_9_948 ();
 DECAPx10_ASAP7_75t_R FILLER_9_970 ();
 DECAPx6_ASAP7_75t_R FILLER_9_992 ();
 FILLER_ASAP7_75t_R FILLER_9_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_9_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_9_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_9_1091 ();
 DECAPx6_ASAP7_75t_R FILLER_9_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_9_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_9_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_10_112 ();
 DECAPx10_ASAP7_75t_R FILLER_10_134 ();
 DECAPx10_ASAP7_75t_R FILLER_10_156 ();
 DECAPx10_ASAP7_75t_R FILLER_10_178 ();
 DECAPx10_ASAP7_75t_R FILLER_10_200 ();
 DECAPx10_ASAP7_75t_R FILLER_10_222 ();
 DECAPx10_ASAP7_75t_R FILLER_10_244 ();
 DECAPx10_ASAP7_75t_R FILLER_10_266 ();
 DECAPx10_ASAP7_75t_R FILLER_10_288 ();
 DECAPx10_ASAP7_75t_R FILLER_10_310 ();
 DECAPx10_ASAP7_75t_R FILLER_10_332 ();
 DECAPx10_ASAP7_75t_R FILLER_10_354 ();
 DECAPx10_ASAP7_75t_R FILLER_10_376 ();
 DECAPx10_ASAP7_75t_R FILLER_10_398 ();
 DECAPx2_ASAP7_75t_R FILLER_10_420 ();
 FILLER_ASAP7_75t_R FILLER_10_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_428 ();
 FILLER_ASAP7_75t_R FILLER_10_451 ();
 FILLER_ASAP7_75t_R FILLER_10_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_461 ();
 DECAPx1_ASAP7_75t_R FILLER_10_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_468 ();
 DECAPx10_ASAP7_75t_R FILLER_10_496 ();
 DECAPx6_ASAP7_75t_R FILLER_10_518 ();
 FILLER_ASAP7_75t_R FILLER_10_532 ();
 FILLER_ASAP7_75t_R FILLER_10_540 ();
 FILLER_ASAP7_75t_R FILLER_10_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_552 ();
 FILLER_ASAP7_75t_R FILLER_10_562 ();
 FILLER_ASAP7_75t_R FILLER_10_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_574 ();
 DECAPx6_ASAP7_75t_R FILLER_10_581 ();
 FILLER_ASAP7_75t_R FILLER_10_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_613 ();
 DECAPx2_ASAP7_75t_R FILLER_10_636 ();
 DECAPx4_ASAP7_75t_R FILLER_10_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_655 ();
 DECAPx10_ASAP7_75t_R FILLER_10_659 ();
 DECAPx4_ASAP7_75t_R FILLER_10_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_691 ();
 DECAPx2_ASAP7_75t_R FILLER_10_698 ();
 FILLER_ASAP7_75t_R FILLER_10_704 ();
 DECAPx10_ASAP7_75t_R FILLER_10_750 ();
 DECAPx10_ASAP7_75t_R FILLER_10_772 ();
 DECAPx10_ASAP7_75t_R FILLER_10_794 ();
 DECAPx6_ASAP7_75t_R FILLER_10_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_830 ();
 DECAPx4_ASAP7_75t_R FILLER_10_834 ();
 FILLER_ASAP7_75t_R FILLER_10_844 ();
 DECAPx10_ASAP7_75t_R FILLER_10_849 ();
 DECAPx10_ASAP7_75t_R FILLER_10_871 ();
 DECAPx10_ASAP7_75t_R FILLER_10_893 ();
 DECAPx10_ASAP7_75t_R FILLER_10_915 ();
 DECAPx4_ASAP7_75t_R FILLER_10_937 ();
 DECAPx10_ASAP7_75t_R FILLER_10_952 ();
 DECAPx10_ASAP7_75t_R FILLER_10_974 ();
 DECAPx10_ASAP7_75t_R FILLER_10_996 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_10_1032 ();
 FILLER_ASAP7_75t_R FILLER_10_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_10_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1112 ();
 FILLER_ASAP7_75t_R FILLER_10_1118 ();
 FILLER_ASAP7_75t_R FILLER_10_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1125 ();
 FILLER_ASAP7_75t_R FILLER_10_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1184 ();
 DECAPx6_ASAP7_75t_R FILLER_10_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_10_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_11_24 ();
 DECAPx10_ASAP7_75t_R FILLER_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_11_68 ();
 DECAPx10_ASAP7_75t_R FILLER_11_90 ();
 DECAPx10_ASAP7_75t_R FILLER_11_112 ();
 DECAPx10_ASAP7_75t_R FILLER_11_134 ();
 DECAPx10_ASAP7_75t_R FILLER_11_156 ();
 DECAPx10_ASAP7_75t_R FILLER_11_178 ();
 DECAPx10_ASAP7_75t_R FILLER_11_200 ();
 DECAPx10_ASAP7_75t_R FILLER_11_222 ();
 DECAPx10_ASAP7_75t_R FILLER_11_244 ();
 DECAPx10_ASAP7_75t_R FILLER_11_266 ();
 DECAPx10_ASAP7_75t_R FILLER_11_288 ();
 DECAPx10_ASAP7_75t_R FILLER_11_310 ();
 DECAPx10_ASAP7_75t_R FILLER_11_332 ();
 DECAPx10_ASAP7_75t_R FILLER_11_354 ();
 DECAPx10_ASAP7_75t_R FILLER_11_376 ();
 DECAPx6_ASAP7_75t_R FILLER_11_398 ();
 FILLER_ASAP7_75t_R FILLER_11_412 ();
 FILLER_ASAP7_75t_R FILLER_11_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_444 ();
 DECAPx10_ASAP7_75t_R FILLER_11_458 ();
 DECAPx1_ASAP7_75t_R FILLER_11_480 ();
 DECAPx6_ASAP7_75t_R FILLER_11_523 ();
 DECAPx1_ASAP7_75t_R FILLER_11_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_541 ();
 DECAPx2_ASAP7_75t_R FILLER_11_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_571 ();
 DECAPx1_ASAP7_75t_R FILLER_11_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_598 ();
 DECAPx1_ASAP7_75t_R FILLER_11_606 ();
 DECAPx2_ASAP7_75t_R FILLER_11_618 ();
 FILLER_ASAP7_75t_R FILLER_11_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_626 ();
 DECAPx6_ASAP7_75t_R FILLER_11_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_664 ();
 DECAPx2_ASAP7_75t_R FILLER_11_668 ();
 DECAPx1_ASAP7_75t_R FILLER_11_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_700 ();
 DECAPx4_ASAP7_75t_R FILLER_11_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_733 ();
 DECAPx10_ASAP7_75t_R FILLER_11_740 ();
 DECAPx10_ASAP7_75t_R FILLER_11_762 ();
 DECAPx4_ASAP7_75t_R FILLER_11_784 ();
 DECAPx10_ASAP7_75t_R FILLER_11_799 ();
 DECAPx10_ASAP7_75t_R FILLER_11_821 ();
 DECAPx10_ASAP7_75t_R FILLER_11_843 ();
 DECAPx10_ASAP7_75t_R FILLER_11_865 ();
 DECAPx10_ASAP7_75t_R FILLER_11_887 ();
 DECAPx6_ASAP7_75t_R FILLER_11_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_923 ();
 DECAPx6_ASAP7_75t_R FILLER_11_926 ();
 DECAPx1_ASAP7_75t_R FILLER_11_940 ();
 DECAPx10_ASAP7_75t_R FILLER_11_947 ();
 DECAPx10_ASAP7_75t_R FILLER_11_969 ();
 DECAPx10_ASAP7_75t_R FILLER_11_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1061 ();
 DECAPx6_ASAP7_75t_R FILLER_11_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_11_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1194 ();
 FILLER_ASAP7_75t_R FILLER_11_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_12_24 ();
 DECAPx10_ASAP7_75t_R FILLER_12_46 ();
 DECAPx10_ASAP7_75t_R FILLER_12_68 ();
 DECAPx10_ASAP7_75t_R FILLER_12_90 ();
 DECAPx10_ASAP7_75t_R FILLER_12_112 ();
 DECAPx10_ASAP7_75t_R FILLER_12_134 ();
 DECAPx10_ASAP7_75t_R FILLER_12_156 ();
 DECAPx10_ASAP7_75t_R FILLER_12_178 ();
 DECAPx10_ASAP7_75t_R FILLER_12_200 ();
 DECAPx10_ASAP7_75t_R FILLER_12_222 ();
 DECAPx10_ASAP7_75t_R FILLER_12_244 ();
 DECAPx10_ASAP7_75t_R FILLER_12_266 ();
 DECAPx10_ASAP7_75t_R FILLER_12_288 ();
 DECAPx10_ASAP7_75t_R FILLER_12_310 ();
 DECAPx10_ASAP7_75t_R FILLER_12_332 ();
 DECAPx10_ASAP7_75t_R FILLER_12_354 ();
 DECAPx10_ASAP7_75t_R FILLER_12_376 ();
 DECAPx10_ASAP7_75t_R FILLER_12_398 ();
 DECAPx4_ASAP7_75t_R FILLER_12_420 ();
 DECAPx10_ASAP7_75t_R FILLER_12_436 ();
 DECAPx1_ASAP7_75t_R FILLER_12_458 ();
 DECAPx2_ASAP7_75t_R FILLER_12_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_470 ();
 DECAPx10_ASAP7_75t_R FILLER_12_493 ();
 DECAPx2_ASAP7_75t_R FILLER_12_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_521 ();
 DECAPx1_ASAP7_75t_R FILLER_12_539 ();
 DECAPx10_ASAP7_75t_R FILLER_12_550 ();
 DECAPx6_ASAP7_75t_R FILLER_12_572 ();
 DECAPx2_ASAP7_75t_R FILLER_12_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_592 ();
 FILLER_ASAP7_75t_R FILLER_12_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_612 ();
 DECAPx1_ASAP7_75t_R FILLER_12_630 ();
 DECAPx4_ASAP7_75t_R FILLER_12_654 ();
 FILLER_ASAP7_75t_R FILLER_12_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_666 ();
 DECAPx1_ASAP7_75t_R FILLER_12_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_676 ();
 DECAPx4_ASAP7_75t_R FILLER_12_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_718 ();
 DECAPx2_ASAP7_75t_R FILLER_12_743 ();
 FILLER_ASAP7_75t_R FILLER_12_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_751 ();
 DECAPx6_ASAP7_75t_R FILLER_12_774 ();
 DECAPx1_ASAP7_75t_R FILLER_12_788 ();
 DECAPx10_ASAP7_75t_R FILLER_12_795 ();
 DECAPx4_ASAP7_75t_R FILLER_12_817 ();
 FILLER_ASAP7_75t_R FILLER_12_827 ();
 DECAPx6_ASAP7_75t_R FILLER_12_851 ();
 DECAPx1_ASAP7_75t_R FILLER_12_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_869 ();
 DECAPx10_ASAP7_75t_R FILLER_12_892 ();
 DECAPx10_ASAP7_75t_R FILLER_12_914 ();
 DECAPx10_ASAP7_75t_R FILLER_12_936 ();
 DECAPx10_ASAP7_75t_R FILLER_12_958 ();
 DECAPx10_ASAP7_75t_R FILLER_12_980 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_12_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_12_1038 ();
 FILLER_ASAP7_75t_R FILLER_12_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_12_1140 ();
 FILLER_ASAP7_75t_R FILLER_12_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_12_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_13_24 ();
 DECAPx10_ASAP7_75t_R FILLER_13_46 ();
 DECAPx10_ASAP7_75t_R FILLER_13_68 ();
 DECAPx10_ASAP7_75t_R FILLER_13_90 ();
 DECAPx10_ASAP7_75t_R FILLER_13_112 ();
 DECAPx10_ASAP7_75t_R FILLER_13_134 ();
 DECAPx10_ASAP7_75t_R FILLER_13_156 ();
 DECAPx10_ASAP7_75t_R FILLER_13_178 ();
 DECAPx10_ASAP7_75t_R FILLER_13_200 ();
 DECAPx10_ASAP7_75t_R FILLER_13_222 ();
 DECAPx10_ASAP7_75t_R FILLER_13_244 ();
 DECAPx10_ASAP7_75t_R FILLER_13_266 ();
 DECAPx10_ASAP7_75t_R FILLER_13_288 ();
 DECAPx10_ASAP7_75t_R FILLER_13_310 ();
 DECAPx10_ASAP7_75t_R FILLER_13_332 ();
 DECAPx10_ASAP7_75t_R FILLER_13_354 ();
 DECAPx10_ASAP7_75t_R FILLER_13_376 ();
 DECAPx2_ASAP7_75t_R FILLER_13_398 ();
 FILLER_ASAP7_75t_R FILLER_13_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_406 ();
 FILLER_ASAP7_75t_R FILLER_13_413 ();
 DECAPx1_ASAP7_75t_R FILLER_13_426 ();
 DECAPx6_ASAP7_75t_R FILLER_13_458 ();
 FILLER_ASAP7_75t_R FILLER_13_472 ();
 DECAPx2_ASAP7_75t_R FILLER_13_480 ();
 DECAPx4_ASAP7_75t_R FILLER_13_506 ();
 FILLER_ASAP7_75t_R FILLER_13_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_540 ();
 DECAPx10_ASAP7_75t_R FILLER_13_569 ();
 DECAPx1_ASAP7_75t_R FILLER_13_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_595 ();
 DECAPx6_ASAP7_75t_R FILLER_13_640 ();
 FILLER_ASAP7_75t_R FILLER_13_654 ();
 FILLER_ASAP7_75t_R FILLER_13_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_692 ();
 DECAPx2_ASAP7_75t_R FILLER_13_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_741 ();
 FILLER_ASAP7_75t_R FILLER_13_753 ();
 DECAPx10_ASAP7_75t_R FILLER_13_761 ();
 DECAPx6_ASAP7_75t_R FILLER_13_783 ();
 DECAPx1_ASAP7_75t_R FILLER_13_797 ();
 DECAPx10_ASAP7_75t_R FILLER_13_835 ();
 DECAPx2_ASAP7_75t_R FILLER_13_857 ();
 FILLER_ASAP7_75t_R FILLER_13_863 ();
 FILLER_ASAP7_75t_R FILLER_13_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_884 ();
 DECAPx6_ASAP7_75t_R FILLER_13_907 ();
 FILLER_ASAP7_75t_R FILLER_13_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_923 ();
 DECAPx10_ASAP7_75t_R FILLER_13_926 ();
 DECAPx10_ASAP7_75t_R FILLER_13_948 ();
 DECAPx10_ASAP7_75t_R FILLER_13_970 ();
 DECAPx10_ASAP7_75t_R FILLER_13_992 ();
 DECAPx4_ASAP7_75t_R FILLER_13_1014 ();
 FILLER_ASAP7_75t_R FILLER_13_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_13_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_13_1041 ();
 FILLER_ASAP7_75t_R FILLER_13_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1060 ();
 FILLER_ASAP7_75t_R FILLER_13_1066 ();
 DECAPx1_ASAP7_75t_R FILLER_13_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1082 ();
 FILLER_ASAP7_75t_R FILLER_13_1086 ();
 DECAPx4_ASAP7_75t_R FILLER_13_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1117 ();
 DECAPx6_ASAP7_75t_R FILLER_13_1139 ();
 FILLER_ASAP7_75t_R FILLER_13_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1155 ();
 FILLER_ASAP7_75t_R FILLER_13_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_13_1186 ();
 FILLER_ASAP7_75t_R FILLER_13_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1194 ();
 FILLER_ASAP7_75t_R FILLER_13_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1205 ();
 FILLER_ASAP7_75t_R FILLER_13_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_14_2 ();
 DECAPx10_ASAP7_75t_R FILLER_14_24 ();
 DECAPx10_ASAP7_75t_R FILLER_14_46 ();
 DECAPx10_ASAP7_75t_R FILLER_14_68 ();
 DECAPx10_ASAP7_75t_R FILLER_14_90 ();
 DECAPx10_ASAP7_75t_R FILLER_14_112 ();
 DECAPx10_ASAP7_75t_R FILLER_14_134 ();
 DECAPx10_ASAP7_75t_R FILLER_14_156 ();
 DECAPx10_ASAP7_75t_R FILLER_14_178 ();
 DECAPx10_ASAP7_75t_R FILLER_14_200 ();
 DECAPx10_ASAP7_75t_R FILLER_14_222 ();
 DECAPx10_ASAP7_75t_R FILLER_14_244 ();
 DECAPx10_ASAP7_75t_R FILLER_14_266 ();
 DECAPx10_ASAP7_75t_R FILLER_14_288 ();
 DECAPx10_ASAP7_75t_R FILLER_14_310 ();
 DECAPx10_ASAP7_75t_R FILLER_14_332 ();
 DECAPx10_ASAP7_75t_R FILLER_14_354 ();
 DECAPx10_ASAP7_75t_R FILLER_14_376 ();
 DECAPx2_ASAP7_75t_R FILLER_14_398 ();
 DECAPx1_ASAP7_75t_R FILLER_14_426 ();
 DECAPx2_ASAP7_75t_R FILLER_14_453 ();
 FILLER_ASAP7_75t_R FILLER_14_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_461 ();
 DECAPx4_ASAP7_75t_R FILLER_14_464 ();
 FILLER_ASAP7_75t_R FILLER_14_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_476 ();
 DECAPx4_ASAP7_75t_R FILLER_14_487 ();
 FILLER_ASAP7_75t_R FILLER_14_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_499 ();
 DECAPx6_ASAP7_75t_R FILLER_14_520 ();
 DECAPx2_ASAP7_75t_R FILLER_14_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_540 ();
 DECAPx2_ASAP7_75t_R FILLER_14_547 ();
 FILLER_ASAP7_75t_R FILLER_14_553 ();
 DECAPx6_ASAP7_75t_R FILLER_14_563 ();
 FILLER_ASAP7_75t_R FILLER_14_577 ();
 DECAPx2_ASAP7_75t_R FILLER_14_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_595 ();
 DECAPx10_ASAP7_75t_R FILLER_14_616 ();
 DECAPx2_ASAP7_75t_R FILLER_14_641 ();
 FILLER_ASAP7_75t_R FILLER_14_647 ();
 DECAPx1_ASAP7_75t_R FILLER_14_655 ();
 DECAPx4_ASAP7_75t_R FILLER_14_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_680 ();
 DECAPx1_ASAP7_75t_R FILLER_14_687 ();
 DECAPx6_ASAP7_75t_R FILLER_14_705 ();
 DECAPx2_ASAP7_75t_R FILLER_14_719 ();
 DECAPx2_ASAP7_75t_R FILLER_14_733 ();
 FILLER_ASAP7_75t_R FILLER_14_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_747 ();
 DECAPx10_ASAP7_75t_R FILLER_14_754 ();
 DECAPx6_ASAP7_75t_R FILLER_14_776 ();
 DECAPx1_ASAP7_75t_R FILLER_14_790 ();
 DECAPx1_ASAP7_75t_R FILLER_14_800 ();
 DECAPx1_ASAP7_75t_R FILLER_14_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_819 ();
 DECAPx4_ASAP7_75t_R FILLER_14_831 ();
 DECAPx4_ASAP7_75t_R FILLER_14_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_873 ();
 DECAPx10_ASAP7_75t_R FILLER_14_891 ();
 DECAPx10_ASAP7_75t_R FILLER_14_913 ();
 DECAPx10_ASAP7_75t_R FILLER_14_935 ();
 DECAPx10_ASAP7_75t_R FILLER_14_957 ();
 DECAPx10_ASAP7_75t_R FILLER_14_979 ();
 DECAPx6_ASAP7_75t_R FILLER_14_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_14_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1023 ();
 DECAPx6_ASAP7_75t_R FILLER_14_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_14_1046 ();
 FILLER_ASAP7_75t_R FILLER_14_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1055 ();
 FILLER_ASAP7_75t_R FILLER_14_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1074 ();
 DECAPx6_ASAP7_75t_R FILLER_14_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1158 ();
 DECAPx6_ASAP7_75t_R FILLER_14_1180 ();
 FILLER_ASAP7_75t_R FILLER_14_1194 ();
 DECAPx4_ASAP7_75t_R FILLER_14_1201 ();
 FILLER_ASAP7_75t_R FILLER_14_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1216 ();
 DECAPx1_ASAP7_75t_R FILLER_14_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_15_2 ();
 DECAPx10_ASAP7_75t_R FILLER_15_24 ();
 DECAPx10_ASAP7_75t_R FILLER_15_46 ();
 DECAPx10_ASAP7_75t_R FILLER_15_68 ();
 DECAPx10_ASAP7_75t_R FILLER_15_90 ();
 DECAPx10_ASAP7_75t_R FILLER_15_112 ();
 DECAPx10_ASAP7_75t_R FILLER_15_134 ();
 DECAPx10_ASAP7_75t_R FILLER_15_156 ();
 DECAPx10_ASAP7_75t_R FILLER_15_178 ();
 DECAPx10_ASAP7_75t_R FILLER_15_200 ();
 DECAPx10_ASAP7_75t_R FILLER_15_222 ();
 DECAPx10_ASAP7_75t_R FILLER_15_244 ();
 DECAPx10_ASAP7_75t_R FILLER_15_266 ();
 DECAPx10_ASAP7_75t_R FILLER_15_288 ();
 DECAPx10_ASAP7_75t_R FILLER_15_310 ();
 DECAPx10_ASAP7_75t_R FILLER_15_332 ();
 DECAPx10_ASAP7_75t_R FILLER_15_354 ();
 DECAPx10_ASAP7_75t_R FILLER_15_376 ();
 DECAPx6_ASAP7_75t_R FILLER_15_398 ();
 DECAPx2_ASAP7_75t_R FILLER_15_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_418 ();
 DECAPx2_ASAP7_75t_R FILLER_15_425 ();
 DECAPx2_ASAP7_75t_R FILLER_15_447 ();
 FILLER_ASAP7_75t_R FILLER_15_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_455 ();
 DECAPx2_ASAP7_75t_R FILLER_15_478 ();
 FILLER_ASAP7_75t_R FILLER_15_484 ();
 DECAPx10_ASAP7_75t_R FILLER_15_511 ();
 DECAPx4_ASAP7_75t_R FILLER_15_533 ();
 FILLER_ASAP7_75t_R FILLER_15_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_545 ();
 DECAPx6_ASAP7_75t_R FILLER_15_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_582 ();
 DECAPx10_ASAP7_75t_R FILLER_15_600 ();
 DECAPx6_ASAP7_75t_R FILLER_15_622 ();
 DECAPx2_ASAP7_75t_R FILLER_15_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_642 ();
 DECAPx2_ASAP7_75t_R FILLER_15_671 ();
 FILLER_ASAP7_75t_R FILLER_15_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_689 ();
 DECAPx6_ASAP7_75t_R FILLER_15_705 ();
 DECAPx2_ASAP7_75t_R FILLER_15_719 ();
 DECAPx2_ASAP7_75t_R FILLER_15_732 ();
 DECAPx2_ASAP7_75t_R FILLER_15_771 ();
 FILLER_ASAP7_75t_R FILLER_15_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_806 ();
 DECAPx6_ASAP7_75t_R FILLER_15_818 ();
 DECAPx6_ASAP7_75t_R FILLER_15_849 ();
 FILLER_ASAP7_75t_R FILLER_15_863 ();
 DECAPx2_ASAP7_75t_R FILLER_15_868 ();
 DECAPx4_ASAP7_75t_R FILLER_15_880 ();
 DECAPx6_ASAP7_75t_R FILLER_15_910 ();
 DECAPx10_ASAP7_75t_R FILLER_15_926 ();
 DECAPx10_ASAP7_75t_R FILLER_15_948 ();
 DECAPx10_ASAP7_75t_R FILLER_15_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_992 ();
 DECAPx10_ASAP7_75t_R FILLER_15_999 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1021 ();
 DECAPx4_ASAP7_75t_R FILLER_15_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_15_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_15_1135 ();
 FILLER_ASAP7_75t_R FILLER_15_1141 ();
 FILLER_ASAP7_75t_R FILLER_15_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1153 ();
 FILLER_ASAP7_75t_R FILLER_15_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1164 ();
 DECAPx4_ASAP7_75t_R FILLER_15_1186 ();
 DECAPx6_ASAP7_75t_R FILLER_15_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_16_2 ();
 DECAPx10_ASAP7_75t_R FILLER_16_24 ();
 DECAPx10_ASAP7_75t_R FILLER_16_46 ();
 DECAPx10_ASAP7_75t_R FILLER_16_68 ();
 DECAPx10_ASAP7_75t_R FILLER_16_90 ();
 DECAPx10_ASAP7_75t_R FILLER_16_112 ();
 DECAPx10_ASAP7_75t_R FILLER_16_134 ();
 DECAPx10_ASAP7_75t_R FILLER_16_156 ();
 DECAPx10_ASAP7_75t_R FILLER_16_178 ();
 DECAPx10_ASAP7_75t_R FILLER_16_200 ();
 DECAPx10_ASAP7_75t_R FILLER_16_222 ();
 DECAPx10_ASAP7_75t_R FILLER_16_244 ();
 DECAPx10_ASAP7_75t_R FILLER_16_266 ();
 DECAPx10_ASAP7_75t_R FILLER_16_288 ();
 DECAPx10_ASAP7_75t_R FILLER_16_310 ();
 DECAPx10_ASAP7_75t_R FILLER_16_332 ();
 DECAPx10_ASAP7_75t_R FILLER_16_354 ();
 DECAPx10_ASAP7_75t_R FILLER_16_376 ();
 DECAPx10_ASAP7_75t_R FILLER_16_398 ();
 DECAPx2_ASAP7_75t_R FILLER_16_420 ();
 FILLER_ASAP7_75t_R FILLER_16_426 ();
 DECAPx6_ASAP7_75t_R FILLER_16_436 ();
 DECAPx2_ASAP7_75t_R FILLER_16_450 ();
 DECAPx2_ASAP7_75t_R FILLER_16_464 ();
 FILLER_ASAP7_75t_R FILLER_16_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_472 ();
 DECAPx2_ASAP7_75t_R FILLER_16_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_501 ();
 DECAPx2_ASAP7_75t_R FILLER_16_524 ();
 FILLER_ASAP7_75t_R FILLER_16_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_550 ();
 DECAPx6_ASAP7_75t_R FILLER_16_559 ();
 DECAPx1_ASAP7_75t_R FILLER_16_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_577 ();
 DECAPx2_ASAP7_75t_R FILLER_16_598 ();
 FILLER_ASAP7_75t_R FILLER_16_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_606 ();
 DECAPx10_ASAP7_75t_R FILLER_16_613 ();
 DECAPx10_ASAP7_75t_R FILLER_16_635 ();
 DECAPx6_ASAP7_75t_R FILLER_16_657 ();
 DECAPx2_ASAP7_75t_R FILLER_16_687 ();
 FILLER_ASAP7_75t_R FILLER_16_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_695 ();
 DECAPx2_ASAP7_75t_R FILLER_16_724 ();
 FILLER_ASAP7_75t_R FILLER_16_743 ();
 DECAPx6_ASAP7_75t_R FILLER_16_779 ();
 FILLER_ASAP7_75t_R FILLER_16_793 ();
 FILLER_ASAP7_75t_R FILLER_16_801 ();
 FILLER_ASAP7_75t_R FILLER_16_815 ();
 DECAPx10_ASAP7_75t_R FILLER_16_825 ();
 DECAPx1_ASAP7_75t_R FILLER_16_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_884 ();
 FILLER_ASAP7_75t_R FILLER_16_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_904 ();
 DECAPx10_ASAP7_75t_R FILLER_16_915 ();
 DECAPx10_ASAP7_75t_R FILLER_16_937 ();
 DECAPx10_ASAP7_75t_R FILLER_16_959 ();
 DECAPx4_ASAP7_75t_R FILLER_16_981 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_16_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1061 ();
 DECAPx6_ASAP7_75t_R FILLER_16_1065 ();
 FILLER_ASAP7_75t_R FILLER_16_1079 ();
 FILLER_ASAP7_75t_R FILLER_16_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_16_1140 ();
 FILLER_ASAP7_75t_R FILLER_16_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_16_1200 ();
 FILLER_ASAP7_75t_R FILLER_16_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1216 ();
 DECAPx1_ASAP7_75t_R FILLER_16_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_17_2 ();
 DECAPx10_ASAP7_75t_R FILLER_17_24 ();
 DECAPx10_ASAP7_75t_R FILLER_17_46 ();
 DECAPx10_ASAP7_75t_R FILLER_17_68 ();
 DECAPx10_ASAP7_75t_R FILLER_17_90 ();
 DECAPx10_ASAP7_75t_R FILLER_17_112 ();
 DECAPx10_ASAP7_75t_R FILLER_17_134 ();
 DECAPx10_ASAP7_75t_R FILLER_17_156 ();
 DECAPx10_ASAP7_75t_R FILLER_17_178 ();
 DECAPx10_ASAP7_75t_R FILLER_17_200 ();
 DECAPx10_ASAP7_75t_R FILLER_17_222 ();
 DECAPx10_ASAP7_75t_R FILLER_17_244 ();
 DECAPx10_ASAP7_75t_R FILLER_17_266 ();
 DECAPx10_ASAP7_75t_R FILLER_17_288 ();
 DECAPx10_ASAP7_75t_R FILLER_17_310 ();
 DECAPx10_ASAP7_75t_R FILLER_17_332 ();
 DECAPx10_ASAP7_75t_R FILLER_17_354 ();
 DECAPx10_ASAP7_75t_R FILLER_17_376 ();
 FILLER_ASAP7_75t_R FILLER_17_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_400 ();
 DECAPx1_ASAP7_75t_R FILLER_17_407 ();
 DECAPx1_ASAP7_75t_R FILLER_17_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_426 ();
 FILLER_ASAP7_75t_R FILLER_17_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_451 ();
 DECAPx1_ASAP7_75t_R FILLER_17_467 ();
 FILLER_ASAP7_75t_R FILLER_17_490 ();
 DECAPx1_ASAP7_75t_R FILLER_17_515 ();
 FILLER_ASAP7_75t_R FILLER_17_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_543 ();
 DECAPx4_ASAP7_75t_R FILLER_17_557 ();
 FILLER_ASAP7_75t_R FILLER_17_567 ();
 DECAPx1_ASAP7_75t_R FILLER_17_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_603 ();
 DECAPx10_ASAP7_75t_R FILLER_17_626 ();
 DECAPx4_ASAP7_75t_R FILLER_17_648 ();
 FILLER_ASAP7_75t_R FILLER_17_658 ();
 DECAPx10_ASAP7_75t_R FILLER_17_694 ();
 DECAPx2_ASAP7_75t_R FILLER_17_716 ();
 DECAPx1_ASAP7_75t_R FILLER_17_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_737 ();
 DECAPx1_ASAP7_75t_R FILLER_17_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_779 ();
 FILLER_ASAP7_75t_R FILLER_17_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_827 ();
 FILLER_ASAP7_75t_R FILLER_17_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_873 ();
 FILLER_ASAP7_75t_R FILLER_17_881 ();
 DECAPx10_ASAP7_75t_R FILLER_17_895 ();
 DECAPx2_ASAP7_75t_R FILLER_17_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_923 ();
 DECAPx10_ASAP7_75t_R FILLER_17_926 ();
 DECAPx10_ASAP7_75t_R FILLER_17_948 ();
 FILLER_ASAP7_75t_R FILLER_17_970 ();
 FILLER_ASAP7_75t_R FILLER_17_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_985 ();
 DECAPx4_ASAP7_75t_R FILLER_17_997 ();
 FILLER_ASAP7_75t_R FILLER_17_1007 ();
 DECAPx6_ASAP7_75t_R FILLER_17_1031 ();
 FILLER_ASAP7_75t_R FILLER_17_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1133 ();
 FILLER_ASAP7_75t_R FILLER_17_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_17_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1172 ();
 DECAPx6_ASAP7_75t_R FILLER_17_1181 ();
 FILLER_ASAP7_75t_R FILLER_17_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_17_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_18_2 ();
 DECAPx10_ASAP7_75t_R FILLER_18_24 ();
 DECAPx10_ASAP7_75t_R FILLER_18_46 ();
 DECAPx10_ASAP7_75t_R FILLER_18_68 ();
 DECAPx10_ASAP7_75t_R FILLER_18_90 ();
 DECAPx10_ASAP7_75t_R FILLER_18_112 ();
 DECAPx10_ASAP7_75t_R FILLER_18_134 ();
 DECAPx10_ASAP7_75t_R FILLER_18_156 ();
 DECAPx10_ASAP7_75t_R FILLER_18_178 ();
 DECAPx10_ASAP7_75t_R FILLER_18_200 ();
 DECAPx10_ASAP7_75t_R FILLER_18_222 ();
 DECAPx10_ASAP7_75t_R FILLER_18_244 ();
 DECAPx10_ASAP7_75t_R FILLER_18_266 ();
 DECAPx10_ASAP7_75t_R FILLER_18_288 ();
 DECAPx10_ASAP7_75t_R FILLER_18_310 ();
 DECAPx10_ASAP7_75t_R FILLER_18_332 ();
 DECAPx10_ASAP7_75t_R FILLER_18_354 ();
 DECAPx6_ASAP7_75t_R FILLER_18_376 ();
 DECAPx2_ASAP7_75t_R FILLER_18_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_396 ();
 DECAPx1_ASAP7_75t_R FILLER_18_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_440 ();
 DECAPx4_ASAP7_75t_R FILLER_18_449 ();
 FILLER_ASAP7_75t_R FILLER_18_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_461 ();
 DECAPx6_ASAP7_75t_R FILLER_18_471 ();
 DECAPx10_ASAP7_75t_R FILLER_18_492 ();
 DECAPx4_ASAP7_75t_R FILLER_18_514 ();
 DECAPx2_ASAP7_75t_R FILLER_18_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_571 ();
 DECAPx10_ASAP7_75t_R FILLER_18_609 ();
 DECAPx6_ASAP7_75t_R FILLER_18_631 ();
 FILLER_ASAP7_75t_R FILLER_18_645 ();
 FILLER_ASAP7_75t_R FILLER_18_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_677 ();
 DECAPx10_ASAP7_75t_R FILLER_18_686 ();
 FILLER_ASAP7_75t_R FILLER_18_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_710 ();
 DECAPx1_ASAP7_75t_R FILLER_18_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_735 ();
 DECAPx1_ASAP7_75t_R FILLER_18_785 ();
 DECAPx4_ASAP7_75t_R FILLER_18_795 ();
 DECAPx2_ASAP7_75t_R FILLER_18_816 ();
 FILLER_ASAP7_75t_R FILLER_18_822 ();
 DECAPx10_ASAP7_75t_R FILLER_18_844 ();
 DECAPx4_ASAP7_75t_R FILLER_18_866 ();
 DECAPx6_ASAP7_75t_R FILLER_18_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_902 ();
 DECAPx10_ASAP7_75t_R FILLER_18_917 ();
 DECAPx6_ASAP7_75t_R FILLER_18_939 ();
 DECAPx1_ASAP7_75t_R FILLER_18_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_957 ();
 FILLER_ASAP7_75t_R FILLER_18_984 ();
 DECAPx2_ASAP7_75t_R FILLER_18_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_998 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_18_1038 ();
 FILLER_ASAP7_75t_R FILLER_18_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_18_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_18_1080 ();
 FILLER_ASAP7_75t_R FILLER_18_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1158 ();
 DECAPx6_ASAP7_75t_R FILLER_18_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1194 ();
 FILLER_ASAP7_75t_R FILLER_18_1198 ();
 FILLER_ASAP7_75t_R FILLER_18_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_19_2 ();
 DECAPx10_ASAP7_75t_R FILLER_19_24 ();
 DECAPx10_ASAP7_75t_R FILLER_19_46 ();
 DECAPx10_ASAP7_75t_R FILLER_19_68 ();
 DECAPx10_ASAP7_75t_R FILLER_19_90 ();
 DECAPx10_ASAP7_75t_R FILLER_19_112 ();
 DECAPx10_ASAP7_75t_R FILLER_19_134 ();
 DECAPx10_ASAP7_75t_R FILLER_19_156 ();
 DECAPx10_ASAP7_75t_R FILLER_19_178 ();
 DECAPx10_ASAP7_75t_R FILLER_19_200 ();
 DECAPx10_ASAP7_75t_R FILLER_19_222 ();
 DECAPx10_ASAP7_75t_R FILLER_19_244 ();
 DECAPx10_ASAP7_75t_R FILLER_19_266 ();
 DECAPx10_ASAP7_75t_R FILLER_19_288 ();
 DECAPx10_ASAP7_75t_R FILLER_19_310 ();
 DECAPx10_ASAP7_75t_R FILLER_19_332 ();
 DECAPx10_ASAP7_75t_R FILLER_19_354 ();
 DECAPx10_ASAP7_75t_R FILLER_19_376 ();
 DECAPx10_ASAP7_75t_R FILLER_19_398 ();
 DECAPx10_ASAP7_75t_R FILLER_19_420 ();
 DECAPx10_ASAP7_75t_R FILLER_19_442 ();
 DECAPx6_ASAP7_75t_R FILLER_19_464 ();
 DECAPx1_ASAP7_75t_R FILLER_19_478 ();
 DECAPx10_ASAP7_75t_R FILLER_19_488 ();
 DECAPx4_ASAP7_75t_R FILLER_19_510 ();
 DECAPx1_ASAP7_75t_R FILLER_19_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_530 ();
 DECAPx10_ASAP7_75t_R FILLER_19_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_564 ();
 DECAPx2_ASAP7_75t_R FILLER_19_580 ();
 FILLER_ASAP7_75t_R FILLER_19_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_588 ();
 DECAPx10_ASAP7_75t_R FILLER_19_629 ();
 DECAPx4_ASAP7_75t_R FILLER_19_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_661 ();
 DECAPx2_ASAP7_75t_R FILLER_19_670 ();
 DECAPx1_ASAP7_75t_R FILLER_19_682 ();
 DECAPx2_ASAP7_75t_R FILLER_19_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_739 ();
 DECAPx1_ASAP7_75t_R FILLER_19_768 ();
 FILLER_ASAP7_75t_R FILLER_19_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_796 ();
 DECAPx1_ASAP7_75t_R FILLER_19_805 ();
 DECAPx1_ASAP7_75t_R FILLER_19_816 ();
 DECAPx1_ASAP7_75t_R FILLER_19_829 ();
 DECAPx2_ASAP7_75t_R FILLER_19_866 ();
 FILLER_ASAP7_75t_R FILLER_19_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_874 ();
 DECAPx1_ASAP7_75t_R FILLER_19_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_901 ();
 DECAPx2_ASAP7_75t_R FILLER_19_926 ();
 FILLER_ASAP7_75t_R FILLER_19_932 ();
 DECAPx4_ASAP7_75t_R FILLER_19_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_978 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1030 ();
 DECAPx6_ASAP7_75t_R FILLER_19_1052 ();
 FILLER_ASAP7_75t_R FILLER_19_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1121 ();
 DECAPx4_ASAP7_75t_R FILLER_19_1143 ();
 FILLER_ASAP7_75t_R FILLER_19_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1155 ();
 FILLER_ASAP7_75t_R FILLER_19_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1166 ();
 FILLER_ASAP7_75t_R FILLER_19_1170 ();
 FILLER_ASAP7_75t_R FILLER_19_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1179 ();
 DECAPx4_ASAP7_75t_R FILLER_19_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_20_2 ();
 DECAPx10_ASAP7_75t_R FILLER_20_24 ();
 DECAPx10_ASAP7_75t_R FILLER_20_46 ();
 DECAPx10_ASAP7_75t_R FILLER_20_68 ();
 DECAPx10_ASAP7_75t_R FILLER_20_90 ();
 DECAPx10_ASAP7_75t_R FILLER_20_112 ();
 DECAPx10_ASAP7_75t_R FILLER_20_134 ();
 DECAPx10_ASAP7_75t_R FILLER_20_156 ();
 DECAPx10_ASAP7_75t_R FILLER_20_178 ();
 DECAPx10_ASAP7_75t_R FILLER_20_200 ();
 DECAPx10_ASAP7_75t_R FILLER_20_222 ();
 DECAPx10_ASAP7_75t_R FILLER_20_244 ();
 DECAPx10_ASAP7_75t_R FILLER_20_266 ();
 DECAPx10_ASAP7_75t_R FILLER_20_288 ();
 DECAPx10_ASAP7_75t_R FILLER_20_310 ();
 DECAPx10_ASAP7_75t_R FILLER_20_332 ();
 DECAPx10_ASAP7_75t_R FILLER_20_354 ();
 DECAPx10_ASAP7_75t_R FILLER_20_376 ();
 DECAPx10_ASAP7_75t_R FILLER_20_398 ();
 DECAPx4_ASAP7_75t_R FILLER_20_420 ();
 FILLER_ASAP7_75t_R FILLER_20_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_461 ();
 DECAPx2_ASAP7_75t_R FILLER_20_476 ();
 DECAPx6_ASAP7_75t_R FILLER_20_496 ();
 DECAPx2_ASAP7_75t_R FILLER_20_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_546 ();
 DECAPx10_ASAP7_75t_R FILLER_20_554 ();
 DECAPx4_ASAP7_75t_R FILLER_20_576 ();
 DECAPx10_ASAP7_75t_R FILLER_20_625 ();
 DECAPx4_ASAP7_75t_R FILLER_20_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_657 ();
 FILLER_ASAP7_75t_R FILLER_20_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_680 ();
 DECAPx4_ASAP7_75t_R FILLER_20_690 ();
 FILLER_ASAP7_75t_R FILLER_20_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_702 ();
 DECAPx10_ASAP7_75t_R FILLER_20_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_747 ();
 DECAPx6_ASAP7_75t_R FILLER_20_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_795 ();
 FILLER_ASAP7_75t_R FILLER_20_802 ();
 FILLER_ASAP7_75t_R FILLER_20_811 ();
 DECAPx2_ASAP7_75t_R FILLER_20_833 ();
 DECAPx1_ASAP7_75t_R FILLER_20_852 ();
 DECAPx2_ASAP7_75t_R FILLER_20_878 ();
 FILLER_ASAP7_75t_R FILLER_20_884 ();
 DECAPx4_ASAP7_75t_R FILLER_20_892 ();
 DECAPx1_ASAP7_75t_R FILLER_20_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_912 ();
 DECAPx6_ASAP7_75t_R FILLER_20_946 ();
 DECAPx4_ASAP7_75t_R FILLER_20_967 ();
 FILLER_ASAP7_75t_R FILLER_20_977 ();
 DECAPx2_ASAP7_75t_R FILLER_20_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_997 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1111 ();
 FILLER_ASAP7_75t_R FILLER_20_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1191 ();
 FILLER_ASAP7_75t_R FILLER_20_1197 ();
 FILLER_ASAP7_75t_R FILLER_20_1204 ();
 FILLER_ASAP7_75t_R FILLER_20_1209 ();
 DECAPx1_ASAP7_75t_R FILLER_20_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_21_2 ();
 DECAPx10_ASAP7_75t_R FILLER_21_24 ();
 DECAPx10_ASAP7_75t_R FILLER_21_46 ();
 DECAPx10_ASAP7_75t_R FILLER_21_68 ();
 DECAPx10_ASAP7_75t_R FILLER_21_90 ();
 DECAPx10_ASAP7_75t_R FILLER_21_112 ();
 DECAPx10_ASAP7_75t_R FILLER_21_134 ();
 DECAPx10_ASAP7_75t_R FILLER_21_156 ();
 DECAPx10_ASAP7_75t_R FILLER_21_178 ();
 DECAPx10_ASAP7_75t_R FILLER_21_200 ();
 DECAPx10_ASAP7_75t_R FILLER_21_222 ();
 DECAPx10_ASAP7_75t_R FILLER_21_244 ();
 DECAPx10_ASAP7_75t_R FILLER_21_266 ();
 DECAPx10_ASAP7_75t_R FILLER_21_288 ();
 DECAPx4_ASAP7_75t_R FILLER_21_310 ();
 DECAPx10_ASAP7_75t_R FILLER_21_326 ();
 DECAPx10_ASAP7_75t_R FILLER_21_348 ();
 DECAPx10_ASAP7_75t_R FILLER_21_370 ();
 DECAPx6_ASAP7_75t_R FILLER_21_392 ();
 FILLER_ASAP7_75t_R FILLER_21_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_408 ();
 FILLER_ASAP7_75t_R FILLER_21_437 ();
 DECAPx2_ASAP7_75t_R FILLER_21_461 ();
 FILLER_ASAP7_75t_R FILLER_21_479 ();
 FILLER_ASAP7_75t_R FILLER_21_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_523 ();
 FILLER_ASAP7_75t_R FILLER_21_546 ();
 FILLER_ASAP7_75t_R FILLER_21_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_566 ();
 FILLER_ASAP7_75t_R FILLER_21_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_591 ();
 DECAPx2_ASAP7_75t_R FILLER_21_600 ();
 DECAPx10_ASAP7_75t_R FILLER_21_612 ();
 DECAPx10_ASAP7_75t_R FILLER_21_634 ();
 DECAPx1_ASAP7_75t_R FILLER_21_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_660 ();
 DECAPx4_ASAP7_75t_R FILLER_21_667 ();
 DECAPx2_ASAP7_75t_R FILLER_21_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_708 ();
 DECAPx10_ASAP7_75t_R FILLER_21_715 ();
 DECAPx6_ASAP7_75t_R FILLER_21_737 ();
 DECAPx2_ASAP7_75t_R FILLER_21_751 ();
 DECAPx10_ASAP7_75t_R FILLER_21_763 ();
 DECAPx4_ASAP7_75t_R FILLER_21_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_795 ();
 DECAPx10_ASAP7_75t_R FILLER_21_803 ();
 DECAPx2_ASAP7_75t_R FILLER_21_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_831 ();
 DECAPx4_ASAP7_75t_R FILLER_21_843 ();
 DECAPx6_ASAP7_75t_R FILLER_21_861 ();
 DECAPx2_ASAP7_75t_R FILLER_21_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_881 ();
 DECAPx6_ASAP7_75t_R FILLER_21_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_904 ();
 DECAPx4_ASAP7_75t_R FILLER_21_912 ();
 FILLER_ASAP7_75t_R FILLER_21_922 ();
 DECAPx2_ASAP7_75t_R FILLER_21_926 ();
 DECAPx1_ASAP7_75t_R FILLER_21_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_958 ();
 DECAPx1_ASAP7_75t_R FILLER_21_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_977 ();
 DECAPx2_ASAP7_75t_R FILLER_21_986 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_21_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_21_1205 ();
 FILLER_ASAP7_75t_R FILLER_21_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1213 ();
 FILLER_ASAP7_75t_R FILLER_21_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_22_2 ();
 DECAPx10_ASAP7_75t_R FILLER_22_24 ();
 DECAPx10_ASAP7_75t_R FILLER_22_46 ();
 DECAPx10_ASAP7_75t_R FILLER_22_68 ();
 DECAPx10_ASAP7_75t_R FILLER_22_90 ();
 DECAPx10_ASAP7_75t_R FILLER_22_112 ();
 DECAPx10_ASAP7_75t_R FILLER_22_134 ();
 DECAPx10_ASAP7_75t_R FILLER_22_156 ();
 DECAPx10_ASAP7_75t_R FILLER_22_178 ();
 DECAPx10_ASAP7_75t_R FILLER_22_200 ();
 DECAPx10_ASAP7_75t_R FILLER_22_222 ();
 DECAPx10_ASAP7_75t_R FILLER_22_244 ();
 DECAPx10_ASAP7_75t_R FILLER_22_266 ();
 DECAPx10_ASAP7_75t_R FILLER_22_288 ();
 DECAPx2_ASAP7_75t_R FILLER_22_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_316 ();
 DECAPx6_ASAP7_75t_R FILLER_22_339 ();
 DECAPx1_ASAP7_75t_R FILLER_22_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_357 ();
 FILLER_ASAP7_75t_R FILLER_22_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_382 ();
 DECAPx6_ASAP7_75t_R FILLER_22_405 ();
 DECAPx1_ASAP7_75t_R FILLER_22_419 ();
 DECAPx1_ASAP7_75t_R FILLER_22_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_445 ();
 DECAPx2_ASAP7_75t_R FILLER_22_454 ();
 FILLER_ASAP7_75t_R FILLER_22_460 ();
 DECAPx6_ASAP7_75t_R FILLER_22_464 ();
 FILLER_ASAP7_75t_R FILLER_22_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_480 ();
 DECAPx6_ASAP7_75t_R FILLER_22_509 ();
 DECAPx1_ASAP7_75t_R FILLER_22_523 ();
 DECAPx1_ASAP7_75t_R FILLER_22_533 ();
 FILLER_ASAP7_75t_R FILLER_22_588 ();
 DECAPx10_ASAP7_75t_R FILLER_22_602 ();
 DECAPx4_ASAP7_75t_R FILLER_22_624 ();
 FILLER_ASAP7_75t_R FILLER_22_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_636 ();
 DECAPx4_ASAP7_75t_R FILLER_22_670 ();
 DECAPx6_ASAP7_75t_R FILLER_22_687 ();
 DECAPx2_ASAP7_75t_R FILLER_22_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_707 ();
 DECAPx4_ASAP7_75t_R FILLER_22_726 ();
 DECAPx10_ASAP7_75t_R FILLER_22_764 ();
 DECAPx2_ASAP7_75t_R FILLER_22_786 ();
 FILLER_ASAP7_75t_R FILLER_22_792 ();
 DECAPx10_ASAP7_75t_R FILLER_22_809 ();
 DECAPx10_ASAP7_75t_R FILLER_22_831 ();
 DECAPx10_ASAP7_75t_R FILLER_22_853 ();
 DECAPx1_ASAP7_75t_R FILLER_22_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_889 ();
 DECAPx2_ASAP7_75t_R FILLER_22_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_902 ();
 DECAPx4_ASAP7_75t_R FILLER_22_920 ();
 FILLER_ASAP7_75t_R FILLER_22_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_932 ();
 FILLER_ASAP7_75t_R FILLER_22_945 ();
 FILLER_ASAP7_75t_R FILLER_22_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_957 ();
 DECAPx10_ASAP7_75t_R FILLER_22_987 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1163 ();
 DECAPx6_ASAP7_75t_R FILLER_22_1185 ();
 DECAPx1_ASAP7_75t_R FILLER_22_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_22_1215 ();
 FILLER_ASAP7_75t_R FILLER_22_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_23_2 ();
 DECAPx10_ASAP7_75t_R FILLER_23_24 ();
 DECAPx10_ASAP7_75t_R FILLER_23_46 ();
 DECAPx10_ASAP7_75t_R FILLER_23_68 ();
 DECAPx10_ASAP7_75t_R FILLER_23_90 ();
 DECAPx10_ASAP7_75t_R FILLER_23_112 ();
 DECAPx10_ASAP7_75t_R FILLER_23_134 ();
 DECAPx10_ASAP7_75t_R FILLER_23_156 ();
 DECAPx10_ASAP7_75t_R FILLER_23_178 ();
 DECAPx10_ASAP7_75t_R FILLER_23_200 ();
 DECAPx10_ASAP7_75t_R FILLER_23_222 ();
 DECAPx10_ASAP7_75t_R FILLER_23_244 ();
 DECAPx10_ASAP7_75t_R FILLER_23_266 ();
 DECAPx10_ASAP7_75t_R FILLER_23_288 ();
 DECAPx1_ASAP7_75t_R FILLER_23_310 ();
 DECAPx10_ASAP7_75t_R FILLER_23_325 ();
 DECAPx2_ASAP7_75t_R FILLER_23_347 ();
 FILLER_ASAP7_75t_R FILLER_23_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_373 ();
 DECAPx10_ASAP7_75t_R FILLER_23_391 ();
 FILLER_ASAP7_75t_R FILLER_23_413 ();
 DECAPx2_ASAP7_75t_R FILLER_23_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_427 ();
 FILLER_ASAP7_75t_R FILLER_23_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_444 ();
 DECAPx1_ASAP7_75t_R FILLER_23_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_455 ();
 DECAPx2_ASAP7_75t_R FILLER_23_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_473 ();
 FILLER_ASAP7_75t_R FILLER_23_486 ();
 DECAPx6_ASAP7_75t_R FILLER_23_516 ();
 DECAPx10_ASAP7_75t_R FILLER_23_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_592 ();
 DECAPx4_ASAP7_75t_R FILLER_23_599 ();
 FILLER_ASAP7_75t_R FILLER_23_609 ();
 DECAPx2_ASAP7_75t_R FILLER_23_633 ();
 FILLER_ASAP7_75t_R FILLER_23_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_641 ();
 DECAPx6_ASAP7_75t_R FILLER_23_648 ();
 DECAPx2_ASAP7_75t_R FILLER_23_668 ();
 FILLER_ASAP7_75t_R FILLER_23_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_682 ();
 DECAPx1_ASAP7_75t_R FILLER_23_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_694 ();
 DECAPx1_ASAP7_75t_R FILLER_23_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_715 ();
 FILLER_ASAP7_75t_R FILLER_23_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_727 ();
 DECAPx6_ASAP7_75t_R FILLER_23_761 ();
 DECAPx1_ASAP7_75t_R FILLER_23_775 ();
 DECAPx1_ASAP7_75t_R FILLER_23_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_800 ();
 DECAPx2_ASAP7_75t_R FILLER_23_808 ();
 FILLER_ASAP7_75t_R FILLER_23_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_816 ();
 DECAPx2_ASAP7_75t_R FILLER_23_834 ();
 DECAPx10_ASAP7_75t_R FILLER_23_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_923 ();
 DECAPx2_ASAP7_75t_R FILLER_23_926 ();
 FILLER_ASAP7_75t_R FILLER_23_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_956 ();
 DECAPx6_ASAP7_75t_R FILLER_23_964 ();
 FILLER_ASAP7_75t_R FILLER_23_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_980 ();
 FILLER_ASAP7_75t_R FILLER_23_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1117 ();
 DECAPx4_ASAP7_75t_R FILLER_23_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_23_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_23_1187 ();
 FILLER_ASAP7_75t_R FILLER_23_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_23_1206 ();
 DECAPx2_ASAP7_75t_R FILLER_23_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_24_2 ();
 DECAPx10_ASAP7_75t_R FILLER_24_24 ();
 DECAPx10_ASAP7_75t_R FILLER_24_46 ();
 DECAPx10_ASAP7_75t_R FILLER_24_68 ();
 DECAPx10_ASAP7_75t_R FILLER_24_90 ();
 DECAPx10_ASAP7_75t_R FILLER_24_112 ();
 DECAPx10_ASAP7_75t_R FILLER_24_134 ();
 DECAPx10_ASAP7_75t_R FILLER_24_156 ();
 DECAPx10_ASAP7_75t_R FILLER_24_178 ();
 DECAPx10_ASAP7_75t_R FILLER_24_200 ();
 DECAPx10_ASAP7_75t_R FILLER_24_222 ();
 DECAPx10_ASAP7_75t_R FILLER_24_244 ();
 DECAPx10_ASAP7_75t_R FILLER_24_266 ();
 DECAPx10_ASAP7_75t_R FILLER_24_288 ();
 DECAPx1_ASAP7_75t_R FILLER_24_310 ();
 DECAPx1_ASAP7_75t_R FILLER_24_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_324 ();
 DECAPx6_ASAP7_75t_R FILLER_24_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_378 ();
 DECAPx2_ASAP7_75t_R FILLER_24_407 ();
 DECAPx1_ASAP7_75t_R FILLER_24_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_439 ();
 DECAPx1_ASAP7_75t_R FILLER_24_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_461 ();
 DECAPx2_ASAP7_75t_R FILLER_24_464 ();
 DECAPx1_ASAP7_75t_R FILLER_24_498 ();
 DECAPx10_ASAP7_75t_R FILLER_24_508 ();
 DECAPx4_ASAP7_75t_R FILLER_24_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_540 ();
 DECAPx6_ASAP7_75t_R FILLER_24_558 ();
 DECAPx1_ASAP7_75t_R FILLER_24_572 ();
 FILLER_ASAP7_75t_R FILLER_24_582 ();
 DECAPx1_ASAP7_75t_R FILLER_24_600 ();
 DECAPx10_ASAP7_75t_R FILLER_24_621 ();
 DECAPx6_ASAP7_75t_R FILLER_24_643 ();
 DECAPx2_ASAP7_75t_R FILLER_24_657 ();
 FILLER_ASAP7_75t_R FILLER_24_669 ();
 DECAPx2_ASAP7_75t_R FILLER_24_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_691 ();
 DECAPx2_ASAP7_75t_R FILLER_24_707 ();
 FILLER_ASAP7_75t_R FILLER_24_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_715 ();
 FILLER_ASAP7_75t_R FILLER_24_724 ();
 DECAPx1_ASAP7_75t_R FILLER_24_738 ();
 DECAPx10_ASAP7_75t_R FILLER_24_748 ();
 DECAPx2_ASAP7_75t_R FILLER_24_770 ();
 FILLER_ASAP7_75t_R FILLER_24_798 ();
 DECAPx2_ASAP7_75t_R FILLER_24_807 ();
 FILLER_ASAP7_75t_R FILLER_24_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_815 ();
 DECAPx2_ASAP7_75t_R FILLER_24_822 ();
 DECAPx10_ASAP7_75t_R FILLER_24_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_878 ();
 DECAPx4_ASAP7_75t_R FILLER_24_887 ();
 DECAPx4_ASAP7_75t_R FILLER_24_919 ();
 DECAPx1_ASAP7_75t_R FILLER_24_952 ();
 DECAPx6_ASAP7_75t_R FILLER_24_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_977 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_24_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_24_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_24_1211 ();
 FILLER_ASAP7_75t_R FILLER_24_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_25_2 ();
 DECAPx10_ASAP7_75t_R FILLER_25_24 ();
 DECAPx10_ASAP7_75t_R FILLER_25_46 ();
 DECAPx10_ASAP7_75t_R FILLER_25_68 ();
 DECAPx10_ASAP7_75t_R FILLER_25_90 ();
 DECAPx10_ASAP7_75t_R FILLER_25_112 ();
 DECAPx10_ASAP7_75t_R FILLER_25_134 ();
 DECAPx10_ASAP7_75t_R FILLER_25_156 ();
 DECAPx10_ASAP7_75t_R FILLER_25_178 ();
 DECAPx10_ASAP7_75t_R FILLER_25_200 ();
 DECAPx10_ASAP7_75t_R FILLER_25_222 ();
 DECAPx10_ASAP7_75t_R FILLER_25_244 ();
 DECAPx10_ASAP7_75t_R FILLER_25_266 ();
 DECAPx2_ASAP7_75t_R FILLER_25_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_316 ();
 DECAPx1_ASAP7_75t_R FILLER_25_323 ();
 DECAPx10_ASAP7_75t_R FILLER_25_334 ();
 DECAPx1_ASAP7_75t_R FILLER_25_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_376 ();
 DECAPx10_ASAP7_75t_R FILLER_25_392 ();
 DECAPx6_ASAP7_75t_R FILLER_25_414 ();
 FILLER_ASAP7_75t_R FILLER_25_438 ();
 FILLER_ASAP7_75t_R FILLER_25_462 ();
 DECAPx4_ASAP7_75t_R FILLER_25_474 ();
 FILLER_ASAP7_75t_R FILLER_25_484 ();
 DECAPx10_ASAP7_75t_R FILLER_25_504 ();
 DECAPx10_ASAP7_75t_R FILLER_25_526 ();
 DECAPx10_ASAP7_75t_R FILLER_25_548 ();
 FILLER_ASAP7_75t_R FILLER_25_570 ();
 DECAPx6_ASAP7_75t_R FILLER_25_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_614 ();
 DECAPx10_ASAP7_75t_R FILLER_25_638 ();
 DECAPx1_ASAP7_75t_R FILLER_25_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_719 ();
 DECAPx2_ASAP7_75t_R FILLER_25_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_740 ();
 DECAPx1_ASAP7_75t_R FILLER_25_758 ();
 DECAPx6_ASAP7_75t_R FILLER_25_768 ();
 DECAPx1_ASAP7_75t_R FILLER_25_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_786 ();
 FILLER_ASAP7_75t_R FILLER_25_797 ();
 DECAPx4_ASAP7_75t_R FILLER_25_833 ();
 DECAPx10_ASAP7_75t_R FILLER_25_854 ();
 DECAPx1_ASAP7_75t_R FILLER_25_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_880 ();
 DECAPx2_ASAP7_75t_R FILLER_25_889 ();
 FILLER_ASAP7_75t_R FILLER_25_895 ();
 DECAPx6_ASAP7_75t_R FILLER_25_903 ();
 DECAPx2_ASAP7_75t_R FILLER_25_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_923 ();
 DECAPx10_ASAP7_75t_R FILLER_25_926 ();
 DECAPx2_ASAP7_75t_R FILLER_25_948 ();
 FILLER_ASAP7_75t_R FILLER_25_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_967 ();
 FILLER_ASAP7_75t_R FILLER_25_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_25_1133 ();
 FILLER_ASAP7_75t_R FILLER_25_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1150 ();
 DECAPx6_ASAP7_75t_R FILLER_25_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_25_1186 ();
 DECAPx6_ASAP7_75t_R FILLER_25_1195 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_26_2 ();
 DECAPx10_ASAP7_75t_R FILLER_26_24 ();
 DECAPx10_ASAP7_75t_R FILLER_26_46 ();
 DECAPx10_ASAP7_75t_R FILLER_26_68 ();
 DECAPx10_ASAP7_75t_R FILLER_26_90 ();
 DECAPx10_ASAP7_75t_R FILLER_26_112 ();
 DECAPx10_ASAP7_75t_R FILLER_26_134 ();
 DECAPx10_ASAP7_75t_R FILLER_26_156 ();
 DECAPx10_ASAP7_75t_R FILLER_26_178 ();
 DECAPx10_ASAP7_75t_R FILLER_26_200 ();
 DECAPx10_ASAP7_75t_R FILLER_26_222 ();
 DECAPx10_ASAP7_75t_R FILLER_26_244 ();
 DECAPx10_ASAP7_75t_R FILLER_26_266 ();
 DECAPx1_ASAP7_75t_R FILLER_26_337 ();
 FILLER_ASAP7_75t_R FILLER_26_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_387 ();
 DECAPx4_ASAP7_75t_R FILLER_26_394 ();
 FILLER_ASAP7_75t_R FILLER_26_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_406 ();
 DECAPx6_ASAP7_75t_R FILLER_26_413 ();
 FILLER_ASAP7_75t_R FILLER_26_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_464 ();
 DECAPx6_ASAP7_75t_R FILLER_26_471 ();
 DECAPx1_ASAP7_75t_R FILLER_26_485 ();
 DECAPx10_ASAP7_75t_R FILLER_26_498 ();
 DECAPx4_ASAP7_75t_R FILLER_26_520 ();
 DECAPx1_ASAP7_75t_R FILLER_26_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_566 ();
 FILLER_ASAP7_75t_R FILLER_26_583 ();
 DECAPx4_ASAP7_75t_R FILLER_26_607 ();
 DECAPx6_ASAP7_75t_R FILLER_26_620 ();
 DECAPx1_ASAP7_75t_R FILLER_26_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_679 ();
 DECAPx4_ASAP7_75t_R FILLER_26_690 ();
 FILLER_ASAP7_75t_R FILLER_26_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_702 ();
 DECAPx2_ASAP7_75t_R FILLER_26_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_731 ();
 DECAPx6_ASAP7_75t_R FILLER_26_738 ();
 DECAPx10_ASAP7_75t_R FILLER_26_772 ();
 DECAPx4_ASAP7_75t_R FILLER_26_794 ();
 DECAPx10_ASAP7_75t_R FILLER_26_812 ();
 DECAPx1_ASAP7_75t_R FILLER_26_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_838 ();
 DECAPx10_ASAP7_75t_R FILLER_26_851 ();
 FILLER_ASAP7_75t_R FILLER_26_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_875 ();
 DECAPx6_ASAP7_75t_R FILLER_26_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_909 ();
 DECAPx10_ASAP7_75t_R FILLER_26_932 ();
 FILLER_ASAP7_75t_R FILLER_26_954 ();
 DECAPx10_ASAP7_75t_R FILLER_26_964 ();
 DECAPx6_ASAP7_75t_R FILLER_26_986 ();
 DECAPx1_ASAP7_75t_R FILLER_26_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1032 ();
 DECAPx6_ASAP7_75t_R FILLER_26_1054 ();
 FILLER_ASAP7_75t_R FILLER_26_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1142 ();
 FILLER_ASAP7_75t_R FILLER_26_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1166 ();
 DECAPx6_ASAP7_75t_R FILLER_26_1172 ();
 FILLER_ASAP7_75t_R FILLER_26_1189 ();
 DECAPx2_ASAP7_75t_R FILLER_26_1196 ();
 FILLER_ASAP7_75t_R FILLER_26_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1204 ();
 DECAPx1_ASAP7_75t_R FILLER_26_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_27_2 ();
 DECAPx10_ASAP7_75t_R FILLER_27_24 ();
 DECAPx10_ASAP7_75t_R FILLER_27_46 ();
 DECAPx10_ASAP7_75t_R FILLER_27_68 ();
 DECAPx10_ASAP7_75t_R FILLER_27_90 ();
 DECAPx10_ASAP7_75t_R FILLER_27_112 ();
 DECAPx10_ASAP7_75t_R FILLER_27_134 ();
 DECAPx10_ASAP7_75t_R FILLER_27_156 ();
 DECAPx10_ASAP7_75t_R FILLER_27_178 ();
 DECAPx10_ASAP7_75t_R FILLER_27_200 ();
 DECAPx10_ASAP7_75t_R FILLER_27_222 ();
 DECAPx10_ASAP7_75t_R FILLER_27_244 ();
 DECAPx10_ASAP7_75t_R FILLER_27_266 ();
 DECAPx4_ASAP7_75t_R FILLER_27_288 ();
 FILLER_ASAP7_75t_R FILLER_27_298 ();
 FILLER_ASAP7_75t_R FILLER_27_306 ();
 DECAPx1_ASAP7_75t_R FILLER_27_319 ();
 FILLER_ASAP7_75t_R FILLER_27_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_340 ();
 DECAPx1_ASAP7_75t_R FILLER_27_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_351 ();
 FILLER_ASAP7_75t_R FILLER_27_372 ();
 DECAPx1_ASAP7_75t_R FILLER_27_381 ();
 DECAPx1_ASAP7_75t_R FILLER_27_391 ();
 FILLER_ASAP7_75t_R FILLER_27_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_403 ();
 FILLER_ASAP7_75t_R FILLER_27_448 ();
 DECAPx4_ASAP7_75t_R FILLER_27_470 ();
 FILLER_ASAP7_75t_R FILLER_27_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_482 ();
 FILLER_ASAP7_75t_R FILLER_27_501 ();
 DECAPx10_ASAP7_75t_R FILLER_27_513 ();
 DECAPx10_ASAP7_75t_R FILLER_27_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_557 ();
 FILLER_ASAP7_75t_R FILLER_27_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_569 ();
 FILLER_ASAP7_75t_R FILLER_27_582 ();
 FILLER_ASAP7_75t_R FILLER_27_601 ();
 DECAPx10_ASAP7_75t_R FILLER_27_613 ();
 DECAPx10_ASAP7_75t_R FILLER_27_635 ();
 DECAPx4_ASAP7_75t_R FILLER_27_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_667 ();
 DECAPx6_ASAP7_75t_R FILLER_27_688 ();
 DECAPx2_ASAP7_75t_R FILLER_27_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_708 ();
 DECAPx1_ASAP7_75t_R FILLER_27_715 ();
 DECAPx1_ASAP7_75t_R FILLER_27_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_729 ();
 DECAPx1_ASAP7_75t_R FILLER_27_745 ();
 DECAPx4_ASAP7_75t_R FILLER_27_771 ();
 DECAPx2_ASAP7_75t_R FILLER_27_787 ();
 DECAPx2_ASAP7_75t_R FILLER_27_804 ();
 DECAPx2_ASAP7_75t_R FILLER_27_817 ();
 FILLER_ASAP7_75t_R FILLER_27_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_825 ();
 FILLER_ASAP7_75t_R FILLER_27_853 ();
 FILLER_ASAP7_75t_R FILLER_27_884 ();
 DECAPx6_ASAP7_75t_R FILLER_27_908 ();
 FILLER_ASAP7_75t_R FILLER_27_922 ();
 DECAPx2_ASAP7_75t_R FILLER_27_926 ();
 DECAPx6_ASAP7_75t_R FILLER_27_960 ();
 FILLER_ASAP7_75t_R FILLER_27_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_976 ();
 DECAPx4_ASAP7_75t_R FILLER_27_987 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_27_1149 ();
 FILLER_ASAP7_75t_R FILLER_27_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_27_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_27_1204 ();
 FILLER_ASAP7_75t_R FILLER_27_1210 ();
 FILLER_ASAP7_75t_R FILLER_27_1215 ();
 FILLER_ASAP7_75t_R FILLER_27_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_28_24 ();
 DECAPx10_ASAP7_75t_R FILLER_28_46 ();
 DECAPx10_ASAP7_75t_R FILLER_28_68 ();
 DECAPx10_ASAP7_75t_R FILLER_28_90 ();
 DECAPx10_ASAP7_75t_R FILLER_28_112 ();
 DECAPx10_ASAP7_75t_R FILLER_28_134 ();
 DECAPx10_ASAP7_75t_R FILLER_28_156 ();
 DECAPx10_ASAP7_75t_R FILLER_28_178 ();
 DECAPx10_ASAP7_75t_R FILLER_28_200 ();
 DECAPx10_ASAP7_75t_R FILLER_28_222 ();
 DECAPx10_ASAP7_75t_R FILLER_28_244 ();
 DECAPx10_ASAP7_75t_R FILLER_28_266 ();
 DECAPx10_ASAP7_75t_R FILLER_28_288 ();
 DECAPx6_ASAP7_75t_R FILLER_28_310 ();
 DECAPx2_ASAP7_75t_R FILLER_28_324 ();
 DECAPx6_ASAP7_75t_R FILLER_28_341 ();
 DECAPx1_ASAP7_75t_R FILLER_28_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_367 ();
 DECAPx6_ASAP7_75t_R FILLER_28_386 ();
 DECAPx2_ASAP7_75t_R FILLER_28_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_431 ();
 DECAPx1_ASAP7_75t_R FILLER_28_438 ();
 DECAPx4_ASAP7_75t_R FILLER_28_452 ();
 DECAPx2_ASAP7_75t_R FILLER_28_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_494 ();
 DECAPx4_ASAP7_75t_R FILLER_28_534 ();
 FILLER_ASAP7_75t_R FILLER_28_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_552 ();
 DECAPx2_ASAP7_75t_R FILLER_28_576 ();
 DECAPx10_ASAP7_75t_R FILLER_28_604 ();
 DECAPx4_ASAP7_75t_R FILLER_28_626 ();
 FILLER_ASAP7_75t_R FILLER_28_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_638 ();
 FILLER_ASAP7_75t_R FILLER_28_667 ();
 DECAPx4_ASAP7_75t_R FILLER_28_675 ();
 FILLER_ASAP7_75t_R FILLER_28_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_687 ();
 DECAPx10_ASAP7_75t_R FILLER_28_691 ();
 FILLER_ASAP7_75t_R FILLER_28_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_715 ();
 FILLER_ASAP7_75t_R FILLER_28_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_740 ();
 DECAPx6_ASAP7_75t_R FILLER_28_758 ();
 DECAPx1_ASAP7_75t_R FILLER_28_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_776 ();
 FILLER_ASAP7_75t_R FILLER_28_805 ();
 DECAPx2_ASAP7_75t_R FILLER_28_835 ();
 FILLER_ASAP7_75t_R FILLER_28_856 ();
 FILLER_ASAP7_75t_R FILLER_28_864 ();
 FILLER_ASAP7_75t_R FILLER_28_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_876 ();
 FILLER_ASAP7_75t_R FILLER_28_884 ();
 DECAPx10_ASAP7_75t_R FILLER_28_892 ();
 DECAPx10_ASAP7_75t_R FILLER_28_955 ();
 DECAPx4_ASAP7_75t_R FILLER_28_977 ();
 FILLER_ASAP7_75t_R FILLER_28_987 ();
 FILLER_ASAP7_75t_R FILLER_28_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1120 ();
 DECAPx6_ASAP7_75t_R FILLER_28_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1160 ();
 DECAPx4_ASAP7_75t_R FILLER_28_1182 ();
 FILLER_ASAP7_75t_R FILLER_28_1192 ();
 DECAPx1_ASAP7_75t_R FILLER_28_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1212 ();
 FILLER_ASAP7_75t_R FILLER_28_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_29_2 ();
 DECAPx10_ASAP7_75t_R FILLER_29_24 ();
 DECAPx10_ASAP7_75t_R FILLER_29_46 ();
 DECAPx10_ASAP7_75t_R FILLER_29_68 ();
 DECAPx10_ASAP7_75t_R FILLER_29_90 ();
 DECAPx10_ASAP7_75t_R FILLER_29_112 ();
 DECAPx10_ASAP7_75t_R FILLER_29_134 ();
 DECAPx10_ASAP7_75t_R FILLER_29_156 ();
 DECAPx10_ASAP7_75t_R FILLER_29_178 ();
 DECAPx10_ASAP7_75t_R FILLER_29_200 ();
 DECAPx10_ASAP7_75t_R FILLER_29_222 ();
 DECAPx10_ASAP7_75t_R FILLER_29_244 ();
 DECAPx10_ASAP7_75t_R FILLER_29_266 ();
 DECAPx2_ASAP7_75t_R FILLER_29_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_324 ();
 DECAPx1_ASAP7_75t_R FILLER_29_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_337 ();
 DECAPx10_ASAP7_75t_R FILLER_29_358 ();
 DECAPx2_ASAP7_75t_R FILLER_29_380 ();
 DECAPx2_ASAP7_75t_R FILLER_29_392 ();
 DECAPx1_ASAP7_75t_R FILLER_29_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_408 ();
 DECAPx2_ASAP7_75t_R FILLER_29_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_445 ();
 DECAPx4_ASAP7_75t_R FILLER_29_466 ();
 FILLER_ASAP7_75t_R FILLER_29_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_484 ();
 DECAPx10_ASAP7_75t_R FILLER_29_491 ();
 DECAPx10_ASAP7_75t_R FILLER_29_513 ();
 DECAPx1_ASAP7_75t_R FILLER_29_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_539 ();
 DECAPx10_ASAP7_75t_R FILLER_29_588 ();
 DECAPx2_ASAP7_75t_R FILLER_29_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_616 ();
 FILLER_ASAP7_75t_R FILLER_29_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_691 ();
 DECAPx10_ASAP7_75t_R FILLER_29_708 ();
 DECAPx1_ASAP7_75t_R FILLER_29_730 ();
 DECAPx6_ASAP7_75t_R FILLER_29_747 ();
 DECAPx1_ASAP7_75t_R FILLER_29_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_765 ();
 DECAPx2_ASAP7_75t_R FILLER_29_769 ();
 FILLER_ASAP7_75t_R FILLER_29_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_777 ();
 DECAPx1_ASAP7_75t_R FILLER_29_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_792 ();
 FILLER_ASAP7_75t_R FILLER_29_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_817 ();
 FILLER_ASAP7_75t_R FILLER_29_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_827 ();
 FILLER_ASAP7_75t_R FILLER_29_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_840 ();
 DECAPx2_ASAP7_75t_R FILLER_29_852 ();
 DECAPx2_ASAP7_75t_R FILLER_29_864 ();
 DECAPx10_ASAP7_75t_R FILLER_29_892 ();
 DECAPx4_ASAP7_75t_R FILLER_29_914 ();
 DECAPx2_ASAP7_75t_R FILLER_29_926 ();
 FILLER_ASAP7_75t_R FILLER_29_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_947 ();
 DECAPx10_ASAP7_75t_R FILLER_29_956 ();
 DECAPx2_ASAP7_75t_R FILLER_29_978 ();
 DECAPx1_ASAP7_75t_R FILLER_29_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1056 ();
 DECAPx4_ASAP7_75t_R FILLER_29_1078 ();
 FILLER_ASAP7_75t_R FILLER_29_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1140 ();
 FILLER_ASAP7_75t_R FILLER_29_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1164 ();
 DECAPx6_ASAP7_75t_R FILLER_29_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_29_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_30_2 ();
 DECAPx10_ASAP7_75t_R FILLER_30_24 ();
 DECAPx10_ASAP7_75t_R FILLER_30_46 ();
 DECAPx10_ASAP7_75t_R FILLER_30_68 ();
 DECAPx10_ASAP7_75t_R FILLER_30_90 ();
 DECAPx10_ASAP7_75t_R FILLER_30_112 ();
 DECAPx10_ASAP7_75t_R FILLER_30_134 ();
 DECAPx10_ASAP7_75t_R FILLER_30_156 ();
 DECAPx10_ASAP7_75t_R FILLER_30_178 ();
 DECAPx10_ASAP7_75t_R FILLER_30_200 ();
 DECAPx10_ASAP7_75t_R FILLER_30_222 ();
 DECAPx10_ASAP7_75t_R FILLER_30_244 ();
 DECAPx10_ASAP7_75t_R FILLER_30_266 ();
 DECAPx10_ASAP7_75t_R FILLER_30_288 ();
 FILLER_ASAP7_75t_R FILLER_30_310 ();
 FILLER_ASAP7_75t_R FILLER_30_318 ();
 DECAPx2_ASAP7_75t_R FILLER_30_326 ();
 FILLER_ASAP7_75t_R FILLER_30_332 ();
 DECAPx10_ASAP7_75t_R FILLER_30_351 ();
 DECAPx1_ASAP7_75t_R FILLER_30_373 ();
 DECAPx1_ASAP7_75t_R FILLER_30_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_388 ();
 DECAPx4_ASAP7_75t_R FILLER_30_420 ();
 FILLER_ASAP7_75t_R FILLER_30_460 ();
 DECAPx4_ASAP7_75t_R FILLER_30_464 ();
 FILLER_ASAP7_75t_R FILLER_30_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_476 ();
 DECAPx6_ASAP7_75t_R FILLER_30_499 ();
 DECAPx1_ASAP7_75t_R FILLER_30_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_517 ();
 DECAPx10_ASAP7_75t_R FILLER_30_521 ();
 DECAPx10_ASAP7_75t_R FILLER_30_543 ();
 DECAPx10_ASAP7_75t_R FILLER_30_565 ();
 DECAPx4_ASAP7_75t_R FILLER_30_587 ();
 FILLER_ASAP7_75t_R FILLER_30_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_599 ();
 FILLER_ASAP7_75t_R FILLER_30_620 ();
 DECAPx6_ASAP7_75t_R FILLER_30_645 ();
 FILLER_ASAP7_75t_R FILLER_30_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_661 ();
 DECAPx10_ASAP7_75t_R FILLER_30_665 ();
 DECAPx4_ASAP7_75t_R FILLER_30_687 ();
 FILLER_ASAP7_75t_R FILLER_30_697 ();
 DECAPx6_ASAP7_75t_R FILLER_30_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_735 ();
 DECAPx6_ASAP7_75t_R FILLER_30_742 ();
 DECAPx10_ASAP7_75t_R FILLER_30_776 ();
 DECAPx2_ASAP7_75t_R FILLER_30_798 ();
 FILLER_ASAP7_75t_R FILLER_30_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_823 ();
 DECAPx2_ASAP7_75t_R FILLER_30_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_844 ();
 DECAPx4_ASAP7_75t_R FILLER_30_862 ();
 FILLER_ASAP7_75t_R FILLER_30_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_874 ();
 FILLER_ASAP7_75t_R FILLER_30_881 ();
 DECAPx10_ASAP7_75t_R FILLER_30_889 ();
 DECAPx2_ASAP7_75t_R FILLER_30_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_917 ();
 DECAPx2_ASAP7_75t_R FILLER_30_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_935 ();
 DECAPx4_ASAP7_75t_R FILLER_30_944 ();
 FILLER_ASAP7_75t_R FILLER_30_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_956 ();
 FILLER_ASAP7_75t_R FILLER_30_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_981 ();
 DECAPx10_ASAP7_75t_R FILLER_30_993 ();
 DECAPx6_ASAP7_75t_R FILLER_30_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_30_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1037 ();
 DECAPx2_ASAP7_75t_R FILLER_30_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1179 ();
 DECAPx6_ASAP7_75t_R FILLER_30_1183 ();
 FILLER_ASAP7_75t_R FILLER_30_1197 ();
 FILLER_ASAP7_75t_R FILLER_30_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_30_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1214 ();
 DECAPx2_ASAP7_75t_R FILLER_30_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_31_2 ();
 DECAPx10_ASAP7_75t_R FILLER_31_24 ();
 DECAPx10_ASAP7_75t_R FILLER_31_46 ();
 DECAPx10_ASAP7_75t_R FILLER_31_68 ();
 DECAPx10_ASAP7_75t_R FILLER_31_90 ();
 DECAPx10_ASAP7_75t_R FILLER_31_112 ();
 DECAPx10_ASAP7_75t_R FILLER_31_134 ();
 DECAPx10_ASAP7_75t_R FILLER_31_156 ();
 DECAPx10_ASAP7_75t_R FILLER_31_178 ();
 DECAPx10_ASAP7_75t_R FILLER_31_200 ();
 DECAPx10_ASAP7_75t_R FILLER_31_222 ();
 DECAPx10_ASAP7_75t_R FILLER_31_244 ();
 DECAPx10_ASAP7_75t_R FILLER_31_266 ();
 DECAPx10_ASAP7_75t_R FILLER_31_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_322 ();
 DECAPx10_ASAP7_75t_R FILLER_31_345 ();
 DECAPx2_ASAP7_75t_R FILLER_31_367 ();
 FILLER_ASAP7_75t_R FILLER_31_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_375 ();
 FILLER_ASAP7_75t_R FILLER_31_383 ();
 DECAPx4_ASAP7_75t_R FILLER_31_402 ();
 FILLER_ASAP7_75t_R FILLER_31_412 ();
 DECAPx2_ASAP7_75t_R FILLER_31_436 ();
 DECAPx1_ASAP7_75t_R FILLER_31_448 ();
 DECAPx10_ASAP7_75t_R FILLER_31_457 ();
 DECAPx6_ASAP7_75t_R FILLER_31_479 ();
 DECAPx2_ASAP7_75t_R FILLER_31_542 ();
 DECAPx10_ASAP7_75t_R FILLER_31_558 ();
 DECAPx10_ASAP7_75t_R FILLER_31_580 ();
 DECAPx6_ASAP7_75t_R FILLER_31_602 ();
 DECAPx1_ASAP7_75t_R FILLER_31_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_620 ();
 DECAPx6_ASAP7_75t_R FILLER_31_627 ();
 FILLER_ASAP7_75t_R FILLER_31_641 ();
 DECAPx2_ASAP7_75t_R FILLER_31_663 ();
 FILLER_ASAP7_75t_R FILLER_31_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_671 ();
 DECAPx6_ASAP7_75t_R FILLER_31_695 ();
 DECAPx1_ASAP7_75t_R FILLER_31_709 ();
 DECAPx10_ASAP7_75t_R FILLER_31_757 ();
 DECAPx2_ASAP7_75t_R FILLER_31_779 ();
 FILLER_ASAP7_75t_R FILLER_31_785 ();
 DECAPx6_ASAP7_75t_R FILLER_31_797 ();
 FILLER_ASAP7_75t_R FILLER_31_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_827 ();
 DECAPx6_ASAP7_75t_R FILLER_31_834 ();
 FILLER_ASAP7_75t_R FILLER_31_848 ();
 FILLER_ASAP7_75t_R FILLER_31_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_855 ();
 DECAPx10_ASAP7_75t_R FILLER_31_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_900 ();
 FILLER_ASAP7_75t_R FILLER_31_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_923 ();
 FILLER_ASAP7_75t_R FILLER_31_932 ();
 DECAPx2_ASAP7_75t_R FILLER_31_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_952 ();
 DECAPx6_ASAP7_75t_R FILLER_31_966 ();
 FILLER_ASAP7_75t_R FILLER_31_980 ();
 DECAPx4_ASAP7_75t_R FILLER_31_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_998 ();
 FILLER_ASAP7_75t_R FILLER_31_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1053 ();
 FILLER_ASAP7_75t_R FILLER_31_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_31_1138 ();
 DECAPx1_ASAP7_75t_R FILLER_31_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1161 ();
 FILLER_ASAP7_75t_R FILLER_31_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1193 ();
 FILLER_ASAP7_75t_R FILLER_31_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_31_1204 ();
 FILLER_ASAP7_75t_R FILLER_31_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_32_2 ();
 DECAPx10_ASAP7_75t_R FILLER_32_24 ();
 DECAPx10_ASAP7_75t_R FILLER_32_46 ();
 DECAPx10_ASAP7_75t_R FILLER_32_68 ();
 DECAPx10_ASAP7_75t_R FILLER_32_90 ();
 DECAPx10_ASAP7_75t_R FILLER_32_112 ();
 DECAPx10_ASAP7_75t_R FILLER_32_134 ();
 DECAPx10_ASAP7_75t_R FILLER_32_156 ();
 DECAPx10_ASAP7_75t_R FILLER_32_178 ();
 DECAPx10_ASAP7_75t_R FILLER_32_200 ();
 DECAPx10_ASAP7_75t_R FILLER_32_222 ();
 DECAPx10_ASAP7_75t_R FILLER_32_244 ();
 DECAPx10_ASAP7_75t_R FILLER_32_266 ();
 DECAPx2_ASAP7_75t_R FILLER_32_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_294 ();
 FILLER_ASAP7_75t_R FILLER_32_317 ();
 DECAPx1_ASAP7_75t_R FILLER_32_325 ();
 FILLER_ASAP7_75t_R FILLER_32_351 ();
 DECAPx1_ASAP7_75t_R FILLER_32_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_369 ();
 FILLER_ASAP7_75t_R FILLER_32_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_392 ();
 DECAPx1_ASAP7_75t_R FILLER_32_421 ();
 DECAPx2_ASAP7_75t_R FILLER_32_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_461 ();
 DECAPx2_ASAP7_75t_R FILLER_32_464 ();
 FILLER_ASAP7_75t_R FILLER_32_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_495 ();
 DECAPx10_ASAP7_75t_R FILLER_32_499 ();
 DECAPx2_ASAP7_75t_R FILLER_32_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_551 ();
 DECAPx10_ASAP7_75t_R FILLER_32_558 ();
 DECAPx10_ASAP7_75t_R FILLER_32_580 ();
 DECAPx2_ASAP7_75t_R FILLER_32_622 ();
 FILLER_ASAP7_75t_R FILLER_32_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_630 ();
 DECAPx1_ASAP7_75t_R FILLER_32_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_681 ();
 DECAPx4_ASAP7_75t_R FILLER_32_714 ();
 FILLER_ASAP7_75t_R FILLER_32_724 ();
 FILLER_ASAP7_75t_R FILLER_32_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_737 ();
 DECAPx10_ASAP7_75t_R FILLER_32_766 ();
 DECAPx2_ASAP7_75t_R FILLER_32_788 ();
 FILLER_ASAP7_75t_R FILLER_32_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_796 ();
 DECAPx1_ASAP7_75t_R FILLER_32_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_823 ();
 DECAPx10_ASAP7_75t_R FILLER_32_849 ();
 DECAPx10_ASAP7_75t_R FILLER_32_871 ();
 DECAPx10_ASAP7_75t_R FILLER_32_893 ();
 DECAPx1_ASAP7_75t_R FILLER_32_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_930 ();
 DECAPx4_ASAP7_75t_R FILLER_32_966 ();
 FILLER_ASAP7_75t_R FILLER_32_976 ();
 FILLER_ASAP7_75t_R FILLER_32_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1057 ();
 DECAPx1_ASAP7_75t_R FILLER_32_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1083 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_32_1117 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1138 ();
 FILLER_ASAP7_75t_R FILLER_32_1152 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_32_1171 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1183 ();
 FILLER_ASAP7_75t_R FILLER_32_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_33_2 ();
 DECAPx10_ASAP7_75t_R FILLER_33_24 ();
 DECAPx10_ASAP7_75t_R FILLER_33_46 ();
 DECAPx10_ASAP7_75t_R FILLER_33_68 ();
 DECAPx10_ASAP7_75t_R FILLER_33_90 ();
 DECAPx10_ASAP7_75t_R FILLER_33_112 ();
 DECAPx10_ASAP7_75t_R FILLER_33_134 ();
 DECAPx10_ASAP7_75t_R FILLER_33_156 ();
 DECAPx6_ASAP7_75t_R FILLER_33_178 ();
 FILLER_ASAP7_75t_R FILLER_33_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_194 ();
 DECAPx10_ASAP7_75t_R FILLER_33_205 ();
 DECAPx10_ASAP7_75t_R FILLER_33_227 ();
 DECAPx10_ASAP7_75t_R FILLER_33_249 ();
 DECAPx10_ASAP7_75t_R FILLER_33_271 ();
 DECAPx4_ASAP7_75t_R FILLER_33_293 ();
 FILLER_ASAP7_75t_R FILLER_33_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_305 ();
 FILLER_ASAP7_75t_R FILLER_33_329 ();
 DECAPx2_ASAP7_75t_R FILLER_33_337 ();
 FILLER_ASAP7_75t_R FILLER_33_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_345 ();
 FILLER_ASAP7_75t_R FILLER_33_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_370 ();
 DECAPx10_ASAP7_75t_R FILLER_33_402 ();
 DECAPx6_ASAP7_75t_R FILLER_33_424 ();
 DECAPx2_ASAP7_75t_R FILLER_33_438 ();
 DECAPx2_ASAP7_75t_R FILLER_33_447 ();
 DECAPx10_ASAP7_75t_R FILLER_33_479 ();
 FILLER_ASAP7_75t_R FILLER_33_501 ();
 DECAPx6_ASAP7_75t_R FILLER_33_506 ();
 DECAPx2_ASAP7_75t_R FILLER_33_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_526 ();
 DECAPx10_ASAP7_75t_R FILLER_33_581 ();
 DECAPx2_ASAP7_75t_R FILLER_33_603 ();
 FILLER_ASAP7_75t_R FILLER_33_629 ();
 DECAPx10_ASAP7_75t_R FILLER_33_637 ();
 DECAPx1_ASAP7_75t_R FILLER_33_659 ();
 DECAPx6_ASAP7_75t_R FILLER_33_666 ();
 DECAPx10_ASAP7_75t_R FILLER_33_705 ();
 DECAPx1_ASAP7_75t_R FILLER_33_727 ();
 DECAPx6_ASAP7_75t_R FILLER_33_740 ();
 DECAPx1_ASAP7_75t_R FILLER_33_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_758 ();
 DECAPx10_ASAP7_75t_R FILLER_33_762 ();
 DECAPx2_ASAP7_75t_R FILLER_33_784 ();
 DECAPx6_ASAP7_75t_R FILLER_33_793 ();
 DECAPx2_ASAP7_75t_R FILLER_33_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_813 ();
 DECAPx10_ASAP7_75t_R FILLER_33_820 ();
 DECAPx10_ASAP7_75t_R FILLER_33_842 ();
 DECAPx6_ASAP7_75t_R FILLER_33_864 ();
 DECAPx1_ASAP7_75t_R FILLER_33_878 ();
 DECAPx6_ASAP7_75t_R FILLER_33_905 ();
 DECAPx1_ASAP7_75t_R FILLER_33_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_923 ();
 DECAPx10_ASAP7_75t_R FILLER_33_926 ();
 DECAPx1_ASAP7_75t_R FILLER_33_948 ();
 DECAPx4_ASAP7_75t_R FILLER_33_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_982 ();
 FILLER_ASAP7_75t_R FILLER_33_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_991 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1001 ();
 FILLER_ASAP7_75t_R FILLER_33_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_33_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1041 ();
 FILLER_ASAP7_75t_R FILLER_33_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_33_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_33_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1096 ();
 FILLER_ASAP7_75t_R FILLER_33_1102 ();
 FILLER_ASAP7_75t_R FILLER_33_1116 ();
 FILLER_ASAP7_75t_R FILLER_33_1132 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1156 ();
 FILLER_ASAP7_75t_R FILLER_33_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1177 ();
 FILLER_ASAP7_75t_R FILLER_33_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1185 ();
 FILLER_ASAP7_75t_R FILLER_33_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1204 ();
 FILLER_ASAP7_75t_R FILLER_33_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_34_2 ();
 DECAPx10_ASAP7_75t_R FILLER_34_24 ();
 DECAPx10_ASAP7_75t_R FILLER_34_46 ();
 DECAPx10_ASAP7_75t_R FILLER_34_68 ();
 DECAPx10_ASAP7_75t_R FILLER_34_90 ();
 DECAPx10_ASAP7_75t_R FILLER_34_112 ();
 DECAPx10_ASAP7_75t_R FILLER_34_134 ();
 DECAPx10_ASAP7_75t_R FILLER_34_156 ();
 DECAPx10_ASAP7_75t_R FILLER_34_178 ();
 DECAPx10_ASAP7_75t_R FILLER_34_200 ();
 DECAPx10_ASAP7_75t_R FILLER_34_222 ();
 DECAPx10_ASAP7_75t_R FILLER_34_244 ();
 DECAPx10_ASAP7_75t_R FILLER_34_266 ();
 DECAPx10_ASAP7_75t_R FILLER_34_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_310 ();
 FILLER_ASAP7_75t_R FILLER_34_329 ();
 DECAPx10_ASAP7_75t_R FILLER_34_338 ();
 DECAPx1_ASAP7_75t_R FILLER_34_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_364 ();
 DECAPx10_ASAP7_75t_R FILLER_34_379 ();
 DECAPx6_ASAP7_75t_R FILLER_34_401 ();
 FILLER_ASAP7_75t_R FILLER_34_415 ();
 DECAPx1_ASAP7_75t_R FILLER_34_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_427 ();
 DECAPx6_ASAP7_75t_R FILLER_34_448 ();
 DECAPx10_ASAP7_75t_R FILLER_34_464 ();
 DECAPx2_ASAP7_75t_R FILLER_34_486 ();
 DECAPx1_ASAP7_75t_R FILLER_34_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_519 ();
 FILLER_ASAP7_75t_R FILLER_34_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_528 ();
 DECAPx10_ASAP7_75t_R FILLER_34_532 ();
 DECAPx10_ASAP7_75t_R FILLER_34_554 ();
 DECAPx4_ASAP7_75t_R FILLER_34_576 ();
 FILLER_ASAP7_75t_R FILLER_34_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_588 ();
 DECAPx4_ASAP7_75t_R FILLER_34_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_619 ();
 DECAPx6_ASAP7_75t_R FILLER_34_629 ();
 DECAPx1_ASAP7_75t_R FILLER_34_643 ();
 DECAPx4_ASAP7_75t_R FILLER_34_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_677 ();
 DECAPx10_ASAP7_75t_R FILLER_34_681 ();
 DECAPx6_ASAP7_75t_R FILLER_34_703 ();
 FILLER_ASAP7_75t_R FILLER_34_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_719 ();
 DECAPx6_ASAP7_75t_R FILLER_34_740 ();
 DECAPx1_ASAP7_75t_R FILLER_34_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_758 ();
 DECAPx10_ASAP7_75t_R FILLER_34_782 ();
 DECAPx6_ASAP7_75t_R FILLER_34_804 ();
 DECAPx2_ASAP7_75t_R FILLER_34_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_824 ();
 DECAPx10_ASAP7_75t_R FILLER_34_893 ();
 DECAPx6_ASAP7_75t_R FILLER_34_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_960 ();
 DECAPx2_ASAP7_75t_R FILLER_34_967 ();
 FILLER_ASAP7_75t_R FILLER_34_973 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1026 ();
 FILLER_ASAP7_75t_R FILLER_34_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1071 ();
 FILLER_ASAP7_75t_R FILLER_34_1077 ();
 FILLER_ASAP7_75t_R FILLER_34_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1087 ();
 DECAPx4_ASAP7_75t_R FILLER_34_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1143 ();
 FILLER_ASAP7_75t_R FILLER_34_1165 ();
 DECAPx4_ASAP7_75t_R FILLER_34_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1180 ();
 DECAPx4_ASAP7_75t_R FILLER_34_1187 ();
 FILLER_ASAP7_75t_R FILLER_34_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1217 ();
 FILLER_ASAP7_75t_R FILLER_34_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_35_2 ();
 DECAPx10_ASAP7_75t_R FILLER_35_24 ();
 DECAPx10_ASAP7_75t_R FILLER_35_46 ();
 DECAPx10_ASAP7_75t_R FILLER_35_68 ();
 DECAPx10_ASAP7_75t_R FILLER_35_90 ();
 DECAPx10_ASAP7_75t_R FILLER_35_112 ();
 DECAPx10_ASAP7_75t_R FILLER_35_134 ();
 DECAPx10_ASAP7_75t_R FILLER_35_156 ();
 DECAPx10_ASAP7_75t_R FILLER_35_178 ();
 DECAPx10_ASAP7_75t_R FILLER_35_200 ();
 DECAPx10_ASAP7_75t_R FILLER_35_222 ();
 DECAPx10_ASAP7_75t_R FILLER_35_244 ();
 DECAPx1_ASAP7_75t_R FILLER_35_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_270 ();
 DECAPx1_ASAP7_75t_R FILLER_35_294 ();
 DECAPx4_ASAP7_75t_R FILLER_35_302 ();
 DECAPx10_ASAP7_75t_R FILLER_35_341 ();
 DECAPx1_ASAP7_75t_R FILLER_35_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_367 ();
 DECAPx10_ASAP7_75t_R FILLER_35_390 ();
 FILLER_ASAP7_75t_R FILLER_35_412 ();
 DECAPx4_ASAP7_75t_R FILLER_35_439 ();
 FILLER_ASAP7_75t_R FILLER_35_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_451 ();
 DECAPx2_ASAP7_75t_R FILLER_35_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_484 ();
 DECAPx1_ASAP7_75t_R FILLER_35_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_492 ();
 DECAPx2_ASAP7_75t_R FILLER_35_513 ();
 DECAPx10_ASAP7_75t_R FILLER_35_539 ();
 DECAPx10_ASAP7_75t_R FILLER_35_561 ();
 DECAPx6_ASAP7_75t_R FILLER_35_583 ();
 DECAPx1_ASAP7_75t_R FILLER_35_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_601 ();
 FILLER_ASAP7_75t_R FILLER_35_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_624 ();
 FILLER_ASAP7_75t_R FILLER_35_647 ();
 DECAPx4_ASAP7_75t_R FILLER_35_652 ();
 FILLER_ASAP7_75t_R FILLER_35_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_685 ();
 DECAPx2_ASAP7_75t_R FILLER_35_732 ();
 DECAPx4_ASAP7_75t_R FILLER_35_765 ();
 DECAPx4_ASAP7_75t_R FILLER_35_795 ();
 FILLER_ASAP7_75t_R FILLER_35_805 ();
 DECAPx1_ASAP7_75t_R FILLER_35_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_852 ();
 DECAPx6_ASAP7_75t_R FILLER_35_856 ();
 DECAPx10_ASAP7_75t_R FILLER_35_876 ();
 DECAPx6_ASAP7_75t_R FILLER_35_898 ();
 FILLER_ASAP7_75t_R FILLER_35_912 ();
 DECAPx1_ASAP7_75t_R FILLER_35_959 ();
 DECAPx1_ASAP7_75t_R FILLER_35_969 ();
 FILLER_ASAP7_75t_R FILLER_35_982 ();
 DECAPx6_ASAP7_75t_R FILLER_35_1020 ();
 FILLER_ASAP7_75t_R FILLER_35_1034 ();
 DECAPx1_ASAP7_75t_R FILLER_35_1042 ();
 FILLER_ASAP7_75t_R FILLER_35_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1109 ();
 DECAPx6_ASAP7_75t_R FILLER_35_1116 ();
 FILLER_ASAP7_75t_R FILLER_35_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1166 ();
 DECAPx6_ASAP7_75t_R FILLER_35_1188 ();
 FILLER_ASAP7_75t_R FILLER_35_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1208 ();
 FILLER_ASAP7_75t_R FILLER_35_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_36_2 ();
 DECAPx10_ASAP7_75t_R FILLER_36_24 ();
 DECAPx10_ASAP7_75t_R FILLER_36_46 ();
 DECAPx10_ASAP7_75t_R FILLER_36_68 ();
 DECAPx10_ASAP7_75t_R FILLER_36_90 ();
 DECAPx10_ASAP7_75t_R FILLER_36_112 ();
 DECAPx10_ASAP7_75t_R FILLER_36_134 ();
 DECAPx10_ASAP7_75t_R FILLER_36_156 ();
 DECAPx10_ASAP7_75t_R FILLER_36_178 ();
 DECAPx10_ASAP7_75t_R FILLER_36_200 ();
 DECAPx10_ASAP7_75t_R FILLER_36_222 ();
 DECAPx4_ASAP7_75t_R FILLER_36_244 ();
 FILLER_ASAP7_75t_R FILLER_36_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_256 ();
 DECAPx10_ASAP7_75t_R FILLER_36_280 ();
 DECAPx10_ASAP7_75t_R FILLER_36_302 ();
 FILLER_ASAP7_75t_R FILLER_36_324 ();
 DECAPx2_ASAP7_75t_R FILLER_36_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_344 ();
 DECAPx6_ASAP7_75t_R FILLER_36_367 ();
 DECAPx2_ASAP7_75t_R FILLER_36_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_416 ();
 DECAPx10_ASAP7_75t_R FILLER_36_427 ();
 DECAPx4_ASAP7_75t_R FILLER_36_449 ();
 FILLER_ASAP7_75t_R FILLER_36_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_461 ();
 DECAPx2_ASAP7_75t_R FILLER_36_464 ();
 FILLER_ASAP7_75t_R FILLER_36_492 ();
 DECAPx10_ASAP7_75t_R FILLER_36_497 ();
 DECAPx10_ASAP7_75t_R FILLER_36_519 ();
 DECAPx10_ASAP7_75t_R FILLER_36_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_563 ();
 FILLER_ASAP7_75t_R FILLER_36_590 ();
 DECAPx2_ASAP7_75t_R FILLER_36_615 ();
 DECAPx2_ASAP7_75t_R FILLER_36_624 ();
 FILLER_ASAP7_75t_R FILLER_36_630 ();
 DECAPx4_ASAP7_75t_R FILLER_36_654 ();
 FILLER_ASAP7_75t_R FILLER_36_664 ();
 DECAPx10_ASAP7_75t_R FILLER_36_698 ();
 DECAPx2_ASAP7_75t_R FILLER_36_720 ();
 FILLER_ASAP7_75t_R FILLER_36_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_728 ();
 DECAPx1_ASAP7_75t_R FILLER_36_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_756 ();
 DECAPx1_ASAP7_75t_R FILLER_36_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_781 ();
 DECAPx1_ASAP7_75t_R FILLER_36_785 ();
 DECAPx6_ASAP7_75t_R FILLER_36_809 ();
 FILLER_ASAP7_75t_R FILLER_36_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_892 ();
 DECAPx10_ASAP7_75t_R FILLER_36_899 ();
 DECAPx10_ASAP7_75t_R FILLER_36_921 ();
 DECAPx2_ASAP7_75t_R FILLER_36_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_972 ();
 FILLER_ASAP7_75t_R FILLER_36_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1008 ();
 FILLER_ASAP7_75t_R FILLER_36_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1080 ();
 FILLER_ASAP7_75t_R FILLER_36_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1096 ();
 FILLER_ASAP7_75t_R FILLER_36_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_37_2 ();
 DECAPx10_ASAP7_75t_R FILLER_37_24 ();
 DECAPx10_ASAP7_75t_R FILLER_37_46 ();
 DECAPx10_ASAP7_75t_R FILLER_37_68 ();
 DECAPx10_ASAP7_75t_R FILLER_37_90 ();
 DECAPx10_ASAP7_75t_R FILLER_37_112 ();
 DECAPx10_ASAP7_75t_R FILLER_37_134 ();
 DECAPx10_ASAP7_75t_R FILLER_37_156 ();
 DECAPx10_ASAP7_75t_R FILLER_37_178 ();
 DECAPx10_ASAP7_75t_R FILLER_37_200 ();
 DECAPx10_ASAP7_75t_R FILLER_37_222 ();
 DECAPx10_ASAP7_75t_R FILLER_37_244 ();
 DECAPx10_ASAP7_75t_R FILLER_37_266 ();
 DECAPx10_ASAP7_75t_R FILLER_37_288 ();
 DECAPx6_ASAP7_75t_R FILLER_37_310 ();
 DECAPx2_ASAP7_75t_R FILLER_37_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_337 ();
 FILLER_ASAP7_75t_R FILLER_37_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_357 ();
 DECAPx2_ASAP7_75t_R FILLER_37_364 ();
 FILLER_ASAP7_75t_R FILLER_37_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_372 ();
 FILLER_ASAP7_75t_R FILLER_37_381 ();
 DECAPx2_ASAP7_75t_R FILLER_37_398 ();
 DECAPx10_ASAP7_75t_R FILLER_37_424 ();
 DECAPx2_ASAP7_75t_R FILLER_37_446 ();
 DECAPx1_ASAP7_75t_R FILLER_37_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_482 ();
 DECAPx6_ASAP7_75t_R FILLER_37_505 ();
 DECAPx10_ASAP7_75t_R FILLER_37_539 ();
 DECAPx6_ASAP7_75t_R FILLER_37_561 ();
 DECAPx1_ASAP7_75t_R FILLER_37_575 ();
 DECAPx2_ASAP7_75t_R FILLER_37_604 ();
 FILLER_ASAP7_75t_R FILLER_37_610 ();
 DECAPx2_ASAP7_75t_R FILLER_37_638 ();
 FILLER_ASAP7_75t_R FILLER_37_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_646 ();
 DECAPx10_ASAP7_75t_R FILLER_37_669 ();
 FILLER_ASAP7_75t_R FILLER_37_691 ();
 DECAPx10_ASAP7_75t_R FILLER_37_703 ();
 DECAPx2_ASAP7_75t_R FILLER_37_725 ();
 FILLER_ASAP7_75t_R FILLER_37_731 ();
 DECAPx10_ASAP7_75t_R FILLER_37_739 ();
 DECAPx6_ASAP7_75t_R FILLER_37_784 ();
 DECAPx1_ASAP7_75t_R FILLER_37_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_802 ();
 DECAPx4_ASAP7_75t_R FILLER_37_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_833 ();
 DECAPx4_ASAP7_75t_R FILLER_37_837 ();
 FILLER_ASAP7_75t_R FILLER_37_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_849 ();
 DECAPx10_ASAP7_75t_R FILLER_37_856 ();
 DECAPx4_ASAP7_75t_R FILLER_37_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_888 ();
 DECAPx4_ASAP7_75t_R FILLER_37_912 ();
 FILLER_ASAP7_75t_R FILLER_37_922 ();
 DECAPx10_ASAP7_75t_R FILLER_37_926 ();
 DECAPx1_ASAP7_75t_R FILLER_37_948 ();
 DECAPx10_ASAP7_75t_R FILLER_37_958 ();
 FILLER_ASAP7_75t_R FILLER_37_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1031 ();
 DECAPx4_ASAP7_75t_R FILLER_37_1053 ();
 FILLER_ASAP7_75t_R FILLER_37_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1065 ();
 DECAPx6_ASAP7_75t_R FILLER_37_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1086 ();
 DECAPx4_ASAP7_75t_R FILLER_37_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_37_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_38_2 ();
 DECAPx10_ASAP7_75t_R FILLER_38_24 ();
 DECAPx10_ASAP7_75t_R FILLER_38_46 ();
 DECAPx10_ASAP7_75t_R FILLER_38_68 ();
 DECAPx10_ASAP7_75t_R FILLER_38_90 ();
 DECAPx10_ASAP7_75t_R FILLER_38_112 ();
 DECAPx10_ASAP7_75t_R FILLER_38_134 ();
 DECAPx10_ASAP7_75t_R FILLER_38_156 ();
 DECAPx10_ASAP7_75t_R FILLER_38_178 ();
 DECAPx10_ASAP7_75t_R FILLER_38_200 ();
 DECAPx10_ASAP7_75t_R FILLER_38_222 ();
 DECAPx10_ASAP7_75t_R FILLER_38_244 ();
 DECAPx10_ASAP7_75t_R FILLER_38_266 ();
 DECAPx10_ASAP7_75t_R FILLER_38_288 ();
 DECAPx2_ASAP7_75t_R FILLER_38_310 ();
 DECAPx2_ASAP7_75t_R FILLER_38_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_350 ();
 DECAPx2_ASAP7_75t_R FILLER_38_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_385 ();
 DECAPx2_ASAP7_75t_R FILLER_38_402 ();
 FILLER_ASAP7_75t_R FILLER_38_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_410 ();
 DECAPx1_ASAP7_75t_R FILLER_38_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_461 ();
 DECAPx10_ASAP7_75t_R FILLER_38_464 ();
 DECAPx1_ASAP7_75t_R FILLER_38_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_496 ();
 DECAPx10_ASAP7_75t_R FILLER_38_552 ();
 DECAPx10_ASAP7_75t_R FILLER_38_574 ();
 DECAPx2_ASAP7_75t_R FILLER_38_596 ();
 DECAPx1_ASAP7_75t_R FILLER_38_608 ();
 DECAPx10_ASAP7_75t_R FILLER_38_618 ();
 DECAPx2_ASAP7_75t_R FILLER_38_640 ();
 FILLER_ASAP7_75t_R FILLER_38_646 ();
 DECAPx4_ASAP7_75t_R FILLER_38_654 ();
 FILLER_ASAP7_75t_R FILLER_38_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_672 ();
 DECAPx2_ASAP7_75t_R FILLER_38_681 ();
 FILLER_ASAP7_75t_R FILLER_38_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_709 ();
 FILLER_ASAP7_75t_R FILLER_38_713 ();
 DECAPx10_ASAP7_75t_R FILLER_38_735 ();
 DECAPx4_ASAP7_75t_R FILLER_38_757 ();
 FILLER_ASAP7_75t_R FILLER_38_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_773 ();
 DECAPx2_ASAP7_75t_R FILLER_38_797 ();
 FILLER_ASAP7_75t_R FILLER_38_803 ();
 DECAPx4_ASAP7_75t_R FILLER_38_811 ();
 DECAPx1_ASAP7_75t_R FILLER_38_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_842 ();
 DECAPx6_ASAP7_75t_R FILLER_38_849 ();
 DECAPx2_ASAP7_75t_R FILLER_38_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_869 ();
 DECAPx1_ASAP7_75t_R FILLER_38_932 ();
 DECAPx1_ASAP7_75t_R FILLER_38_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_944 ();
 DECAPx2_ASAP7_75t_R FILLER_38_960 ();
 FILLER_ASAP7_75t_R FILLER_38_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_968 ();
 FILLER_ASAP7_75t_R FILLER_38_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_977 ();
 DECAPx2_ASAP7_75t_R FILLER_38_981 ();
 FILLER_ASAP7_75t_R FILLER_38_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_998 ();
 DECAPx6_ASAP7_75t_R FILLER_38_1021 ();
 FILLER_ASAP7_75t_R FILLER_38_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1099 ();
 DECAPx4_ASAP7_75t_R FILLER_38_1112 ();
 DECAPx4_ASAP7_75t_R FILLER_38_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1187 ();
 FILLER_ASAP7_75t_R FILLER_38_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_39_2 ();
 DECAPx10_ASAP7_75t_R FILLER_39_24 ();
 DECAPx10_ASAP7_75t_R FILLER_39_46 ();
 DECAPx10_ASAP7_75t_R FILLER_39_68 ();
 DECAPx10_ASAP7_75t_R FILLER_39_90 ();
 DECAPx10_ASAP7_75t_R FILLER_39_112 ();
 DECAPx10_ASAP7_75t_R FILLER_39_134 ();
 DECAPx10_ASAP7_75t_R FILLER_39_156 ();
 DECAPx10_ASAP7_75t_R FILLER_39_178 ();
 DECAPx10_ASAP7_75t_R FILLER_39_200 ();
 DECAPx10_ASAP7_75t_R FILLER_39_222 ();
 DECAPx10_ASAP7_75t_R FILLER_39_244 ();
 DECAPx10_ASAP7_75t_R FILLER_39_266 ();
 DECAPx10_ASAP7_75t_R FILLER_39_288 ();
 DECAPx6_ASAP7_75t_R FILLER_39_310 ();
 DECAPx2_ASAP7_75t_R FILLER_39_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_330 ();
 DECAPx6_ASAP7_75t_R FILLER_39_339 ();
 DECAPx1_ASAP7_75t_R FILLER_39_353 ();
 DECAPx2_ASAP7_75t_R FILLER_39_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_371 ();
 DECAPx2_ASAP7_75t_R FILLER_39_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_385 ();
 DECAPx6_ASAP7_75t_R FILLER_39_400 ();
 FILLER_ASAP7_75t_R FILLER_39_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_416 ();
 DECAPx10_ASAP7_75t_R FILLER_39_420 ();
 DECAPx1_ASAP7_75t_R FILLER_39_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_470 ();
 FILLER_ASAP7_75t_R FILLER_39_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_495 ();
 FILLER_ASAP7_75t_R FILLER_39_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_514 ();
 DECAPx4_ASAP7_75t_R FILLER_39_518 ();
 DECAPx1_ASAP7_75t_R FILLER_39_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_535 ();
 FILLER_ASAP7_75t_R FILLER_39_539 ();
 FILLER_ASAP7_75t_R FILLER_39_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_563 ();
 FILLER_ASAP7_75t_R FILLER_39_576 ();
 DECAPx4_ASAP7_75t_R FILLER_39_584 ();
 FILLER_ASAP7_75t_R FILLER_39_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_616 ();
 DECAPx2_ASAP7_75t_R FILLER_39_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_629 ();
 DECAPx2_ASAP7_75t_R FILLER_39_650 ();
 FILLER_ASAP7_75t_R FILLER_39_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_658 ();
 DECAPx4_ASAP7_75t_R FILLER_39_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_680 ();
 DECAPx4_ASAP7_75t_R FILLER_39_708 ();
 FILLER_ASAP7_75t_R FILLER_39_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_720 ();
 DECAPx1_ASAP7_75t_R FILLER_39_743 ();
 DECAPx6_ASAP7_75t_R FILLER_39_751 ();
 DECAPx6_ASAP7_75t_R FILLER_39_785 ();
 FILLER_ASAP7_75t_R FILLER_39_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_846 ();
 FILLER_ASAP7_75t_R FILLER_39_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_855 ();
 DECAPx4_ASAP7_75t_R FILLER_39_912 ();
 FILLER_ASAP7_75t_R FILLER_39_922 ();
 DECAPx6_ASAP7_75t_R FILLER_39_926 ();
 FILLER_ASAP7_75t_R FILLER_39_940 ();
 FILLER_ASAP7_75t_R FILLER_39_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_966 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1012 ();
 DECAPx4_ASAP7_75t_R FILLER_39_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1051 ();
 FILLER_ASAP7_75t_R FILLER_39_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1059 ();
 FILLER_ASAP7_75t_R FILLER_39_1066 ();
 DECAPx4_ASAP7_75t_R FILLER_39_1085 ();
 FILLER_ASAP7_75t_R FILLER_39_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1108 ();
 FILLER_ASAP7_75t_R FILLER_39_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_39_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1185 ();
 FILLER_ASAP7_75t_R FILLER_39_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1199 ();
 FILLER_ASAP7_75t_R FILLER_39_1205 ();
 FILLER_ASAP7_75t_R FILLER_39_1215 ();
 FILLER_ASAP7_75t_R FILLER_39_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_40_2 ();
 DECAPx10_ASAP7_75t_R FILLER_40_24 ();
 DECAPx10_ASAP7_75t_R FILLER_40_46 ();
 DECAPx10_ASAP7_75t_R FILLER_40_68 ();
 DECAPx10_ASAP7_75t_R FILLER_40_90 ();
 DECAPx10_ASAP7_75t_R FILLER_40_112 ();
 DECAPx10_ASAP7_75t_R FILLER_40_134 ();
 DECAPx10_ASAP7_75t_R FILLER_40_156 ();
 DECAPx10_ASAP7_75t_R FILLER_40_178 ();
 DECAPx10_ASAP7_75t_R FILLER_40_200 ();
 DECAPx10_ASAP7_75t_R FILLER_40_222 ();
 DECAPx10_ASAP7_75t_R FILLER_40_244 ();
 DECAPx10_ASAP7_75t_R FILLER_40_266 ();
 DECAPx10_ASAP7_75t_R FILLER_40_288 ();
 DECAPx10_ASAP7_75t_R FILLER_40_310 ();
 DECAPx4_ASAP7_75t_R FILLER_40_332 ();
 DECAPx2_ASAP7_75t_R FILLER_40_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_365 ();
 DECAPx1_ASAP7_75t_R FILLER_40_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_383 ();
 DECAPx10_ASAP7_75t_R FILLER_40_418 ();
 DECAPx10_ASAP7_75t_R FILLER_40_440 ();
 DECAPx10_ASAP7_75t_R FILLER_40_464 ();
 DECAPx2_ASAP7_75t_R FILLER_40_486 ();
 FILLER_ASAP7_75t_R FILLER_40_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_511 ();
 DECAPx6_ASAP7_75t_R FILLER_40_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_532 ();
 DECAPx1_ASAP7_75t_R FILLER_40_553 ();
 DECAPx1_ASAP7_75t_R FILLER_40_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_609 ();
 FILLER_ASAP7_75t_R FILLER_40_616 ();
 DECAPx2_ASAP7_75t_R FILLER_40_640 ();
 FILLER_ASAP7_75t_R FILLER_40_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_648 ();
 DECAPx1_ASAP7_75t_R FILLER_40_659 ();
 FILLER_ASAP7_75t_R FILLER_40_674 ();
 DECAPx10_ASAP7_75t_R FILLER_40_691 ();
 DECAPx4_ASAP7_75t_R FILLER_40_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_723 ();
 DECAPx2_ASAP7_75t_R FILLER_40_727 ();
 FILLER_ASAP7_75t_R FILLER_40_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_735 ();
 FILLER_ASAP7_75t_R FILLER_40_765 ();
 FILLER_ASAP7_75t_R FILLER_40_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_772 ();
 DECAPx1_ASAP7_75t_R FILLER_40_779 ();
 DECAPx10_ASAP7_75t_R FILLER_40_786 ();
 FILLER_ASAP7_75t_R FILLER_40_808 ();
 DECAPx4_ASAP7_75t_R FILLER_40_839 ();
 FILLER_ASAP7_75t_R FILLER_40_849 ();
 DECAPx4_ASAP7_75t_R FILLER_40_861 ();
 FILLER_ASAP7_75t_R FILLER_40_871 ();
 DECAPx4_ASAP7_75t_R FILLER_40_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_903 ();
 FILLER_ASAP7_75t_R FILLER_40_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_913 ();
 DECAPx6_ASAP7_75t_R FILLER_40_917 ();
 FILLER_ASAP7_75t_R FILLER_40_951 ();
 FILLER_ASAP7_75t_R FILLER_40_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_977 ();
 FILLER_ASAP7_75t_R FILLER_40_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_992 ();
 DECAPx6_ASAP7_75t_R FILLER_40_999 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1013 ();
 DECAPx4_ASAP7_75t_R FILLER_40_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1037 ();
 FILLER_ASAP7_75t_R FILLER_40_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1078 ();
 FILLER_ASAP7_75t_R FILLER_40_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1119 ();
 FILLER_ASAP7_75t_R FILLER_40_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1155 ();
 DECAPx6_ASAP7_75t_R FILLER_40_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1191 ();
 FILLER_ASAP7_75t_R FILLER_40_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_41_2 ();
 DECAPx10_ASAP7_75t_R FILLER_41_24 ();
 DECAPx10_ASAP7_75t_R FILLER_41_46 ();
 DECAPx10_ASAP7_75t_R FILLER_41_68 ();
 DECAPx10_ASAP7_75t_R FILLER_41_90 ();
 DECAPx10_ASAP7_75t_R FILLER_41_112 ();
 DECAPx10_ASAP7_75t_R FILLER_41_134 ();
 DECAPx10_ASAP7_75t_R FILLER_41_156 ();
 DECAPx10_ASAP7_75t_R FILLER_41_178 ();
 DECAPx10_ASAP7_75t_R FILLER_41_200 ();
 DECAPx10_ASAP7_75t_R FILLER_41_222 ();
 DECAPx10_ASAP7_75t_R FILLER_41_244 ();
 DECAPx4_ASAP7_75t_R FILLER_41_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_276 ();
 DECAPx6_ASAP7_75t_R FILLER_41_321 ();
 FILLER_ASAP7_75t_R FILLER_41_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_337 ();
 FILLER_ASAP7_75t_R FILLER_41_366 ();
 DECAPx10_ASAP7_75t_R FILLER_41_376 ();
 DECAPx6_ASAP7_75t_R FILLER_41_398 ();
 FILLER_ASAP7_75t_R FILLER_41_412 ();
 DECAPx6_ASAP7_75t_R FILLER_41_444 ();
 DECAPx1_ASAP7_75t_R FILLER_41_458 ();
 DECAPx6_ASAP7_75t_R FILLER_41_482 ();
 DECAPx1_ASAP7_75t_R FILLER_41_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_500 ();
 DECAPx10_ASAP7_75t_R FILLER_41_522 ();
 DECAPx4_ASAP7_75t_R FILLER_41_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_554 ();
 DECAPx10_ASAP7_75t_R FILLER_41_558 ();
 DECAPx4_ASAP7_75t_R FILLER_41_580 ();
 FILLER_ASAP7_75t_R FILLER_41_590 ();
 FILLER_ASAP7_75t_R FILLER_41_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_600 ();
 DECAPx10_ASAP7_75t_R FILLER_41_613 ();
 DECAPx2_ASAP7_75t_R FILLER_41_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_641 ();
 DECAPx6_ASAP7_75t_R FILLER_41_655 ();
 DECAPx2_ASAP7_75t_R FILLER_41_669 ();
 DECAPx10_ASAP7_75t_R FILLER_41_687 ();
 DECAPx6_ASAP7_75t_R FILLER_41_709 ();
 DECAPx2_ASAP7_75t_R FILLER_41_729 ();
 FILLER_ASAP7_75t_R FILLER_41_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_737 ();
 DECAPx6_ASAP7_75t_R FILLER_41_741 ();
 DECAPx6_ASAP7_75t_R FILLER_41_795 ();
 DECAPx1_ASAP7_75t_R FILLER_41_809 ();
 DECAPx6_ASAP7_75t_R FILLER_41_819 ();
 DECAPx10_ASAP7_75t_R FILLER_41_851 ();
 FILLER_ASAP7_75t_R FILLER_41_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_885 ();
 DECAPx6_ASAP7_75t_R FILLER_41_892 ();
 DECAPx2_ASAP7_75t_R FILLER_41_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_912 ();
 DECAPx2_ASAP7_75t_R FILLER_41_916 ();
 FILLER_ASAP7_75t_R FILLER_41_922 ();
 DECAPx1_ASAP7_75t_R FILLER_41_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_950 ();
 DECAPx1_ASAP7_75t_R FILLER_41_955 ();
 FILLER_ASAP7_75t_R FILLER_41_979 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_41_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1046 ();
 FILLER_ASAP7_75t_R FILLER_41_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1141 ();
 DECAPx6_ASAP7_75t_R FILLER_41_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_41_1177 ();
 FILLER_ASAP7_75t_R FILLER_41_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1186 ();
 DECAPx4_ASAP7_75t_R FILLER_41_1192 ();
 FILLER_ASAP7_75t_R FILLER_41_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_42_2 ();
 DECAPx10_ASAP7_75t_R FILLER_42_24 ();
 DECAPx10_ASAP7_75t_R FILLER_42_46 ();
 DECAPx10_ASAP7_75t_R FILLER_42_68 ();
 DECAPx10_ASAP7_75t_R FILLER_42_90 ();
 DECAPx10_ASAP7_75t_R FILLER_42_112 ();
 DECAPx10_ASAP7_75t_R FILLER_42_134 ();
 DECAPx10_ASAP7_75t_R FILLER_42_156 ();
 DECAPx10_ASAP7_75t_R FILLER_42_178 ();
 DECAPx10_ASAP7_75t_R FILLER_42_200 ();
 DECAPx10_ASAP7_75t_R FILLER_42_248 ();
 DECAPx1_ASAP7_75t_R FILLER_42_270 ();
 DECAPx4_ASAP7_75t_R FILLER_42_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_301 ();
 DECAPx6_ASAP7_75t_R FILLER_42_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_356 ();
 FILLER_ASAP7_75t_R FILLER_42_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_392 ();
 DECAPx10_ASAP7_75t_R FILLER_42_415 ();
 FILLER_ASAP7_75t_R FILLER_42_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_461 ();
 DECAPx4_ASAP7_75t_R FILLER_42_464 ();
 DECAPx1_ASAP7_75t_R FILLER_42_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_514 ();
 DECAPx4_ASAP7_75t_R FILLER_42_560 ();
 DECAPx4_ASAP7_75t_R FILLER_42_610 ();
 FILLER_ASAP7_75t_R FILLER_42_620 ();
 FILLER_ASAP7_75t_R FILLER_42_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_650 ();
 FILLER_ASAP7_75t_R FILLER_42_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_656 ();
 DECAPx1_ASAP7_75t_R FILLER_42_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_679 ();
 DECAPx4_ASAP7_75t_R FILLER_42_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_703 ();
 DECAPx4_ASAP7_75t_R FILLER_42_746 ();
 DECAPx6_ASAP7_75t_R FILLER_42_759 ();
 DECAPx1_ASAP7_75t_R FILLER_42_773 ();
 DECAPx10_ASAP7_75t_R FILLER_42_780 ();
 DECAPx1_ASAP7_75t_R FILLER_42_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_841 ();
 FILLER_ASAP7_75t_R FILLER_42_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_858 ();
 DECAPx4_ASAP7_75t_R FILLER_42_862 ();
 DECAPx2_ASAP7_75t_R FILLER_42_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_891 ();
 DECAPx10_ASAP7_75t_R FILLER_42_912 ();
 DECAPx10_ASAP7_75t_R FILLER_42_934 ();
 DECAPx10_ASAP7_75t_R FILLER_42_956 ();
 DECAPx10_ASAP7_75t_R FILLER_42_978 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1022 ();
 FILLER_ASAP7_75t_R FILLER_42_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1078 ();
 DECAPx6_ASAP7_75t_R FILLER_42_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1136 ();
 DECAPx4_ASAP7_75t_R FILLER_42_1158 ();
 FILLER_ASAP7_75t_R FILLER_42_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_42_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1208 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_43_2 ();
 DECAPx10_ASAP7_75t_R FILLER_43_24 ();
 DECAPx10_ASAP7_75t_R FILLER_43_46 ();
 DECAPx10_ASAP7_75t_R FILLER_43_68 ();
 DECAPx10_ASAP7_75t_R FILLER_43_90 ();
 DECAPx10_ASAP7_75t_R FILLER_43_112 ();
 DECAPx10_ASAP7_75t_R FILLER_43_134 ();
 DECAPx4_ASAP7_75t_R FILLER_43_156 ();
 DECAPx2_ASAP7_75t_R FILLER_43_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_189 ();
 DECAPx6_ASAP7_75t_R FILLER_43_200 ();
 DECAPx2_ASAP7_75t_R FILLER_43_220 ();
 FILLER_ASAP7_75t_R FILLER_43_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_239 ();
 DECAPx6_ASAP7_75t_R FILLER_43_256 ();
 DECAPx2_ASAP7_75t_R FILLER_43_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_276 ();
 DECAPx4_ASAP7_75t_R FILLER_43_348 ();
 FILLER_ASAP7_75t_R FILLER_43_358 ();
 DECAPx6_ASAP7_75t_R FILLER_43_399 ();
 DECAPx2_ASAP7_75t_R FILLER_43_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_419 ();
 FILLER_ASAP7_75t_R FILLER_43_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_440 ();
 DECAPx2_ASAP7_75t_R FILLER_43_447 ();
 FILLER_ASAP7_75t_R FILLER_43_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_455 ();
 DECAPx1_ASAP7_75t_R FILLER_43_480 ();
 DECAPx6_ASAP7_75t_R FILLER_43_487 ();
 FILLER_ASAP7_75t_R FILLER_43_501 ();
 FILLER_ASAP7_75t_R FILLER_43_512 ();
 DECAPx4_ASAP7_75t_R FILLER_43_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_536 ();
 DECAPx2_ASAP7_75t_R FILLER_43_560 ();
 FILLER_ASAP7_75t_R FILLER_43_566 ();
 DECAPx1_ASAP7_75t_R FILLER_43_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_584 ();
 FILLER_ASAP7_75t_R FILLER_43_591 ();
 DECAPx1_ASAP7_75t_R FILLER_43_613 ();
 DECAPx6_ASAP7_75t_R FILLER_43_640 ();
 DECAPx1_ASAP7_75t_R FILLER_43_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_671 ();
 DECAPx1_ASAP7_75t_R FILLER_43_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_723 ();
 FILLER_ASAP7_75t_R FILLER_43_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_769 ();
 DECAPx10_ASAP7_75t_R FILLER_43_790 ();
 DECAPx1_ASAP7_75t_R FILLER_43_812 ();
 FILLER_ASAP7_75t_R FILLER_43_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_834 ();
 DECAPx1_ASAP7_75t_R FILLER_43_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_856 ();
 DECAPx1_ASAP7_75t_R FILLER_43_863 ();
 DECAPx6_ASAP7_75t_R FILLER_43_907 ();
 FILLER_ASAP7_75t_R FILLER_43_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_923 ();
 FILLER_ASAP7_75t_R FILLER_43_926 ();
 FILLER_ASAP7_75t_R FILLER_43_952 ();
 FILLER_ASAP7_75t_R FILLER_43_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_980 ();
 DECAPx6_ASAP7_75t_R FILLER_43_987 ();
 FILLER_ASAP7_75t_R FILLER_43_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1047 ();
 FILLER_ASAP7_75t_R FILLER_43_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1121 ();
 FILLER_ASAP7_75t_R FILLER_43_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_43_1149 ();
 FILLER_ASAP7_75t_R FILLER_43_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1167 ();
 FILLER_ASAP7_75t_R FILLER_43_1173 ();
 FILLER_ASAP7_75t_R FILLER_43_1191 ();
 FILLER_ASAP7_75t_R FILLER_43_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_44_2 ();
 DECAPx10_ASAP7_75t_R FILLER_44_24 ();
 DECAPx10_ASAP7_75t_R FILLER_44_46 ();
 DECAPx10_ASAP7_75t_R FILLER_44_68 ();
 DECAPx10_ASAP7_75t_R FILLER_44_90 ();
 DECAPx10_ASAP7_75t_R FILLER_44_112 ();
 DECAPx10_ASAP7_75t_R FILLER_44_134 ();
 DECAPx6_ASAP7_75t_R FILLER_44_156 ();
 FILLER_ASAP7_75t_R FILLER_44_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_172 ();
 DECAPx6_ASAP7_75t_R FILLER_44_193 ();
 DECAPx10_ASAP7_75t_R FILLER_44_262 ();
 DECAPx1_ASAP7_75t_R FILLER_44_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_294 ();
 FILLER_ASAP7_75t_R FILLER_44_303 ();
 DECAPx10_ASAP7_75t_R FILLER_44_335 ();
 FILLER_ASAP7_75t_R FILLER_44_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_359 ();
 DECAPx10_ASAP7_75t_R FILLER_44_366 ();
 DECAPx10_ASAP7_75t_R FILLER_44_388 ();
 DECAPx10_ASAP7_75t_R FILLER_44_410 ();
 FILLER_ASAP7_75t_R FILLER_44_432 ();
 DECAPx1_ASAP7_75t_R FILLER_44_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_458 ();
 DECAPx6_ASAP7_75t_R FILLER_44_464 ();
 DECAPx2_ASAP7_75t_R FILLER_44_478 ();
 DECAPx4_ASAP7_75t_R FILLER_44_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_506 ();
 DECAPx2_ASAP7_75t_R FILLER_44_529 ();
 FILLER_ASAP7_75t_R FILLER_44_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_537 ();
 DECAPx6_ASAP7_75t_R FILLER_44_544 ();
 DECAPx2_ASAP7_75t_R FILLER_44_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_564 ();
 DECAPx6_ASAP7_75t_R FILLER_44_638 ();
 DECAPx1_ASAP7_75t_R FILLER_44_652 ();
 DECAPx2_ASAP7_75t_R FILLER_44_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_680 ();
 DECAPx4_ASAP7_75t_R FILLER_44_689 ();
 DECAPx2_ASAP7_75t_R FILLER_44_732 ();
 FILLER_ASAP7_75t_R FILLER_44_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_740 ();
 DECAPx4_ASAP7_75t_R FILLER_44_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_757 ();
 DECAPx1_ASAP7_75t_R FILLER_44_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_768 ();
 FILLER_ASAP7_75t_R FILLER_44_775 ();
 DECAPx10_ASAP7_75t_R FILLER_44_800 ();
 FILLER_ASAP7_75t_R FILLER_44_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_824 ();
 FILLER_ASAP7_75t_R FILLER_44_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_845 ();
 FILLER_ASAP7_75t_R FILLER_44_852 ();
 DECAPx4_ASAP7_75t_R FILLER_44_857 ();
 FILLER_ASAP7_75t_R FILLER_44_867 ();
 DECAPx6_ASAP7_75t_R FILLER_44_895 ();
 DECAPx2_ASAP7_75t_R FILLER_44_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_915 ();
 DECAPx1_ASAP7_75t_R FILLER_44_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_923 ();
 DECAPx2_ASAP7_75t_R FILLER_44_927 ();
 FILLER_ASAP7_75t_R FILLER_44_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_935 ();
 FILLER_ASAP7_75t_R FILLER_44_980 ();
 FILLER_ASAP7_75t_R FILLER_44_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1037 ();
 DECAPx4_ASAP7_75t_R FILLER_44_1102 ();
 FILLER_ASAP7_75t_R FILLER_44_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1122 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1144 ();
 FILLER_ASAP7_75t_R FILLER_44_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1160 ();
 FILLER_ASAP7_75t_R FILLER_44_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1174 ();
 FILLER_ASAP7_75t_R FILLER_44_1178 ();
 FILLER_ASAP7_75t_R FILLER_44_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1216 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_45_2 ();
 DECAPx10_ASAP7_75t_R FILLER_45_24 ();
 DECAPx10_ASAP7_75t_R FILLER_45_46 ();
 DECAPx10_ASAP7_75t_R FILLER_45_68 ();
 DECAPx10_ASAP7_75t_R FILLER_45_90 ();
 DECAPx10_ASAP7_75t_R FILLER_45_112 ();
 DECAPx10_ASAP7_75t_R FILLER_45_134 ();
 DECAPx6_ASAP7_75t_R FILLER_45_156 ();
 DECAPx6_ASAP7_75t_R FILLER_45_192 ();
 DECAPx2_ASAP7_75t_R FILLER_45_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_223 ();
 DECAPx10_ASAP7_75t_R FILLER_45_238 ();
 DECAPx2_ASAP7_75t_R FILLER_45_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_301 ();
 FILLER_ASAP7_75t_R FILLER_45_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_319 ();
 DECAPx10_ASAP7_75t_R FILLER_45_334 ();
 DECAPx10_ASAP7_75t_R FILLER_45_356 ();
 DECAPx10_ASAP7_75t_R FILLER_45_378 ();
 DECAPx10_ASAP7_75t_R FILLER_45_400 ();
 DECAPx4_ASAP7_75t_R FILLER_45_422 ();
 FILLER_ASAP7_75t_R FILLER_45_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_454 ();
 DECAPx1_ASAP7_75t_R FILLER_45_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_498 ();
 FILLER_ASAP7_75t_R FILLER_45_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_507 ();
 DECAPx2_ASAP7_75t_R FILLER_45_531 ();
 FILLER_ASAP7_75t_R FILLER_45_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_539 ();
 DECAPx4_ASAP7_75t_R FILLER_45_548 ();
 DECAPx10_ASAP7_75t_R FILLER_45_561 ();
 DECAPx10_ASAP7_75t_R FILLER_45_583 ();
 DECAPx4_ASAP7_75t_R FILLER_45_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_644 ();
 FILLER_ASAP7_75t_R FILLER_45_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_659 ();
 FILLER_ASAP7_75t_R FILLER_45_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_676 ();
 DECAPx10_ASAP7_75t_R FILLER_45_690 ();
 DECAPx2_ASAP7_75t_R FILLER_45_734 ();
 FILLER_ASAP7_75t_R FILLER_45_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_742 ();
 DECAPx1_ASAP7_75t_R FILLER_45_755 ();
 FILLER_ASAP7_75t_R FILLER_45_775 ();
 DECAPx10_ASAP7_75t_R FILLER_45_800 ();
 FILLER_ASAP7_75t_R FILLER_45_822 ();
 FILLER_ASAP7_75t_R FILLER_45_839 ();
 DECAPx2_ASAP7_75t_R FILLER_45_847 ();
 FILLER_ASAP7_75t_R FILLER_45_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_855 ();
 DECAPx1_ASAP7_75t_R FILLER_45_866 ();
 DECAPx10_ASAP7_75t_R FILLER_45_876 ();
 DECAPx1_ASAP7_75t_R FILLER_45_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_902 ();
 DECAPx1_ASAP7_75t_R FILLER_45_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_920 ();
 DECAPx4_ASAP7_75t_R FILLER_45_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_936 ();
 FILLER_ASAP7_75t_R FILLER_45_957 ();
 DECAPx4_ASAP7_75t_R FILLER_45_963 ();
 FILLER_ASAP7_75t_R FILLER_45_973 ();
 DECAPx10_ASAP7_75t_R FILLER_45_981 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_45_1033 ();
 FILLER_ASAP7_75t_R FILLER_45_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1051 ();
 FILLER_ASAP7_75t_R FILLER_45_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_45_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_45_1157 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_45_1193 ();
 FILLER_ASAP7_75t_R FILLER_45_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_46_2 ();
 DECAPx10_ASAP7_75t_R FILLER_46_24 ();
 DECAPx10_ASAP7_75t_R FILLER_46_46 ();
 DECAPx10_ASAP7_75t_R FILLER_46_68 ();
 DECAPx10_ASAP7_75t_R FILLER_46_90 ();
 DECAPx10_ASAP7_75t_R FILLER_46_112 ();
 DECAPx10_ASAP7_75t_R FILLER_46_134 ();
 DECAPx6_ASAP7_75t_R FILLER_46_156 ();
 DECAPx1_ASAP7_75t_R FILLER_46_170 ();
 DECAPx2_ASAP7_75t_R FILLER_46_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_186 ();
 DECAPx6_ASAP7_75t_R FILLER_46_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_232 ();
 DECAPx10_ASAP7_75t_R FILLER_46_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_266 ();
 FILLER_ASAP7_75t_R FILLER_46_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_320 ();
 DECAPx10_ASAP7_75t_R FILLER_46_338 ();
 DECAPx10_ASAP7_75t_R FILLER_46_360 ();
 DECAPx10_ASAP7_75t_R FILLER_46_382 ();
 DECAPx6_ASAP7_75t_R FILLER_46_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_418 ();
 DECAPx4_ASAP7_75t_R FILLER_46_425 ();
 FILLER_ASAP7_75t_R FILLER_46_435 ();
 DECAPx2_ASAP7_75t_R FILLER_46_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_449 ();
 FILLER_ASAP7_75t_R FILLER_46_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_464 ();
 DECAPx2_ASAP7_75t_R FILLER_46_468 ();
 FILLER_ASAP7_75t_R FILLER_46_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_476 ();
 DECAPx2_ASAP7_75t_R FILLER_46_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_486 ();
 DECAPx1_ASAP7_75t_R FILLER_46_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_497 ();
 FILLER_ASAP7_75t_R FILLER_46_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_512 ();
 DECAPx1_ASAP7_75t_R FILLER_46_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_528 ();
 DECAPx2_ASAP7_75t_R FILLER_46_535 ();
 DECAPx10_ASAP7_75t_R FILLER_46_561 ();
 DECAPx10_ASAP7_75t_R FILLER_46_583 ();
 DECAPx10_ASAP7_75t_R FILLER_46_605 ();
 DECAPx1_ASAP7_75t_R FILLER_46_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_631 ();
 DECAPx10_ASAP7_75t_R FILLER_46_690 ();
 DECAPx1_ASAP7_75t_R FILLER_46_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_716 ();
 DECAPx6_ASAP7_75t_R FILLER_46_723 ();
 DECAPx2_ASAP7_75t_R FILLER_46_752 ();
 FILLER_ASAP7_75t_R FILLER_46_758 ();
 DECAPx1_ASAP7_75t_R FILLER_46_767 ();
 DECAPx10_ASAP7_75t_R FILLER_46_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_796 ();
 DECAPx1_ASAP7_75t_R FILLER_46_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_835 ();
 DECAPx2_ASAP7_75t_R FILLER_46_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_854 ();
 DECAPx2_ASAP7_75t_R FILLER_46_862 ();
 DECAPx2_ASAP7_75t_R FILLER_46_874 ();
 FILLER_ASAP7_75t_R FILLER_46_880 ();
 DECAPx10_ASAP7_75t_R FILLER_46_919 ();
 DECAPx6_ASAP7_75t_R FILLER_46_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_975 ();
 DECAPx10_ASAP7_75t_R FILLER_46_999 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1076 ();
 FILLER_ASAP7_75t_R FILLER_46_1098 ();
 FILLER_ASAP7_75t_R FILLER_46_1122 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1184 ();
 FILLER_ASAP7_75t_R FILLER_46_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_47_2 ();
 DECAPx10_ASAP7_75t_R FILLER_47_24 ();
 DECAPx10_ASAP7_75t_R FILLER_47_46 ();
 DECAPx10_ASAP7_75t_R FILLER_47_68 ();
 DECAPx10_ASAP7_75t_R FILLER_47_90 ();
 DECAPx10_ASAP7_75t_R FILLER_47_112 ();
 DECAPx10_ASAP7_75t_R FILLER_47_134 ();
 DECAPx6_ASAP7_75t_R FILLER_47_156 ();
 DECAPx1_ASAP7_75t_R FILLER_47_170 ();
 FILLER_ASAP7_75t_R FILLER_47_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_197 ();
 DECAPx2_ASAP7_75t_R FILLER_47_204 ();
 DECAPx4_ASAP7_75t_R FILLER_47_232 ();
 DECAPx10_ASAP7_75t_R FILLER_47_248 ();
 DECAPx2_ASAP7_75t_R FILLER_47_270 ();
 FILLER_ASAP7_75t_R FILLER_47_276 ();
 DECAPx6_ASAP7_75t_R FILLER_47_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_313 ();
 DECAPx4_ASAP7_75t_R FILLER_47_320 ();
 FILLER_ASAP7_75t_R FILLER_47_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_332 ();
 DECAPx10_ASAP7_75t_R FILLER_47_355 ();
 DECAPx10_ASAP7_75t_R FILLER_47_377 ();
 DECAPx6_ASAP7_75t_R FILLER_47_399 ();
 DECAPx1_ASAP7_75t_R FILLER_47_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_417 ();
 DECAPx1_ASAP7_75t_R FILLER_47_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_451 ();
 DECAPx2_ASAP7_75t_R FILLER_47_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_464 ();
 DECAPx1_ASAP7_75t_R FILLER_47_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_489 ();
 FILLER_ASAP7_75t_R FILLER_47_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_525 ();
 FILLER_ASAP7_75t_R FILLER_47_538 ();
 DECAPx10_ASAP7_75t_R FILLER_47_546 ();
 DECAPx10_ASAP7_75t_R FILLER_47_568 ();
 DECAPx1_ASAP7_75t_R FILLER_47_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_594 ();
 DECAPx6_ASAP7_75t_R FILLER_47_617 ();
 DECAPx2_ASAP7_75t_R FILLER_47_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_653 ();
 FILLER_ASAP7_75t_R FILLER_47_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_664 ();
 DECAPx4_ASAP7_75t_R FILLER_47_687 ();
 FILLER_ASAP7_75t_R FILLER_47_697 ();
 DECAPx4_ASAP7_75t_R FILLER_47_719 ();
 DECAPx2_ASAP7_75t_R FILLER_47_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_741 ();
 FILLER_ASAP7_75t_R FILLER_47_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_753 ();
 DECAPx6_ASAP7_75t_R FILLER_47_763 ();
 FILLER_ASAP7_75t_R FILLER_47_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_779 ();
 DECAPx4_ASAP7_75t_R FILLER_47_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_829 ();
 DECAPx1_ASAP7_75t_R FILLER_47_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_841 ();
 DECAPx2_ASAP7_75t_R FILLER_47_852 ();
 FILLER_ASAP7_75t_R FILLER_47_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_866 ();
 DECAPx4_ASAP7_75t_R FILLER_47_873 ();
 DECAPx1_ASAP7_75t_R FILLER_47_889 ();
 DECAPx4_ASAP7_75t_R FILLER_47_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_923 ();
 DECAPx6_ASAP7_75t_R FILLER_47_926 ();
 FILLER_ASAP7_75t_R FILLER_47_940 ();
 FILLER_ASAP7_75t_R FILLER_47_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_974 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1061 ();
 DECAPx6_ASAP7_75t_R FILLER_47_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_47_1097 ();
 FILLER_ASAP7_75t_R FILLER_47_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1150 ();
 FILLER_ASAP7_75t_R FILLER_47_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1182 ();
 FILLER_ASAP7_75t_R FILLER_47_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1215 ();
 FILLER_ASAP7_75t_R FILLER_47_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_48_2 ();
 DECAPx10_ASAP7_75t_R FILLER_48_24 ();
 DECAPx10_ASAP7_75t_R FILLER_48_46 ();
 DECAPx10_ASAP7_75t_R FILLER_48_68 ();
 DECAPx10_ASAP7_75t_R FILLER_48_90 ();
 DECAPx10_ASAP7_75t_R FILLER_48_112 ();
 DECAPx10_ASAP7_75t_R FILLER_48_134 ();
 DECAPx6_ASAP7_75t_R FILLER_48_156 ();
 FILLER_ASAP7_75t_R FILLER_48_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_172 ();
 DECAPx2_ASAP7_75t_R FILLER_48_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_191 ();
 FILLER_ASAP7_75t_R FILLER_48_218 ();
 DECAPx2_ASAP7_75t_R FILLER_48_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_234 ();
 DECAPx1_ASAP7_75t_R FILLER_48_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_268 ();
 DECAPx1_ASAP7_75t_R FILLER_48_280 ();
 DECAPx2_ASAP7_75t_R FILLER_48_291 ();
 DECAPx6_ASAP7_75t_R FILLER_48_304 ();
 DECAPx6_ASAP7_75t_R FILLER_48_326 ();
 DECAPx1_ASAP7_75t_R FILLER_48_340 ();
 DECAPx10_ASAP7_75t_R FILLER_48_374 ();
 DECAPx10_ASAP7_75t_R FILLER_48_396 ();
 DECAPx10_ASAP7_75t_R FILLER_48_418 ();
 FILLER_ASAP7_75t_R FILLER_48_440 ();
 DECAPx6_ASAP7_75t_R FILLER_48_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_478 ();
 DECAPx2_ASAP7_75t_R FILLER_48_493 ();
 DECAPx2_ASAP7_75t_R FILLER_48_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_508 ();
 FILLER_ASAP7_75t_R FILLER_48_521 ();
 FILLER_ASAP7_75t_R FILLER_48_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_541 ();
 FILLER_ASAP7_75t_R FILLER_48_550 ();
 DECAPx2_ASAP7_75t_R FILLER_48_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_586 ();
 DECAPx2_ASAP7_75t_R FILLER_48_609 ();
 DECAPx4_ASAP7_75t_R FILLER_48_659 ();
 DECAPx6_ASAP7_75t_R FILLER_48_683 ();
 DECAPx2_ASAP7_75t_R FILLER_48_697 ();
 DECAPx2_ASAP7_75t_R FILLER_48_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_733 ();
 DECAPx6_ASAP7_75t_R FILLER_48_753 ();
 DECAPx6_ASAP7_75t_R FILLER_48_785 ();
 FILLER_ASAP7_75t_R FILLER_48_799 ();
 DECAPx10_ASAP7_75t_R FILLER_48_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_829 ();
 FILLER_ASAP7_75t_R FILLER_48_838 ();
 DECAPx6_ASAP7_75t_R FILLER_48_846 ();
 DECAPx2_ASAP7_75t_R FILLER_48_860 ();
 DECAPx2_ASAP7_75t_R FILLER_48_886 ();
 DECAPx2_ASAP7_75t_R FILLER_48_912 ();
 FILLER_ASAP7_75t_R FILLER_48_918 ();
 DECAPx4_ASAP7_75t_R FILLER_48_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_933 ();
 DECAPx1_ASAP7_75t_R FILLER_48_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_991 ();
 DECAPx2_ASAP7_75t_R FILLER_48_998 ();
 FILLER_ASAP7_75t_R FILLER_48_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1063 ();
 FILLER_ASAP7_75t_R FILLER_48_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1108 ();
 FILLER_ASAP7_75t_R FILLER_48_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1143 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1173 ();
 FILLER_ASAP7_75t_R FILLER_48_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1204 ();
 FILLER_ASAP7_75t_R FILLER_48_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_49_2 ();
 DECAPx10_ASAP7_75t_R FILLER_49_24 ();
 DECAPx10_ASAP7_75t_R FILLER_49_46 ();
 DECAPx10_ASAP7_75t_R FILLER_49_68 ();
 DECAPx10_ASAP7_75t_R FILLER_49_90 ();
 DECAPx10_ASAP7_75t_R FILLER_49_112 ();
 DECAPx10_ASAP7_75t_R FILLER_49_134 ();
 DECAPx6_ASAP7_75t_R FILLER_49_156 ();
 DECAPx2_ASAP7_75t_R FILLER_49_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_176 ();
 FILLER_ASAP7_75t_R FILLER_49_194 ();
 DECAPx10_ASAP7_75t_R FILLER_49_203 ();
 FILLER_ASAP7_75t_R FILLER_49_225 ();
 DECAPx4_ASAP7_75t_R FILLER_49_249 ();
 DECAPx4_ASAP7_75t_R FILLER_49_287 ();
 FILLER_ASAP7_75t_R FILLER_49_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_319 ();
 DECAPx10_ASAP7_75t_R FILLER_49_348 ();
 DECAPx6_ASAP7_75t_R FILLER_49_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_384 ();
 DECAPx1_ASAP7_75t_R FILLER_49_445 ();
 DECAPx4_ASAP7_75t_R FILLER_49_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_517 ();
 DECAPx1_ASAP7_75t_R FILLER_49_526 ();
 DECAPx1_ASAP7_75t_R FILLER_49_538 ();
 DECAPx10_ASAP7_75t_R FILLER_49_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_567 ();
 DECAPx4_ASAP7_75t_R FILLER_49_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_584 ();
 DECAPx10_ASAP7_75t_R FILLER_49_607 ();
 DECAPx2_ASAP7_75t_R FILLER_49_629 ();
 FILLER_ASAP7_75t_R FILLER_49_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_637 ();
 FILLER_ASAP7_75t_R FILLER_49_657 ();
 DECAPx10_ASAP7_75t_R FILLER_49_677 ();
 DECAPx1_ASAP7_75t_R FILLER_49_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_703 ();
 DECAPx2_ASAP7_75t_R FILLER_49_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_716 ();
 DECAPx2_ASAP7_75t_R FILLER_49_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_743 ();
 DECAPx1_ASAP7_75t_R FILLER_49_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_767 ();
 DECAPx1_ASAP7_75t_R FILLER_49_774 ();
 DECAPx4_ASAP7_75t_R FILLER_49_790 ();
 FILLER_ASAP7_75t_R FILLER_49_800 ();
 DECAPx2_ASAP7_75t_R FILLER_49_824 ();
 FILLER_ASAP7_75t_R FILLER_49_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_835 ();
 DECAPx4_ASAP7_75t_R FILLER_49_863 ();
 FILLER_ASAP7_75t_R FILLER_49_873 ();
 DECAPx10_ASAP7_75t_R FILLER_49_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_923 ();
 DECAPx10_ASAP7_75t_R FILLER_49_926 ();
 DECAPx1_ASAP7_75t_R FILLER_49_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_952 ();
 DECAPx10_ASAP7_75t_R FILLER_49_975 ();
 DECAPx2_ASAP7_75t_R FILLER_49_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1032 ();
 FILLER_ASAP7_75t_R FILLER_49_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1063 ();
 DECAPx4_ASAP7_75t_R FILLER_49_1076 ();
 DECAPx4_ASAP7_75t_R FILLER_49_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1108 ();
 FILLER_ASAP7_75t_R FILLER_49_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1140 ();
 FILLER_ASAP7_75t_R FILLER_49_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_50_2 ();
 DECAPx10_ASAP7_75t_R FILLER_50_24 ();
 DECAPx10_ASAP7_75t_R FILLER_50_46 ();
 DECAPx10_ASAP7_75t_R FILLER_50_68 ();
 DECAPx10_ASAP7_75t_R FILLER_50_90 ();
 DECAPx10_ASAP7_75t_R FILLER_50_112 ();
 DECAPx10_ASAP7_75t_R FILLER_50_134 ();
 DECAPx4_ASAP7_75t_R FILLER_50_156 ();
 FILLER_ASAP7_75t_R FILLER_50_166 ();
 DECAPx10_ASAP7_75t_R FILLER_50_190 ();
 DECAPx4_ASAP7_75t_R FILLER_50_212 ();
 FILLER_ASAP7_75t_R FILLER_50_222 ();
 DECAPx10_ASAP7_75t_R FILLER_50_238 ();
 DECAPx10_ASAP7_75t_R FILLER_50_260 ();
 DECAPx1_ASAP7_75t_R FILLER_50_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_286 ();
 DECAPx2_ASAP7_75t_R FILLER_50_309 ();
 FILLER_ASAP7_75t_R FILLER_50_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_317 ();
 FILLER_ASAP7_75t_R FILLER_50_332 ();
 DECAPx2_ASAP7_75t_R FILLER_50_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_391 ();
 DECAPx10_ASAP7_75t_R FILLER_50_398 ();
 DECAPx6_ASAP7_75t_R FILLER_50_420 ();
 DECAPx2_ASAP7_75t_R FILLER_50_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_453 ();
 FILLER_ASAP7_75t_R FILLER_50_460 ();
 DECAPx1_ASAP7_75t_R FILLER_50_490 ();
 DECAPx4_ASAP7_75t_R FILLER_50_500 ();
 FILLER_ASAP7_75t_R FILLER_50_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_526 ();
 DECAPx4_ASAP7_75t_R FILLER_50_535 ();
 DECAPx2_ASAP7_75t_R FILLER_50_558 ();
 DECAPx10_ASAP7_75t_R FILLER_50_586 ();
 DECAPx4_ASAP7_75t_R FILLER_50_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_618 ();
 DECAPx1_ASAP7_75t_R FILLER_50_647 ();
 FILLER_ASAP7_75t_R FILLER_50_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_671 ();
 DECAPx2_ASAP7_75t_R FILLER_50_682 ();
 DECAPx6_ASAP7_75t_R FILLER_50_708 ();
 FILLER_ASAP7_75t_R FILLER_50_753 ();
 FILLER_ASAP7_75t_R FILLER_50_762 ();
 FILLER_ASAP7_75t_R FILLER_50_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_780 ();
 DECAPx10_ASAP7_75t_R FILLER_50_789 ();
 DECAPx2_ASAP7_75t_R FILLER_50_811 ();
 DECAPx1_ASAP7_75t_R FILLER_50_839 ();
 DECAPx1_ASAP7_75t_R FILLER_50_853 ();
 DECAPx4_ASAP7_75t_R FILLER_50_864 ();
 DECAPx4_ASAP7_75t_R FILLER_50_880 ();
 DECAPx10_ASAP7_75t_R FILLER_50_910 ();
 DECAPx1_ASAP7_75t_R FILLER_50_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_957 ();
 DECAPx6_ASAP7_75t_R FILLER_50_986 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1081 ();
 FILLER_ASAP7_75t_R FILLER_50_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1129 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1151 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_51_2 ();
 DECAPx10_ASAP7_75t_R FILLER_51_24 ();
 DECAPx10_ASAP7_75t_R FILLER_51_46 ();
 DECAPx10_ASAP7_75t_R FILLER_51_68 ();
 DECAPx10_ASAP7_75t_R FILLER_51_90 ();
 DECAPx10_ASAP7_75t_R FILLER_51_112 ();
 DECAPx10_ASAP7_75t_R FILLER_51_134 ();
 DECAPx2_ASAP7_75t_R FILLER_51_156 ();
 FILLER_ASAP7_75t_R FILLER_51_162 ();
 FILLER_ASAP7_75t_R FILLER_51_182 ();
 DECAPx2_ASAP7_75t_R FILLER_51_201 ();
 DECAPx4_ASAP7_75t_R FILLER_51_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_243 ();
 DECAPx1_ASAP7_75t_R FILLER_51_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_278 ();
 FILLER_ASAP7_75t_R FILLER_51_285 ();
 DECAPx10_ASAP7_75t_R FILLER_51_293 ();
 DECAPx2_ASAP7_75t_R FILLER_51_315 ();
 FILLER_ASAP7_75t_R FILLER_51_321 ();
 DECAPx10_ASAP7_75t_R FILLER_51_340 ();
 DECAPx2_ASAP7_75t_R FILLER_51_362 ();
 DECAPx2_ASAP7_75t_R FILLER_51_379 ();
 FILLER_ASAP7_75t_R FILLER_51_396 ();
 DECAPx4_ASAP7_75t_R FILLER_51_408 ();
 FILLER_ASAP7_75t_R FILLER_51_418 ();
 FILLER_ASAP7_75t_R FILLER_51_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_460 ();
 DECAPx1_ASAP7_75t_R FILLER_51_464 ();
 DECAPx2_ASAP7_75t_R FILLER_51_501 ();
 FILLER_ASAP7_75t_R FILLER_51_507 ();
 FILLER_ASAP7_75t_R FILLER_51_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_518 ();
 DECAPx6_ASAP7_75t_R FILLER_51_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_551 ();
 FILLER_ASAP7_75t_R FILLER_51_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_582 ();
 DECAPx6_ASAP7_75t_R FILLER_51_605 ();
 DECAPx2_ASAP7_75t_R FILLER_51_619 ();
 DECAPx6_ASAP7_75t_R FILLER_51_653 ();
 FILLER_ASAP7_75t_R FILLER_51_667 ();
 DECAPx10_ASAP7_75t_R FILLER_51_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_698 ();
 FILLER_ASAP7_75t_R FILLER_51_705 ();
 DECAPx4_ASAP7_75t_R FILLER_51_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_741 ();
 DECAPx2_ASAP7_75t_R FILLER_51_749 ();
 FILLER_ASAP7_75t_R FILLER_51_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_757 ();
 FILLER_ASAP7_75t_R FILLER_51_765 ();
 DECAPx2_ASAP7_75t_R FILLER_51_773 ();
 FILLER_ASAP7_75t_R FILLER_51_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_789 ();
 DECAPx2_ASAP7_75t_R FILLER_51_812 ();
 FILLER_ASAP7_75t_R FILLER_51_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_820 ();
 DECAPx2_ASAP7_75t_R FILLER_51_853 ();
 FILLER_ASAP7_75t_R FILLER_51_862 ();
 FILLER_ASAP7_75t_R FILLER_51_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_892 ();
 DECAPx2_ASAP7_75t_R FILLER_51_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_905 ();
 DECAPx2_ASAP7_75t_R FILLER_51_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_932 ();
 DECAPx10_ASAP7_75t_R FILLER_51_939 ();
 DECAPx6_ASAP7_75t_R FILLER_51_961 ();
 FILLER_ASAP7_75t_R FILLER_51_975 ();
 DECAPx2_ASAP7_75t_R FILLER_51_997 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_51_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1047 ();
 FILLER_ASAP7_75t_R FILLER_51_1053 ();
 FILLER_ASAP7_75t_R FILLER_51_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1120 ();
 DECAPx4_ASAP7_75t_R FILLER_51_1142 ();
 FILLER_ASAP7_75t_R FILLER_51_1152 ();
 FILLER_ASAP7_75t_R FILLER_51_1181 ();
 FILLER_ASAP7_75t_R FILLER_51_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_52_2 ();
 DECAPx10_ASAP7_75t_R FILLER_52_24 ();
 DECAPx10_ASAP7_75t_R FILLER_52_46 ();
 DECAPx10_ASAP7_75t_R FILLER_52_68 ();
 DECAPx10_ASAP7_75t_R FILLER_52_90 ();
 DECAPx10_ASAP7_75t_R FILLER_52_112 ();
 DECAPx6_ASAP7_75t_R FILLER_52_134 ();
 DECAPx1_ASAP7_75t_R FILLER_52_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_152 ();
 FILLER_ASAP7_75t_R FILLER_52_181 ();
 DECAPx10_ASAP7_75t_R FILLER_52_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_222 ();
 DECAPx10_ASAP7_75t_R FILLER_52_235 ();
 DECAPx1_ASAP7_75t_R FILLER_52_257 ();
 DECAPx6_ASAP7_75t_R FILLER_52_300 ();
 DECAPx1_ASAP7_75t_R FILLER_52_314 ();
 DECAPx10_ASAP7_75t_R FILLER_52_343 ();
 DECAPx4_ASAP7_75t_R FILLER_52_365 ();
 FILLER_ASAP7_75t_R FILLER_52_381 ();
 DECAPx10_ASAP7_75t_R FILLER_52_405 ();
 FILLER_ASAP7_75t_R FILLER_52_427 ();
 DECAPx1_ASAP7_75t_R FILLER_52_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_461 ();
 DECAPx1_ASAP7_75t_R FILLER_52_490 ();
 DECAPx10_ASAP7_75t_R FILLER_52_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_543 ();
 DECAPx1_ASAP7_75t_R FILLER_52_588 ();
 DECAPx4_ASAP7_75t_R FILLER_52_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_630 ();
 DECAPx6_ASAP7_75t_R FILLER_52_651 ();
 FILLER_ASAP7_75t_R FILLER_52_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_667 ();
 DECAPx6_ASAP7_75t_R FILLER_52_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_699 ();
 DECAPx2_ASAP7_75t_R FILLER_52_712 ();
 FILLER_ASAP7_75t_R FILLER_52_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_720 ();
 FILLER_ASAP7_75t_R FILLER_52_728 ();
 DECAPx4_ASAP7_75t_R FILLER_52_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_753 ();
 DECAPx6_ASAP7_75t_R FILLER_52_768 ();
 FILLER_ASAP7_75t_R FILLER_52_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_790 ();
 DECAPx6_ASAP7_75t_R FILLER_52_797 ();
 DECAPx1_ASAP7_75t_R FILLER_52_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_859 ();
 DECAPx10_ASAP7_75t_R FILLER_52_867 ();
 DECAPx2_ASAP7_75t_R FILLER_52_889 ();
 DECAPx6_ASAP7_75t_R FILLER_52_917 ();
 FILLER_ASAP7_75t_R FILLER_52_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_953 ();
 DECAPx1_ASAP7_75t_R FILLER_52_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_986 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_52_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1152 ();
 FILLER_ASAP7_75t_R FILLER_52_1158 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_52_1187 ();
 FILLER_ASAP7_75t_R FILLER_52_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_53_2 ();
 DECAPx10_ASAP7_75t_R FILLER_53_24 ();
 DECAPx10_ASAP7_75t_R FILLER_53_46 ();
 DECAPx10_ASAP7_75t_R FILLER_53_68 ();
 DECAPx10_ASAP7_75t_R FILLER_53_90 ();
 DECAPx10_ASAP7_75t_R FILLER_53_112 ();
 DECAPx10_ASAP7_75t_R FILLER_53_134 ();
 DECAPx6_ASAP7_75t_R FILLER_53_156 ();
 DECAPx1_ASAP7_75t_R FILLER_53_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_174 ();
 DECAPx2_ASAP7_75t_R FILLER_53_187 ();
 FILLER_ASAP7_75t_R FILLER_53_193 ();
 FILLER_ASAP7_75t_R FILLER_53_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_219 ();
 FILLER_ASAP7_75t_R FILLER_53_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_228 ();
 DECAPx2_ASAP7_75t_R FILLER_53_251 ();
 DECAPx6_ASAP7_75t_R FILLER_53_293 ();
 DECAPx1_ASAP7_75t_R FILLER_53_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_311 ();
 FILLER_ASAP7_75t_R FILLER_53_323 ();
 FILLER_ASAP7_75t_R FILLER_53_331 ();
 FILLER_ASAP7_75t_R FILLER_53_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_357 ();
 FILLER_ASAP7_75t_R FILLER_53_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_366 ();
 DECAPx2_ASAP7_75t_R FILLER_53_378 ();
 FILLER_ASAP7_75t_R FILLER_53_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_386 ();
 DECAPx4_ASAP7_75t_R FILLER_53_393 ();
 DECAPx10_ASAP7_75t_R FILLER_53_425 ();
 DECAPx10_ASAP7_75t_R FILLER_53_447 ();
 DECAPx2_ASAP7_75t_R FILLER_53_469 ();
 FILLER_ASAP7_75t_R FILLER_53_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_477 ();
 FILLER_ASAP7_75t_R FILLER_53_482 ();
 DECAPx4_ASAP7_75t_R FILLER_53_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_520 ();
 DECAPx6_ASAP7_75t_R FILLER_53_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_569 ();
 DECAPx4_ASAP7_75t_R FILLER_53_576 ();
 FILLER_ASAP7_75t_R FILLER_53_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_588 ();
 DECAPx10_ASAP7_75t_R FILLER_53_611 ();
 DECAPx4_ASAP7_75t_R FILLER_53_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_643 ();
 DECAPx10_ASAP7_75t_R FILLER_53_682 ();
 DECAPx6_ASAP7_75t_R FILLER_53_704 ();
 DECAPx2_ASAP7_75t_R FILLER_53_725 ();
 FILLER_ASAP7_75t_R FILLER_53_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_748 ();
 DECAPx4_ASAP7_75t_R FILLER_53_763 ();
 FILLER_ASAP7_75t_R FILLER_53_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_775 ();
 DECAPx6_ASAP7_75t_R FILLER_53_798 ();
 DECAPx2_ASAP7_75t_R FILLER_53_812 ();
 DECAPx1_ASAP7_75t_R FILLER_53_821 ();
 DECAPx10_ASAP7_75t_R FILLER_53_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_874 ();
 DECAPx4_ASAP7_75t_R FILLER_53_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_891 ();
 DECAPx2_ASAP7_75t_R FILLER_53_898 ();
 FILLER_ASAP7_75t_R FILLER_53_904 ();
 FILLER_ASAP7_75t_R FILLER_53_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_928 ();
 DECAPx10_ASAP7_75t_R FILLER_53_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_957 ();
 DECAPx6_ASAP7_75t_R FILLER_53_964 ();
 FILLER_ASAP7_75t_R FILLER_53_978 ();
 FILLER_ASAP7_75t_R FILLER_53_983 ();
 DECAPx2_ASAP7_75t_R FILLER_53_997 ();
 FILLER_ASAP7_75t_R FILLER_53_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1011 ();
 FILLER_ASAP7_75t_R FILLER_53_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1025 ();
 FILLER_ASAP7_75t_R FILLER_53_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1054 ();
 FILLER_ASAP7_75t_R FILLER_53_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_53_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1095 ();
 FILLER_ASAP7_75t_R FILLER_53_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_53_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1143 ();
 FILLER_ASAP7_75t_R FILLER_53_1185 ();
 DECAPx1_ASAP7_75t_R FILLER_53_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_54_2 ();
 DECAPx10_ASAP7_75t_R FILLER_54_24 ();
 DECAPx10_ASAP7_75t_R FILLER_54_46 ();
 DECAPx10_ASAP7_75t_R FILLER_54_68 ();
 DECAPx10_ASAP7_75t_R FILLER_54_90 ();
 DECAPx10_ASAP7_75t_R FILLER_54_112 ();
 DECAPx10_ASAP7_75t_R FILLER_54_134 ();
 DECAPx6_ASAP7_75t_R FILLER_54_156 ();
 DECAPx2_ASAP7_75t_R FILLER_54_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_185 ();
 FILLER_ASAP7_75t_R FILLER_54_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_199 ();
 FILLER_ASAP7_75t_R FILLER_54_215 ();
 DECAPx2_ASAP7_75t_R FILLER_54_233 ();
 FILLER_ASAP7_75t_R FILLER_54_239 ();
 DECAPx2_ASAP7_75t_R FILLER_54_263 ();
 FILLER_ASAP7_75t_R FILLER_54_269 ();
 DECAPx6_ASAP7_75t_R FILLER_54_299 ();
 FILLER_ASAP7_75t_R FILLER_54_313 ();
 DECAPx4_ASAP7_75t_R FILLER_54_339 ();
 FILLER_ASAP7_75t_R FILLER_54_349 ();
 DECAPx4_ASAP7_75t_R FILLER_54_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_404 ();
 FILLER_ASAP7_75t_R FILLER_54_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_413 ();
 DECAPx2_ASAP7_75t_R FILLER_54_420 ();
 DECAPx6_ASAP7_75t_R FILLER_54_446 ();
 FILLER_ASAP7_75t_R FILLER_54_460 ();
 DECAPx10_ASAP7_75t_R FILLER_54_464 ();
 DECAPx10_ASAP7_75t_R FILLER_54_486 ();
 DECAPx1_ASAP7_75t_R FILLER_54_508 ();
 DECAPx10_ASAP7_75t_R FILLER_54_532 ();
 DECAPx6_ASAP7_75t_R FILLER_54_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_568 ();
 DECAPx4_ASAP7_75t_R FILLER_54_591 ();
 FILLER_ASAP7_75t_R FILLER_54_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_603 ();
 DECAPx4_ASAP7_75t_R FILLER_54_626 ();
 FILLER_ASAP7_75t_R FILLER_54_636 ();
 DECAPx1_ASAP7_75t_R FILLER_54_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_662 ();
 DECAPx1_ASAP7_75t_R FILLER_54_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_680 ();
 DECAPx2_ASAP7_75t_R FILLER_54_701 ();
 FILLER_ASAP7_75t_R FILLER_54_707 ();
 DECAPx4_ASAP7_75t_R FILLER_54_715 ();
 DECAPx2_ASAP7_75t_R FILLER_54_735 ();
 FILLER_ASAP7_75t_R FILLER_54_775 ();
 DECAPx10_ASAP7_75t_R FILLER_54_797 ();
 DECAPx10_ASAP7_75t_R FILLER_54_819 ();
 DECAPx10_ASAP7_75t_R FILLER_54_841 ();
 DECAPx2_ASAP7_75t_R FILLER_54_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_937 ();
 DECAPx2_ASAP7_75t_R FILLER_54_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_986 ();
 DECAPx4_ASAP7_75t_R FILLER_54_993 ();
 FILLER_ASAP7_75t_R FILLER_54_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_54_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1166 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_55_2 ();
 DECAPx10_ASAP7_75t_R FILLER_55_24 ();
 DECAPx10_ASAP7_75t_R FILLER_55_46 ();
 DECAPx10_ASAP7_75t_R FILLER_55_68 ();
 DECAPx10_ASAP7_75t_R FILLER_55_90 ();
 DECAPx10_ASAP7_75t_R FILLER_55_112 ();
 DECAPx10_ASAP7_75t_R FILLER_55_134 ();
 DECAPx1_ASAP7_75t_R FILLER_55_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_160 ();
 FILLER_ASAP7_75t_R FILLER_55_183 ();
 DECAPx6_ASAP7_75t_R FILLER_55_212 ();
 DECAPx1_ASAP7_75t_R FILLER_55_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_230 ();
 DECAPx6_ASAP7_75t_R FILLER_55_256 ();
 DECAPx6_ASAP7_75t_R FILLER_55_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_320 ();
 DECAPx2_ASAP7_75t_R FILLER_55_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_333 ();
 DECAPx6_ASAP7_75t_R FILLER_55_356 ();
 FILLER_ASAP7_75t_R FILLER_55_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_372 ();
 DECAPx10_ASAP7_75t_R FILLER_55_381 ();
 DECAPx6_ASAP7_75t_R FILLER_55_403 ();
 FILLER_ASAP7_75t_R FILLER_55_417 ();
 DECAPx2_ASAP7_75t_R FILLER_55_436 ();
 FILLER_ASAP7_75t_R FILLER_55_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_444 ();
 DECAPx10_ASAP7_75t_R FILLER_55_455 ();
 DECAPx6_ASAP7_75t_R FILLER_55_477 ();
 DECAPx2_ASAP7_75t_R FILLER_55_491 ();
 DECAPx2_ASAP7_75t_R FILLER_55_522 ();
 FILLER_ASAP7_75t_R FILLER_55_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_530 ();
 DECAPx10_ASAP7_75t_R FILLER_55_553 ();
 DECAPx10_ASAP7_75t_R FILLER_55_575 ();
 FILLER_ASAP7_75t_R FILLER_55_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_599 ();
 DECAPx6_ASAP7_75t_R FILLER_55_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_620 ();
 DECAPx2_ASAP7_75t_R FILLER_55_643 ();
 FILLER_ASAP7_75t_R FILLER_55_649 ();
 DECAPx6_ASAP7_75t_R FILLER_55_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_687 ();
 DECAPx6_ASAP7_75t_R FILLER_55_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_708 ();
 DECAPx6_ASAP7_75t_R FILLER_55_731 ();
 FILLER_ASAP7_75t_R FILLER_55_745 ();
 FILLER_ASAP7_75t_R FILLER_55_759 ();
 DECAPx4_ASAP7_75t_R FILLER_55_765 ();
 FILLER_ASAP7_75t_R FILLER_55_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_780 ();
 DECAPx6_ASAP7_75t_R FILLER_55_803 ();
 DECAPx2_ASAP7_75t_R FILLER_55_817 ();
 FILLER_ASAP7_75t_R FILLER_55_871 ();
 DECAPx6_ASAP7_75t_R FILLER_55_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_926 ();
 FILLER_ASAP7_75t_R FILLER_55_933 ();
 DECAPx10_ASAP7_75t_R FILLER_55_941 ();
 DECAPx6_ASAP7_75t_R FILLER_55_963 ();
 FILLER_ASAP7_75t_R FILLER_55_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_992 ();
 DECAPx1_ASAP7_75t_R FILLER_55_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_55_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1069 ();
 FILLER_ASAP7_75t_R FILLER_55_1075 ();
 FILLER_ASAP7_75t_R FILLER_55_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1116 ();
 FILLER_ASAP7_75t_R FILLER_55_1122 ();
 DECAPx6_ASAP7_75t_R FILLER_55_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1195 ();
 FILLER_ASAP7_75t_R FILLER_55_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_56_2 ();
 DECAPx10_ASAP7_75t_R FILLER_56_24 ();
 DECAPx10_ASAP7_75t_R FILLER_56_46 ();
 DECAPx10_ASAP7_75t_R FILLER_56_68 ();
 DECAPx10_ASAP7_75t_R FILLER_56_90 ();
 DECAPx10_ASAP7_75t_R FILLER_56_112 ();
 DECAPx10_ASAP7_75t_R FILLER_56_134 ();
 DECAPx6_ASAP7_75t_R FILLER_56_156 ();
 DECAPx2_ASAP7_75t_R FILLER_56_170 ();
 DECAPx4_ASAP7_75t_R FILLER_56_182 ();
 FILLER_ASAP7_75t_R FILLER_56_192 ();
 DECAPx4_ASAP7_75t_R FILLER_56_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_210 ();
 DECAPx2_ASAP7_75t_R FILLER_56_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_228 ();
 DECAPx2_ASAP7_75t_R FILLER_56_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_241 ();
 DECAPx10_ASAP7_75t_R FILLER_56_248 ();
 DECAPx6_ASAP7_75t_R FILLER_56_270 ();
 DECAPx2_ASAP7_75t_R FILLER_56_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_290 ();
 DECAPx10_ASAP7_75t_R FILLER_56_319 ();
 DECAPx6_ASAP7_75t_R FILLER_56_341 ();
 FILLER_ASAP7_75t_R FILLER_56_355 ();
 DECAPx2_ASAP7_75t_R FILLER_56_383 ();
 FILLER_ASAP7_75t_R FILLER_56_389 ();
 FILLER_ASAP7_75t_R FILLER_56_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_408 ();
 DECAPx10_ASAP7_75t_R FILLER_56_422 ();
 DECAPx6_ASAP7_75t_R FILLER_56_444 ();
 DECAPx1_ASAP7_75t_R FILLER_56_458 ();
 DECAPx2_ASAP7_75t_R FILLER_56_464 ();
 FILLER_ASAP7_75t_R FILLER_56_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_472 ();
 DECAPx10_ASAP7_75t_R FILLER_56_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_517 ();
 DECAPx2_ASAP7_75t_R FILLER_56_540 ();
 FILLER_ASAP7_75t_R FILLER_56_546 ();
 DECAPx4_ASAP7_75t_R FILLER_56_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_584 ();
 DECAPx6_ASAP7_75t_R FILLER_56_605 ();
 DECAPx2_ASAP7_75t_R FILLER_56_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_625 ();
 DECAPx1_ASAP7_75t_R FILLER_56_629 ();
 DECAPx4_ASAP7_75t_R FILLER_56_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_649 ();
 FILLER_ASAP7_75t_R FILLER_56_682 ();
 DECAPx2_ASAP7_75t_R FILLER_56_732 ();
 DECAPx2_ASAP7_75t_R FILLER_56_759 ();
 DECAPx2_ASAP7_75t_R FILLER_56_773 ();
 FILLER_ASAP7_75t_R FILLER_56_799 ();
 FILLER_ASAP7_75t_R FILLER_56_807 ();
 DECAPx10_ASAP7_75t_R FILLER_56_829 ();
 DECAPx10_ASAP7_75t_R FILLER_56_873 ();
 DECAPx10_ASAP7_75t_R FILLER_56_895 ();
 DECAPx6_ASAP7_75t_R FILLER_56_917 ();
 DECAPx1_ASAP7_75t_R FILLER_56_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_935 ();
 DECAPx6_ASAP7_75t_R FILLER_56_964 ();
 FILLER_ASAP7_75t_R FILLER_56_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1063 ();
 FILLER_ASAP7_75t_R FILLER_56_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_56_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1115 ();
 FILLER_ASAP7_75t_R FILLER_56_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1124 ();
 FILLER_ASAP7_75t_R FILLER_56_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1140 ();
 FILLER_ASAP7_75t_R FILLER_56_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1148 ();
 DECAPx1_ASAP7_75t_R FILLER_56_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_57_2 ();
 DECAPx10_ASAP7_75t_R FILLER_57_24 ();
 DECAPx10_ASAP7_75t_R FILLER_57_46 ();
 DECAPx10_ASAP7_75t_R FILLER_57_68 ();
 DECAPx10_ASAP7_75t_R FILLER_57_90 ();
 DECAPx10_ASAP7_75t_R FILLER_57_112 ();
 DECAPx10_ASAP7_75t_R FILLER_57_134 ();
 DECAPx10_ASAP7_75t_R FILLER_57_156 ();
 FILLER_ASAP7_75t_R FILLER_57_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_180 ();
 DECAPx6_ASAP7_75t_R FILLER_57_192 ();
 DECAPx1_ASAP7_75t_R FILLER_57_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_210 ();
 DECAPx2_ASAP7_75t_R FILLER_57_233 ();
 FILLER_ASAP7_75t_R FILLER_57_239 ();
 DECAPx10_ASAP7_75t_R FILLER_57_263 ();
 DECAPx6_ASAP7_75t_R FILLER_57_285 ();
 DECAPx2_ASAP7_75t_R FILLER_57_299 ();
 DECAPx1_ASAP7_75t_R FILLER_57_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_352 ();
 FILLER_ASAP7_75t_R FILLER_57_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_377 ();
 DECAPx2_ASAP7_75t_R FILLER_57_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_426 ();
 DECAPx10_ASAP7_75t_R FILLER_57_449 ();
 DECAPx1_ASAP7_75t_R FILLER_57_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_475 ();
 DECAPx4_ASAP7_75t_R FILLER_57_482 ();
 FILLER_ASAP7_75t_R FILLER_57_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_515 ();
 DECAPx6_ASAP7_75t_R FILLER_57_526 ();
 DECAPx1_ASAP7_75t_R FILLER_57_540 ();
 DECAPx4_ASAP7_75t_R FILLER_57_550 ();
 FILLER_ASAP7_75t_R FILLER_57_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_584 ();
 DECAPx2_ASAP7_75t_R FILLER_57_605 ();
 FILLER_ASAP7_75t_R FILLER_57_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_613 ();
 DECAPx2_ASAP7_75t_R FILLER_57_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_626 ();
 DECAPx1_ASAP7_75t_R FILLER_57_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_645 ();
 DECAPx10_ASAP7_75t_R FILLER_57_655 ();
 DECAPx2_ASAP7_75t_R FILLER_57_677 ();
 FILLER_ASAP7_75t_R FILLER_57_683 ();
 DECAPx10_ASAP7_75t_R FILLER_57_691 ();
 DECAPx10_ASAP7_75t_R FILLER_57_713 ();
 DECAPx2_ASAP7_75t_R FILLER_57_735 ();
 DECAPx2_ASAP7_75t_R FILLER_57_744 ();
 DECAPx4_ASAP7_75t_R FILLER_57_756 ();
 FILLER_ASAP7_75t_R FILLER_57_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_768 ();
 DECAPx10_ASAP7_75t_R FILLER_57_781 ();
 DECAPx4_ASAP7_75t_R FILLER_57_803 ();
 FILLER_ASAP7_75t_R FILLER_57_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_815 ();
 FILLER_ASAP7_75t_R FILLER_57_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_862 ();
 DECAPx10_ASAP7_75t_R FILLER_57_869 ();
 DECAPx10_ASAP7_75t_R FILLER_57_891 ();
 DECAPx4_ASAP7_75t_R FILLER_57_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_923 ();
 DECAPx6_ASAP7_75t_R FILLER_57_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_960 ();
 FILLER_ASAP7_75t_R FILLER_57_968 ();
 FILLER_ASAP7_75t_R FILLER_57_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_986 ();
 DECAPx2_ASAP7_75t_R FILLER_57_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1091 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1178 ();
 FILLER_ASAP7_75t_R FILLER_57_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1203 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1213 ();
 FILLER_ASAP7_75t_R FILLER_57_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_58_2 ();
 DECAPx10_ASAP7_75t_R FILLER_58_24 ();
 DECAPx10_ASAP7_75t_R FILLER_58_46 ();
 DECAPx10_ASAP7_75t_R FILLER_58_68 ();
 DECAPx10_ASAP7_75t_R FILLER_58_90 ();
 DECAPx10_ASAP7_75t_R FILLER_58_112 ();
 DECAPx10_ASAP7_75t_R FILLER_58_134 ();
 DECAPx10_ASAP7_75t_R FILLER_58_156 ();
 DECAPx1_ASAP7_75t_R FILLER_58_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_182 ();
 DECAPx4_ASAP7_75t_R FILLER_58_205 ();
 DECAPx6_ASAP7_75t_R FILLER_58_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_245 ();
 DECAPx2_ASAP7_75t_R FILLER_58_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_273 ();
 FILLER_ASAP7_75t_R FILLER_58_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_286 ();
 FILLER_ASAP7_75t_R FILLER_58_309 ();
 FILLER_ASAP7_75t_R FILLER_58_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_319 ();
 DECAPx1_ASAP7_75t_R FILLER_58_337 ();
 DECAPx10_ASAP7_75t_R FILLER_58_351 ();
 DECAPx10_ASAP7_75t_R FILLER_58_373 ();
 DECAPx4_ASAP7_75t_R FILLER_58_408 ();
 FILLER_ASAP7_75t_R FILLER_58_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_420 ();
 FILLER_ASAP7_75t_R FILLER_58_427 ();
 DECAPx6_ASAP7_75t_R FILLER_58_435 ();
 FILLER_ASAP7_75t_R FILLER_58_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_461 ();
 DECAPx10_ASAP7_75t_R FILLER_58_464 ();
 FILLER_ASAP7_75t_R FILLER_58_486 ();
 DECAPx2_ASAP7_75t_R FILLER_58_516 ();
 DECAPx1_ASAP7_75t_R FILLER_58_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_588 ();
 DECAPx1_ASAP7_75t_R FILLER_58_607 ();
 DECAPx2_ASAP7_75t_R FILLER_58_622 ();
 DECAPx2_ASAP7_75t_R FILLER_58_640 ();
 DECAPx4_ASAP7_75t_R FILLER_58_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_663 ();
 DECAPx6_ASAP7_75t_R FILLER_58_667 ();
 DECAPx1_ASAP7_75t_R FILLER_58_681 ();
 DECAPx1_ASAP7_75t_R FILLER_58_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_695 ();
 DECAPx2_ASAP7_75t_R FILLER_58_702 ();
 FILLER_ASAP7_75t_R FILLER_58_708 ();
 DECAPx6_ASAP7_75t_R FILLER_58_730 ();
 DECAPx2_ASAP7_75t_R FILLER_58_747 ();
 DECAPx4_ASAP7_75t_R FILLER_58_760 ();
 FILLER_ASAP7_75t_R FILLER_58_770 ();
 DECAPx6_ASAP7_75t_R FILLER_58_794 ();
 DECAPx2_ASAP7_75t_R FILLER_58_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_814 ();
 FILLER_ASAP7_75t_R FILLER_58_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_826 ();
 DECAPx4_ASAP7_75t_R FILLER_58_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_859 ();
 DECAPx4_ASAP7_75t_R FILLER_58_878 ();
 DECAPx1_ASAP7_75t_R FILLER_58_912 ();
 DECAPx10_ASAP7_75t_R FILLER_58_936 ();
 DECAPx2_ASAP7_75t_R FILLER_58_958 ();
 FILLER_ASAP7_75t_R FILLER_58_964 ();
 FILLER_ASAP7_75t_R FILLER_58_978 ();
 DECAPx4_ASAP7_75t_R FILLER_58_1002 ();
 FILLER_ASAP7_75t_R FILLER_58_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1050 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1086 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1109 ();
 FILLER_ASAP7_75t_R FILLER_58_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1162 ();
 FILLER_ASAP7_75t_R FILLER_58_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1202 ();
 FILLER_ASAP7_75t_R FILLER_58_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_59_2 ();
 DECAPx10_ASAP7_75t_R FILLER_59_24 ();
 DECAPx10_ASAP7_75t_R FILLER_59_46 ();
 DECAPx10_ASAP7_75t_R FILLER_59_68 ();
 DECAPx10_ASAP7_75t_R FILLER_59_90 ();
 DECAPx10_ASAP7_75t_R FILLER_59_112 ();
 DECAPx10_ASAP7_75t_R FILLER_59_134 ();
 DECAPx10_ASAP7_75t_R FILLER_59_156 ();
 DECAPx4_ASAP7_75t_R FILLER_59_178 ();
 DECAPx1_ASAP7_75t_R FILLER_59_194 ();
 DECAPx6_ASAP7_75t_R FILLER_59_220 ();
 DECAPx2_ASAP7_75t_R FILLER_59_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_260 ();
 DECAPx2_ASAP7_75t_R FILLER_59_283 ();
 DECAPx6_ASAP7_75t_R FILLER_59_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_309 ();
 DECAPx10_ASAP7_75t_R FILLER_59_316 ();
 DECAPx6_ASAP7_75t_R FILLER_59_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_352 ();
 FILLER_ASAP7_75t_R FILLER_59_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_361 ();
 DECAPx1_ASAP7_75t_R FILLER_59_393 ();
 DECAPx6_ASAP7_75t_R FILLER_59_403 ();
 FILLER_ASAP7_75t_R FILLER_59_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_437 ();
 DECAPx1_ASAP7_75t_R FILLER_59_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_462 ();
 DECAPx4_ASAP7_75t_R FILLER_59_485 ();
 FILLER_ASAP7_75t_R FILLER_59_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_497 ();
 FILLER_ASAP7_75t_R FILLER_59_504 ();
 DECAPx2_ASAP7_75t_R FILLER_59_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_554 ();
 DECAPx2_ASAP7_75t_R FILLER_59_567 ();
 FILLER_ASAP7_75t_R FILLER_59_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_575 ();
 DECAPx10_ASAP7_75t_R FILLER_59_585 ();
 DECAPx4_ASAP7_75t_R FILLER_59_607 ();
 FILLER_ASAP7_75t_R FILLER_59_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_619 ();
 DECAPx2_ASAP7_75t_R FILLER_59_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_632 ();
 DECAPx2_ASAP7_75t_R FILLER_59_646 ();
 FILLER_ASAP7_75t_R FILLER_59_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_674 ();
 FILLER_ASAP7_75t_R FILLER_59_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_725 ();
 DECAPx6_ASAP7_75t_R FILLER_59_732 ();
 FILLER_ASAP7_75t_R FILLER_59_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_770 ();
 DECAPx10_ASAP7_75t_R FILLER_59_777 ();
 DECAPx10_ASAP7_75t_R FILLER_59_799 ();
 DECAPx6_ASAP7_75t_R FILLER_59_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_841 ();
 FILLER_ASAP7_75t_R FILLER_59_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_866 ();
 FILLER_ASAP7_75t_R FILLER_59_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_891 ();
 FILLER_ASAP7_75t_R FILLER_59_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_926 ();
 DECAPx6_ASAP7_75t_R FILLER_59_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_947 ();
 FILLER_ASAP7_75t_R FILLER_59_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_985 ();
 DECAPx2_ASAP7_75t_R FILLER_59_990 ();
 FILLER_ASAP7_75t_R FILLER_59_996 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1055 ();
 FILLER_ASAP7_75t_R FILLER_59_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_59_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1149 ();
 FILLER_ASAP7_75t_R FILLER_59_1157 ();
 FILLER_ASAP7_75t_R FILLER_59_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_59_1186 ();
 FILLER_ASAP7_75t_R FILLER_59_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1205 ();
 FILLER_ASAP7_75t_R FILLER_59_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_60_2 ();
 DECAPx10_ASAP7_75t_R FILLER_60_24 ();
 DECAPx10_ASAP7_75t_R FILLER_60_46 ();
 DECAPx10_ASAP7_75t_R FILLER_60_68 ();
 DECAPx10_ASAP7_75t_R FILLER_60_90 ();
 DECAPx10_ASAP7_75t_R FILLER_60_112 ();
 DECAPx10_ASAP7_75t_R FILLER_60_134 ();
 DECAPx10_ASAP7_75t_R FILLER_60_156 ();
 DECAPx10_ASAP7_75t_R FILLER_60_178 ();
 DECAPx1_ASAP7_75t_R FILLER_60_200 ();
 DECAPx1_ASAP7_75t_R FILLER_60_216 ();
 DECAPx2_ASAP7_75t_R FILLER_60_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_233 ();
 DECAPx2_ASAP7_75t_R FILLER_60_253 ();
 DECAPx6_ASAP7_75t_R FILLER_60_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_281 ();
 DECAPx6_ASAP7_75t_R FILLER_60_293 ();
 DECAPx2_ASAP7_75t_R FILLER_60_307 ();
 DECAPx2_ASAP7_75t_R FILLER_60_341 ();
 FILLER_ASAP7_75t_R FILLER_60_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_349 ();
 FILLER_ASAP7_75t_R FILLER_60_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_381 ();
 DECAPx4_ASAP7_75t_R FILLER_60_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_398 ();
 DECAPx4_ASAP7_75t_R FILLER_60_429 ();
 FILLER_ASAP7_75t_R FILLER_60_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_441 ();
 FILLER_ASAP7_75t_R FILLER_60_460 ();
 DECAPx6_ASAP7_75t_R FILLER_60_470 ();
 FILLER_ASAP7_75t_R FILLER_60_484 ();
 DECAPx2_ASAP7_75t_R FILLER_60_506 ();
 FILLER_ASAP7_75t_R FILLER_60_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_520 ();
 DECAPx2_ASAP7_75t_R FILLER_60_527 ();
 DECAPx1_ASAP7_75t_R FILLER_60_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_564 ();
 FILLER_ASAP7_75t_R FILLER_60_577 ();
 DECAPx4_ASAP7_75t_R FILLER_60_593 ();
 FILLER_ASAP7_75t_R FILLER_60_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_612 ();
 DECAPx2_ASAP7_75t_R FILLER_60_623 ();
 FILLER_ASAP7_75t_R FILLER_60_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_639 ();
 DECAPx10_ASAP7_75t_R FILLER_60_656 ();
 DECAPx10_ASAP7_75t_R FILLER_60_678 ();
 DECAPx6_ASAP7_75t_R FILLER_60_700 ();
 DECAPx2_ASAP7_75t_R FILLER_60_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_720 ();
 DECAPx6_ASAP7_75t_R FILLER_60_743 ();
 FILLER_ASAP7_75t_R FILLER_60_757 ();
 FILLER_ASAP7_75t_R FILLER_60_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_782 ();
 DECAPx2_ASAP7_75t_R FILLER_60_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_819 ();
 FILLER_ASAP7_75t_R FILLER_60_826 ();
 DECAPx6_ASAP7_75t_R FILLER_60_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_852 ();
 DECAPx2_ASAP7_75t_R FILLER_60_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_887 ();
 DECAPx4_ASAP7_75t_R FILLER_60_910 ();
 DECAPx6_ASAP7_75t_R FILLER_60_926 ();
 FILLER_ASAP7_75t_R FILLER_60_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_942 ();
 FILLER_ASAP7_75t_R FILLER_60_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_973 ();
 DECAPx6_ASAP7_75t_R FILLER_60_988 ();
 FILLER_ASAP7_75t_R FILLER_60_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1055 ();
 DECAPx4_ASAP7_75t_R FILLER_60_1077 ();
 FILLER_ASAP7_75t_R FILLER_60_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1140 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_60_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1168 ();
 FILLER_ASAP7_75t_R FILLER_60_1214 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_61_2 ();
 DECAPx10_ASAP7_75t_R FILLER_61_24 ();
 DECAPx10_ASAP7_75t_R FILLER_61_46 ();
 DECAPx10_ASAP7_75t_R FILLER_61_68 ();
 DECAPx10_ASAP7_75t_R FILLER_61_90 ();
 DECAPx10_ASAP7_75t_R FILLER_61_112 ();
 DECAPx10_ASAP7_75t_R FILLER_61_134 ();
 DECAPx10_ASAP7_75t_R FILLER_61_156 ();
 DECAPx4_ASAP7_75t_R FILLER_61_178 ();
 FILLER_ASAP7_75t_R FILLER_61_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_190 ();
 DECAPx2_ASAP7_75t_R FILLER_61_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_208 ();
 DECAPx1_ASAP7_75t_R FILLER_61_216 ();
 DECAPx1_ASAP7_75t_R FILLER_61_232 ();
 DECAPx4_ASAP7_75t_R FILLER_61_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_254 ();
 DECAPx10_ASAP7_75t_R FILLER_61_261 ();
 DECAPx1_ASAP7_75t_R FILLER_61_283 ();
 DECAPx4_ASAP7_75t_R FILLER_61_309 ();
 DECAPx10_ASAP7_75t_R FILLER_61_325 ();
 DECAPx10_ASAP7_75t_R FILLER_61_347 ();
 FILLER_ASAP7_75t_R FILLER_61_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_371 ();
 FILLER_ASAP7_75t_R FILLER_61_379 ();
 DECAPx10_ASAP7_75t_R FILLER_61_433 ();
 DECAPx6_ASAP7_75t_R FILLER_61_455 ();
 DECAPx1_ASAP7_75t_R FILLER_61_491 ();
 DECAPx10_ASAP7_75t_R FILLER_61_511 ();
 DECAPx4_ASAP7_75t_R FILLER_61_533 ();
 FILLER_ASAP7_75t_R FILLER_61_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_545 ();
 FILLER_ASAP7_75t_R FILLER_61_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_586 ();
 DECAPx2_ASAP7_75t_R FILLER_61_594 ();
 FILLER_ASAP7_75t_R FILLER_61_616 ();
 DECAPx1_ASAP7_75t_R FILLER_61_625 ();
 DECAPx6_ASAP7_75t_R FILLER_61_635 ();
 DECAPx1_ASAP7_75t_R FILLER_61_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_673 ();
 DECAPx2_ASAP7_75t_R FILLER_61_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_686 ();
 FILLER_ASAP7_75t_R FILLER_61_715 ();
 DECAPx4_ASAP7_75t_R FILLER_61_723 ();
 FILLER_ASAP7_75t_R FILLER_61_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_764 ();
 FILLER_ASAP7_75t_R FILLER_61_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_803 ();
 FILLER_ASAP7_75t_R FILLER_61_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_838 ();
 FILLER_ASAP7_75t_R FILLER_61_847 ();
 DECAPx6_ASAP7_75t_R FILLER_61_857 ();
 DECAPx1_ASAP7_75t_R FILLER_61_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_875 ();
 DECAPx10_ASAP7_75t_R FILLER_61_896 ();
 DECAPx2_ASAP7_75t_R FILLER_61_918 ();
 DECAPx10_ASAP7_75t_R FILLER_61_926 ();
 DECAPx6_ASAP7_75t_R FILLER_61_948 ();
 FILLER_ASAP7_75t_R FILLER_61_962 ();
 DECAPx2_ASAP7_75t_R FILLER_61_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_976 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1043 ();
 FILLER_ASAP7_75t_R FILLER_61_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1074 ();
 FILLER_ASAP7_75t_R FILLER_61_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_61_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1096 ();
 DECAPx6_ASAP7_75t_R FILLER_61_1103 ();
 FILLER_ASAP7_75t_R FILLER_61_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_62_2 ();
 DECAPx10_ASAP7_75t_R FILLER_62_24 ();
 DECAPx10_ASAP7_75t_R FILLER_62_46 ();
 DECAPx10_ASAP7_75t_R FILLER_62_68 ();
 DECAPx10_ASAP7_75t_R FILLER_62_90 ();
 DECAPx10_ASAP7_75t_R FILLER_62_112 ();
 DECAPx10_ASAP7_75t_R FILLER_62_134 ();
 DECAPx10_ASAP7_75t_R FILLER_62_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_207 ();
 DECAPx1_ASAP7_75t_R FILLER_62_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_219 ();
 FILLER_ASAP7_75t_R FILLER_62_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_234 ();
 DECAPx4_ASAP7_75t_R FILLER_62_268 ();
 FILLER_ASAP7_75t_R FILLER_62_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_280 ();
 FILLER_ASAP7_75t_R FILLER_62_306 ();
 DECAPx2_ASAP7_75t_R FILLER_62_329 ();
 DECAPx2_ASAP7_75t_R FILLER_62_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_348 ();
 DECAPx10_ASAP7_75t_R FILLER_62_359 ();
 DECAPx10_ASAP7_75t_R FILLER_62_381 ();
 DECAPx6_ASAP7_75t_R FILLER_62_403 ();
 DECAPx2_ASAP7_75t_R FILLER_62_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_423 ();
 DECAPx1_ASAP7_75t_R FILLER_62_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_461 ();
 DECAPx4_ASAP7_75t_R FILLER_62_464 ();
 FILLER_ASAP7_75t_R FILLER_62_474 ();
 DECAPx10_ASAP7_75t_R FILLER_62_524 ();
 DECAPx10_ASAP7_75t_R FILLER_62_546 ();
 DECAPx1_ASAP7_75t_R FILLER_62_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_572 ();
 FILLER_ASAP7_75t_R FILLER_62_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_578 ();
 FILLER_ASAP7_75t_R FILLER_62_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_587 ();
 FILLER_ASAP7_75t_R FILLER_62_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_607 ();
 DECAPx2_ASAP7_75t_R FILLER_62_618 ();
 DECAPx4_ASAP7_75t_R FILLER_62_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_648 ();
 DECAPx6_ASAP7_75t_R FILLER_62_655 ();
 DECAPx1_ASAP7_75t_R FILLER_62_669 ();
 DECAPx6_ASAP7_75t_R FILLER_62_699 ();
 FILLER_ASAP7_75t_R FILLER_62_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_758 ();
 DECAPx2_ASAP7_75t_R FILLER_62_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_771 ();
 DECAPx6_ASAP7_75t_R FILLER_62_778 ();
 DECAPx1_ASAP7_75t_R FILLER_62_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_796 ();
 DECAPx2_ASAP7_75t_R FILLER_62_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_818 ();
 FILLER_ASAP7_75t_R FILLER_62_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_827 ();
 DECAPx6_ASAP7_75t_R FILLER_62_838 ();
 DECAPx10_ASAP7_75t_R FILLER_62_860 ();
 DECAPx10_ASAP7_75t_R FILLER_62_882 ();
 DECAPx6_ASAP7_75t_R FILLER_62_904 ();
 FILLER_ASAP7_75t_R FILLER_62_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_974 ();
 FILLER_ASAP7_75t_R FILLER_62_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1018 ();
 FILLER_ASAP7_75t_R FILLER_62_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1068 ();
 FILLER_ASAP7_75t_R FILLER_62_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1081 ();
 FILLER_ASAP7_75t_R FILLER_62_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1093 ();
 FILLER_ASAP7_75t_R FILLER_62_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1133 ();
 FILLER_ASAP7_75t_R FILLER_62_1155 ();
 FILLER_ASAP7_75t_R FILLER_62_1171 ();
 FILLER_ASAP7_75t_R FILLER_62_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1200 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_63_2 ();
 DECAPx10_ASAP7_75t_R FILLER_63_24 ();
 DECAPx10_ASAP7_75t_R FILLER_63_46 ();
 DECAPx10_ASAP7_75t_R FILLER_63_68 ();
 DECAPx10_ASAP7_75t_R FILLER_63_90 ();
 DECAPx10_ASAP7_75t_R FILLER_63_112 ();
 DECAPx10_ASAP7_75t_R FILLER_63_134 ();
 DECAPx10_ASAP7_75t_R FILLER_63_156 ();
 DECAPx10_ASAP7_75t_R FILLER_63_178 ();
 DECAPx10_ASAP7_75t_R FILLER_63_218 ();
 DECAPx10_ASAP7_75t_R FILLER_63_240 ();
 DECAPx2_ASAP7_75t_R FILLER_63_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_296 ();
 DECAPx1_ASAP7_75t_R FILLER_63_304 ();
 DECAPx4_ASAP7_75t_R FILLER_63_315 ();
 DECAPx6_ASAP7_75t_R FILLER_63_342 ();
 DECAPx1_ASAP7_75t_R FILLER_63_356 ();
 DECAPx6_ASAP7_75t_R FILLER_63_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_433 ();
 DECAPx10_ASAP7_75t_R FILLER_63_440 ();
 DECAPx6_ASAP7_75t_R FILLER_63_462 ();
 FILLER_ASAP7_75t_R FILLER_63_476 ();
 DECAPx10_ASAP7_75t_R FILLER_63_500 ();
 DECAPx1_ASAP7_75t_R FILLER_63_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_526 ();
 DECAPx4_ASAP7_75t_R FILLER_63_532 ();
 FILLER_ASAP7_75t_R FILLER_63_542 ();
 DECAPx1_ASAP7_75t_R FILLER_63_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_564 ();
 FILLER_ASAP7_75t_R FILLER_63_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_592 ();
 DECAPx1_ASAP7_75t_R FILLER_63_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_609 ();
 DECAPx2_ASAP7_75t_R FILLER_63_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_633 ();
 DECAPx2_ASAP7_75t_R FILLER_63_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_682 ();
 DECAPx6_ASAP7_75t_R FILLER_63_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_739 ();
 DECAPx10_ASAP7_75t_R FILLER_63_746 ();
 DECAPx10_ASAP7_75t_R FILLER_63_768 ();
 DECAPx2_ASAP7_75t_R FILLER_63_790 ();
 FILLER_ASAP7_75t_R FILLER_63_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_817 ();
 DECAPx2_ASAP7_75t_R FILLER_63_824 ();
 FILLER_ASAP7_75t_R FILLER_63_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_849 ();
 DECAPx10_ASAP7_75t_R FILLER_63_888 ();
 DECAPx6_ASAP7_75t_R FILLER_63_910 ();
 FILLER_ASAP7_75t_R FILLER_63_926 ();
 FILLER_ASAP7_75t_R FILLER_63_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_950 ();
 FILLER_ASAP7_75t_R FILLER_63_971 ();
 DECAPx2_ASAP7_75t_R FILLER_63_995 ();
 FILLER_ASAP7_75t_R FILLER_63_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1017 ();
 FILLER_ASAP7_75t_R FILLER_63_1039 ();
 FILLER_ASAP7_75t_R FILLER_63_1075 ();
 FILLER_ASAP7_75t_R FILLER_63_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1112 ();
 FILLER_ASAP7_75t_R FILLER_63_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1171 ();
 DECAPx4_ASAP7_75t_R FILLER_63_1179 ();
 FILLER_ASAP7_75t_R FILLER_63_1189 ();
 FILLER_ASAP7_75t_R FILLER_63_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_64_2 ();
 DECAPx10_ASAP7_75t_R FILLER_64_24 ();
 DECAPx10_ASAP7_75t_R FILLER_64_46 ();
 DECAPx10_ASAP7_75t_R FILLER_64_68 ();
 DECAPx2_ASAP7_75t_R FILLER_64_90 ();
 FILLER_ASAP7_75t_R FILLER_64_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_98 ();
 DECAPx10_ASAP7_75t_R FILLER_64_133 ();
 DECAPx10_ASAP7_75t_R FILLER_64_155 ();
 DECAPx10_ASAP7_75t_R FILLER_64_177 ();
 DECAPx2_ASAP7_75t_R FILLER_64_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_205 ();
 DECAPx6_ASAP7_75t_R FILLER_64_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_228 ();
 DECAPx2_ASAP7_75t_R FILLER_64_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_282 ();
 DECAPx2_ASAP7_75t_R FILLER_64_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_297 ();
 DECAPx1_ASAP7_75t_R FILLER_64_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_308 ();
 FILLER_ASAP7_75t_R FILLER_64_321 ();
 DECAPx1_ASAP7_75t_R FILLER_64_329 ();
 FILLER_ASAP7_75t_R FILLER_64_355 ();
 DECAPx1_ASAP7_75t_R FILLER_64_377 ();
 DECAPx1_ASAP7_75t_R FILLER_64_392 ();
 DECAPx6_ASAP7_75t_R FILLER_64_408 ();
 DECAPx2_ASAP7_75t_R FILLER_64_422 ();
 DECAPx2_ASAP7_75t_R FILLER_64_456 ();
 DECAPx10_ASAP7_75t_R FILLER_64_464 ();
 DECAPx1_ASAP7_75t_R FILLER_64_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_490 ();
 FILLER_ASAP7_75t_R FILLER_64_517 ();
 DECAPx6_ASAP7_75t_R FILLER_64_525 ();
 FILLER_ASAP7_75t_R FILLER_64_539 ();
 DECAPx6_ASAP7_75t_R FILLER_64_558 ();
 DECAPx2_ASAP7_75t_R FILLER_64_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_578 ();
 DECAPx1_ASAP7_75t_R FILLER_64_597 ();
 DECAPx2_ASAP7_75t_R FILLER_64_607 ();
 FILLER_ASAP7_75t_R FILLER_64_613 ();
 DECAPx6_ASAP7_75t_R FILLER_64_623 ();
 DECAPx1_ASAP7_75t_R FILLER_64_657 ();
 DECAPx2_ASAP7_75t_R FILLER_64_695 ();
 FILLER_ASAP7_75t_R FILLER_64_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_703 ();
 FILLER_ASAP7_75t_R FILLER_64_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_712 ();
 DECAPx6_ASAP7_75t_R FILLER_64_751 ();
 FILLER_ASAP7_75t_R FILLER_64_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_767 ();
 FILLER_ASAP7_75t_R FILLER_64_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_805 ();
 DECAPx1_ASAP7_75t_R FILLER_64_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_819 ();
 FILLER_ASAP7_75t_R FILLER_64_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_828 ();
 DECAPx2_ASAP7_75t_R FILLER_64_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_853 ();
 DECAPx1_ASAP7_75t_R FILLER_64_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_880 ();
 DECAPx10_ASAP7_75t_R FILLER_64_887 ();
 FILLER_ASAP7_75t_R FILLER_64_909 ();
 DECAPx2_ASAP7_75t_R FILLER_64_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_939 ();
 DECAPx2_ASAP7_75t_R FILLER_64_965 ();
 FILLER_ASAP7_75t_R FILLER_64_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_973 ();
 DECAPx6_ASAP7_75t_R FILLER_64_988 ();
 DECAPx1_ASAP7_75t_R FILLER_64_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1020 ();
 FILLER_ASAP7_75t_R FILLER_64_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1059 ();
 FILLER_ASAP7_75t_R FILLER_64_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_64_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1152 ();
 FILLER_ASAP7_75t_R FILLER_64_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1176 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1183 ();
 FILLER_ASAP7_75t_R FILLER_64_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1212 ();
 FILLER_ASAP7_75t_R FILLER_64_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_65_2 ();
 DECAPx10_ASAP7_75t_R FILLER_65_24 ();
 DECAPx10_ASAP7_75t_R FILLER_65_46 ();
 DECAPx10_ASAP7_75t_R FILLER_65_68 ();
 DECAPx6_ASAP7_75t_R FILLER_65_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_104 ();
 DECAPx2_ASAP7_75t_R FILLER_65_116 ();
 FILLER_ASAP7_75t_R FILLER_65_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_124 ();
 DECAPx1_ASAP7_75t_R FILLER_65_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_151 ();
 DECAPx4_ASAP7_75t_R FILLER_65_158 ();
 FILLER_ASAP7_75t_R FILLER_65_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_170 ();
 DECAPx2_ASAP7_75t_R FILLER_65_177 ();
 FILLER_ASAP7_75t_R FILLER_65_183 ();
 DECAPx1_ASAP7_75t_R FILLER_65_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_217 ();
 DECAPx6_ASAP7_75t_R FILLER_65_224 ();
 FILLER_ASAP7_75t_R FILLER_65_238 ();
 DECAPx2_ASAP7_75t_R FILLER_65_273 ();
 FILLER_ASAP7_75t_R FILLER_65_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_281 ();
 DECAPx6_ASAP7_75t_R FILLER_65_288 ();
 FILLER_ASAP7_75t_R FILLER_65_302 ();
 FILLER_ASAP7_75t_R FILLER_65_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_318 ();
 DECAPx6_ASAP7_75t_R FILLER_65_333 ();
 DECAPx2_ASAP7_75t_R FILLER_65_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_353 ();
 DECAPx6_ASAP7_75t_R FILLER_65_364 ();
 FILLER_ASAP7_75t_R FILLER_65_378 ();
 DECAPx4_ASAP7_75t_R FILLER_65_409 ();
 DECAPx10_ASAP7_75t_R FILLER_65_427 ();
 DECAPx10_ASAP7_75t_R FILLER_65_449 ();
 FILLER_ASAP7_75t_R FILLER_65_471 ();
 DECAPx6_ASAP7_75t_R FILLER_65_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_514 ();
 FILLER_ASAP7_75t_R FILLER_65_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_549 ();
 FILLER_ASAP7_75t_R FILLER_65_563 ();
 DECAPx2_ASAP7_75t_R FILLER_65_577 ();
 FILLER_ASAP7_75t_R FILLER_65_583 ();
 FILLER_ASAP7_75t_R FILLER_65_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_596 ();
 DECAPx6_ASAP7_75t_R FILLER_65_600 ();
 DECAPx6_ASAP7_75t_R FILLER_65_624 ();
 FILLER_ASAP7_75t_R FILLER_65_638 ();
 DECAPx10_ASAP7_75t_R FILLER_65_648 ();
 DECAPx10_ASAP7_75t_R FILLER_65_670 ();
 DECAPx4_ASAP7_75t_R FILLER_65_692 ();
 FILLER_ASAP7_75t_R FILLER_65_702 ();
 DECAPx6_ASAP7_75t_R FILLER_65_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_730 ();
 DECAPx10_ASAP7_75t_R FILLER_65_753 ();
 DECAPx6_ASAP7_75t_R FILLER_65_775 ();
 DECAPx1_ASAP7_75t_R FILLER_65_789 ();
 FILLER_ASAP7_75t_R FILLER_65_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_809 ();
 DECAPx4_ASAP7_75t_R FILLER_65_836 ();
 FILLER_ASAP7_75t_R FILLER_65_846 ();
 DECAPx2_ASAP7_75t_R FILLER_65_876 ();
 FILLER_ASAP7_75t_R FILLER_65_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_884 ();
 DECAPx6_ASAP7_75t_R FILLER_65_903 ();
 DECAPx2_ASAP7_75t_R FILLER_65_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_923 ();
 DECAPx6_ASAP7_75t_R FILLER_65_932 ();
 FILLER_ASAP7_75t_R FILLER_65_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_948 ();
 DECAPx10_ASAP7_75t_R FILLER_65_986 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1024 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1050 ();
 FILLER_ASAP7_75t_R FILLER_65_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_65_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1115 ();
 FILLER_ASAP7_75t_R FILLER_65_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1161 ();
 FILLER_ASAP7_75t_R FILLER_65_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1208 ();
 FILLER_ASAP7_75t_R FILLER_65_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_66_2 ();
 DECAPx10_ASAP7_75t_R FILLER_66_24 ();
 DECAPx10_ASAP7_75t_R FILLER_66_46 ();
 DECAPx6_ASAP7_75t_R FILLER_66_68 ();
 DECAPx1_ASAP7_75t_R FILLER_66_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_109 ();
 FILLER_ASAP7_75t_R FILLER_66_117 ();
 DECAPx6_ASAP7_75t_R FILLER_66_130 ();
 FILLER_ASAP7_75t_R FILLER_66_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_146 ();
 DECAPx10_ASAP7_75t_R FILLER_66_191 ();
 FILLER_ASAP7_75t_R FILLER_66_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_215 ();
 FILLER_ASAP7_75t_R FILLER_66_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_240 ();
 DECAPx6_ASAP7_75t_R FILLER_66_247 ();
 DECAPx2_ASAP7_75t_R FILLER_66_261 ();
 DECAPx1_ASAP7_75t_R FILLER_66_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_310 ();
 FILLER_ASAP7_75t_R FILLER_66_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_324 ();
 DECAPx2_ASAP7_75t_R FILLER_66_347 ();
 FILLER_ASAP7_75t_R FILLER_66_353 ();
 DECAPx2_ASAP7_75t_R FILLER_66_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_383 ();
 DECAPx2_ASAP7_75t_R FILLER_66_390 ();
 DECAPx1_ASAP7_75t_R FILLER_66_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_461 ();
 DECAPx6_ASAP7_75t_R FILLER_66_464 ();
 FILLER_ASAP7_75t_R FILLER_66_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_533 ();
 FILLER_ASAP7_75t_R FILLER_66_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_557 ();
 DECAPx6_ASAP7_75t_R FILLER_66_565 ();
 DECAPx1_ASAP7_75t_R FILLER_66_579 ();
 FILLER_ASAP7_75t_R FILLER_66_589 ();
 DECAPx2_ASAP7_75t_R FILLER_66_610 ();
 FILLER_ASAP7_75t_R FILLER_66_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_626 ();
 DECAPx2_ASAP7_75t_R FILLER_66_633 ();
 FILLER_ASAP7_75t_R FILLER_66_639 ();
 DECAPx1_ASAP7_75t_R FILLER_66_647 ();
 DECAPx10_ASAP7_75t_R FILLER_66_657 ();
 DECAPx10_ASAP7_75t_R FILLER_66_679 ();
 DECAPx10_ASAP7_75t_R FILLER_66_723 ();
 DECAPx2_ASAP7_75t_R FILLER_66_745 ();
 FILLER_ASAP7_75t_R FILLER_66_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_776 ();
 DECAPx2_ASAP7_75t_R FILLER_66_807 ();
 FILLER_ASAP7_75t_R FILLER_66_813 ();
 DECAPx10_ASAP7_75t_R FILLER_66_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_843 ();
 DECAPx2_ASAP7_75t_R FILLER_66_852 ();
 FILLER_ASAP7_75t_R FILLER_66_858 ();
 DECAPx4_ASAP7_75t_R FILLER_66_890 ();
 DECAPx1_ASAP7_75t_R FILLER_66_918 ();
 DECAPx10_ASAP7_75t_R FILLER_66_944 ();
 DECAPx1_ASAP7_75t_R FILLER_66_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_970 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1041 ();
 FILLER_ASAP7_75t_R FILLER_66_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1069 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1091 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1137 ();
 FILLER_ASAP7_75t_R FILLER_66_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1171 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_67_2 ();
 DECAPx10_ASAP7_75t_R FILLER_67_24 ();
 DECAPx10_ASAP7_75t_R FILLER_67_46 ();
 DECAPx10_ASAP7_75t_R FILLER_67_68 ();
 DECAPx6_ASAP7_75t_R FILLER_67_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_110 ();
 DECAPx2_ASAP7_75t_R FILLER_67_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_142 ();
 DECAPx2_ASAP7_75t_R FILLER_67_154 ();
 FILLER_ASAP7_75t_R FILLER_67_160 ();
 DECAPx10_ASAP7_75t_R FILLER_67_173 ();
 FILLER_ASAP7_75t_R FILLER_67_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_219 ();
 DECAPx2_ASAP7_75t_R FILLER_67_233 ();
 FILLER_ASAP7_75t_R FILLER_67_239 ();
 DECAPx4_ASAP7_75t_R FILLER_67_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_262 ();
 DECAPx10_ASAP7_75t_R FILLER_67_285 ();
 DECAPx10_ASAP7_75t_R FILLER_67_307 ();
 DECAPx2_ASAP7_75t_R FILLER_67_329 ();
 DECAPx4_ASAP7_75t_R FILLER_67_345 ();
 DECAPx10_ASAP7_75t_R FILLER_67_378 ();
 DECAPx6_ASAP7_75t_R FILLER_67_423 ();
 FILLER_ASAP7_75t_R FILLER_67_437 ();
 DECAPx10_ASAP7_75t_R FILLER_67_456 ();
 DECAPx4_ASAP7_75t_R FILLER_67_478 ();
 FILLER_ASAP7_75t_R FILLER_67_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_490 ();
 DECAPx6_ASAP7_75t_R FILLER_67_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_518 ();
 FILLER_ASAP7_75t_R FILLER_67_529 ();
 DECAPx10_ASAP7_75t_R FILLER_67_555 ();
 DECAPx1_ASAP7_75t_R FILLER_67_577 ();
 DECAPx2_ASAP7_75t_R FILLER_67_591 ();
 FILLER_ASAP7_75t_R FILLER_67_597 ();
 DECAPx10_ASAP7_75t_R FILLER_67_611 ();
 DECAPx6_ASAP7_75t_R FILLER_67_633 ();
 DECAPx1_ASAP7_75t_R FILLER_67_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_692 ();
 DECAPx10_ASAP7_75t_R FILLER_67_715 ();
 DECAPx4_ASAP7_75t_R FILLER_67_737 ();
 FILLER_ASAP7_75t_R FILLER_67_747 ();
 DECAPx6_ASAP7_75t_R FILLER_67_793 ();
 DECAPx2_ASAP7_75t_R FILLER_67_807 ();
 FILLER_ASAP7_75t_R FILLER_67_824 ();
 DECAPx1_ASAP7_75t_R FILLER_67_838 ();
 DECAPx10_ASAP7_75t_R FILLER_67_885 ();
 DECAPx6_ASAP7_75t_R FILLER_67_907 ();
 FILLER_ASAP7_75t_R FILLER_67_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_923 ();
 DECAPx1_ASAP7_75t_R FILLER_67_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_930 ();
 DECAPx6_ASAP7_75t_R FILLER_67_937 ();
 FILLER_ASAP7_75t_R FILLER_67_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_977 ();
 DECAPx2_ASAP7_75t_R FILLER_67_981 ();
 FILLER_ASAP7_75t_R FILLER_67_987 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_67_1036 ();
 FILLER_ASAP7_75t_R FILLER_67_1046 ();
 FILLER_ASAP7_75t_R FILLER_67_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1086 ();
 FILLER_ASAP7_75t_R FILLER_67_1109 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1166 ();
 FILLER_ASAP7_75t_R FILLER_67_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1174 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1182 ();
 FILLER_ASAP7_75t_R FILLER_67_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1190 ();
 DECAPx4_ASAP7_75t_R FILLER_67_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_68_2 ();
 DECAPx10_ASAP7_75t_R FILLER_68_24 ();
 DECAPx10_ASAP7_75t_R FILLER_68_46 ();
 DECAPx10_ASAP7_75t_R FILLER_68_68 ();
 DECAPx4_ASAP7_75t_R FILLER_68_90 ();
 FILLER_ASAP7_75t_R FILLER_68_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_102 ();
 FILLER_ASAP7_75t_R FILLER_68_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_117 ();
 DECAPx1_ASAP7_75t_R FILLER_68_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_130 ();
 FILLER_ASAP7_75t_R FILLER_68_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_139 ();
 DECAPx2_ASAP7_75t_R FILLER_68_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_174 ();
 DECAPx1_ASAP7_75t_R FILLER_68_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_224 ();
 FILLER_ASAP7_75t_R FILLER_68_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_233 ();
 DECAPx1_ASAP7_75t_R FILLER_68_243 ();
 DECAPx4_ASAP7_75t_R FILLER_68_269 ();
 FILLER_ASAP7_75t_R FILLER_68_279 ();
 DECAPx2_ASAP7_75t_R FILLER_68_303 ();
 FILLER_ASAP7_75t_R FILLER_68_309 ();
 DECAPx6_ASAP7_75t_R FILLER_68_317 ();
 DECAPx2_ASAP7_75t_R FILLER_68_337 ();
 FILLER_ASAP7_75t_R FILLER_68_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_367 ();
 DECAPx6_ASAP7_75t_R FILLER_68_401 ();
 DECAPx1_ASAP7_75t_R FILLER_68_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_426 ();
 DECAPx10_ASAP7_75t_R FILLER_68_434 ();
 DECAPx2_ASAP7_75t_R FILLER_68_456 ();
 DECAPx2_ASAP7_75t_R FILLER_68_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_496 ();
 DECAPx1_ASAP7_75t_R FILLER_68_517 ();
 DECAPx6_ASAP7_75t_R FILLER_68_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_539 ();
 DECAPx2_ASAP7_75t_R FILLER_68_554 ();
 FILLER_ASAP7_75t_R FILLER_68_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_568 ();
 DECAPx2_ASAP7_75t_R FILLER_68_609 ();
 FILLER_ASAP7_75t_R FILLER_68_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_617 ();
 FILLER_ASAP7_75t_R FILLER_68_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_636 ();
 DECAPx1_ASAP7_75t_R FILLER_68_665 ();
 DECAPx2_ASAP7_75t_R FILLER_68_691 ();
 FILLER_ASAP7_75t_R FILLER_68_697 ();
 DECAPx4_ASAP7_75t_R FILLER_68_705 ();
 FILLER_ASAP7_75t_R FILLER_68_715 ();
 DECAPx2_ASAP7_75t_R FILLER_68_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_751 ();
 DECAPx2_ASAP7_75t_R FILLER_68_772 ();
 DECAPx1_ASAP7_75t_R FILLER_68_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_796 ();
 FILLER_ASAP7_75t_R FILLER_68_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_815 ();
 DECAPx2_ASAP7_75t_R FILLER_68_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_845 ();
 DECAPx6_ASAP7_75t_R FILLER_68_854 ();
 DECAPx2_ASAP7_75t_R FILLER_68_868 ();
 DECAPx2_ASAP7_75t_R FILLER_68_904 ();
 FILLER_ASAP7_75t_R FILLER_68_910 ();
 DECAPx1_ASAP7_75t_R FILLER_68_956 ();
 FILLER_ASAP7_75t_R FILLER_68_982 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1102 ();
 FILLER_ASAP7_75t_R FILLER_68_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_68_1130 ();
 FILLER_ASAP7_75t_R FILLER_68_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1166 ();
 FILLER_ASAP7_75t_R FILLER_68_1174 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1182 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_69_2 ();
 DECAPx10_ASAP7_75t_R FILLER_69_24 ();
 DECAPx10_ASAP7_75t_R FILLER_69_46 ();
 DECAPx6_ASAP7_75t_R FILLER_69_68 ();
 DECAPx2_ASAP7_75t_R FILLER_69_82 ();
 DECAPx2_ASAP7_75t_R FILLER_69_110 ();
 FILLER_ASAP7_75t_R FILLER_69_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_126 ();
 DECAPx2_ASAP7_75t_R FILLER_69_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_153 ();
 FILLER_ASAP7_75t_R FILLER_69_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_181 ();
 DECAPx10_ASAP7_75t_R FILLER_69_190 ();
 DECAPx1_ASAP7_75t_R FILLER_69_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_216 ();
 DECAPx1_ASAP7_75t_R FILLER_69_245 ();
 DECAPx10_ASAP7_75t_R FILLER_69_255 ();
 DECAPx1_ASAP7_75t_R FILLER_69_277 ();
 DECAPx2_ASAP7_75t_R FILLER_69_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_312 ();
 DECAPx2_ASAP7_75t_R FILLER_69_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_339 ();
 FILLER_ASAP7_75t_R FILLER_69_356 ();
 FILLER_ASAP7_75t_R FILLER_69_372 ();
 DECAPx4_ASAP7_75t_R FILLER_69_380 ();
 FILLER_ASAP7_75t_R FILLER_69_390 ();
 DECAPx4_ASAP7_75t_R FILLER_69_404 ();
 FILLER_ASAP7_75t_R FILLER_69_414 ();
 FILLER_ASAP7_75t_R FILLER_69_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_449 ();
 FILLER_ASAP7_75t_R FILLER_69_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_458 ();
 DECAPx2_ASAP7_75t_R FILLER_69_481 ();
 FILLER_ASAP7_75t_R FILLER_69_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_496 ();
 FILLER_ASAP7_75t_R FILLER_69_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_521 ();
 DECAPx2_ASAP7_75t_R FILLER_69_537 ();
 FILLER_ASAP7_75t_R FILLER_69_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_545 ();
 FILLER_ASAP7_75t_R FILLER_69_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_569 ();
 DECAPx10_ASAP7_75t_R FILLER_69_580 ();
 DECAPx6_ASAP7_75t_R FILLER_69_602 ();
 DECAPx2_ASAP7_75t_R FILLER_69_643 ();
 FILLER_ASAP7_75t_R FILLER_69_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_651 ();
 DECAPx10_ASAP7_75t_R FILLER_69_655 ();
 DECAPx10_ASAP7_75t_R FILLER_69_677 ();
 FILLER_ASAP7_75t_R FILLER_69_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_701 ();
 DECAPx4_ASAP7_75t_R FILLER_69_708 ();
 DECAPx10_ASAP7_75t_R FILLER_69_724 ();
 DECAPx2_ASAP7_75t_R FILLER_69_746 ();
 FILLER_ASAP7_75t_R FILLER_69_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_754 ();
 DECAPx1_ASAP7_75t_R FILLER_69_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_781 ();
 DECAPx10_ASAP7_75t_R FILLER_69_786 ();
 FILLER_ASAP7_75t_R FILLER_69_808 ();
 DECAPx2_ASAP7_75t_R FILLER_69_822 ();
 DECAPx4_ASAP7_75t_R FILLER_69_838 ();
 FILLER_ASAP7_75t_R FILLER_69_848 ();
 DECAPx6_ASAP7_75t_R FILLER_69_866 ();
 DECAPx10_ASAP7_75t_R FILLER_69_926 ();
 DECAPx1_ASAP7_75t_R FILLER_69_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_952 ();
 FILLER_ASAP7_75t_R FILLER_69_973 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1019 ();
 FILLER_ASAP7_75t_R FILLER_69_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1048 ();
 FILLER_ASAP7_75t_R FILLER_69_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1063 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1095 ();
 DECAPx6_ASAP7_75t_R FILLER_69_1107 ();
 FILLER_ASAP7_75t_R FILLER_69_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1123 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1141 ();
 FILLER_ASAP7_75t_R FILLER_69_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1153 ();
 FILLER_ASAP7_75t_R FILLER_69_1162 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1184 ();
 DECAPx1_ASAP7_75t_R FILLER_69_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1209 ();
 FILLER_ASAP7_75t_R FILLER_69_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_70_2 ();
 DECAPx10_ASAP7_75t_R FILLER_70_24 ();
 DECAPx10_ASAP7_75t_R FILLER_70_46 ();
 DECAPx6_ASAP7_75t_R FILLER_70_68 ();
 FILLER_ASAP7_75t_R FILLER_70_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_95 ();
 FILLER_ASAP7_75t_R FILLER_70_111 ();
 DECAPx10_ASAP7_75t_R FILLER_70_122 ();
 FILLER_ASAP7_75t_R FILLER_70_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_160 ();
 DECAPx10_ASAP7_75t_R FILLER_70_168 ();
 DECAPx4_ASAP7_75t_R FILLER_70_190 ();
 FILLER_ASAP7_75t_R FILLER_70_200 ();
 DECAPx4_ASAP7_75t_R FILLER_70_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_218 ();
 DECAPx2_ASAP7_75t_R FILLER_70_236 ();
 DECAPx6_ASAP7_75t_R FILLER_70_264 ();
 DECAPx1_ASAP7_75t_R FILLER_70_278 ();
 DECAPx1_ASAP7_75t_R FILLER_70_307 ();
 DECAPx4_ASAP7_75t_R FILLER_70_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_343 ();
 DECAPx10_ASAP7_75t_R FILLER_70_377 ();
 DECAPx2_ASAP7_75t_R FILLER_70_399 ();
 DECAPx4_ASAP7_75t_R FILLER_70_413 ();
 FILLER_ASAP7_75t_R FILLER_70_423 ();
 DECAPx1_ASAP7_75t_R FILLER_70_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_450 ();
 DECAPx10_ASAP7_75t_R FILLER_70_464 ();
 DECAPx2_ASAP7_75t_R FILLER_70_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_492 ();
 DECAPx4_ASAP7_75t_R FILLER_70_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_525 ();
 DECAPx6_ASAP7_75t_R FILLER_70_541 ();
 DECAPx1_ASAP7_75t_R FILLER_70_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_569 ();
 FILLER_ASAP7_75t_R FILLER_70_594 ();
 DECAPx2_ASAP7_75t_R FILLER_70_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_641 ();
 DECAPx10_ASAP7_75t_R FILLER_70_648 ();
 DECAPx10_ASAP7_75t_R FILLER_70_670 ();
 DECAPx1_ASAP7_75t_R FILLER_70_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_696 ();
 DECAPx10_ASAP7_75t_R FILLER_70_763 ();
 DECAPx2_ASAP7_75t_R FILLER_70_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_791 ();
 DECAPx2_ASAP7_75t_R FILLER_70_804 ();
 FILLER_ASAP7_75t_R FILLER_70_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_826 ();
 FILLER_ASAP7_75t_R FILLER_70_837 ();
 DECAPx2_ASAP7_75t_R FILLER_70_847 ();
 FILLER_ASAP7_75t_R FILLER_70_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_855 ();
 DECAPx10_ASAP7_75t_R FILLER_70_876 ();
 DECAPx6_ASAP7_75t_R FILLER_70_898 ();
 DECAPx2_ASAP7_75t_R FILLER_70_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_918 ();
 DECAPx10_ASAP7_75t_R FILLER_70_949 ();
 DECAPx10_ASAP7_75t_R FILLER_70_971 ();
 DECAPx10_ASAP7_75t_R FILLER_70_993 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1088 ();
 FILLER_ASAP7_75t_R FILLER_70_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1163 ();
 FILLER_ASAP7_75t_R FILLER_70_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1171 ();
 FILLER_ASAP7_75t_R FILLER_70_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_71_2 ();
 DECAPx10_ASAP7_75t_R FILLER_71_24 ();
 DECAPx10_ASAP7_75t_R FILLER_71_46 ();
 DECAPx1_ASAP7_75t_R FILLER_71_68 ();
 DECAPx1_ASAP7_75t_R FILLER_71_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_98 ();
 DECAPx1_ASAP7_75t_R FILLER_71_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_109 ();
 FILLER_ASAP7_75t_R FILLER_71_135 ();
 DECAPx2_ASAP7_75t_R FILLER_71_157 ();
 DECAPx6_ASAP7_75t_R FILLER_71_181 ();
 DECAPx1_ASAP7_75t_R FILLER_71_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_199 ();
 DECAPx2_ASAP7_75t_R FILLER_71_222 ();
 FILLER_ASAP7_75t_R FILLER_71_228 ();
 FILLER_ASAP7_75t_R FILLER_71_245 ();
 DECAPx10_ASAP7_75t_R FILLER_71_253 ();
 DECAPx1_ASAP7_75t_R FILLER_71_275 ();
 DECAPx1_ASAP7_75t_R FILLER_71_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_289 ();
 DECAPx10_ASAP7_75t_R FILLER_71_318 ();
 DECAPx10_ASAP7_75t_R FILLER_71_340 ();
 FILLER_ASAP7_75t_R FILLER_71_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_364 ();
 DECAPx6_ASAP7_75t_R FILLER_71_387 ();
 DECAPx2_ASAP7_75t_R FILLER_71_429 ();
 FILLER_ASAP7_75t_R FILLER_71_435 ();
 FILLER_ASAP7_75t_R FILLER_71_449 ();
 DECAPx10_ASAP7_75t_R FILLER_71_487 ();
 DECAPx1_ASAP7_75t_R FILLER_71_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_537 ();
 DECAPx6_ASAP7_75t_R FILLER_71_558 ();
 FILLER_ASAP7_75t_R FILLER_71_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_574 ();
 DECAPx2_ASAP7_75t_R FILLER_71_589 ();
 FILLER_ASAP7_75t_R FILLER_71_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_597 ();
 DECAPx10_ASAP7_75t_R FILLER_71_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_637 ();
 FILLER_ASAP7_75t_R FILLER_71_650 ();
 DECAPx2_ASAP7_75t_R FILLER_71_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_665 ();
 DECAPx2_ASAP7_75t_R FILLER_71_696 ();
 DECAPx1_ASAP7_75t_R FILLER_71_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_728 ();
 DECAPx4_ASAP7_75t_R FILLER_71_755 ();
 FILLER_ASAP7_75t_R FILLER_71_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_767 ();
 DECAPx6_ASAP7_75t_R FILLER_71_785 ();
 FILLER_ASAP7_75t_R FILLER_71_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_801 ();
 FILLER_ASAP7_75t_R FILLER_71_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_807 ();
 DECAPx6_ASAP7_75t_R FILLER_71_814 ();
 DECAPx2_ASAP7_75t_R FILLER_71_838 ();
 FILLER_ASAP7_75t_R FILLER_71_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_846 ();
 DECAPx2_ASAP7_75t_R FILLER_71_875 ();
 FILLER_ASAP7_75t_R FILLER_71_881 ();
 DECAPx4_ASAP7_75t_R FILLER_71_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_932 ();
 DECAPx2_ASAP7_75t_R FILLER_71_955 ();
 DECAPx10_ASAP7_75t_R FILLER_71_967 ();
 DECAPx6_ASAP7_75t_R FILLER_71_989 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1051 ();
 FILLER_ASAP7_75t_R FILLER_71_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_71_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1157 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_71_1215 ();
 FILLER_ASAP7_75t_R FILLER_71_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_72_2 ();
 DECAPx10_ASAP7_75t_R FILLER_72_24 ();
 DECAPx10_ASAP7_75t_R FILLER_72_46 ();
 DECAPx6_ASAP7_75t_R FILLER_72_68 ();
 DECAPx2_ASAP7_75t_R FILLER_72_82 ();
 DECAPx2_ASAP7_75t_R FILLER_72_94 ();
 DECAPx2_ASAP7_75t_R FILLER_72_106 ();
 FILLER_ASAP7_75t_R FILLER_72_112 ();
 DECAPx1_ASAP7_75t_R FILLER_72_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_125 ();
 DECAPx10_ASAP7_75t_R FILLER_72_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_176 ();
 DECAPx1_ASAP7_75t_R FILLER_72_190 ();
 DECAPx4_ASAP7_75t_R FILLER_72_205 ();
 DECAPx10_ASAP7_75t_R FILLER_72_241 ();
 DECAPx4_ASAP7_75t_R FILLER_72_263 ();
 DECAPx1_ASAP7_75t_R FILLER_72_295 ();
 DECAPx10_ASAP7_75t_R FILLER_72_308 ();
 DECAPx6_ASAP7_75t_R FILLER_72_330 ();
 FILLER_ASAP7_75t_R FILLER_72_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_346 ();
 DECAPx1_ASAP7_75t_R FILLER_72_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_373 ();
 DECAPx1_ASAP7_75t_R FILLER_72_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_398 ();
 FILLER_ASAP7_75t_R FILLER_72_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_410 ();
 DECAPx2_ASAP7_75t_R FILLER_72_418 ();
 FILLER_ASAP7_75t_R FILLER_72_424 ();
 DECAPx4_ASAP7_75t_R FILLER_72_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_464 ();
 DECAPx10_ASAP7_75t_R FILLER_72_487 ();
 DECAPx2_ASAP7_75t_R FILLER_72_509 ();
 FILLER_ASAP7_75t_R FILLER_72_515 ();
 DECAPx2_ASAP7_75t_R FILLER_72_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_555 ();
 DECAPx2_ASAP7_75t_R FILLER_72_563 ();
 FILLER_ASAP7_75t_R FILLER_72_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_571 ();
 DECAPx10_ASAP7_75t_R FILLER_72_578 ();
 DECAPx6_ASAP7_75t_R FILLER_72_600 ();
 FILLER_ASAP7_75t_R FILLER_72_626 ();
 DECAPx6_ASAP7_75t_R FILLER_72_640 ();
 FILLER_ASAP7_75t_R FILLER_72_682 ();
 DECAPx4_ASAP7_75t_R FILLER_72_694 ();
 FILLER_ASAP7_75t_R FILLER_72_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_706 ();
 DECAPx2_ASAP7_75t_R FILLER_72_713 ();
 DECAPx4_ASAP7_75t_R FILLER_72_752 ();
 FILLER_ASAP7_75t_R FILLER_72_762 ();
 FILLER_ASAP7_75t_R FILLER_72_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_776 ();
 DECAPx1_ASAP7_75t_R FILLER_72_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_791 ();
 FILLER_ASAP7_75t_R FILLER_72_804 ();
 DECAPx1_ASAP7_75t_R FILLER_72_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_816 ();
 DECAPx1_ASAP7_75t_R FILLER_72_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_827 ();
 DECAPx2_ASAP7_75t_R FILLER_72_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_852 ();
 DECAPx1_ASAP7_75t_R FILLER_72_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_865 ();
 DECAPx10_ASAP7_75t_R FILLER_72_872 ();
 DECAPx6_ASAP7_75t_R FILLER_72_894 ();
 DECAPx1_ASAP7_75t_R FILLER_72_908 ();
 DECAPx2_ASAP7_75t_R FILLER_72_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_934 ();
 DECAPx2_ASAP7_75t_R FILLER_72_951 ();
 DECAPx4_ASAP7_75t_R FILLER_72_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_989 ();
 DECAPx4_ASAP7_75t_R FILLER_72_1013 ();
 FILLER_ASAP7_75t_R FILLER_72_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1025 ();
 FILLER_ASAP7_75t_R FILLER_72_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1048 ();
 FILLER_ASAP7_75t_R FILLER_72_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_72_1146 ();
 FILLER_ASAP7_75t_R FILLER_72_1156 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1166 ();
 FILLER_ASAP7_75t_R FILLER_72_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_73_2 ();
 FILLER_ASAP7_75t_R FILLER_73_24 ();
 DECAPx10_ASAP7_75t_R FILLER_73_38 ();
 DECAPx10_ASAP7_75t_R FILLER_73_60 ();
 DECAPx2_ASAP7_75t_R FILLER_73_82 ();
 DECAPx10_ASAP7_75t_R FILLER_73_105 ();
 DECAPx10_ASAP7_75t_R FILLER_73_127 ();
 DECAPx6_ASAP7_75t_R FILLER_73_149 ();
 DECAPx1_ASAP7_75t_R FILLER_73_163 ();
 DECAPx4_ASAP7_75t_R FILLER_73_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_205 ();
 DECAPx10_ASAP7_75t_R FILLER_73_217 ();
 DECAPx10_ASAP7_75t_R FILLER_73_239 ();
 DECAPx10_ASAP7_75t_R FILLER_73_261 ();
 DECAPx1_ASAP7_75t_R FILLER_73_283 ();
 DECAPx1_ASAP7_75t_R FILLER_73_305 ();
 DECAPx6_ASAP7_75t_R FILLER_73_337 ();
 FILLER_ASAP7_75t_R FILLER_73_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_359 ();
 DECAPx2_ASAP7_75t_R FILLER_73_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_390 ();
 DECAPx10_ASAP7_75t_R FILLER_73_409 ();
 DECAPx1_ASAP7_75t_R FILLER_73_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_435 ();
 FILLER_ASAP7_75t_R FILLER_73_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_456 ();
 DECAPx4_ASAP7_75t_R FILLER_73_507 ();
 FILLER_ASAP7_75t_R FILLER_73_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_523 ();
 DECAPx2_ASAP7_75t_R FILLER_73_541 ();
 FILLER_ASAP7_75t_R FILLER_73_547 ();
 DECAPx2_ASAP7_75t_R FILLER_73_564 ();
 DECAPx10_ASAP7_75t_R FILLER_73_581 ();
 DECAPx6_ASAP7_75t_R FILLER_73_603 ();
 DECAPx4_ASAP7_75t_R FILLER_73_625 ();
 FILLER_ASAP7_75t_R FILLER_73_635 ();
 DECAPx2_ASAP7_75t_R FILLER_73_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_651 ();
 DECAPx2_ASAP7_75t_R FILLER_73_658 ();
 FILLER_ASAP7_75t_R FILLER_73_664 ();
 DECAPx10_ASAP7_75t_R FILLER_73_686 ();
 DECAPx1_ASAP7_75t_R FILLER_73_708 ();
 DECAPx1_ASAP7_75t_R FILLER_73_760 ();
 FILLER_ASAP7_75t_R FILLER_73_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_781 ();
 DECAPx1_ASAP7_75t_R FILLER_73_792 ();
 FILLER_ASAP7_75t_R FILLER_73_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_801 ();
 DECAPx1_ASAP7_75t_R FILLER_73_816 ();
 DECAPx6_ASAP7_75t_R FILLER_73_826 ();
 FILLER_ASAP7_75t_R FILLER_73_840 ();
 DECAPx6_ASAP7_75t_R FILLER_73_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_886 ();
 DECAPx10_ASAP7_75t_R FILLER_73_895 ();
 DECAPx2_ASAP7_75t_R FILLER_73_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_923 ();
 DECAPx2_ASAP7_75t_R FILLER_73_926 ();
 FILLER_ASAP7_75t_R FILLER_73_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_934 ();
 DECAPx2_ASAP7_75t_R FILLER_73_963 ();
 FILLER_ASAP7_75t_R FILLER_73_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_971 ();
 DECAPx10_ASAP7_75t_R FILLER_73_994 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1022 ();
 DECAPx1_ASAP7_75t_R FILLER_73_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_73_1120 ();
 FILLER_ASAP7_75t_R FILLER_73_1134 ();
 FILLER_ASAP7_75t_R FILLER_73_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1168 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1186 ();
 FILLER_ASAP7_75t_R FILLER_73_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1209 ();
 DECAPx6_ASAP7_75t_R FILLER_74_8 ();
 FILLER_ASAP7_75t_R FILLER_74_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_24 ();
 DECAPx10_ASAP7_75t_R FILLER_74_31 ();
 DECAPx10_ASAP7_75t_R FILLER_74_53 ();
 DECAPx2_ASAP7_75t_R FILLER_74_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_104 ();
 DECAPx1_ASAP7_75t_R FILLER_74_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_131 ();
 DECAPx4_ASAP7_75t_R FILLER_74_164 ();
 FILLER_ASAP7_75t_R FILLER_74_192 ();
 DECAPx10_ASAP7_75t_R FILLER_74_218 ();
 DECAPx10_ASAP7_75t_R FILLER_74_240 ();
 DECAPx10_ASAP7_75t_R FILLER_74_262 ();
 DECAPx10_ASAP7_75t_R FILLER_74_304 ();
 DECAPx10_ASAP7_75t_R FILLER_74_326 ();
 DECAPx6_ASAP7_75t_R FILLER_74_348 ();
 DECAPx2_ASAP7_75t_R FILLER_74_362 ();
 DECAPx2_ASAP7_75t_R FILLER_74_372 ();
 FILLER_ASAP7_75t_R FILLER_74_378 ();
 DECAPx1_ASAP7_75t_R FILLER_74_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_388 ();
 FILLER_ASAP7_75t_R FILLER_74_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_402 ();
 DECAPx10_ASAP7_75t_R FILLER_74_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_431 ();
 DECAPx2_ASAP7_75t_R FILLER_74_454 ();
 FILLER_ASAP7_75t_R FILLER_74_460 ();
 FILLER_ASAP7_75t_R FILLER_74_475 ();
 DECAPx4_ASAP7_75t_R FILLER_74_495 ();
 FILLER_ASAP7_75t_R FILLER_74_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_507 ();
 FILLER_ASAP7_75t_R FILLER_74_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_542 ();
 DECAPx1_ASAP7_75t_R FILLER_74_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_557 ();
 DECAPx1_ASAP7_75t_R FILLER_74_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_568 ();
 FILLER_ASAP7_75t_R FILLER_74_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_589 ();
 DECAPx6_ASAP7_75t_R FILLER_74_600 ();
 FILLER_ASAP7_75t_R FILLER_74_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_645 ();
 FILLER_ASAP7_75t_R FILLER_74_658 ();
 DECAPx10_ASAP7_75t_R FILLER_74_688 ();
 DECAPx4_ASAP7_75t_R FILLER_74_710 ();
 FILLER_ASAP7_75t_R FILLER_74_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_722 ();
 DECAPx10_ASAP7_75t_R FILLER_74_747 ();
 DECAPx1_ASAP7_75t_R FILLER_74_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_773 ();
 DECAPx2_ASAP7_75t_R FILLER_74_787 ();
 FILLER_ASAP7_75t_R FILLER_74_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_795 ();
 FILLER_ASAP7_75t_R FILLER_74_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_812 ();
 FILLER_ASAP7_75t_R FILLER_74_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_837 ();
 DECAPx2_ASAP7_75t_R FILLER_74_863 ();
 FILLER_ASAP7_75t_R FILLER_74_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_871 ();
 DECAPx4_ASAP7_75t_R FILLER_74_892 ();
 FILLER_ASAP7_75t_R FILLER_74_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_904 ();
 DECAPx4_ASAP7_75t_R FILLER_74_931 ();
 DECAPx10_ASAP7_75t_R FILLER_74_985 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1028 ();
 FILLER_ASAP7_75t_R FILLER_74_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1059 ();
 FILLER_ASAP7_75t_R FILLER_74_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1110 ();
 FILLER_ASAP7_75t_R FILLER_74_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1169 ();
 FILLER_ASAP7_75t_R FILLER_74_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1181 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1204 ();
 FILLER_ASAP7_75t_R FILLER_74_1214 ();
 FILLER_ASAP7_75t_R FILLER_74_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_75_2 ();
 DECAPx10_ASAP7_75t_R FILLER_75_24 ();
 DECAPx10_ASAP7_75t_R FILLER_75_46 ();
 DECAPx10_ASAP7_75t_R FILLER_75_68 ();
 DECAPx6_ASAP7_75t_R FILLER_75_90 ();
 FILLER_ASAP7_75t_R FILLER_75_104 ();
 DECAPx6_ASAP7_75t_R FILLER_75_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_132 ();
 FILLER_ASAP7_75t_R FILLER_75_155 ();
 DECAPx6_ASAP7_75t_R FILLER_75_176 ();
 FILLER_ASAP7_75t_R FILLER_75_190 ();
 DECAPx6_ASAP7_75t_R FILLER_75_234 ();
 DECAPx1_ASAP7_75t_R FILLER_75_248 ();
 DECAPx4_ASAP7_75t_R FILLER_75_270 ();
 FILLER_ASAP7_75t_R FILLER_75_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_301 ();
 DECAPx10_ASAP7_75t_R FILLER_75_326 ();
 DECAPx10_ASAP7_75t_R FILLER_75_348 ();
 DECAPx10_ASAP7_75t_R FILLER_75_370 ();
 DECAPx1_ASAP7_75t_R FILLER_75_392 ();
 DECAPx6_ASAP7_75t_R FILLER_75_421 ();
 FILLER_ASAP7_75t_R FILLER_75_435 ();
 DECAPx10_ASAP7_75t_R FILLER_75_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_477 ();
 FILLER_ASAP7_75t_R FILLER_75_490 ();
 DECAPx1_ASAP7_75t_R FILLER_75_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_557 ();
 FILLER_ASAP7_75t_R FILLER_75_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_567 ();
 DECAPx2_ASAP7_75t_R FILLER_75_588 ();
 FILLER_ASAP7_75t_R FILLER_75_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_602 ();
 DECAPx2_ASAP7_75t_R FILLER_75_611 ();
 DECAPx1_ASAP7_75t_R FILLER_75_623 ();
 DECAPx2_ASAP7_75t_R FILLER_75_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_639 ();
 DECAPx10_ASAP7_75t_R FILLER_75_684 ();
 DECAPx6_ASAP7_75t_R FILLER_75_706 ();
 FILLER_ASAP7_75t_R FILLER_75_720 ();
 DECAPx2_ASAP7_75t_R FILLER_75_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_746 ();
 DECAPx1_ASAP7_75t_R FILLER_75_753 ();
 DECAPx2_ASAP7_75t_R FILLER_75_763 ();
 FILLER_ASAP7_75t_R FILLER_75_769 ();
 DECAPx2_ASAP7_75t_R FILLER_75_781 ();
 FILLER_ASAP7_75t_R FILLER_75_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_801 ();
 DECAPx2_ASAP7_75t_R FILLER_75_812 ();
 FILLER_ASAP7_75t_R FILLER_75_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_820 ();
 DECAPx2_ASAP7_75t_R FILLER_75_824 ();
 DECAPx1_ASAP7_75t_R FILLER_75_837 ();
 DECAPx1_ASAP7_75t_R FILLER_75_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_856 ();
 DECAPx2_ASAP7_75t_R FILLER_75_875 ();
 FILLER_ASAP7_75t_R FILLER_75_881 ();
 DECAPx6_ASAP7_75t_R FILLER_75_905 ();
 DECAPx1_ASAP7_75t_R FILLER_75_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_923 ();
 DECAPx10_ASAP7_75t_R FILLER_75_948 ();
 DECAPx2_ASAP7_75t_R FILLER_75_970 ();
 FILLER_ASAP7_75t_R FILLER_75_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_978 ();
 DECAPx6_ASAP7_75t_R FILLER_75_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1015 ();
 FILLER_ASAP7_75t_R FILLER_75_1041 ();
 DECAPx4_ASAP7_75t_R FILLER_75_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_75_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1163 ();
 DECAPx4_ASAP7_75t_R FILLER_75_1181 ();
 FILLER_ASAP7_75t_R FILLER_75_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1220 ();
 DECAPx6_ASAP7_75t_R FILLER_76_2 ();
 FILLER_ASAP7_75t_R FILLER_76_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_18 ();
 DECAPx10_ASAP7_75t_R FILLER_76_25 ();
 DECAPx10_ASAP7_75t_R FILLER_76_47 ();
 DECAPx10_ASAP7_75t_R FILLER_76_69 ();
 DECAPx6_ASAP7_75t_R FILLER_76_91 ();
 DECAPx2_ASAP7_75t_R FILLER_76_105 ();
 FILLER_ASAP7_75t_R FILLER_76_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_132 ();
 DECAPx2_ASAP7_75t_R FILLER_76_139 ();
 FILLER_ASAP7_75t_R FILLER_76_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_147 ();
 DECAPx6_ASAP7_75t_R FILLER_76_175 ();
 DECAPx1_ASAP7_75t_R FILLER_76_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_193 ();
 DECAPx10_ASAP7_75t_R FILLER_76_200 ();
 DECAPx10_ASAP7_75t_R FILLER_76_222 ();
 DECAPx10_ASAP7_75t_R FILLER_76_244 ();
 DECAPx6_ASAP7_75t_R FILLER_76_266 ();
 FILLER_ASAP7_75t_R FILLER_76_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_282 ();
 DECAPx1_ASAP7_75t_R FILLER_76_305 ();
 DECAPx6_ASAP7_75t_R FILLER_76_312 ();
 FILLER_ASAP7_75t_R FILLER_76_326 ();
 DECAPx6_ASAP7_75t_R FILLER_76_368 ();
 DECAPx2_ASAP7_75t_R FILLER_76_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_408 ();
 DECAPx2_ASAP7_75t_R FILLER_76_431 ();
 FILLER_ASAP7_75t_R FILLER_76_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_439 ();
 DECAPx2_ASAP7_75t_R FILLER_76_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_470 ();
 DECAPx1_ASAP7_75t_R FILLER_76_478 ();
 DECAPx1_ASAP7_75t_R FILLER_76_488 ();
 DECAPx6_ASAP7_75t_R FILLER_76_498 ();
 FILLER_ASAP7_75t_R FILLER_76_512 ();
 DECAPx2_ASAP7_75t_R FILLER_76_517 ();
 FILLER_ASAP7_75t_R FILLER_76_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_559 ();
 DECAPx1_ASAP7_75t_R FILLER_76_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_579 ();
 DECAPx2_ASAP7_75t_R FILLER_76_606 ();
 DECAPx2_ASAP7_75t_R FILLER_76_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_648 ();
 DECAPx10_ASAP7_75t_R FILLER_76_655 ();
 DECAPx10_ASAP7_75t_R FILLER_76_677 ();
 DECAPx6_ASAP7_75t_R FILLER_76_699 ();
 FILLER_ASAP7_75t_R FILLER_76_713 ();
 DECAPx6_ASAP7_75t_R FILLER_76_733 ();
 DECAPx1_ASAP7_75t_R FILLER_76_747 ();
 DECAPx2_ASAP7_75t_R FILLER_76_763 ();
 DECAPx2_ASAP7_75t_R FILLER_76_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_784 ();
 DECAPx1_ASAP7_75t_R FILLER_76_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_796 ();
 DECAPx4_ASAP7_75t_R FILLER_76_800 ();
 FILLER_ASAP7_75t_R FILLER_76_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_812 ();
 DECAPx2_ASAP7_75t_R FILLER_76_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_828 ();
 DECAPx10_ASAP7_75t_R FILLER_76_857 ();
 DECAPx10_ASAP7_75t_R FILLER_76_879 ();
 DECAPx1_ASAP7_75t_R FILLER_76_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_905 ();
 FILLER_ASAP7_75t_R FILLER_76_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_914 ();
 FILLER_ASAP7_75t_R FILLER_76_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_937 ();
 DECAPx2_ASAP7_75t_R FILLER_76_946 ();
 DECAPx2_ASAP7_75t_R FILLER_76_958 ();
 FILLER_ASAP7_75t_R FILLER_76_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_966 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1001 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1043 ();
 FILLER_ASAP7_75t_R FILLER_76_1052 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1153 ();
 DECAPx4_ASAP7_75t_R FILLER_76_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1197 ();
 FILLER_ASAP7_75t_R FILLER_76_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1205 ();
 DECAPx6_ASAP7_75t_R FILLER_77_2 ();
 DECAPx10_ASAP7_75t_R FILLER_77_22 ();
 DECAPx10_ASAP7_75t_R FILLER_77_44 ();
 DECAPx10_ASAP7_75t_R FILLER_77_66 ();
 DECAPx4_ASAP7_75t_R FILLER_77_88 ();
 FILLER_ASAP7_75t_R FILLER_77_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_100 ();
 FILLER_ASAP7_75t_R FILLER_77_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_114 ();
 DECAPx2_ASAP7_75t_R FILLER_77_123 ();
 FILLER_ASAP7_75t_R FILLER_77_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_131 ();
 DECAPx10_ASAP7_75t_R FILLER_77_140 ();
 DECAPx1_ASAP7_75t_R FILLER_77_162 ();
 DECAPx10_ASAP7_75t_R FILLER_77_194 ();
 DECAPx10_ASAP7_75t_R FILLER_77_216 ();
 DECAPx2_ASAP7_75t_R FILLER_77_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_264 ();
 DECAPx6_ASAP7_75t_R FILLER_77_271 ();
 DECAPx1_ASAP7_75t_R FILLER_77_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_315 ();
 DECAPx4_ASAP7_75t_R FILLER_77_320 ();
 FILLER_ASAP7_75t_R FILLER_77_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_336 ();
 DECAPx6_ASAP7_75t_R FILLER_77_357 ();
 DECAPx1_ASAP7_75t_R FILLER_77_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_375 ();
 DECAPx2_ASAP7_75t_R FILLER_77_416 ();
 FILLER_ASAP7_75t_R FILLER_77_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_430 ();
 DECAPx2_ASAP7_75t_R FILLER_77_450 ();
 FILLER_ASAP7_75t_R FILLER_77_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_484 ();
 DECAPx1_ASAP7_75t_R FILLER_77_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_500 ();
 DECAPx10_ASAP7_75t_R FILLER_77_523 ();
 FILLER_ASAP7_75t_R FILLER_77_545 ();
 FILLER_ASAP7_75t_R FILLER_77_561 ();
 DECAPx6_ASAP7_75t_R FILLER_77_576 ();
 DECAPx2_ASAP7_75t_R FILLER_77_590 ();
 DECAPx10_ASAP7_75t_R FILLER_77_604 ();
 DECAPx2_ASAP7_75t_R FILLER_77_626 ();
 FILLER_ASAP7_75t_R FILLER_77_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_634 ();
 DECAPx6_ASAP7_75t_R FILLER_77_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_655 ();
 DECAPx1_ASAP7_75t_R FILLER_77_670 ();
 DECAPx10_ASAP7_75t_R FILLER_77_694 ();
 DECAPx6_ASAP7_75t_R FILLER_77_734 ();
 FILLER_ASAP7_75t_R FILLER_77_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_750 ();
 FILLER_ASAP7_75t_R FILLER_77_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_784 ();
 DECAPx2_ASAP7_75t_R FILLER_77_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_825 ();
 DECAPx10_ASAP7_75t_R FILLER_77_844 ();
 DECAPx10_ASAP7_75t_R FILLER_77_866 ();
 DECAPx4_ASAP7_75t_R FILLER_77_888 ();
 FILLER_ASAP7_75t_R FILLER_77_898 ();
 DECAPx2_ASAP7_75t_R FILLER_77_918 ();
 DECAPx2_ASAP7_75t_R FILLER_77_939 ();
 FILLER_ASAP7_75t_R FILLER_77_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_954 ();
 DECAPx4_ASAP7_75t_R FILLER_77_961 ();
 DECAPx2_ASAP7_75t_R FILLER_77_974 ();
 FILLER_ASAP7_75t_R FILLER_77_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_982 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_77_1129 ();
 FILLER_ASAP7_75t_R FILLER_77_1139 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1180 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1202 ();
 FILLER_ASAP7_75t_R FILLER_77_1216 ();
 FILLER_ASAP7_75t_R FILLER_78_2 ();
 DECAPx10_ASAP7_75t_R FILLER_78_10 ();
 DECAPx10_ASAP7_75t_R FILLER_78_32 ();
 DECAPx10_ASAP7_75t_R FILLER_78_54 ();
 DECAPx2_ASAP7_75t_R FILLER_78_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_82 ();
 DECAPx10_ASAP7_75t_R FILLER_78_124 ();
 DECAPx1_ASAP7_75t_R FILLER_78_146 ();
 DECAPx4_ASAP7_75t_R FILLER_78_160 ();
 DECAPx2_ASAP7_75t_R FILLER_78_178 ();
 FILLER_ASAP7_75t_R FILLER_78_184 ();
 DECAPx10_ASAP7_75t_R FILLER_78_214 ();
 DECAPx1_ASAP7_75t_R FILLER_78_236 ();
 DECAPx2_ASAP7_75t_R FILLER_78_266 ();
 DECAPx4_ASAP7_75t_R FILLER_78_294 ();
 FILLER_ASAP7_75t_R FILLER_78_304 ();
 DECAPx2_ASAP7_75t_R FILLER_78_326 ();
 DECAPx4_ASAP7_75t_R FILLER_78_335 ();
 DECAPx10_ASAP7_75t_R FILLER_78_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_393 ();
 DECAPx6_ASAP7_75t_R FILLER_78_405 ();
 DECAPx2_ASAP7_75t_R FILLER_78_453 ();
 FILLER_ASAP7_75t_R FILLER_78_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_461 ();
 DECAPx1_ASAP7_75t_R FILLER_78_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_490 ();
 DECAPx2_ASAP7_75t_R FILLER_78_497 ();
 DECAPx10_ASAP7_75t_R FILLER_78_509 ();
 DECAPx6_ASAP7_75t_R FILLER_78_531 ();
 FILLER_ASAP7_75t_R FILLER_78_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_553 ();
 DECAPx6_ASAP7_75t_R FILLER_78_576 ();
 FILLER_ASAP7_75t_R FILLER_78_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_592 ();
 FILLER_ASAP7_75t_R FILLER_78_599 ();
 DECAPx2_ASAP7_75t_R FILLER_78_623 ();
 FILLER_ASAP7_75t_R FILLER_78_629 ();
 FILLER_ASAP7_75t_R FILLER_78_653 ();
 DECAPx10_ASAP7_75t_R FILLER_78_711 ();
 FILLER_ASAP7_75t_R FILLER_78_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_768 ();
 DECAPx1_ASAP7_75t_R FILLER_78_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_779 ();
 DECAPx1_ASAP7_75t_R FILLER_78_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_798 ();
 DECAPx2_ASAP7_75t_R FILLER_78_830 ();
 FILLER_ASAP7_75t_R FILLER_78_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_838 ();
 DECAPx10_ASAP7_75t_R FILLER_78_843 ();
 DECAPx1_ASAP7_75t_R FILLER_78_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_893 ();
 FILLER_ASAP7_75t_R FILLER_78_900 ();
 DECAPx1_ASAP7_75t_R FILLER_78_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_912 ();
 DECAPx2_ASAP7_75t_R FILLER_78_923 ();
 FILLER_ASAP7_75t_R FILLER_78_939 ();
 FILLER_ASAP7_75t_R FILLER_78_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_957 ();
 DECAPx2_ASAP7_75t_R FILLER_78_979 ();
 DECAPx4_ASAP7_75t_R FILLER_78_1013 ();
 FILLER_ASAP7_75t_R FILLER_78_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_78_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1117 ();
 FILLER_ASAP7_75t_R FILLER_78_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_78_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1169 ();
 FILLER_ASAP7_75t_R FILLER_78_1176 ();
 FILLER_ASAP7_75t_R FILLER_78_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_79_2 ();
 DECAPx10_ASAP7_75t_R FILLER_79_24 ();
 DECAPx10_ASAP7_75t_R FILLER_79_46 ();
 DECAPx10_ASAP7_75t_R FILLER_79_68 ();
 DECAPx6_ASAP7_75t_R FILLER_79_90 ();
 DECAPx2_ASAP7_75t_R FILLER_79_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_110 ();
 DECAPx2_ASAP7_75t_R FILLER_79_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_123 ();
 FILLER_ASAP7_75t_R FILLER_79_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_132 ();
 DECAPx6_ASAP7_75t_R FILLER_79_148 ();
 FILLER_ASAP7_75t_R FILLER_79_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_164 ();
 DECAPx10_ASAP7_75t_R FILLER_79_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_203 ();
 DECAPx10_ASAP7_75t_R FILLER_79_234 ();
 DECAPx6_ASAP7_75t_R FILLER_79_256 ();
 FILLER_ASAP7_75t_R FILLER_79_270 ();
 DECAPx6_ASAP7_75t_R FILLER_79_278 ();
 DECAPx2_ASAP7_75t_R FILLER_79_292 ();
 DECAPx1_ASAP7_75t_R FILLER_79_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_305 ();
 DECAPx6_ASAP7_75t_R FILLER_79_318 ();
 DECAPx1_ASAP7_75t_R FILLER_79_332 ();
 DECAPx2_ASAP7_75t_R FILLER_79_343 ();
 FILLER_ASAP7_75t_R FILLER_79_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_390 ();
 DECAPx6_ASAP7_75t_R FILLER_79_417 ();
 FILLER_ASAP7_75t_R FILLER_79_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_433 ();
 FILLER_ASAP7_75t_R FILLER_79_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_453 ();
 DECAPx10_ASAP7_75t_R FILLER_79_461 ();
 DECAPx2_ASAP7_75t_R FILLER_79_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_489 ();
 DECAPx10_ASAP7_75t_R FILLER_79_510 ();
 DECAPx6_ASAP7_75t_R FILLER_79_532 ();
 DECAPx2_ASAP7_75t_R FILLER_79_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_559 ();
 DECAPx1_ASAP7_75t_R FILLER_79_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_569 ();
 DECAPx1_ASAP7_75t_R FILLER_79_590 ();
 DECAPx10_ASAP7_75t_R FILLER_79_602 ();
 DECAPx4_ASAP7_75t_R FILLER_79_624 ();
 DECAPx10_ASAP7_75t_R FILLER_79_656 ();
 DECAPx10_ASAP7_75t_R FILLER_79_678 ();
 DECAPx6_ASAP7_75t_R FILLER_79_700 ();
 DECAPx2_ASAP7_75t_R FILLER_79_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_720 ();
 DECAPx2_ASAP7_75t_R FILLER_79_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_749 ();
 FILLER_ASAP7_75t_R FILLER_79_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_758 ();
 DECAPx10_ASAP7_75t_R FILLER_79_762 ();
 DECAPx4_ASAP7_75t_R FILLER_79_784 ();
 FILLER_ASAP7_75t_R FILLER_79_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_796 ();
 DECAPx2_ASAP7_75t_R FILLER_79_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_817 ();
 FILLER_ASAP7_75t_R FILLER_79_826 ();
 DECAPx4_ASAP7_75t_R FILLER_79_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_858 ();
 DECAPx4_ASAP7_75t_R FILLER_79_877 ();
 FILLER_ASAP7_75t_R FILLER_79_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_923 ();
 DECAPx6_ASAP7_75t_R FILLER_79_926 ();
 FILLER_ASAP7_75t_R FILLER_79_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_942 ();
 FILLER_ASAP7_75t_R FILLER_79_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_966 ();
 DECAPx2_ASAP7_75t_R FILLER_79_980 ();
 FILLER_ASAP7_75t_R FILLER_79_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_988 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1011 ();
 DECAPx6_ASAP7_75t_R FILLER_79_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1073 ();
 DECAPx6_ASAP7_75t_R FILLER_79_1105 ();
 FILLER_ASAP7_75t_R FILLER_79_1119 ();
 FILLER_ASAP7_75t_R FILLER_79_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1162 ();
 FILLER_ASAP7_75t_R FILLER_79_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1170 ();
 FILLER_ASAP7_75t_R FILLER_79_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_80_8 ();
 DECAPx10_ASAP7_75t_R FILLER_80_30 ();
 DECAPx10_ASAP7_75t_R FILLER_80_52 ();
 DECAPx10_ASAP7_75t_R FILLER_80_74 ();
 DECAPx4_ASAP7_75t_R FILLER_80_96 ();
 FILLER_ASAP7_75t_R FILLER_80_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_143 ();
 DECAPx2_ASAP7_75t_R FILLER_80_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_175 ();
 FILLER_ASAP7_75t_R FILLER_80_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_186 ();
 DECAPx1_ASAP7_75t_R FILLER_80_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_197 ();
 DECAPx10_ASAP7_75t_R FILLER_80_215 ();
 DECAPx6_ASAP7_75t_R FILLER_80_237 ();
 FILLER_ASAP7_75t_R FILLER_80_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_332 ();
 DECAPx2_ASAP7_75t_R FILLER_80_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_354 ();
 DECAPx6_ASAP7_75t_R FILLER_80_387 ();
 FILLER_ASAP7_75t_R FILLER_80_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_448 ();
 DECAPx10_ASAP7_75t_R FILLER_80_464 ();
 DECAPx4_ASAP7_75t_R FILLER_80_497 ();
 DECAPx10_ASAP7_75t_R FILLER_80_513 ();
 FILLER_ASAP7_75t_R FILLER_80_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_591 ();
 DECAPx1_ASAP7_75t_R FILLER_80_614 ();
 DECAPx4_ASAP7_75t_R FILLER_80_650 ();
 FILLER_ASAP7_75t_R FILLER_80_660 ();
 DECAPx10_ASAP7_75t_R FILLER_80_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_747 ();
 DECAPx4_ASAP7_75t_R FILLER_80_774 ();
 DECAPx4_ASAP7_75t_R FILLER_80_794 ();
 FILLER_ASAP7_75t_R FILLER_80_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_806 ();
 FILLER_ASAP7_75t_R FILLER_80_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_839 ();
 DECAPx4_ASAP7_75t_R FILLER_80_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_902 ();
 DECAPx2_ASAP7_75t_R FILLER_80_943 ();
 FILLER_ASAP7_75t_R FILLER_80_949 ();
 DECAPx2_ASAP7_75t_R FILLER_80_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_963 ();
 DECAPx6_ASAP7_75t_R FILLER_80_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_981 ();
 DECAPx4_ASAP7_75t_R FILLER_80_1004 ();
 FILLER_ASAP7_75t_R FILLER_80_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1038 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1060 ();
 FILLER_ASAP7_75t_R FILLER_80_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1080 ();
 DECAPx4_ASAP7_75t_R FILLER_80_1102 ();
 FILLER_ASAP7_75t_R FILLER_80_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1114 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_80_1184 ();
 FILLER_ASAP7_75t_R FILLER_80_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1213 ();
 DECAPx6_ASAP7_75t_R FILLER_81_2 ();
 FILLER_ASAP7_75t_R FILLER_81_16 ();
 DECAPx10_ASAP7_75t_R FILLER_81_24 ();
 DECAPx10_ASAP7_75t_R FILLER_81_46 ();
 DECAPx10_ASAP7_75t_R FILLER_81_68 ();
 DECAPx2_ASAP7_75t_R FILLER_81_90 ();
 DECAPx4_ASAP7_75t_R FILLER_81_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_134 ();
 FILLER_ASAP7_75t_R FILLER_81_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_185 ();
 DECAPx10_ASAP7_75t_R FILLER_81_197 ();
 DECAPx10_ASAP7_75t_R FILLER_81_219 ();
 DECAPx10_ASAP7_75t_R FILLER_81_241 ();
 DECAPx10_ASAP7_75t_R FILLER_81_263 ();
 DECAPx4_ASAP7_75t_R FILLER_81_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_295 ();
 DECAPx6_ASAP7_75t_R FILLER_81_302 ();
 FILLER_ASAP7_75t_R FILLER_81_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_318 ();
 DECAPx2_ASAP7_75t_R FILLER_81_325 ();
 DECAPx6_ASAP7_75t_R FILLER_81_338 ();
 FILLER_ASAP7_75t_R FILLER_81_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_354 ();
 DECAPx10_ASAP7_75t_R FILLER_81_361 ();
 DECAPx6_ASAP7_75t_R FILLER_81_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_397 ();
 FILLER_ASAP7_75t_R FILLER_81_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_416 ();
 DECAPx6_ASAP7_75t_R FILLER_81_428 ();
 DECAPx1_ASAP7_75t_R FILLER_81_442 ();
 DECAPx4_ASAP7_75t_R FILLER_81_468 ();
 FILLER_ASAP7_75t_R FILLER_81_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_480 ();
 DECAPx2_ASAP7_75t_R FILLER_81_487 ();
 FILLER_ASAP7_75t_R FILLER_81_493 ();
 DECAPx2_ASAP7_75t_R FILLER_81_513 ();
 FILLER_ASAP7_75t_R FILLER_81_519 ();
 DECAPx10_ASAP7_75t_R FILLER_81_543 ();
 DECAPx2_ASAP7_75t_R FILLER_81_565 ();
 FILLER_ASAP7_75t_R FILLER_81_571 ();
 FILLER_ASAP7_75t_R FILLER_81_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_639 ();
 DECAPx4_ASAP7_75t_R FILLER_81_648 ();
 FILLER_ASAP7_75t_R FILLER_81_658 ();
 DECAPx2_ASAP7_75t_R FILLER_81_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_675 ();
 DECAPx10_ASAP7_75t_R FILLER_81_690 ();
 DECAPx6_ASAP7_75t_R FILLER_81_712 ();
 FILLER_ASAP7_75t_R FILLER_81_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_728 ();
 DECAPx4_ASAP7_75t_R FILLER_81_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_761 ();
 FILLER_ASAP7_75t_R FILLER_81_770 ();
 FILLER_ASAP7_75t_R FILLER_81_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_831 ();
 FILLER_ASAP7_75t_R FILLER_81_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_840 ();
 DECAPx10_ASAP7_75t_R FILLER_81_863 ();
 DECAPx4_ASAP7_75t_R FILLER_81_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_901 ();
 DECAPx1_ASAP7_75t_R FILLER_81_908 ();
 DECAPx2_ASAP7_75t_R FILLER_81_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_932 ();
 DECAPx1_ASAP7_75t_R FILLER_81_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_947 ();
 DECAPx1_ASAP7_75t_R FILLER_81_954 ();
 FILLER_ASAP7_75t_R FILLER_81_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_975 ();
 DECAPx6_ASAP7_75t_R FILLER_81_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1050 ();
 DECAPx6_ASAP7_75t_R FILLER_81_1057 ();
 FILLER_ASAP7_75t_R FILLER_81_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_81_1116 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1130 ();
 DECAPx6_ASAP7_75t_R FILLER_81_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1161 ();
 FILLER_ASAP7_75t_R FILLER_81_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_82_2 ();
 DECAPx10_ASAP7_75t_R FILLER_82_24 ();
 DECAPx10_ASAP7_75t_R FILLER_82_46 ();
 DECAPx10_ASAP7_75t_R FILLER_82_68 ();
 DECAPx4_ASAP7_75t_R FILLER_82_90 ();
 FILLER_ASAP7_75t_R FILLER_82_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_102 ();
 DECAPx6_ASAP7_75t_R FILLER_82_120 ();
 DECAPx2_ASAP7_75t_R FILLER_82_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_140 ();
 FILLER_ASAP7_75t_R FILLER_82_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_150 ();
 DECAPx6_ASAP7_75t_R FILLER_82_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_173 ();
 DECAPx2_ASAP7_75t_R FILLER_82_180 ();
 FILLER_ASAP7_75t_R FILLER_82_186 ();
 DECAPx10_ASAP7_75t_R FILLER_82_194 ();
 DECAPx10_ASAP7_75t_R FILLER_82_216 ();
 DECAPx10_ASAP7_75t_R FILLER_82_238 ();
 DECAPx6_ASAP7_75t_R FILLER_82_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_274 ();
 FILLER_ASAP7_75t_R FILLER_82_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_299 ();
 DECAPx4_ASAP7_75t_R FILLER_82_332 ();
 FILLER_ASAP7_75t_R FILLER_82_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_350 ();
 DECAPx10_ASAP7_75t_R FILLER_82_365 ();
 DECAPx6_ASAP7_75t_R FILLER_82_387 ();
 DECAPx1_ASAP7_75t_R FILLER_82_401 ();
 DECAPx10_ASAP7_75t_R FILLER_82_427 ();
 FILLER_ASAP7_75t_R FILLER_82_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_451 ();
 DECAPx1_ASAP7_75t_R FILLER_82_458 ();
 DECAPx2_ASAP7_75t_R FILLER_82_464 ();
 DECAPx1_ASAP7_75t_R FILLER_82_496 ();
 FILLER_ASAP7_75t_R FILLER_82_508 ();
 DECAPx10_ASAP7_75t_R FILLER_82_527 ();
 DECAPx6_ASAP7_75t_R FILLER_82_549 ();
 DECAPx2_ASAP7_75t_R FILLER_82_563 ();
 DECAPx1_ASAP7_75t_R FILLER_82_591 ();
 DECAPx4_ASAP7_75t_R FILLER_82_603 ();
 FILLER_ASAP7_75t_R FILLER_82_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_623 ();
 FILLER_ASAP7_75t_R FILLER_82_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_642 ();
 DECAPx10_ASAP7_75t_R FILLER_82_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_673 ();
 DECAPx4_ASAP7_75t_R FILLER_82_684 ();
 FILLER_ASAP7_75t_R FILLER_82_694 ();
 DECAPx2_ASAP7_75t_R FILLER_82_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_746 ();
 FILLER_ASAP7_75t_R FILLER_82_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_755 ();
 DECAPx1_ASAP7_75t_R FILLER_82_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_783 ();
 DECAPx1_ASAP7_75t_R FILLER_82_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_800 ();
 DECAPx10_ASAP7_75t_R FILLER_82_807 ();
 DECAPx2_ASAP7_75t_R FILLER_82_829 ();
 FILLER_ASAP7_75t_R FILLER_82_835 ();
 DECAPx10_ASAP7_75t_R FILLER_82_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_890 ();
 FILLER_ASAP7_75t_R FILLER_82_897 ();
 FILLER_ASAP7_75t_R FILLER_82_908 ();
 FILLER_ASAP7_75t_R FILLER_82_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_918 ();
 DECAPx2_ASAP7_75t_R FILLER_82_926 ();
 FILLER_ASAP7_75t_R FILLER_82_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_934 ();
 DECAPx1_ASAP7_75t_R FILLER_82_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_949 ();
 FILLER_ASAP7_75t_R FILLER_82_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_958 ();
 DECAPx6_ASAP7_75t_R FILLER_82_978 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1036 ();
 FILLER_ASAP7_75t_R FILLER_82_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1078 ();
 FILLER_ASAP7_75t_R FILLER_82_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1090 ();
 DECAPx4_ASAP7_75t_R FILLER_82_1114 ();
 FILLER_ASAP7_75t_R FILLER_82_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1156 ();
 FILLER_ASAP7_75t_R FILLER_82_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_82_1185 ();
 FILLER_ASAP7_75t_R FILLER_82_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1210 ();
 FILLER_ASAP7_75t_R FILLER_82_1216 ();
 DECAPx2_ASAP7_75t_R FILLER_83_2 ();
 FILLER_ASAP7_75t_R FILLER_83_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_10 ();
 DECAPx10_ASAP7_75t_R FILLER_83_17 ();
 DECAPx10_ASAP7_75t_R FILLER_83_39 ();
 DECAPx10_ASAP7_75t_R FILLER_83_61 ();
 DECAPx10_ASAP7_75t_R FILLER_83_83 ();
 FILLER_ASAP7_75t_R FILLER_83_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_138 ();
 DECAPx6_ASAP7_75t_R FILLER_83_151 ();
 FILLER_ASAP7_75t_R FILLER_83_165 ();
 DECAPx2_ASAP7_75t_R FILLER_83_178 ();
 DECAPx4_ASAP7_75t_R FILLER_83_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_263 ();
 DECAPx6_ASAP7_75t_R FILLER_83_270 ();
 FILLER_ASAP7_75t_R FILLER_83_313 ();
 FILLER_ASAP7_75t_R FILLER_83_321 ();
 DECAPx2_ASAP7_75t_R FILLER_83_329 ();
 DECAPx1_ASAP7_75t_R FILLER_83_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_349 ();
 DECAPx10_ASAP7_75t_R FILLER_83_383 ();
 DECAPx10_ASAP7_75t_R FILLER_83_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_427 ();
 FILLER_ASAP7_75t_R FILLER_83_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_441 ();
 DECAPx4_ASAP7_75t_R FILLER_83_448 ();
 DECAPx2_ASAP7_75t_R FILLER_83_466 ();
 FILLER_ASAP7_75t_R FILLER_83_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_474 ();
 FILLER_ASAP7_75t_R FILLER_83_502 ();
 DECAPx10_ASAP7_75t_R FILLER_83_526 ();
 DECAPx10_ASAP7_75t_R FILLER_83_548 ();
 DECAPx4_ASAP7_75t_R FILLER_83_570 ();
 FILLER_ASAP7_75t_R FILLER_83_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_622 ();
 DECAPx6_ASAP7_75t_R FILLER_83_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_653 ();
 DECAPx2_ASAP7_75t_R FILLER_83_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_670 ();
 DECAPx6_ASAP7_75t_R FILLER_83_691 ();
 DECAPx6_ASAP7_75t_R FILLER_83_727 ();
 FILLER_ASAP7_75t_R FILLER_83_741 ();
 DECAPx2_ASAP7_75t_R FILLER_83_759 ();
 FILLER_ASAP7_75t_R FILLER_83_765 ();
 DECAPx2_ASAP7_75t_R FILLER_83_773 ();
 FILLER_ASAP7_75t_R FILLER_83_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_781 ();
 FILLER_ASAP7_75t_R FILLER_83_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_790 ();
 FILLER_ASAP7_75t_R FILLER_83_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_818 ();
 DECAPx10_ASAP7_75t_R FILLER_83_826 ();
 DECAPx2_ASAP7_75t_R FILLER_83_848 ();
 FILLER_ASAP7_75t_R FILLER_83_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_856 ();
 DECAPx2_ASAP7_75t_R FILLER_83_879 ();
 FILLER_ASAP7_75t_R FILLER_83_885 ();
 DECAPx4_ASAP7_75t_R FILLER_83_899 ();
 FILLER_ASAP7_75t_R FILLER_83_922 ();
 DECAPx6_ASAP7_75t_R FILLER_83_926 ();
 DECAPx1_ASAP7_75t_R FILLER_83_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_951 ();
 DECAPx1_ASAP7_75t_R FILLER_83_963 ();
 DECAPx10_ASAP7_75t_R FILLER_83_985 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_83_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1052 ();
 DECAPx4_ASAP7_75t_R FILLER_83_1059 ();
 FILLER_ASAP7_75t_R FILLER_83_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1071 ();
 DECAPx4_ASAP7_75t_R FILLER_83_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1207 ();
 FILLER_ASAP7_75t_R FILLER_83_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1223 ();
 DECAPx4_ASAP7_75t_R FILLER_84_2 ();
 DECAPx10_ASAP7_75t_R FILLER_84_18 ();
 DECAPx10_ASAP7_75t_R FILLER_84_40 ();
 DECAPx10_ASAP7_75t_R FILLER_84_62 ();
 DECAPx10_ASAP7_75t_R FILLER_84_84 ();
 DECAPx10_ASAP7_75t_R FILLER_84_106 ();
 FILLER_ASAP7_75t_R FILLER_84_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_130 ();
 DECAPx6_ASAP7_75t_R FILLER_84_153 ();
 DECAPx1_ASAP7_75t_R FILLER_84_167 ();
 DECAPx6_ASAP7_75t_R FILLER_84_193 ();
 FILLER_ASAP7_75t_R FILLER_84_207 ();
 DECAPx1_ASAP7_75t_R FILLER_84_212 ();
 DECAPx6_ASAP7_75t_R FILLER_84_222 ();
 DECAPx1_ASAP7_75t_R FILLER_84_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_240 ();
 FILLER_ASAP7_75t_R FILLER_84_281 ();
 DECAPx10_ASAP7_75t_R FILLER_84_289 ();
 DECAPx6_ASAP7_75t_R FILLER_84_329 ();
 DECAPx1_ASAP7_75t_R FILLER_84_343 ();
 DECAPx2_ASAP7_75t_R FILLER_84_364 ();
 DECAPx2_ASAP7_75t_R FILLER_84_397 ();
 FILLER_ASAP7_75t_R FILLER_84_403 ();
 FILLER_ASAP7_75t_R FILLER_84_422 ();
 FILLER_ASAP7_75t_R FILLER_84_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_461 ();
 DECAPx4_ASAP7_75t_R FILLER_84_464 ();
 FILLER_ASAP7_75t_R FILLER_84_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_476 ();
 DECAPx10_ASAP7_75t_R FILLER_84_499 ();
 DECAPx6_ASAP7_75t_R FILLER_84_521 ();
 DECAPx10_ASAP7_75t_R FILLER_84_571 ();
 DECAPx6_ASAP7_75t_R FILLER_84_593 ();
 FILLER_ASAP7_75t_R FILLER_84_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_616 ();
 FILLER_ASAP7_75t_R FILLER_84_624 ();
 FILLER_ASAP7_75t_R FILLER_84_633 ();
 DECAPx1_ASAP7_75t_R FILLER_84_641 ();
 FILLER_ASAP7_75t_R FILLER_84_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_653 ();
 DECAPx2_ASAP7_75t_R FILLER_84_661 ();
 FILLER_ASAP7_75t_R FILLER_84_667 ();
 FILLER_ASAP7_75t_R FILLER_84_676 ();
 DECAPx10_ASAP7_75t_R FILLER_84_692 ();
 DECAPx10_ASAP7_75t_R FILLER_84_714 ();
 DECAPx6_ASAP7_75t_R FILLER_84_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_750 ();
 DECAPx2_ASAP7_75t_R FILLER_84_771 ();
 FILLER_ASAP7_75t_R FILLER_84_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_790 ();
 DECAPx2_ASAP7_75t_R FILLER_84_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_804 ();
 DECAPx2_ASAP7_75t_R FILLER_84_812 ();
 FILLER_ASAP7_75t_R FILLER_84_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_820 ();
 DECAPx2_ASAP7_75t_R FILLER_84_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_866 ();
 DECAPx1_ASAP7_75t_R FILLER_84_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_915 ();
 DECAPx6_ASAP7_75t_R FILLER_84_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_956 ();
 FILLER_ASAP7_75t_R FILLER_84_963 ();
 DECAPx1_ASAP7_75t_R FILLER_84_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_997 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1062 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1084 ();
 FILLER_ASAP7_75t_R FILLER_84_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1136 ();
 FILLER_ASAP7_75t_R FILLER_84_1147 ();
 FILLER_ASAP7_75t_R FILLER_84_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1168 ();
 FILLER_ASAP7_75t_R FILLER_84_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1191 ();
 FILLER_ASAP7_75t_R FILLER_84_1201 ();
 FILLER_ASAP7_75t_R FILLER_84_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_85_2 ();
 DECAPx10_ASAP7_75t_R FILLER_85_24 ();
 DECAPx10_ASAP7_75t_R FILLER_85_46 ();
 DECAPx10_ASAP7_75t_R FILLER_85_68 ();
 DECAPx10_ASAP7_75t_R FILLER_85_90 ();
 DECAPx6_ASAP7_75t_R FILLER_85_112 ();
 DECAPx6_ASAP7_75t_R FILLER_85_159 ();
 DECAPx10_ASAP7_75t_R FILLER_85_179 ();
 DECAPx1_ASAP7_75t_R FILLER_85_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_205 ();
 DECAPx10_ASAP7_75t_R FILLER_85_212 ();
 DECAPx4_ASAP7_75t_R FILLER_85_234 ();
 FILLER_ASAP7_75t_R FILLER_85_244 ();
 FILLER_ASAP7_75t_R FILLER_85_252 ();
 DECAPx2_ASAP7_75t_R FILLER_85_260 ();
 FILLER_ASAP7_75t_R FILLER_85_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_268 ();
 DECAPx1_ASAP7_75t_R FILLER_85_291 ();
 FILLER_ASAP7_75t_R FILLER_85_315 ();
 DECAPx1_ASAP7_75t_R FILLER_85_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_331 ();
 FILLER_ASAP7_75t_R FILLER_85_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_344 ();
 DECAPx4_ASAP7_75t_R FILLER_85_358 ();
 FILLER_ASAP7_75t_R FILLER_85_368 ();
 DECAPx10_ASAP7_75t_R FILLER_85_377 ();
 FILLER_ASAP7_75t_R FILLER_85_421 ();
 DECAPx10_ASAP7_75t_R FILLER_85_437 ();
 DECAPx10_ASAP7_75t_R FILLER_85_459 ();
 DECAPx6_ASAP7_75t_R FILLER_85_487 ();
 DECAPx2_ASAP7_75t_R FILLER_85_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_507 ();
 DECAPx6_ASAP7_75t_R FILLER_85_537 ();
 DECAPx6_ASAP7_75t_R FILLER_85_557 ();
 DECAPx1_ASAP7_75t_R FILLER_85_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_575 ();
 DECAPx1_ASAP7_75t_R FILLER_85_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_612 ();
 DECAPx2_ASAP7_75t_R FILLER_85_621 ();
 FILLER_ASAP7_75t_R FILLER_85_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_629 ();
 FILLER_ASAP7_75t_R FILLER_85_640 ();
 DECAPx2_ASAP7_75t_R FILLER_85_656 ();
 FILLER_ASAP7_75t_R FILLER_85_662 ();
 DECAPx6_ASAP7_75t_R FILLER_85_703 ();
 DECAPx1_ASAP7_75t_R FILLER_85_717 ();
 DECAPx4_ASAP7_75t_R FILLER_85_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_753 ();
 DECAPx2_ASAP7_75t_R FILLER_85_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_766 ();
 FILLER_ASAP7_75t_R FILLER_85_774 ();
 DECAPx2_ASAP7_75t_R FILLER_85_788 ();
 FILLER_ASAP7_75t_R FILLER_85_794 ();
 DECAPx1_ASAP7_75t_R FILLER_85_802 ();
 DECAPx10_ASAP7_75t_R FILLER_85_835 ();
 DECAPx10_ASAP7_75t_R FILLER_85_857 ();
 DECAPx6_ASAP7_75t_R FILLER_85_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_893 ();
 DECAPx2_ASAP7_75t_R FILLER_85_916 ();
 FILLER_ASAP7_75t_R FILLER_85_922 ();
 DECAPx4_ASAP7_75t_R FILLER_85_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_957 ();
 DECAPx1_ASAP7_75t_R FILLER_85_973 ();
 DECAPx10_ASAP7_75t_R FILLER_85_999 ();
 FILLER_ASAP7_75t_R FILLER_85_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1046 ();
 FILLER_ASAP7_75t_R FILLER_85_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1135 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1182 ();
 FILLER_ASAP7_75t_R FILLER_85_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1190 ();
 FILLER_ASAP7_75t_R FILLER_85_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_86_2 ();
 DECAPx10_ASAP7_75t_R FILLER_86_24 ();
 DECAPx10_ASAP7_75t_R FILLER_86_46 ();
 DECAPx10_ASAP7_75t_R FILLER_86_68 ();
 DECAPx10_ASAP7_75t_R FILLER_86_90 ();
 FILLER_ASAP7_75t_R FILLER_86_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_114 ();
 DECAPx1_ASAP7_75t_R FILLER_86_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_162 ();
 DECAPx2_ASAP7_75t_R FILLER_86_169 ();
 DECAPx10_ASAP7_75t_R FILLER_86_185 ();
 DECAPx10_ASAP7_75t_R FILLER_86_207 ();
 DECAPx4_ASAP7_75t_R FILLER_86_229 ();
 DECAPx1_ASAP7_75t_R FILLER_86_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_261 ();
 DECAPx2_ASAP7_75t_R FILLER_86_268 ();
 DECAPx2_ASAP7_75t_R FILLER_86_280 ();
 FILLER_ASAP7_75t_R FILLER_86_296 ();
 FILLER_ASAP7_75t_R FILLER_86_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_343 ();
 FILLER_ASAP7_75t_R FILLER_86_364 ();
 DECAPx2_ASAP7_75t_R FILLER_86_374 ();
 DECAPx10_ASAP7_75t_R FILLER_86_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_424 ();
 FILLER_ASAP7_75t_R FILLER_86_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_441 ();
 DECAPx4_ASAP7_75t_R FILLER_86_449 ();
 FILLER_ASAP7_75t_R FILLER_86_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_461 ();
 DECAPx6_ASAP7_75t_R FILLER_86_484 ();
 DECAPx2_ASAP7_75t_R FILLER_86_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_504 ();
 FILLER_ASAP7_75t_R FILLER_86_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_517 ();
 FILLER_ASAP7_75t_R FILLER_86_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_526 ();
 FILLER_ASAP7_75t_R FILLER_86_530 ();
 DECAPx10_ASAP7_75t_R FILLER_86_537 ();
 DECAPx2_ASAP7_75t_R FILLER_86_559 ();
 FILLER_ASAP7_75t_R FILLER_86_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_567 ();
 DECAPx1_ASAP7_75t_R FILLER_86_598 ();
 DECAPx1_ASAP7_75t_R FILLER_86_612 ();
 DECAPx6_ASAP7_75t_R FILLER_86_630 ();
 DECAPx1_ASAP7_75t_R FILLER_86_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_648 ();
 DECAPx6_ASAP7_75t_R FILLER_86_652 ();
 DECAPx2_ASAP7_75t_R FILLER_86_672 ();
 DECAPx2_ASAP7_75t_R FILLER_86_688 ();
 FILLER_ASAP7_75t_R FILLER_86_694 ();
 DECAPx10_ASAP7_75t_R FILLER_86_713 ();
 DECAPx10_ASAP7_75t_R FILLER_86_735 ();
 DECAPx6_ASAP7_75t_R FILLER_86_757 ();
 DECAPx1_ASAP7_75t_R FILLER_86_771 ();
 DECAPx6_ASAP7_75t_R FILLER_86_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_807 ();
 DECAPx1_ASAP7_75t_R FILLER_86_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_818 ();
 DECAPx6_ASAP7_75t_R FILLER_86_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_839 ();
 DECAPx2_ASAP7_75t_R FILLER_86_884 ();
 DECAPx1_ASAP7_75t_R FILLER_86_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_914 ();
 DECAPx4_ASAP7_75t_R FILLER_86_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_949 ();
 DECAPx1_ASAP7_75t_R FILLER_86_969 ();
 DECAPx6_ASAP7_75t_R FILLER_86_993 ();
 FILLER_ASAP7_75t_R FILLER_86_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1012 ();
 FILLER_ASAP7_75t_R FILLER_86_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1050 ();
 FILLER_ASAP7_75t_R FILLER_86_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_86_1115 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_86_1149 ();
 FILLER_ASAP7_75t_R FILLER_86_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_86_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1215 ();
 FILLER_ASAP7_75t_R FILLER_86_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_87_2 ();
 DECAPx10_ASAP7_75t_R FILLER_87_24 ();
 DECAPx10_ASAP7_75t_R FILLER_87_46 ();
 DECAPx10_ASAP7_75t_R FILLER_87_68 ();
 DECAPx10_ASAP7_75t_R FILLER_87_90 ();
 DECAPx6_ASAP7_75t_R FILLER_87_112 ();
 DECAPx2_ASAP7_75t_R FILLER_87_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_149 ();
 DECAPx1_ASAP7_75t_R FILLER_87_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_197 ();
 DECAPx10_ASAP7_75t_R FILLER_87_204 ();
 DECAPx6_ASAP7_75t_R FILLER_87_226 ();
 DECAPx2_ASAP7_75t_R FILLER_87_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_272 ();
 DECAPx1_ASAP7_75t_R FILLER_87_296 ();
 DECAPx4_ASAP7_75t_R FILLER_87_307 ();
 FILLER_ASAP7_75t_R FILLER_87_317 ();
 DECAPx2_ASAP7_75t_R FILLER_87_322 ();
 FILLER_ASAP7_75t_R FILLER_87_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_330 ();
 DECAPx4_ASAP7_75t_R FILLER_87_337 ();
 DECAPx1_ASAP7_75t_R FILLER_87_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_368 ();
 DECAPx1_ASAP7_75t_R FILLER_87_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_435 ();
 DECAPx1_ASAP7_75t_R FILLER_87_447 ();
 DECAPx6_ASAP7_75t_R FILLER_87_475 ();
 DECAPx2_ASAP7_75t_R FILLER_87_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_517 ();
 DECAPx10_ASAP7_75t_R FILLER_87_538 ();
 DECAPx1_ASAP7_75t_R FILLER_87_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_564 ();
 FILLER_ASAP7_75t_R FILLER_87_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_589 ();
 DECAPx1_ASAP7_75t_R FILLER_87_598 ();
 DECAPx2_ASAP7_75t_R FILLER_87_612 ();
 FILLER_ASAP7_75t_R FILLER_87_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_620 ();
 DECAPx4_ASAP7_75t_R FILLER_87_624 ();
 DECAPx1_ASAP7_75t_R FILLER_87_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_648 ();
 DECAPx2_ASAP7_75t_R FILLER_87_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_665 ();
 DECAPx2_ASAP7_75t_R FILLER_87_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_705 ();
 DECAPx4_ASAP7_75t_R FILLER_87_716 ();
 FILLER_ASAP7_75t_R FILLER_87_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_728 ();
 DECAPx10_ASAP7_75t_R FILLER_87_751 ();
 DECAPx4_ASAP7_75t_R FILLER_87_773 ();
 DECAPx1_ASAP7_75t_R FILLER_87_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_810 ();
 DECAPx1_ASAP7_75t_R FILLER_87_818 ();
 DECAPx10_ASAP7_75t_R FILLER_87_851 ();
 DECAPx6_ASAP7_75t_R FILLER_87_873 ();
 DECAPx1_ASAP7_75t_R FILLER_87_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_891 ();
 DECAPx1_ASAP7_75t_R FILLER_87_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_923 ();
 DECAPx6_ASAP7_75t_R FILLER_87_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_940 ();
 DECAPx10_ASAP7_75t_R FILLER_87_956 ();
 DECAPx2_ASAP7_75t_R FILLER_87_978 ();
 FILLER_ASAP7_75t_R FILLER_87_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_986 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1009 ();
 FILLER_ASAP7_75t_R FILLER_87_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1075 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1153 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1201 ();
 FILLER_ASAP7_75t_R FILLER_87_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_88_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_24 ();
 DECAPx10_ASAP7_75t_R FILLER_88_31 ();
 DECAPx10_ASAP7_75t_R FILLER_88_53 ();
 DECAPx10_ASAP7_75t_R FILLER_88_75 ();
 DECAPx10_ASAP7_75t_R FILLER_88_97 ();
 DECAPx6_ASAP7_75t_R FILLER_88_119 ();
 FILLER_ASAP7_75t_R FILLER_88_133 ();
 DECAPx4_ASAP7_75t_R FILLER_88_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_151 ();
 DECAPx6_ASAP7_75t_R FILLER_88_158 ();
 DECAPx1_ASAP7_75t_R FILLER_88_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_176 ();
 DECAPx2_ASAP7_75t_R FILLER_88_180 ();
 FILLER_ASAP7_75t_R FILLER_88_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_188 ();
 DECAPx10_ASAP7_75t_R FILLER_88_213 ();
 DECAPx6_ASAP7_75t_R FILLER_88_235 ();
 DECAPx2_ASAP7_75t_R FILLER_88_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_255 ();
 DECAPx4_ASAP7_75t_R FILLER_88_284 ();
 FILLER_ASAP7_75t_R FILLER_88_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_296 ();
 DECAPx4_ASAP7_75t_R FILLER_88_303 ();
 FILLER_ASAP7_75t_R FILLER_88_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_315 ();
 DECAPx4_ASAP7_75t_R FILLER_88_336 ();
 FILLER_ASAP7_75t_R FILLER_88_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_348 ();
 DECAPx6_ASAP7_75t_R FILLER_88_352 ();
 DECAPx6_ASAP7_75t_R FILLER_88_385 ();
 DECAPx1_ASAP7_75t_R FILLER_88_421 ();
 FILLER_ASAP7_75t_R FILLER_88_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_464 ();
 DECAPx4_ASAP7_75t_R FILLER_88_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_509 ();
 DECAPx10_ASAP7_75t_R FILLER_88_527 ();
 DECAPx6_ASAP7_75t_R FILLER_88_549 ();
 DECAPx2_ASAP7_75t_R FILLER_88_595 ();
 FILLER_ASAP7_75t_R FILLER_88_601 ();
 FILLER_ASAP7_75t_R FILLER_88_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_617 ();
 DECAPx2_ASAP7_75t_R FILLER_88_633 ();
 FILLER_ASAP7_75t_R FILLER_88_639 ();
 DECAPx6_ASAP7_75t_R FILLER_88_644 ();
 DECAPx1_ASAP7_75t_R FILLER_88_658 ();
 DECAPx2_ASAP7_75t_R FILLER_88_676 ();
 FILLER_ASAP7_75t_R FILLER_88_682 ();
 DECAPx2_ASAP7_75t_R FILLER_88_690 ();
 FILLER_ASAP7_75t_R FILLER_88_696 ();
 DECAPx10_ASAP7_75t_R FILLER_88_718 ();
 DECAPx4_ASAP7_75t_R FILLER_88_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_750 ();
 DECAPx1_ASAP7_75t_R FILLER_88_795 ();
 FILLER_ASAP7_75t_R FILLER_88_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_814 ();
 DECAPx10_ASAP7_75t_R FILLER_88_822 ();
 DECAPx10_ASAP7_75t_R FILLER_88_844 ();
 DECAPx6_ASAP7_75t_R FILLER_88_866 ();
 DECAPx2_ASAP7_75t_R FILLER_88_880 ();
 DECAPx2_ASAP7_75t_R FILLER_88_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_898 ();
 DECAPx6_ASAP7_75t_R FILLER_88_917 ();
 DECAPx1_ASAP7_75t_R FILLER_88_931 ();
 DECAPx4_ASAP7_75t_R FILLER_88_950 ();
 FILLER_ASAP7_75t_R FILLER_88_960 ();
 DECAPx10_ASAP7_75t_R FILLER_88_972 ();
 DECAPx10_ASAP7_75t_R FILLER_88_994 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1016 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1068 ();
 FILLER_ASAP7_75t_R FILLER_88_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1115 ();
 FILLER_ASAP7_75t_R FILLER_88_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1131 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1138 ();
 FILLER_ASAP7_75t_R FILLER_88_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1157 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1170 ();
 FILLER_ASAP7_75t_R FILLER_88_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1182 ();
 FILLER_ASAP7_75t_R FILLER_88_1189 ();
 FILLER_ASAP7_75t_R FILLER_88_1197 ();
 FILLER_ASAP7_75t_R FILLER_88_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_89_2 ();
 FILLER_ASAP7_75t_R FILLER_89_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_10 ();
 DECAPx10_ASAP7_75t_R FILLER_89_17 ();
 DECAPx10_ASAP7_75t_R FILLER_89_39 ();
 DECAPx10_ASAP7_75t_R FILLER_89_61 ();
 DECAPx10_ASAP7_75t_R FILLER_89_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_105 ();
 DECAPx4_ASAP7_75t_R FILLER_89_112 ();
 DECAPx4_ASAP7_75t_R FILLER_89_144 ();
 FILLER_ASAP7_75t_R FILLER_89_154 ();
 DECAPx2_ASAP7_75t_R FILLER_89_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_168 ();
 DECAPx10_ASAP7_75t_R FILLER_89_180 ();
 DECAPx10_ASAP7_75t_R FILLER_89_202 ();
 DECAPx4_ASAP7_75t_R FILLER_89_224 ();
 FILLER_ASAP7_75t_R FILLER_89_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_277 ();
 FILLER_ASAP7_75t_R FILLER_89_284 ();
 DECAPx1_ASAP7_75t_R FILLER_89_306 ();
 FILLER_ASAP7_75t_R FILLER_89_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_321 ();
 DECAPx4_ASAP7_75t_R FILLER_89_337 ();
 FILLER_ASAP7_75t_R FILLER_89_347 ();
 DECAPx6_ASAP7_75t_R FILLER_89_355 ();
 DECAPx1_ASAP7_75t_R FILLER_89_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_373 ();
 DECAPx10_ASAP7_75t_R FILLER_89_394 ();
 DECAPx10_ASAP7_75t_R FILLER_89_416 ();
 DECAPx2_ASAP7_75t_R FILLER_89_438 ();
 DECAPx2_ASAP7_75t_R FILLER_89_450 ();
 DECAPx10_ASAP7_75t_R FILLER_89_463 ();
 DECAPx2_ASAP7_75t_R FILLER_89_485 ();
 FILLER_ASAP7_75t_R FILLER_89_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_493 ();
 DECAPx4_ASAP7_75t_R FILLER_89_502 ();
 FILLER_ASAP7_75t_R FILLER_89_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_514 ();
 DECAPx4_ASAP7_75t_R FILLER_89_541 ();
 FILLER_ASAP7_75t_R FILLER_89_551 ();
 DECAPx6_ASAP7_75t_R FILLER_89_573 ();
 DECAPx2_ASAP7_75t_R FILLER_89_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_593 ();
 FILLER_ASAP7_75t_R FILLER_89_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_602 ();
 FILLER_ASAP7_75t_R FILLER_89_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_633 ();
 DECAPx6_ASAP7_75t_R FILLER_89_648 ();
 DECAPx2_ASAP7_75t_R FILLER_89_671 ();
 FILLER_ASAP7_75t_R FILLER_89_677 ();
 DECAPx10_ASAP7_75t_R FILLER_89_706 ();
 DECAPx6_ASAP7_75t_R FILLER_89_728 ();
 FILLER_ASAP7_75t_R FILLER_89_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_744 ();
 DECAPx6_ASAP7_75t_R FILLER_89_767 ();
 DECAPx1_ASAP7_75t_R FILLER_89_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_785 ();
 DECAPx4_ASAP7_75t_R FILLER_89_796 ();
 DECAPx10_ASAP7_75t_R FILLER_89_819 ();
 DECAPx2_ASAP7_75t_R FILLER_89_841 ();
 FILLER_ASAP7_75t_R FILLER_89_847 ();
 FILLER_ASAP7_75t_R FILLER_89_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_883 ();
 DECAPx2_ASAP7_75t_R FILLER_89_916 ();
 FILLER_ASAP7_75t_R FILLER_89_922 ();
 DECAPx1_ASAP7_75t_R FILLER_89_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_942 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1001 ();
 FILLER_ASAP7_75t_R FILLER_89_1015 ();
 FILLER_ASAP7_75t_R FILLER_89_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1022 ();
 DECAPx1_ASAP7_75t_R FILLER_89_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1047 ();
 FILLER_ASAP7_75t_R FILLER_89_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_89_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1143 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1168 ();
 FILLER_ASAP7_75t_R FILLER_89_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_90_2 ();
 DECAPx10_ASAP7_75t_R FILLER_90_24 ();
 DECAPx10_ASAP7_75t_R FILLER_90_46 ();
 DECAPx10_ASAP7_75t_R FILLER_90_68 ();
 DECAPx1_ASAP7_75t_R FILLER_90_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_131 ();
 FILLER_ASAP7_75t_R FILLER_90_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_150 ();
 FILLER_ASAP7_75t_R FILLER_90_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_175 ();
 FILLER_ASAP7_75t_R FILLER_90_198 ();
 DECAPx10_ASAP7_75t_R FILLER_90_220 ();
 DECAPx10_ASAP7_75t_R FILLER_90_248 ();
 DECAPx10_ASAP7_75t_R FILLER_90_270 ();
 DECAPx6_ASAP7_75t_R FILLER_90_292 ();
 DECAPx4_ASAP7_75t_R FILLER_90_318 ();
 FILLER_ASAP7_75t_R FILLER_90_328 ();
 DECAPx2_ASAP7_75t_R FILLER_90_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_342 ();
 FILLER_ASAP7_75t_R FILLER_90_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_375 ();
 FILLER_ASAP7_75t_R FILLER_90_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_397 ();
 FILLER_ASAP7_75t_R FILLER_90_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_410 ();
 DECAPx1_ASAP7_75t_R FILLER_90_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_440 ();
 DECAPx2_ASAP7_75t_R FILLER_90_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_461 ();
 DECAPx4_ASAP7_75t_R FILLER_90_464 ();
 FILLER_ASAP7_75t_R FILLER_90_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_476 ();
 DECAPx2_ASAP7_75t_R FILLER_90_485 ();
 DECAPx10_ASAP7_75t_R FILLER_90_507 ();
 DECAPx10_ASAP7_75t_R FILLER_90_529 ();
 DECAPx2_ASAP7_75t_R FILLER_90_551 ();
 DECAPx2_ASAP7_75t_R FILLER_90_563 ();
 DECAPx4_ASAP7_75t_R FILLER_90_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_599 ();
 DECAPx2_ASAP7_75t_R FILLER_90_610 ();
 DECAPx6_ASAP7_75t_R FILLER_90_622 ();
 DECAPx1_ASAP7_75t_R FILLER_90_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_646 ();
 DECAPx2_ASAP7_75t_R FILLER_90_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_660 ();
 DECAPx1_ASAP7_75t_R FILLER_90_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_673 ();
 FILLER_ASAP7_75t_R FILLER_90_677 ();
 DECAPx4_ASAP7_75t_R FILLER_90_685 ();
 FILLER_ASAP7_75t_R FILLER_90_695 ();
 FILLER_ASAP7_75t_R FILLER_90_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_705 ();
 DECAPx6_ASAP7_75t_R FILLER_90_718 ();
 DECAPx1_ASAP7_75t_R FILLER_90_732 ();
 DECAPx2_ASAP7_75t_R FILLER_90_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_762 ();
 DECAPx4_ASAP7_75t_R FILLER_90_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_813 ();
 DECAPx4_ASAP7_75t_R FILLER_90_827 ();
 FILLER_ASAP7_75t_R FILLER_90_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_839 ();
 DECAPx4_ASAP7_75t_R FILLER_90_890 ();
 FILLER_ASAP7_75t_R FILLER_90_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_902 ();
 DECAPx1_ASAP7_75t_R FILLER_90_917 ();
 DECAPx2_ASAP7_75t_R FILLER_90_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_941 ();
 DECAPx1_ASAP7_75t_R FILLER_90_948 ();
 DECAPx2_ASAP7_75t_R FILLER_90_959 ();
 FILLER_ASAP7_75t_R FILLER_90_965 ();
 DECAPx2_ASAP7_75t_R FILLER_90_973 ();
 FILLER_ASAP7_75t_R FILLER_90_979 ();
 DECAPx6_ASAP7_75t_R FILLER_90_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1026 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1056 ();
 FILLER_ASAP7_75t_R FILLER_90_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1064 ();
 FILLER_ASAP7_75t_R FILLER_90_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1103 ();
 FILLER_ASAP7_75t_R FILLER_90_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1155 ();
 FILLER_ASAP7_75t_R FILLER_90_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1189 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1196 ();
 FILLER_ASAP7_75t_R FILLER_90_1202 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_91_2 ();
 DECAPx10_ASAP7_75t_R FILLER_91_24 ();
 DECAPx10_ASAP7_75t_R FILLER_91_46 ();
 DECAPx10_ASAP7_75t_R FILLER_91_68 ();
 FILLER_ASAP7_75t_R FILLER_91_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_92 ();
 FILLER_ASAP7_75t_R FILLER_91_116 ();
 FILLER_ASAP7_75t_R FILLER_91_129 ();
 DECAPx2_ASAP7_75t_R FILLER_91_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_170 ();
 DECAPx1_ASAP7_75t_R FILLER_91_183 ();
 DECAPx6_ASAP7_75t_R FILLER_91_204 ();
 FILLER_ASAP7_75t_R FILLER_91_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_220 ();
 DECAPx6_ASAP7_75t_R FILLER_91_231 ();
 DECAPx2_ASAP7_75t_R FILLER_91_251 ();
 FILLER_ASAP7_75t_R FILLER_91_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_285 ();
 FILLER_ASAP7_75t_R FILLER_91_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_292 ();
 DECAPx1_ASAP7_75t_R FILLER_91_327 ();
 DECAPx6_ASAP7_75t_R FILLER_91_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_367 ();
 DECAPx2_ASAP7_75t_R FILLER_91_390 ();
 FILLER_ASAP7_75t_R FILLER_91_406 ();
 DECAPx2_ASAP7_75t_R FILLER_91_465 ();
 FILLER_ASAP7_75t_R FILLER_91_471 ();
 DECAPx10_ASAP7_75t_R FILLER_91_517 ();
 DECAPx10_ASAP7_75t_R FILLER_91_539 ();
 DECAPx10_ASAP7_75t_R FILLER_91_561 ();
 FILLER_ASAP7_75t_R FILLER_91_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_594 ();
 DECAPx2_ASAP7_75t_R FILLER_91_611 ();
 FILLER_ASAP7_75t_R FILLER_91_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_619 ();
 FILLER_ASAP7_75t_R FILLER_91_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_638 ();
 DECAPx2_ASAP7_75t_R FILLER_91_655 ();
 FILLER_ASAP7_75t_R FILLER_91_661 ();
 DECAPx1_ASAP7_75t_R FILLER_91_669 ();
 FILLER_ASAP7_75t_R FILLER_91_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_696 ();
 FILLER_ASAP7_75t_R FILLER_91_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_725 ();
 DECAPx6_ASAP7_75t_R FILLER_91_736 ();
 DECAPx6_ASAP7_75t_R FILLER_91_772 ();
 DECAPx1_ASAP7_75t_R FILLER_91_786 ();
 DECAPx1_ASAP7_75t_R FILLER_91_812 ();
 FILLER_ASAP7_75t_R FILLER_91_838 ();
 DECAPx10_ASAP7_75t_R FILLER_91_850 ();
 DECAPx4_ASAP7_75t_R FILLER_91_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_882 ();
 FILLER_ASAP7_75t_R FILLER_91_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_911 ();
 DECAPx2_ASAP7_75t_R FILLER_91_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_934 ();
 DECAPx1_ASAP7_75t_R FILLER_91_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_961 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1016 ();
 FILLER_ASAP7_75t_R FILLER_91_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1058 ();
 FILLER_ASAP7_75t_R FILLER_91_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1081 ();
 FILLER_ASAP7_75t_R FILLER_91_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1115 ();
 DECAPx6_ASAP7_75t_R FILLER_91_1131 ();
 FILLER_ASAP7_75t_R FILLER_91_1145 ();
 FILLER_ASAP7_75t_R FILLER_91_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1166 ();
 FILLER_ASAP7_75t_R FILLER_91_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1174 ();
 DECAPx6_ASAP7_75t_R FILLER_91_1197 ();
 FILLER_ASAP7_75t_R FILLER_91_1211 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1223 ();
 FILLER_ASAP7_75t_R FILLER_92_2 ();
 DECAPx10_ASAP7_75t_R FILLER_92_16 ();
 DECAPx10_ASAP7_75t_R FILLER_92_38 ();
 DECAPx10_ASAP7_75t_R FILLER_92_60 ();
 DECAPx10_ASAP7_75t_R FILLER_92_82 ();
 FILLER_ASAP7_75t_R FILLER_92_112 ();
 DECAPx1_ASAP7_75t_R FILLER_92_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_134 ();
 DECAPx4_ASAP7_75t_R FILLER_92_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_167 ();
 FILLER_ASAP7_75t_R FILLER_92_175 ();
 DECAPx10_ASAP7_75t_R FILLER_92_185 ();
 DECAPx10_ASAP7_75t_R FILLER_92_207 ();
 FILLER_ASAP7_75t_R FILLER_92_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_231 ();
 DECAPx1_ASAP7_75t_R FILLER_92_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_256 ();
 DECAPx10_ASAP7_75t_R FILLER_92_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_285 ();
 FILLER_ASAP7_75t_R FILLER_92_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_308 ();
 DECAPx10_ASAP7_75t_R FILLER_92_321 ();
 DECAPx2_ASAP7_75t_R FILLER_92_343 ();
 FILLER_ASAP7_75t_R FILLER_92_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_359 ();
 DECAPx10_ASAP7_75t_R FILLER_92_372 ();
 DECAPx10_ASAP7_75t_R FILLER_92_394 ();
 DECAPx4_ASAP7_75t_R FILLER_92_416 ();
 DECAPx2_ASAP7_75t_R FILLER_92_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_454 ();
 FILLER_ASAP7_75t_R FILLER_92_464 ();
 DECAPx1_ASAP7_75t_R FILLER_92_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_490 ();
 DECAPx10_ASAP7_75t_R FILLER_92_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_566 ();
 DECAPx1_ASAP7_75t_R FILLER_92_597 ();
 DECAPx1_ASAP7_75t_R FILLER_92_629 ();
 DECAPx1_ASAP7_75t_R FILLER_92_639 ();
 DECAPx4_ASAP7_75t_R FILLER_92_651 ();
 FILLER_ASAP7_75t_R FILLER_92_673 ();
 DECAPx4_ASAP7_75t_R FILLER_92_678 ();
 FILLER_ASAP7_75t_R FILLER_92_688 ();
 FILLER_ASAP7_75t_R FILLER_92_709 ();
 DECAPx10_ASAP7_75t_R FILLER_92_728 ();
 DECAPx10_ASAP7_75t_R FILLER_92_750 ();
 DECAPx1_ASAP7_75t_R FILLER_92_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_776 ();
 DECAPx2_ASAP7_75t_R FILLER_92_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_827 ();
 DECAPx2_ASAP7_75t_R FILLER_92_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_856 ();
 DECAPx6_ASAP7_75t_R FILLER_92_879 ();
 FILLER_ASAP7_75t_R FILLER_92_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_895 ();
 DECAPx10_ASAP7_75t_R FILLER_92_916 ();
 DECAPx2_ASAP7_75t_R FILLER_92_950 ();
 DECAPx10_ASAP7_75t_R FILLER_92_969 ();
 DECAPx10_ASAP7_75t_R FILLER_92_991 ();
 FILLER_ASAP7_75t_R FILLER_92_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1026 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1059 ();
 FILLER_ASAP7_75t_R FILLER_92_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1099 ();
 FILLER_ASAP7_75t_R FILLER_92_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1181 ();
 FILLER_ASAP7_75t_R FILLER_92_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1196 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1208 ();
 FILLER_ASAP7_75t_R FILLER_92_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_93_2 ();
 DECAPx10_ASAP7_75t_R FILLER_93_24 ();
 DECAPx10_ASAP7_75t_R FILLER_93_46 ();
 DECAPx6_ASAP7_75t_R FILLER_93_68 ();
 DECAPx2_ASAP7_75t_R FILLER_93_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_88 ();
 DECAPx2_ASAP7_75t_R FILLER_93_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_123 ();
 DECAPx6_ASAP7_75t_R FILLER_93_141 ();
 FILLER_ASAP7_75t_R FILLER_93_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_157 ();
 FILLER_ASAP7_75t_R FILLER_93_168 ();
 DECAPx10_ASAP7_75t_R FILLER_93_182 ();
 DECAPx10_ASAP7_75t_R FILLER_93_204 ();
 DECAPx10_ASAP7_75t_R FILLER_93_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_248 ();
 FILLER_ASAP7_75t_R FILLER_93_277 ();
 DECAPx2_ASAP7_75t_R FILLER_93_282 ();
 DECAPx4_ASAP7_75t_R FILLER_93_329 ();
 DECAPx2_ASAP7_75t_R FILLER_93_345 ();
 FILLER_ASAP7_75t_R FILLER_93_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_353 ();
 DECAPx6_ASAP7_75t_R FILLER_93_376 ();
 DECAPx2_ASAP7_75t_R FILLER_93_390 ();
 DECAPx6_ASAP7_75t_R FILLER_93_408 ();
 DECAPx2_ASAP7_75t_R FILLER_93_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_428 ();
 DECAPx10_ASAP7_75t_R FILLER_93_435 ();
 FILLER_ASAP7_75t_R FILLER_93_457 ();
 DECAPx10_ASAP7_75t_R FILLER_93_485 ();
 DECAPx6_ASAP7_75t_R FILLER_93_507 ();
 DECAPx10_ASAP7_75t_R FILLER_93_527 ();
 DECAPx4_ASAP7_75t_R FILLER_93_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_559 ();
 DECAPx4_ASAP7_75t_R FILLER_93_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_610 ();
 DECAPx4_ASAP7_75t_R FILLER_93_617 ();
 FILLER_ASAP7_75t_R FILLER_93_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_629 ();
 DECAPx10_ASAP7_75t_R FILLER_93_636 ();
 DECAPx1_ASAP7_75t_R FILLER_93_658 ();
 FILLER_ASAP7_75t_R FILLER_93_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_679 ();
 DECAPx4_ASAP7_75t_R FILLER_93_692 ();
 FILLER_ASAP7_75t_R FILLER_93_702 ();
 DECAPx2_ASAP7_75t_R FILLER_93_715 ();
 FILLER_ASAP7_75t_R FILLER_93_721 ();
 DECAPx10_ASAP7_75t_R FILLER_93_726 ();
 DECAPx10_ASAP7_75t_R FILLER_93_770 ();
 DECAPx6_ASAP7_75t_R FILLER_93_814 ();
 DECAPx2_ASAP7_75t_R FILLER_93_828 ();
 DECAPx10_ASAP7_75t_R FILLER_93_856 ();
 DECAPx6_ASAP7_75t_R FILLER_93_878 ();
 FILLER_ASAP7_75t_R FILLER_93_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_915 ();
 FILLER_ASAP7_75t_R FILLER_93_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_926 ();
 FILLER_ASAP7_75t_R FILLER_93_933 ();
 DECAPx4_ASAP7_75t_R FILLER_93_941 ();
 FILLER_ASAP7_75t_R FILLER_93_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_956 ();
 FILLER_ASAP7_75t_R FILLER_93_965 ();
 DECAPx6_ASAP7_75t_R FILLER_93_987 ();
 FILLER_ASAP7_75t_R FILLER_93_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1034 ();
 FILLER_ASAP7_75t_R FILLER_93_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_93_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_93_1078 ();
 FILLER_ASAP7_75t_R FILLER_93_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1090 ();
 FILLER_ASAP7_75t_R FILLER_93_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1127 ();
 FILLER_ASAP7_75t_R FILLER_93_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1176 ();
 FILLER_ASAP7_75t_R FILLER_93_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_93_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_94_2 ();
 DECAPx10_ASAP7_75t_R FILLER_94_24 ();
 DECAPx10_ASAP7_75t_R FILLER_94_46 ();
 DECAPx10_ASAP7_75t_R FILLER_94_68 ();
 DECAPx6_ASAP7_75t_R FILLER_94_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_104 ();
 FILLER_ASAP7_75t_R FILLER_94_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_113 ();
 DECAPx6_ASAP7_75t_R FILLER_94_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_164 ();
 DECAPx2_ASAP7_75t_R FILLER_94_187 ();
 FILLER_ASAP7_75t_R FILLER_94_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_195 ();
 DECAPx10_ASAP7_75t_R FILLER_94_218 ();
 FILLER_ASAP7_75t_R FILLER_94_240 ();
 DECAPx10_ASAP7_75t_R FILLER_94_248 ();
 FILLER_ASAP7_75t_R FILLER_94_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_272 ();
 DECAPx1_ASAP7_75t_R FILLER_94_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_320 ();
 DECAPx2_ASAP7_75t_R FILLER_94_367 ();
 FILLER_ASAP7_75t_R FILLER_94_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_393 ();
 DECAPx10_ASAP7_75t_R FILLER_94_417 ();
 DECAPx1_ASAP7_75t_R FILLER_94_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_450 ();
 DECAPx2_ASAP7_75t_R FILLER_94_464 ();
 FILLER_ASAP7_75t_R FILLER_94_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_472 ();
 DECAPx2_ASAP7_75t_R FILLER_94_481 ();
 FILLER_ASAP7_75t_R FILLER_94_487 ();
 DECAPx4_ASAP7_75t_R FILLER_94_500 ();
 DECAPx6_ASAP7_75t_R FILLER_94_543 ();
 FILLER_ASAP7_75t_R FILLER_94_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_559 ();
 DECAPx2_ASAP7_75t_R FILLER_94_578 ();
 FILLER_ASAP7_75t_R FILLER_94_584 ();
 DECAPx6_ASAP7_75t_R FILLER_94_616 ();
 FILLER_ASAP7_75t_R FILLER_94_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_652 ();
 DECAPx2_ASAP7_75t_R FILLER_94_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_705 ();
 DECAPx1_ASAP7_75t_R FILLER_94_712 ();
 DECAPx10_ASAP7_75t_R FILLER_94_747 ();
 FILLER_ASAP7_75t_R FILLER_94_769 ();
 DECAPx2_ASAP7_75t_R FILLER_94_793 ();
 DECAPx6_ASAP7_75t_R FILLER_94_841 ();
 DECAPx1_ASAP7_75t_R FILLER_94_855 ();
 FILLER_ASAP7_75t_R FILLER_94_877 ();
 DECAPx6_ASAP7_75t_R FILLER_94_893 ();
 FILLER_ASAP7_75t_R FILLER_94_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_933 ();
 DECAPx1_ASAP7_75t_R FILLER_94_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_947 ();
 DECAPx6_ASAP7_75t_R FILLER_94_964 ();
 FILLER_ASAP7_75t_R FILLER_94_978 ();
 DECAPx10_ASAP7_75t_R FILLER_94_986 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1008 ();
 FILLER_ASAP7_75t_R FILLER_94_1018 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_94_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1073 ();
 DECAPx6_ASAP7_75t_R FILLER_94_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1126 ();
 FILLER_ASAP7_75t_R FILLER_94_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1167 ();
 FILLER_ASAP7_75t_R FILLER_94_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1185 ();
 FILLER_ASAP7_75t_R FILLER_94_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_95_2 ();
 DECAPx10_ASAP7_75t_R FILLER_95_24 ();
 DECAPx10_ASAP7_75t_R FILLER_95_46 ();
 DECAPx6_ASAP7_75t_R FILLER_95_68 ();
 FILLER_ASAP7_75t_R FILLER_95_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_84 ();
 DECAPx2_ASAP7_75t_R FILLER_95_96 ();
 FILLER_ASAP7_75t_R FILLER_95_108 ();
 DECAPx10_ASAP7_75t_R FILLER_95_118 ();
 DECAPx10_ASAP7_75t_R FILLER_95_140 ();
 DECAPx2_ASAP7_75t_R FILLER_95_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_168 ();
 DECAPx2_ASAP7_75t_R FILLER_95_183 ();
 DECAPx10_ASAP7_75t_R FILLER_95_206 ();
 DECAPx2_ASAP7_75t_R FILLER_95_228 ();
 FILLER_ASAP7_75t_R FILLER_95_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_236 ();
 DECAPx6_ASAP7_75t_R FILLER_95_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_295 ();
 DECAPx10_ASAP7_75t_R FILLER_95_300 ();
 DECAPx1_ASAP7_75t_R FILLER_95_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_326 ();
 DECAPx10_ASAP7_75t_R FILLER_95_347 ();
 DECAPx2_ASAP7_75t_R FILLER_95_369 ();
 FILLER_ASAP7_75t_R FILLER_95_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_377 ();
 DECAPx2_ASAP7_75t_R FILLER_95_403 ();
 FILLER_ASAP7_75t_R FILLER_95_409 ();
 DECAPx6_ASAP7_75t_R FILLER_95_424 ();
 FILLER_ASAP7_75t_R FILLER_95_438 ();
 FILLER_ASAP7_75t_R FILLER_95_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_470 ();
 DECAPx1_ASAP7_75t_R FILLER_95_515 ();
 DECAPx2_ASAP7_75t_R FILLER_95_525 ();
 FILLER_ASAP7_75t_R FILLER_95_531 ();
 DECAPx2_ASAP7_75t_R FILLER_95_559 ();
 FILLER_ASAP7_75t_R FILLER_95_565 ();
 DECAPx6_ASAP7_75t_R FILLER_95_611 ();
 DECAPx1_ASAP7_75t_R FILLER_95_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_629 ();
 DECAPx6_ASAP7_75t_R FILLER_95_638 ();
 FILLER_ASAP7_75t_R FILLER_95_652 ();
 DECAPx1_ASAP7_75t_R FILLER_95_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_664 ();
 DECAPx1_ASAP7_75t_R FILLER_95_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_675 ();
 FILLER_ASAP7_75t_R FILLER_95_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_695 ();
 DECAPx10_ASAP7_75t_R FILLER_95_738 ();
 DECAPx10_ASAP7_75t_R FILLER_95_760 ();
 DECAPx6_ASAP7_75t_R FILLER_95_782 ();
 DECAPx2_ASAP7_75t_R FILLER_95_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_825 ();
 DECAPx10_ASAP7_75t_R FILLER_95_848 ();
 DECAPx10_ASAP7_75t_R FILLER_95_870 ();
 DECAPx2_ASAP7_75t_R FILLER_95_892 ();
 FILLER_ASAP7_75t_R FILLER_95_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_900 ();
 DECAPx2_ASAP7_75t_R FILLER_95_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_947 ();
 DECAPx2_ASAP7_75t_R FILLER_95_954 ();
 FILLER_ASAP7_75t_R FILLER_95_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_962 ();
 DECAPx6_ASAP7_75t_R FILLER_95_985 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1059 ();
 FILLER_ASAP7_75t_R FILLER_95_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1111 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1143 ();
 FILLER_ASAP7_75t_R FILLER_95_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_96_2 ();
 DECAPx10_ASAP7_75t_R FILLER_96_24 ();
 DECAPx10_ASAP7_75t_R FILLER_96_46 ();
 DECAPx1_ASAP7_75t_R FILLER_96_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_72 ();
 DECAPx1_ASAP7_75t_R FILLER_96_95 ();
 FILLER_ASAP7_75t_R FILLER_96_133 ();
 DECAPx1_ASAP7_75t_R FILLER_96_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_167 ();
 DECAPx2_ASAP7_75t_R FILLER_96_183 ();
 FILLER_ASAP7_75t_R FILLER_96_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_191 ();
 DECAPx2_ASAP7_75t_R FILLER_96_204 ();
 FILLER_ASAP7_75t_R FILLER_96_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_212 ();
 DECAPx6_ASAP7_75t_R FILLER_96_235 ();
 DECAPx1_ASAP7_75t_R FILLER_96_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_253 ();
 FILLER_ASAP7_75t_R FILLER_96_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_262 ();
 DECAPx6_ASAP7_75t_R FILLER_96_285 ();
 DECAPx1_ASAP7_75t_R FILLER_96_299 ();
 DECAPx6_ASAP7_75t_R FILLER_96_325 ();
 DECAPx1_ASAP7_75t_R FILLER_96_339 ();
 DECAPx1_ASAP7_75t_R FILLER_96_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_367 ();
 DECAPx4_ASAP7_75t_R FILLER_96_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_396 ();
 FILLER_ASAP7_75t_R FILLER_96_403 ();
 DECAPx6_ASAP7_75t_R FILLER_96_431 ();
 DECAPx4_ASAP7_75t_R FILLER_96_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_474 ();
 DECAPx4_ASAP7_75t_R FILLER_96_486 ();
 FILLER_ASAP7_75t_R FILLER_96_496 ();
 DECAPx10_ASAP7_75t_R FILLER_96_504 ();
 DECAPx6_ASAP7_75t_R FILLER_96_526 ();
 DECAPx10_ASAP7_75t_R FILLER_96_550 ();
 DECAPx4_ASAP7_75t_R FILLER_96_572 ();
 FILLER_ASAP7_75t_R FILLER_96_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_584 ();
 DECAPx2_ASAP7_75t_R FILLER_96_629 ();
 FILLER_ASAP7_75t_R FILLER_96_643 ();
 DECAPx1_ASAP7_75t_R FILLER_96_655 ();
 DECAPx1_ASAP7_75t_R FILLER_96_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_682 ();
 DECAPx4_ASAP7_75t_R FILLER_96_707 ();
 FILLER_ASAP7_75t_R FILLER_96_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_719 ();
 DECAPx10_ASAP7_75t_R FILLER_96_740 ();
 DECAPx2_ASAP7_75t_R FILLER_96_762 ();
 FILLER_ASAP7_75t_R FILLER_96_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_770 ();
 DECAPx6_ASAP7_75t_R FILLER_96_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_837 ();
 DECAPx10_ASAP7_75t_R FILLER_96_858 ();
 DECAPx6_ASAP7_75t_R FILLER_96_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_894 ();
 DECAPx2_ASAP7_75t_R FILLER_96_909 ();
 FILLER_ASAP7_75t_R FILLER_96_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_931 ();
 FILLER_ASAP7_75t_R FILLER_96_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_941 ();
 FILLER_ASAP7_75t_R FILLER_96_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_957 ();
 FILLER_ASAP7_75t_R FILLER_96_964 ();
 DECAPx1_ASAP7_75t_R FILLER_96_972 ();
 DECAPx10_ASAP7_75t_R FILLER_96_984 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1028 ();
 FILLER_ASAP7_75t_R FILLER_96_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1042 ();
 FILLER_ASAP7_75t_R FILLER_96_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1050 ();
 DECAPx6_ASAP7_75t_R FILLER_96_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1120 ();
 FILLER_ASAP7_75t_R FILLER_96_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_96_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1178 ();
 FILLER_ASAP7_75t_R FILLER_96_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1186 ();
 FILLER_ASAP7_75t_R FILLER_96_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1203 ();
 FILLER_ASAP7_75t_R FILLER_96_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_97_2 ();
 DECAPx10_ASAP7_75t_R FILLER_97_24 ();
 DECAPx10_ASAP7_75t_R FILLER_97_46 ();
 DECAPx6_ASAP7_75t_R FILLER_97_68 ();
 FILLER_ASAP7_75t_R FILLER_97_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_96 ();
 DECAPx2_ASAP7_75t_R FILLER_97_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_121 ();
 DECAPx2_ASAP7_75t_R FILLER_97_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_136 ();
 DECAPx10_ASAP7_75t_R FILLER_97_143 ();
 DECAPx1_ASAP7_75t_R FILLER_97_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_169 ();
 DECAPx2_ASAP7_75t_R FILLER_97_184 ();
 DECAPx1_ASAP7_75t_R FILLER_97_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_201 ();
 DECAPx10_ASAP7_75t_R FILLER_97_219 ();
 DECAPx10_ASAP7_75t_R FILLER_97_241 ();
 DECAPx10_ASAP7_75t_R FILLER_97_263 ();
 DECAPx2_ASAP7_75t_R FILLER_97_285 ();
 FILLER_ASAP7_75t_R FILLER_97_291 ();
 DECAPx4_ASAP7_75t_R FILLER_97_303 ();
 DECAPx10_ASAP7_75t_R FILLER_97_319 ();
 DECAPx2_ASAP7_75t_R FILLER_97_341 ();
 FILLER_ASAP7_75t_R FILLER_97_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_423 ();
 DECAPx10_ASAP7_75t_R FILLER_97_430 ();
 DECAPx2_ASAP7_75t_R FILLER_97_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_458 ();
 FILLER_ASAP7_75t_R FILLER_97_481 ();
 DECAPx10_ASAP7_75t_R FILLER_97_511 ();
 DECAPx6_ASAP7_75t_R FILLER_97_533 ();
 FILLER_ASAP7_75t_R FILLER_97_547 ();
 DECAPx4_ASAP7_75t_R FILLER_97_567 ();
 DECAPx2_ASAP7_75t_R FILLER_97_643 ();
 DECAPx2_ASAP7_75t_R FILLER_97_656 ();
 DECAPx2_ASAP7_75t_R FILLER_97_672 ();
 FILLER_ASAP7_75t_R FILLER_97_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_695 ();
 DECAPx2_ASAP7_75t_R FILLER_97_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_708 ();
 DECAPx10_ASAP7_75t_R FILLER_97_733 ();
 DECAPx2_ASAP7_75t_R FILLER_97_755 ();
 DECAPx6_ASAP7_75t_R FILLER_97_803 ();
 DECAPx2_ASAP7_75t_R FILLER_97_839 ();
 FILLER_ASAP7_75t_R FILLER_97_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_847 ();
 DECAPx6_ASAP7_75t_R FILLER_97_870 ();
 DECAPx1_ASAP7_75t_R FILLER_97_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_888 ();
 DECAPx2_ASAP7_75t_R FILLER_97_895 ();
 FILLER_ASAP7_75t_R FILLER_97_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_903 ();
 DECAPx1_ASAP7_75t_R FILLER_97_911 ();
 FILLER_ASAP7_75t_R FILLER_97_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_923 ();
 DECAPx1_ASAP7_75t_R FILLER_97_926 ();
 DECAPx1_ASAP7_75t_R FILLER_97_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_940 ();
 DECAPx6_ASAP7_75t_R FILLER_97_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_963 ();
 DECAPx6_ASAP7_75t_R FILLER_97_982 ();
 DECAPx1_ASAP7_75t_R FILLER_97_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1021 ();
 FILLER_ASAP7_75t_R FILLER_97_1027 ();
 FILLER_ASAP7_75t_R FILLER_97_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1132 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1155 ();
 FILLER_ASAP7_75t_R FILLER_97_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1215 ();
 FILLER_ASAP7_75t_R FILLER_97_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_98_2 ();
 DECAPx10_ASAP7_75t_R FILLER_98_24 ();
 DECAPx10_ASAP7_75t_R FILLER_98_46 ();
 DECAPx6_ASAP7_75t_R FILLER_98_68 ();
 DECAPx1_ASAP7_75t_R FILLER_98_82 ();
 DECAPx6_ASAP7_75t_R FILLER_98_108 ();
 FILLER_ASAP7_75t_R FILLER_98_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_131 ();
 DECAPx4_ASAP7_75t_R FILLER_98_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_153 ();
 FILLER_ASAP7_75t_R FILLER_98_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_209 ();
 DECAPx6_ASAP7_75t_R FILLER_98_216 ();
 DECAPx2_ASAP7_75t_R FILLER_98_230 ();
 DECAPx10_ASAP7_75t_R FILLER_98_264 ();
 FILLER_ASAP7_75t_R FILLER_98_286 ();
 FILLER_ASAP7_75t_R FILLER_98_296 ();
 DECAPx2_ASAP7_75t_R FILLER_98_318 ();
 FILLER_ASAP7_75t_R FILLER_98_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_326 ();
 DECAPx1_ASAP7_75t_R FILLER_98_349 ();
 DECAPx6_ASAP7_75t_R FILLER_98_361 ();
 DECAPx6_ASAP7_75t_R FILLER_98_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_392 ();
 FILLER_ASAP7_75t_R FILLER_98_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_402 ();
 FILLER_ASAP7_75t_R FILLER_98_409 ();
 FILLER_ASAP7_75t_R FILLER_98_423 ();
 DECAPx10_ASAP7_75t_R FILLER_98_431 ();
 DECAPx2_ASAP7_75t_R FILLER_98_453 ();
 FILLER_ASAP7_75t_R FILLER_98_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_461 ();
 DECAPx10_ASAP7_75t_R FILLER_98_464 ();
 DECAPx2_ASAP7_75t_R FILLER_98_486 ();
 FILLER_ASAP7_75t_R FILLER_98_492 ();
 DECAPx6_ASAP7_75t_R FILLER_98_512 ();
 DECAPx2_ASAP7_75t_R FILLER_98_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_532 ();
 DECAPx6_ASAP7_75t_R FILLER_98_543 ();
 FILLER_ASAP7_75t_R FILLER_98_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_578 ();
 DECAPx10_ASAP7_75t_R FILLER_98_585 ();
 DECAPx1_ASAP7_75t_R FILLER_98_607 ();
 FILLER_ASAP7_75t_R FILLER_98_633 ();
 DECAPx2_ASAP7_75t_R FILLER_98_672 ();
 FILLER_ASAP7_75t_R FILLER_98_678 ();
 FILLER_ASAP7_75t_R FILLER_98_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_698 ();
 DECAPx2_ASAP7_75t_R FILLER_98_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_714 ();
 DECAPx6_ASAP7_75t_R FILLER_98_737 ();
 DECAPx1_ASAP7_75t_R FILLER_98_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_755 ();
 DECAPx10_ASAP7_75t_R FILLER_98_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_800 ();
 FILLER_ASAP7_75t_R FILLER_98_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_825 ();
 DECAPx4_ASAP7_75t_R FILLER_98_848 ();
 FILLER_ASAP7_75t_R FILLER_98_858 ();
 FILLER_ASAP7_75t_R FILLER_98_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_884 ();
 DECAPx4_ASAP7_75t_R FILLER_98_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_898 ();
 DECAPx1_ASAP7_75t_R FILLER_98_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_934 ();
 FILLER_ASAP7_75t_R FILLER_98_949 ();
 DECAPx10_ASAP7_75t_R FILLER_98_957 ();
 DECAPx6_ASAP7_75t_R FILLER_98_979 ();
 DECAPx1_ASAP7_75t_R FILLER_98_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_997 ();
 DECAPx4_ASAP7_75t_R FILLER_98_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1029 ();
 FILLER_ASAP7_75t_R FILLER_98_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_98_1044 ();
 FILLER_ASAP7_75t_R FILLER_98_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1124 ();
 FILLER_ASAP7_75t_R FILLER_98_1130 ();
 FILLER_ASAP7_75t_R FILLER_98_1186 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_99_2 ();
 DECAPx10_ASAP7_75t_R FILLER_99_24 ();
 DECAPx10_ASAP7_75t_R FILLER_99_46 ();
 DECAPx10_ASAP7_75t_R FILLER_99_68 ();
 DECAPx10_ASAP7_75t_R FILLER_99_90 ();
 FILLER_ASAP7_75t_R FILLER_99_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_114 ();
 DECAPx4_ASAP7_75t_R FILLER_99_129 ();
 DECAPx10_ASAP7_75t_R FILLER_99_147 ();
 DECAPx6_ASAP7_75t_R FILLER_99_169 ();
 DECAPx2_ASAP7_75t_R FILLER_99_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_189 ();
 FILLER_ASAP7_75t_R FILLER_99_196 ();
 DECAPx10_ASAP7_75t_R FILLER_99_210 ();
 DECAPx10_ASAP7_75t_R FILLER_99_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_254 ();
 DECAPx4_ASAP7_75t_R FILLER_99_277 ();
 DECAPx2_ASAP7_75t_R FILLER_99_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_309 ();
 DECAPx6_ASAP7_75t_R FILLER_99_332 ();
 FILLER_ASAP7_75t_R FILLER_99_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_348 ();
 DECAPx6_ASAP7_75t_R FILLER_99_359 ();
 FILLER_ASAP7_75t_R FILLER_99_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_375 ();
 DECAPx6_ASAP7_75t_R FILLER_99_391 ();
 FILLER_ASAP7_75t_R FILLER_99_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_407 ();
 DECAPx1_ASAP7_75t_R FILLER_99_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_415 ();
 FILLER_ASAP7_75t_R FILLER_99_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_426 ();
 DECAPx10_ASAP7_75t_R FILLER_99_448 ();
 DECAPx10_ASAP7_75t_R FILLER_99_470 ();
 DECAPx4_ASAP7_75t_R FILLER_99_492 ();
 FILLER_ASAP7_75t_R FILLER_99_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_504 ();
 DECAPx2_ASAP7_75t_R FILLER_99_511 ();
 FILLER_ASAP7_75t_R FILLER_99_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_519 ();
 DECAPx10_ASAP7_75t_R FILLER_99_538 ();
 DECAPx6_ASAP7_75t_R FILLER_99_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_574 ();
 DECAPx2_ASAP7_75t_R FILLER_99_586 ();
 FILLER_ASAP7_75t_R FILLER_99_592 ();
 DECAPx2_ASAP7_75t_R FILLER_99_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_622 ();
 DECAPx6_ASAP7_75t_R FILLER_99_645 ();
 FILLER_ASAP7_75t_R FILLER_99_659 ();
 FILLER_ASAP7_75t_R FILLER_99_669 ();
 DECAPx6_ASAP7_75t_R FILLER_99_679 ();
 FILLER_ASAP7_75t_R FILLER_99_693 ();
 FILLER_ASAP7_75t_R FILLER_99_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_711 ();
 DECAPx1_ASAP7_75t_R FILLER_99_721 ();
 DECAPx1_ASAP7_75t_R FILLER_99_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_741 ();
 FILLER_ASAP7_75t_R FILLER_99_748 ();
 DECAPx4_ASAP7_75t_R FILLER_99_790 ();
 DECAPx10_ASAP7_75t_R FILLER_99_822 ();
 DECAPx10_ASAP7_75t_R FILLER_99_844 ();
 DECAPx4_ASAP7_75t_R FILLER_99_866 ();
 FILLER_ASAP7_75t_R FILLER_99_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_878 ();
 DECAPx1_ASAP7_75t_R FILLER_99_903 ();
 FILLER_ASAP7_75t_R FILLER_99_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_923 ();
 FILLER_ASAP7_75t_R FILLER_99_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_948 ();
 FILLER_ASAP7_75t_R FILLER_99_955 ();
 FILLER_ASAP7_75t_R FILLER_99_963 ();
 FILLER_ASAP7_75t_R FILLER_99_972 ();
 DECAPx10_ASAP7_75t_R FILLER_99_980 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1002 ();
 DECAPx4_ASAP7_75t_R FILLER_99_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1057 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1079 ();
 FILLER_ASAP7_75t_R FILLER_99_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1133 ();
 FILLER_ASAP7_75t_R FILLER_99_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1170 ();
 FILLER_ASAP7_75t_R FILLER_99_1176 ();
 DECAPx4_ASAP7_75t_R FILLER_99_1190 ();
 FILLER_ASAP7_75t_R FILLER_99_1200 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1216 ();
 FILLER_ASAP7_75t_R FILLER_99_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_100_2 ();
 DECAPx10_ASAP7_75t_R FILLER_100_24 ();
 DECAPx10_ASAP7_75t_R FILLER_100_46 ();
 DECAPx10_ASAP7_75t_R FILLER_100_68 ();
 DECAPx6_ASAP7_75t_R FILLER_100_90 ();
 DECAPx1_ASAP7_75t_R FILLER_100_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_108 ();
 DECAPx2_ASAP7_75t_R FILLER_100_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_168 ();
 DECAPx6_ASAP7_75t_R FILLER_100_183 ();
 DECAPx10_ASAP7_75t_R FILLER_100_206 ();
 DECAPx10_ASAP7_75t_R FILLER_100_228 ();
 DECAPx10_ASAP7_75t_R FILLER_100_256 ();
 DECAPx1_ASAP7_75t_R FILLER_100_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_282 ();
 FILLER_ASAP7_75t_R FILLER_100_293 ();
 DECAPx6_ASAP7_75t_R FILLER_100_315 ();
 DECAPx4_ASAP7_75t_R FILLER_100_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_367 ();
 DECAPx2_ASAP7_75t_R FILLER_100_384 ();
 DECAPx2_ASAP7_75t_R FILLER_100_403 ();
 FILLER_ASAP7_75t_R FILLER_100_416 ();
 DECAPx1_ASAP7_75t_R FILLER_100_426 ();
 DECAPx1_ASAP7_75t_R FILLER_100_436 ();
 DECAPx10_ASAP7_75t_R FILLER_100_464 ();
 DECAPx1_ASAP7_75t_R FILLER_100_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_490 ();
 DECAPx10_ASAP7_75t_R FILLER_100_513 ();
 FILLER_ASAP7_75t_R FILLER_100_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_537 ();
 DECAPx10_ASAP7_75t_R FILLER_100_548 ();
 DECAPx1_ASAP7_75t_R FILLER_100_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_574 ();
 DECAPx10_ASAP7_75t_R FILLER_100_599 ();
 DECAPx4_ASAP7_75t_R FILLER_100_621 ();
 FILLER_ASAP7_75t_R FILLER_100_631 ();
 DECAPx1_ASAP7_75t_R FILLER_100_666 ();
 DECAPx4_ASAP7_75t_R FILLER_100_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_704 ();
 DECAPx1_ASAP7_75t_R FILLER_100_726 ();
 DECAPx10_ASAP7_75t_R FILLER_100_736 ();
 FILLER_ASAP7_75t_R FILLER_100_758 ();
 DECAPx10_ASAP7_75t_R FILLER_100_780 ();
 DECAPx10_ASAP7_75t_R FILLER_100_802 ();
 FILLER_ASAP7_75t_R FILLER_100_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_826 ();
 DECAPx2_ASAP7_75t_R FILLER_100_889 ();
 DECAPx2_ASAP7_75t_R FILLER_100_917 ();
 FILLER_ASAP7_75t_R FILLER_100_961 ();
 FILLER_ASAP7_75t_R FILLER_100_969 ();
 DECAPx10_ASAP7_75t_R FILLER_100_999 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1021 ();
 FILLER_ASAP7_75t_R FILLER_100_1043 ();
 DECAPx4_ASAP7_75t_R FILLER_100_1065 ();
 FILLER_ASAP7_75t_R FILLER_100_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1103 ();
 FILLER_ASAP7_75t_R FILLER_100_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_101_2 ();
 DECAPx10_ASAP7_75t_R FILLER_101_24 ();
 DECAPx10_ASAP7_75t_R FILLER_101_46 ();
 DECAPx10_ASAP7_75t_R FILLER_101_68 ();
 DECAPx4_ASAP7_75t_R FILLER_101_90 ();
 DECAPx10_ASAP7_75t_R FILLER_101_131 ();
 DECAPx2_ASAP7_75t_R FILLER_101_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_159 ();
 DECAPx6_ASAP7_75t_R FILLER_101_182 ();
 FILLER_ASAP7_75t_R FILLER_101_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_198 ();
 DECAPx4_ASAP7_75t_R FILLER_101_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_229 ();
 DECAPx2_ASAP7_75t_R FILLER_101_274 ();
 FILLER_ASAP7_75t_R FILLER_101_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_282 ();
 DECAPx1_ASAP7_75t_R FILLER_101_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_343 ();
 FILLER_ASAP7_75t_R FILLER_101_359 ();
 DECAPx1_ASAP7_75t_R FILLER_101_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_421 ();
 DECAPx10_ASAP7_75t_R FILLER_101_426 ();
 DECAPx1_ASAP7_75t_R FILLER_101_448 ();
 DECAPx6_ASAP7_75t_R FILLER_101_482 ();
 DECAPx1_ASAP7_75t_R FILLER_101_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_500 ();
 FILLER_ASAP7_75t_R FILLER_101_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_516 ();
 DECAPx10_ASAP7_75t_R FILLER_101_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_620 ();
 DECAPx4_ASAP7_75t_R FILLER_101_643 ();
 FILLER_ASAP7_75t_R FILLER_101_653 ();
 DECAPx1_ASAP7_75t_R FILLER_101_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_669 ();
 DECAPx2_ASAP7_75t_R FILLER_101_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_701 ();
 DECAPx10_ASAP7_75t_R FILLER_101_727 ();
 DECAPx10_ASAP7_75t_R FILLER_101_749 ();
 DECAPx4_ASAP7_75t_R FILLER_101_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_790 ();
 FILLER_ASAP7_75t_R FILLER_101_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_799 ();
 DECAPx10_ASAP7_75t_R FILLER_101_806 ();
 DECAPx1_ASAP7_75t_R FILLER_101_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_832 ();
 DECAPx1_ASAP7_75t_R FILLER_101_845 ();
 DECAPx1_ASAP7_75t_R FILLER_101_861 ();
 DECAPx4_ASAP7_75t_R FILLER_101_883 ();
 FILLER_ASAP7_75t_R FILLER_101_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_901 ();
 FILLER_ASAP7_75t_R FILLER_101_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_917 ();
 FILLER_ASAP7_75t_R FILLER_101_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_970 ();
 DECAPx2_ASAP7_75t_R FILLER_101_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_987 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1038 ();
 FILLER_ASAP7_75t_R FILLER_101_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1183 ();
 FILLER_ASAP7_75t_R FILLER_101_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_102_2 ();
 DECAPx10_ASAP7_75t_R FILLER_102_24 ();
 DECAPx10_ASAP7_75t_R FILLER_102_46 ();
 DECAPx10_ASAP7_75t_R FILLER_102_68 ();
 DECAPx10_ASAP7_75t_R FILLER_102_90 ();
 DECAPx10_ASAP7_75t_R FILLER_102_112 ();
 FILLER_ASAP7_75t_R FILLER_102_134 ();
 DECAPx2_ASAP7_75t_R FILLER_102_142 ();
 DECAPx2_ASAP7_75t_R FILLER_102_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_162 ();
 FILLER_ASAP7_75t_R FILLER_102_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_171 ();
 DECAPx2_ASAP7_75t_R FILLER_102_189 ();
 FILLER_ASAP7_75t_R FILLER_102_195 ();
 DECAPx10_ASAP7_75t_R FILLER_102_219 ();
 DECAPx10_ASAP7_75t_R FILLER_102_241 ();
 DECAPx6_ASAP7_75t_R FILLER_102_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_277 ();
 DECAPx2_ASAP7_75t_R FILLER_102_294 ();
 FILLER_ASAP7_75t_R FILLER_102_300 ();
 DECAPx6_ASAP7_75t_R FILLER_102_320 ();
 DECAPx2_ASAP7_75t_R FILLER_102_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_340 ();
 DECAPx4_ASAP7_75t_R FILLER_102_355 ();
 FILLER_ASAP7_75t_R FILLER_102_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_384 ();
 DECAPx6_ASAP7_75t_R FILLER_102_412 ();
 FILLER_ASAP7_75t_R FILLER_102_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_428 ();
 FILLER_ASAP7_75t_R FILLER_102_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_461 ();
 DECAPx6_ASAP7_75t_R FILLER_102_464 ();
 DECAPx1_ASAP7_75t_R FILLER_102_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_505 ();
 FILLER_ASAP7_75t_R FILLER_102_513 ();
 DECAPx1_ASAP7_75t_R FILLER_102_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_553 ();
 FILLER_ASAP7_75t_R FILLER_102_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_574 ();
 DECAPx10_ASAP7_75t_R FILLER_102_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_618 ();
 DECAPx10_ASAP7_75t_R FILLER_102_649 ();
 FILLER_ASAP7_75t_R FILLER_102_671 ();
 FILLER_ASAP7_75t_R FILLER_102_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_682 ();
 FILLER_ASAP7_75t_R FILLER_102_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_692 ();
 DECAPx6_ASAP7_75t_R FILLER_102_701 ();
 DECAPx1_ASAP7_75t_R FILLER_102_715 ();
 DECAPx10_ASAP7_75t_R FILLER_102_725 ();
 DECAPx6_ASAP7_75t_R FILLER_102_747 ();
 DECAPx2_ASAP7_75t_R FILLER_102_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_767 ();
 DECAPx2_ASAP7_75t_R FILLER_102_775 ();
 FILLER_ASAP7_75t_R FILLER_102_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_790 ();
 FILLER_ASAP7_75t_R FILLER_102_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_807 ();
 DECAPx1_ASAP7_75t_R FILLER_102_832 ();
 DECAPx1_ASAP7_75t_R FILLER_102_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_864 ();
 DECAPx10_ASAP7_75t_R FILLER_102_875 ();
 DECAPx6_ASAP7_75t_R FILLER_102_897 ();
 DECAPx1_ASAP7_75t_R FILLER_102_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_915 ();
 FILLER_ASAP7_75t_R FILLER_102_922 ();
 FILLER_ASAP7_75t_R FILLER_102_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_934 ();
 DECAPx6_ASAP7_75t_R FILLER_102_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_959 ();
 DECAPx10_ASAP7_75t_R FILLER_102_970 ();
 DECAPx4_ASAP7_75t_R FILLER_102_992 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1060 ();
 FILLER_ASAP7_75t_R FILLER_102_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1074 ();
 FILLER_ASAP7_75t_R FILLER_102_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1107 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1114 ();
 FILLER_ASAP7_75t_R FILLER_102_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1130 ();
 FILLER_ASAP7_75t_R FILLER_102_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1199 ();
 FILLER_ASAP7_75t_R FILLER_102_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1207 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_103_2 ();
 DECAPx10_ASAP7_75t_R FILLER_103_24 ();
 DECAPx10_ASAP7_75t_R FILLER_103_46 ();
 DECAPx10_ASAP7_75t_R FILLER_103_68 ();
 DECAPx6_ASAP7_75t_R FILLER_103_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_104 ();
 DECAPx1_ASAP7_75t_R FILLER_103_127 ();
 DECAPx6_ASAP7_75t_R FILLER_103_160 ();
 FILLER_ASAP7_75t_R FILLER_103_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_176 ();
 DECAPx10_ASAP7_75t_R FILLER_103_205 ();
 DECAPx2_ASAP7_75t_R FILLER_103_227 ();
 DECAPx6_ASAP7_75t_R FILLER_103_283 ();
 FILLER_ASAP7_75t_R FILLER_103_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_305 ();
 DECAPx2_ASAP7_75t_R FILLER_103_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_318 ();
 DECAPx4_ASAP7_75t_R FILLER_103_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_337 ();
 DECAPx1_ASAP7_75t_R FILLER_103_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_359 ();
 DECAPx4_ASAP7_75t_R FILLER_103_366 ();
 FILLER_ASAP7_75t_R FILLER_103_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_378 ();
 DECAPx2_ASAP7_75t_R FILLER_103_385 ();
 DECAPx1_ASAP7_75t_R FILLER_103_409 ();
 DECAPx2_ASAP7_75t_R FILLER_103_423 ();
 FILLER_ASAP7_75t_R FILLER_103_436 ();
 DECAPx2_ASAP7_75t_R FILLER_103_441 ();
 FILLER_ASAP7_75t_R FILLER_103_447 ();
 DECAPx10_ASAP7_75t_R FILLER_103_471 ();
 DECAPx2_ASAP7_75t_R FILLER_103_493 ();
 FILLER_ASAP7_75t_R FILLER_103_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_501 ();
 FILLER_ASAP7_75t_R FILLER_103_524 ();
 DECAPx2_ASAP7_75t_R FILLER_103_548 ();
 FILLER_ASAP7_75t_R FILLER_103_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_571 ();
 FILLER_ASAP7_75t_R FILLER_103_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_595 ();
 DECAPx4_ASAP7_75t_R FILLER_103_608 ();
 DECAPx10_ASAP7_75t_R FILLER_103_640 ();
 DECAPx10_ASAP7_75t_R FILLER_103_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_692 ();
 DECAPx2_ASAP7_75t_R FILLER_103_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_719 ();
 DECAPx2_ASAP7_75t_R FILLER_103_734 ();
 FILLER_ASAP7_75t_R FILLER_103_740 ();
 FILLER_ASAP7_75t_R FILLER_103_790 ();
 DECAPx6_ASAP7_75t_R FILLER_103_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_836 ();
 DECAPx4_ASAP7_75t_R FILLER_103_843 ();
 FILLER_ASAP7_75t_R FILLER_103_859 ();
 DECAPx6_ASAP7_75t_R FILLER_103_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_881 ();
 DECAPx6_ASAP7_75t_R FILLER_103_908 ();
 FILLER_ASAP7_75t_R FILLER_103_922 ();
 DECAPx10_ASAP7_75t_R FILLER_103_926 ();
 DECAPx2_ASAP7_75t_R FILLER_103_948 ();
 FILLER_ASAP7_75t_R FILLER_103_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_956 ();
 DECAPx4_ASAP7_75t_R FILLER_103_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1022 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1057 ();
 FILLER_ASAP7_75t_R FILLER_103_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1081 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1104 ();
 FILLER_ASAP7_75t_R FILLER_103_1118 ();
 DECAPx4_ASAP7_75t_R FILLER_103_1142 ();
 FILLER_ASAP7_75t_R FILLER_103_1152 ();
 DECAPx4_ASAP7_75t_R FILLER_103_1160 ();
 FILLER_ASAP7_75t_R FILLER_103_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1216 ();
 FILLER_ASAP7_75t_R FILLER_103_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_104_2 ();
 DECAPx10_ASAP7_75t_R FILLER_104_24 ();
 DECAPx10_ASAP7_75t_R FILLER_104_46 ();
 DECAPx10_ASAP7_75t_R FILLER_104_68 ();
 DECAPx10_ASAP7_75t_R FILLER_104_90 ();
 DECAPx2_ASAP7_75t_R FILLER_104_112 ();
 DECAPx2_ASAP7_75t_R FILLER_104_135 ();
 FILLER_ASAP7_75t_R FILLER_104_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_143 ();
 FILLER_ASAP7_75t_R FILLER_104_179 ();
 DECAPx6_ASAP7_75t_R FILLER_104_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_201 ();
 DECAPx10_ASAP7_75t_R FILLER_104_224 ();
 DECAPx2_ASAP7_75t_R FILLER_104_246 ();
 FILLER_ASAP7_75t_R FILLER_104_258 ();
 DECAPx6_ASAP7_75t_R FILLER_104_266 ();
 DECAPx1_ASAP7_75t_R FILLER_104_280 ();
 DECAPx1_ASAP7_75t_R FILLER_104_308 ();
 FILLER_ASAP7_75t_R FILLER_104_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_341 ();
 DECAPx6_ASAP7_75t_R FILLER_104_348 ();
 DECAPx2_ASAP7_75t_R FILLER_104_362 ();
 DECAPx1_ASAP7_75t_R FILLER_104_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_379 ();
 FILLER_ASAP7_75t_R FILLER_104_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_393 ();
 FILLER_ASAP7_75t_R FILLER_104_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_425 ();
 DECAPx6_ASAP7_75t_R FILLER_104_448 ();
 FILLER_ASAP7_75t_R FILLER_104_464 ();
 DECAPx10_ASAP7_75t_R FILLER_104_476 ();
 FILLER_ASAP7_75t_R FILLER_104_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_514 ();
 DECAPx10_ASAP7_75t_R FILLER_104_537 ();
 FILLER_ASAP7_75t_R FILLER_104_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_571 ();
 DECAPx1_ASAP7_75t_R FILLER_104_590 ();
 DECAPx2_ASAP7_75t_R FILLER_104_600 ();
 FILLER_ASAP7_75t_R FILLER_104_606 ();
 DECAPx1_ASAP7_75t_R FILLER_104_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_628 ();
 FILLER_ASAP7_75t_R FILLER_104_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_653 ();
 DECAPx4_ASAP7_75t_R FILLER_104_674 ();
 DECAPx2_ASAP7_75t_R FILLER_104_693 ();
 FILLER_ASAP7_75t_R FILLER_104_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_701 ();
 DECAPx10_ASAP7_75t_R FILLER_104_708 ();
 DECAPx4_ASAP7_75t_R FILLER_104_730 ();
 FILLER_ASAP7_75t_R FILLER_104_740 ();
 FILLER_ASAP7_75t_R FILLER_104_752 ();
 FILLER_ASAP7_75t_R FILLER_104_766 ();
 FILLER_ASAP7_75t_R FILLER_104_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_776 ();
 FILLER_ASAP7_75t_R FILLER_104_787 ();
 FILLER_ASAP7_75t_R FILLER_104_797 ();
 DECAPx1_ASAP7_75t_R FILLER_104_805 ();
 FILLER_ASAP7_75t_R FILLER_104_815 ();
 DECAPx1_ASAP7_75t_R FILLER_104_823 ();
 FILLER_ASAP7_75t_R FILLER_104_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_835 ();
 DECAPx2_ASAP7_75t_R FILLER_104_842 ();
 FILLER_ASAP7_75t_R FILLER_104_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_857 ();
 DECAPx2_ASAP7_75t_R FILLER_104_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_876 ();
 DECAPx10_ASAP7_75t_R FILLER_104_895 ();
 DECAPx6_ASAP7_75t_R FILLER_104_917 ();
 DECAPx1_ASAP7_75t_R FILLER_104_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_935 ();
 DECAPx10_ASAP7_75t_R FILLER_104_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_976 ();
 DECAPx4_ASAP7_75t_R FILLER_104_983 ();
 FILLER_ASAP7_75t_R FILLER_104_993 ();
 FILLER_ASAP7_75t_R FILLER_104_1001 ();
 FILLER_ASAP7_75t_R FILLER_104_1025 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1055 ();
 DECAPx4_ASAP7_75t_R FILLER_104_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1086 ();
 FILLER_ASAP7_75t_R FILLER_104_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1150 ();
 FILLER_ASAP7_75t_R FILLER_104_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_105_2 ();
 DECAPx10_ASAP7_75t_R FILLER_105_24 ();
 DECAPx10_ASAP7_75t_R FILLER_105_46 ();
 DECAPx10_ASAP7_75t_R FILLER_105_68 ();
 DECAPx10_ASAP7_75t_R FILLER_105_90 ();
 DECAPx4_ASAP7_75t_R FILLER_105_112 ();
 FILLER_ASAP7_75t_R FILLER_105_122 ();
 DECAPx6_ASAP7_75t_R FILLER_105_130 ();
 DECAPx2_ASAP7_75t_R FILLER_105_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_185 ();
 DECAPx10_ASAP7_75t_R FILLER_105_211 ();
 DECAPx1_ASAP7_75t_R FILLER_105_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_237 ();
 DECAPx2_ASAP7_75t_R FILLER_105_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_288 ();
 DECAPx2_ASAP7_75t_R FILLER_105_313 ();
 DECAPx2_ASAP7_75t_R FILLER_105_325 ();
 DECAPx2_ASAP7_75t_R FILLER_105_339 ();
 FILLER_ASAP7_75t_R FILLER_105_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_347 ();
 DECAPx2_ASAP7_75t_R FILLER_105_356 ();
 FILLER_ASAP7_75t_R FILLER_105_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_380 ();
 DECAPx2_ASAP7_75t_R FILLER_105_389 ();
 FILLER_ASAP7_75t_R FILLER_105_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_397 ();
 DECAPx10_ASAP7_75t_R FILLER_105_405 ();
 DECAPx1_ASAP7_75t_R FILLER_105_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_431 ();
 DECAPx10_ASAP7_75t_R FILLER_105_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_461 ();
 DECAPx6_ASAP7_75t_R FILLER_105_482 ();
 DECAPx1_ASAP7_75t_R FILLER_105_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_537 ();
 FILLER_ASAP7_75t_R FILLER_105_550 ();
 FILLER_ASAP7_75t_R FILLER_105_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_562 ();
 DECAPx1_ASAP7_75t_R FILLER_105_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_573 ();
 DECAPx6_ASAP7_75t_R FILLER_105_580 ();
 DECAPx2_ASAP7_75t_R FILLER_105_594 ();
 DECAPx4_ASAP7_75t_R FILLER_105_630 ();
 DECAPx1_ASAP7_75t_R FILLER_105_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_666 ();
 DECAPx6_ASAP7_75t_R FILLER_105_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_701 ();
 DECAPx1_ASAP7_75t_R FILLER_105_712 ();
 DECAPx6_ASAP7_75t_R FILLER_105_740 ();
 DECAPx1_ASAP7_75t_R FILLER_105_754 ();
 DECAPx1_ASAP7_75t_R FILLER_105_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_769 ();
 FILLER_ASAP7_75t_R FILLER_105_790 ();
 DECAPx2_ASAP7_75t_R FILLER_105_804 ();
 FILLER_ASAP7_75t_R FILLER_105_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_863 ();
 DECAPx2_ASAP7_75t_R FILLER_105_870 ();
 FILLER_ASAP7_75t_R FILLER_105_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_878 ();
 FILLER_ASAP7_75t_R FILLER_105_897 ();
 DECAPx1_ASAP7_75t_R FILLER_105_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_923 ();
 DECAPx10_ASAP7_75t_R FILLER_105_926 ();
 DECAPx6_ASAP7_75t_R FILLER_105_948 ();
 FILLER_ASAP7_75t_R FILLER_105_962 ();
 DECAPx2_ASAP7_75t_R FILLER_105_982 ();
 FILLER_ASAP7_75t_R FILLER_105_988 ();
 FILLER_ASAP7_75t_R FILLER_105_993 ();
 FILLER_ASAP7_75t_R FILLER_105_998 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1009 ();
 FILLER_ASAP7_75t_R FILLER_105_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1033 ();
 FILLER_ASAP7_75t_R FILLER_105_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1087 ();
 FILLER_ASAP7_75t_R FILLER_105_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1121 ();
 FILLER_ASAP7_75t_R FILLER_105_1135 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1154 ();
 FILLER_ASAP7_75t_R FILLER_105_1164 ();
 DECAPx6_ASAP7_75t_R FILLER_105_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1193 ();
 FILLER_ASAP7_75t_R FILLER_105_1208 ();
 FILLER_ASAP7_75t_R FILLER_105_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_106_2 ();
 DECAPx10_ASAP7_75t_R FILLER_106_24 ();
 DECAPx10_ASAP7_75t_R FILLER_106_46 ();
 DECAPx10_ASAP7_75t_R FILLER_106_68 ();
 DECAPx10_ASAP7_75t_R FILLER_106_90 ();
 DECAPx2_ASAP7_75t_R FILLER_106_112 ();
 DECAPx1_ASAP7_75t_R FILLER_106_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_133 ();
 DECAPx6_ASAP7_75t_R FILLER_106_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_158 ();
 DECAPx1_ASAP7_75t_R FILLER_106_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_175 ();
 DECAPx10_ASAP7_75t_R FILLER_106_183 ();
 DECAPx10_ASAP7_75t_R FILLER_106_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_227 ();
 DECAPx4_ASAP7_75t_R FILLER_106_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_282 ();
 DECAPx6_ASAP7_75t_R FILLER_106_313 ();
 DECAPx2_ASAP7_75t_R FILLER_106_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_343 ();
 DECAPx2_ASAP7_75t_R FILLER_106_354 ();
 FILLER_ASAP7_75t_R FILLER_106_360 ();
 DECAPx4_ASAP7_75t_R FILLER_106_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_394 ();
 DECAPx2_ASAP7_75t_R FILLER_106_418 ();
 FILLER_ASAP7_75t_R FILLER_106_424 ();
 DECAPx10_ASAP7_75t_R FILLER_106_432 ();
 DECAPx2_ASAP7_75t_R FILLER_106_454 ();
 FILLER_ASAP7_75t_R FILLER_106_460 ();
 FILLER_ASAP7_75t_R FILLER_106_464 ();
 DECAPx10_ASAP7_75t_R FILLER_106_469 ();
 DECAPx4_ASAP7_75t_R FILLER_106_491 ();
 FILLER_ASAP7_75t_R FILLER_106_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_503 ();
 DECAPx10_ASAP7_75t_R FILLER_106_526 ();
 DECAPx6_ASAP7_75t_R FILLER_106_548 ();
 DECAPx1_ASAP7_75t_R FILLER_106_562 ();
 DECAPx2_ASAP7_75t_R FILLER_106_572 ();
 FILLER_ASAP7_75t_R FILLER_106_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_580 ();
 DECAPx10_ASAP7_75t_R FILLER_106_594 ();
 DECAPx10_ASAP7_75t_R FILLER_106_616 ();
 DECAPx10_ASAP7_75t_R FILLER_106_638 ();
 DECAPx4_ASAP7_75t_R FILLER_106_660 ();
 DECAPx6_ASAP7_75t_R FILLER_106_692 ();
 DECAPx2_ASAP7_75t_R FILLER_106_706 ();
 DECAPx6_ASAP7_75t_R FILLER_106_732 ();
 DECAPx1_ASAP7_75t_R FILLER_106_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_750 ();
 DECAPx10_ASAP7_75t_R FILLER_106_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_793 ();
 DECAPx4_ASAP7_75t_R FILLER_106_800 ();
 FILLER_ASAP7_75t_R FILLER_106_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_819 ();
 DECAPx2_ASAP7_75t_R FILLER_106_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_844 ();
 DECAPx4_ASAP7_75t_R FILLER_106_869 ();
 FILLER_ASAP7_75t_R FILLER_106_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_881 ();
 FILLER_ASAP7_75t_R FILLER_106_886 ();
 DECAPx2_ASAP7_75t_R FILLER_106_908 ();
 FILLER_ASAP7_75t_R FILLER_106_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_916 ();
 DECAPx6_ASAP7_75t_R FILLER_106_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_963 ();
 DECAPx1_ASAP7_75t_R FILLER_106_982 ();
 DECAPx1_ASAP7_75t_R FILLER_106_995 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_106_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1085 ();
 DECAPx4_ASAP7_75t_R FILLER_106_1092 ();
 FILLER_ASAP7_75t_R FILLER_106_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1111 ();
 FILLER_ASAP7_75t_R FILLER_106_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1146 ();
 FILLER_ASAP7_75t_R FILLER_106_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1171 ();
 DECAPx4_ASAP7_75t_R FILLER_106_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1209 ();
 FILLER_ASAP7_75t_R FILLER_106_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_107_2 ();
 DECAPx10_ASAP7_75t_R FILLER_107_24 ();
 DECAPx10_ASAP7_75t_R FILLER_107_46 ();
 DECAPx10_ASAP7_75t_R FILLER_107_68 ();
 DECAPx10_ASAP7_75t_R FILLER_107_90 ();
 DECAPx1_ASAP7_75t_R FILLER_107_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_116 ();
 DECAPx4_ASAP7_75t_R FILLER_107_167 ();
 FILLER_ASAP7_75t_R FILLER_107_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_196 ();
 DECAPx10_ASAP7_75t_R FILLER_107_225 ();
 DECAPx10_ASAP7_75t_R FILLER_107_247 ();
 DECAPx6_ASAP7_75t_R FILLER_107_269 ();
 DECAPx6_ASAP7_75t_R FILLER_107_289 ();
 DECAPx1_ASAP7_75t_R FILLER_107_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_307 ();
 DECAPx1_ASAP7_75t_R FILLER_107_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_324 ();
 FILLER_ASAP7_75t_R FILLER_107_331 ();
 DECAPx1_ASAP7_75t_R FILLER_107_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_349 ();
 DECAPx6_ASAP7_75t_R FILLER_107_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_370 ();
 DECAPx4_ASAP7_75t_R FILLER_107_389 ();
 DECAPx1_ASAP7_75t_R FILLER_107_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_431 ();
 DECAPx10_ASAP7_75t_R FILLER_107_478 ();
 DECAPx2_ASAP7_75t_R FILLER_107_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_506 ();
 FILLER_ASAP7_75t_R FILLER_107_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_516 ();
 DECAPx4_ASAP7_75t_R FILLER_107_539 ();
 FILLER_ASAP7_75t_R FILLER_107_549 ();
 DECAPx1_ASAP7_75t_R FILLER_107_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_563 ();
 DECAPx1_ASAP7_75t_R FILLER_107_573 ();
 DECAPx2_ASAP7_75t_R FILLER_107_594 ();
 DECAPx6_ASAP7_75t_R FILLER_107_624 ();
 DECAPx1_ASAP7_75t_R FILLER_107_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_642 ();
 FILLER_ASAP7_75t_R FILLER_107_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_698 ();
 DECAPx6_ASAP7_75t_R FILLER_107_717 ();
 DECAPx1_ASAP7_75t_R FILLER_107_731 ();
 DECAPx2_ASAP7_75t_R FILLER_107_752 ();
 DECAPx6_ASAP7_75t_R FILLER_107_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_786 ();
 DECAPx10_ASAP7_75t_R FILLER_107_801 ();
 DECAPx2_ASAP7_75t_R FILLER_107_823 ();
 FILLER_ASAP7_75t_R FILLER_107_829 ();
 DECAPx10_ASAP7_75t_R FILLER_107_870 ();
 DECAPx10_ASAP7_75t_R FILLER_107_892 ();
 DECAPx4_ASAP7_75t_R FILLER_107_914 ();
 DECAPx2_ASAP7_75t_R FILLER_107_926 ();
 FILLER_ASAP7_75t_R FILLER_107_932 ();
 DECAPx2_ASAP7_75t_R FILLER_107_944 ();
 DECAPx4_ASAP7_75t_R FILLER_107_968 ();
 FILLER_ASAP7_75t_R FILLER_107_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_980 ();
 FILLER_ASAP7_75t_R FILLER_107_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_107_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1085 ();
 FILLER_ASAP7_75t_R FILLER_107_1094 ();
 DECAPx1_ASAP7_75t_R FILLER_107_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1124 ();
 FILLER_ASAP7_75t_R FILLER_107_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1189 ();
 FILLER_ASAP7_75t_R FILLER_107_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_108_2 ();
 DECAPx10_ASAP7_75t_R FILLER_108_24 ();
 DECAPx10_ASAP7_75t_R FILLER_108_46 ();
 DECAPx10_ASAP7_75t_R FILLER_108_68 ();
 DECAPx10_ASAP7_75t_R FILLER_108_90 ();
 DECAPx4_ASAP7_75t_R FILLER_108_112 ();
 FILLER_ASAP7_75t_R FILLER_108_122 ();
 DECAPx10_ASAP7_75t_R FILLER_108_130 ();
 DECAPx2_ASAP7_75t_R FILLER_108_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_158 ();
 DECAPx6_ASAP7_75t_R FILLER_108_165 ();
 DECAPx2_ASAP7_75t_R FILLER_108_179 ();
 DECAPx10_ASAP7_75t_R FILLER_108_196 ();
 DECAPx10_ASAP7_75t_R FILLER_108_218 ();
 DECAPx2_ASAP7_75t_R FILLER_108_240 ();
 FILLER_ASAP7_75t_R FILLER_108_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_248 ();
 FILLER_ASAP7_75t_R FILLER_108_271 ();
 DECAPx10_ASAP7_75t_R FILLER_108_279 ();
 DECAPx6_ASAP7_75t_R FILLER_108_301 ();
 DECAPx10_ASAP7_75t_R FILLER_108_321 ();
 DECAPx2_ASAP7_75t_R FILLER_108_343 ();
 DECAPx1_ASAP7_75t_R FILLER_108_368 ();
 FILLER_ASAP7_75t_R FILLER_108_382 ();
 DECAPx6_ASAP7_75t_R FILLER_108_396 ();
 DECAPx4_ASAP7_75t_R FILLER_108_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_423 ();
 FILLER_ASAP7_75t_R FILLER_108_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_461 ();
 DECAPx6_ASAP7_75t_R FILLER_108_464 ();
 DECAPx1_ASAP7_75t_R FILLER_108_478 ();
 DECAPx1_ASAP7_75t_R FILLER_108_504 ();
 FILLER_ASAP7_75t_R FILLER_108_515 ();
 FILLER_ASAP7_75t_R FILLER_108_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_583 ();
 DECAPx4_ASAP7_75t_R FILLER_108_590 ();
 DECAPx1_ASAP7_75t_R FILLER_108_610 ();
 DECAPx10_ASAP7_75t_R FILLER_108_670 ();
 DECAPx10_ASAP7_75t_R FILLER_108_692 ();
 DECAPx10_ASAP7_75t_R FILLER_108_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_736 ();
 DECAPx2_ASAP7_75t_R FILLER_108_745 ();
 FILLER_ASAP7_75t_R FILLER_108_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_771 ();
 DECAPx4_ASAP7_75t_R FILLER_108_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_799 ();
 DECAPx4_ASAP7_75t_R FILLER_108_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_816 ();
 FILLER_ASAP7_75t_R FILLER_108_823 ();
 DECAPx1_ASAP7_75t_R FILLER_108_831 ();
 FILLER_ASAP7_75t_R FILLER_108_841 ();
 DECAPx1_ASAP7_75t_R FILLER_108_849 ();
 DECAPx4_ASAP7_75t_R FILLER_108_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_877 ();
 DECAPx10_ASAP7_75t_R FILLER_108_924 ();
 DECAPx6_ASAP7_75t_R FILLER_108_946 ();
 FILLER_ASAP7_75t_R FILLER_108_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1043 ();
 FILLER_ASAP7_75t_R FILLER_108_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1119 ();
 FILLER_ASAP7_75t_R FILLER_108_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_109_2 ();
 DECAPx10_ASAP7_75t_R FILLER_109_24 ();
 DECAPx10_ASAP7_75t_R FILLER_109_46 ();
 DECAPx10_ASAP7_75t_R FILLER_109_68 ();
 DECAPx10_ASAP7_75t_R FILLER_109_90 ();
 DECAPx10_ASAP7_75t_R FILLER_109_112 ();
 DECAPx4_ASAP7_75t_R FILLER_109_134 ();
 FILLER_ASAP7_75t_R FILLER_109_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_146 ();
 FILLER_ASAP7_75t_R FILLER_109_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_187 ();
 DECAPx2_ASAP7_75t_R FILLER_109_218 ();
 FILLER_ASAP7_75t_R FILLER_109_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_226 ();
 DECAPx6_ASAP7_75t_R FILLER_109_253 ();
 DECAPx2_ASAP7_75t_R FILLER_109_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_273 ();
 FILLER_ASAP7_75t_R FILLER_109_280 ();
 DECAPx4_ASAP7_75t_R FILLER_109_301 ();
 FILLER_ASAP7_75t_R FILLER_109_311 ();
 DECAPx2_ASAP7_75t_R FILLER_109_321 ();
 DECAPx10_ASAP7_75t_R FILLER_109_343 ();
 DECAPx6_ASAP7_75t_R FILLER_109_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_379 ();
 DECAPx1_ASAP7_75t_R FILLER_109_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_411 ();
 DECAPx6_ASAP7_75t_R FILLER_109_425 ();
 DECAPx2_ASAP7_75t_R FILLER_109_439 ();
 DECAPx2_ASAP7_75t_R FILLER_109_473 ();
 FILLER_ASAP7_75t_R FILLER_109_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_481 ();
 DECAPx10_ASAP7_75t_R FILLER_109_510 ();
 DECAPx1_ASAP7_75t_R FILLER_109_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_536 ();
 DECAPx10_ASAP7_75t_R FILLER_109_549 ();
 DECAPx6_ASAP7_75t_R FILLER_109_571 ();
 DECAPx2_ASAP7_75t_R FILLER_109_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_622 ();
 DECAPx10_ASAP7_75t_R FILLER_109_636 ();
 DECAPx10_ASAP7_75t_R FILLER_109_658 ();
 DECAPx2_ASAP7_75t_R FILLER_109_702 ();
 DECAPx6_ASAP7_75t_R FILLER_109_718 ();
 FILLER_ASAP7_75t_R FILLER_109_732 ();
 FILLER_ASAP7_75t_R FILLER_109_764 ();
 DECAPx6_ASAP7_75t_R FILLER_109_773 ();
 DECAPx1_ASAP7_75t_R FILLER_109_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_791 ();
 DECAPx2_ASAP7_75t_R FILLER_109_808 ();
 FILLER_ASAP7_75t_R FILLER_109_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_816 ();
 FILLER_ASAP7_75t_R FILLER_109_823 ();
 FILLER_ASAP7_75t_R FILLER_109_833 ();
 DECAPx1_ASAP7_75t_R FILLER_109_841 ();
 FILLER_ASAP7_75t_R FILLER_109_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_853 ();
 DECAPx1_ASAP7_75t_R FILLER_109_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_872 ();
 FILLER_ASAP7_75t_R FILLER_109_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_897 ();
 DECAPx1_ASAP7_75t_R FILLER_109_920 ();
 DECAPx6_ASAP7_75t_R FILLER_109_926 ();
 FILLER_ASAP7_75t_R FILLER_109_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_942 ();
 DECAPx1_ASAP7_75t_R FILLER_109_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_965 ();
 DECAPx6_ASAP7_75t_R FILLER_109_984 ();
 DECAPx1_ASAP7_75t_R FILLER_109_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1070 ();
 FILLER_ASAP7_75t_R FILLER_109_1084 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1155 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1172 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_110_2 ();
 DECAPx10_ASAP7_75t_R FILLER_110_24 ();
 DECAPx10_ASAP7_75t_R FILLER_110_46 ();
 DECAPx10_ASAP7_75t_R FILLER_110_68 ();
 DECAPx10_ASAP7_75t_R FILLER_110_90 ();
 DECAPx10_ASAP7_75t_R FILLER_110_112 ();
 DECAPx4_ASAP7_75t_R FILLER_110_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_144 ();
 DECAPx1_ASAP7_75t_R FILLER_110_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_171 ();
 DECAPx6_ASAP7_75t_R FILLER_110_200 ();
 DECAPx2_ASAP7_75t_R FILLER_110_214 ();
 FILLER_ASAP7_75t_R FILLER_110_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_266 ();
 DECAPx1_ASAP7_75t_R FILLER_110_281 ();
 DECAPx4_ASAP7_75t_R FILLER_110_304 ();
 FILLER_ASAP7_75t_R FILLER_110_314 ();
 DECAPx2_ASAP7_75t_R FILLER_110_322 ();
 DECAPx6_ASAP7_75t_R FILLER_110_347 ();
 FILLER_ASAP7_75t_R FILLER_110_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_363 ();
 DECAPx10_ASAP7_75t_R FILLER_110_382 ();
 FILLER_ASAP7_75t_R FILLER_110_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_419 ();
 DECAPx10_ASAP7_75t_R FILLER_110_464 ();
 DECAPx6_ASAP7_75t_R FILLER_110_486 ();
 FILLER_ASAP7_75t_R FILLER_110_500 ();
 DECAPx6_ASAP7_75t_R FILLER_110_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_542 ();
 DECAPx2_ASAP7_75t_R FILLER_110_575 ();
 FILLER_ASAP7_75t_R FILLER_110_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_583 ();
 DECAPx10_ASAP7_75t_R FILLER_110_587 ();
 DECAPx4_ASAP7_75t_R FILLER_110_612 ();
 FILLER_ASAP7_75t_R FILLER_110_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_624 ();
 DECAPx10_ASAP7_75t_R FILLER_110_631 ();
 DECAPx6_ASAP7_75t_R FILLER_110_653 ();
 DECAPx2_ASAP7_75t_R FILLER_110_667 ();
 FILLER_ASAP7_75t_R FILLER_110_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_730 ();
 DECAPx1_ASAP7_75t_R FILLER_110_746 ();
 DECAPx6_ASAP7_75t_R FILLER_110_764 ();
 DECAPx1_ASAP7_75t_R FILLER_110_778 ();
 DECAPx1_ASAP7_75t_R FILLER_110_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_814 ();
 DECAPx2_ASAP7_75t_R FILLER_110_829 ();
 DECAPx2_ASAP7_75t_R FILLER_110_851 ();
 DECAPx10_ASAP7_75t_R FILLER_110_863 ();
 DECAPx10_ASAP7_75t_R FILLER_110_885 ();
 DECAPx10_ASAP7_75t_R FILLER_110_907 ();
 DECAPx10_ASAP7_75t_R FILLER_110_929 ();
 DECAPx2_ASAP7_75t_R FILLER_110_951 ();
 FILLER_ASAP7_75t_R FILLER_110_957 ();
 DECAPx10_ASAP7_75t_R FILLER_110_977 ();
 FILLER_ASAP7_75t_R FILLER_110_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1078 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1121 ();
 FILLER_ASAP7_75t_R FILLER_110_1135 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1187 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1197 ();
 FILLER_ASAP7_75t_R FILLER_110_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_111_2 ();
 DECAPx10_ASAP7_75t_R FILLER_111_24 ();
 DECAPx10_ASAP7_75t_R FILLER_111_46 ();
 DECAPx10_ASAP7_75t_R FILLER_111_68 ();
 DECAPx4_ASAP7_75t_R FILLER_111_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_100 ();
 DECAPx10_ASAP7_75t_R FILLER_111_107 ();
 DECAPx10_ASAP7_75t_R FILLER_111_129 ();
 DECAPx1_ASAP7_75t_R FILLER_111_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_155 ();
 DECAPx4_ASAP7_75t_R FILLER_111_162 ();
 FILLER_ASAP7_75t_R FILLER_111_172 ();
 DECAPx10_ASAP7_75t_R FILLER_111_184 ();
 DECAPx4_ASAP7_75t_R FILLER_111_206 ();
 FILLER_ASAP7_75t_R FILLER_111_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_218 ();
 DECAPx6_ASAP7_75t_R FILLER_111_253 ();
 DECAPx10_ASAP7_75t_R FILLER_111_281 ();
 DECAPx2_ASAP7_75t_R FILLER_111_303 ();
 DECAPx6_ASAP7_75t_R FILLER_111_315 ();
 DECAPx1_ASAP7_75t_R FILLER_111_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_339 ();
 DECAPx1_ASAP7_75t_R FILLER_111_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_366 ();
 FILLER_ASAP7_75t_R FILLER_111_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_386 ();
 DECAPx10_ASAP7_75t_R FILLER_111_410 ();
 DECAPx10_ASAP7_75t_R FILLER_111_432 ();
 FILLER_ASAP7_75t_R FILLER_111_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_456 ();
 DECAPx10_ASAP7_75t_R FILLER_111_465 ();
 DECAPx6_ASAP7_75t_R FILLER_111_487 ();
 DECAPx2_ASAP7_75t_R FILLER_111_501 ();
 DECAPx1_ASAP7_75t_R FILLER_111_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_517 ();
 DECAPx10_ASAP7_75t_R FILLER_111_528 ();
 DECAPx10_ASAP7_75t_R FILLER_111_550 ();
 DECAPx1_ASAP7_75t_R FILLER_111_578 ();
 FILLER_ASAP7_75t_R FILLER_111_588 ();
 DECAPx2_ASAP7_75t_R FILLER_111_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_619 ();
 DECAPx10_ASAP7_75t_R FILLER_111_626 ();
 FILLER_ASAP7_75t_R FILLER_111_648 ();
 DECAPx6_ASAP7_75t_R FILLER_111_672 ();
 FILLER_ASAP7_75t_R FILLER_111_686 ();
 DECAPx6_ASAP7_75t_R FILLER_111_706 ();
 DECAPx1_ASAP7_75t_R FILLER_111_720 ();
 FILLER_ASAP7_75t_R FILLER_111_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_751 ();
 FILLER_ASAP7_75t_R FILLER_111_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_760 ();
 DECAPx4_ASAP7_75t_R FILLER_111_775 ();
 FILLER_ASAP7_75t_R FILLER_111_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_787 ();
 DECAPx2_ASAP7_75t_R FILLER_111_804 ();
 FILLER_ASAP7_75t_R FILLER_111_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_823 ();
 DECAPx6_ASAP7_75t_R FILLER_111_830 ();
 FILLER_ASAP7_75t_R FILLER_111_844 ();
 FILLER_ASAP7_75t_R FILLER_111_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_854 ();
 DECAPx6_ASAP7_75t_R FILLER_111_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_875 ();
 DECAPx1_ASAP7_75t_R FILLER_111_880 ();
 DECAPx6_ASAP7_75t_R FILLER_111_904 ();
 DECAPx2_ASAP7_75t_R FILLER_111_918 ();
 DECAPx6_ASAP7_75t_R FILLER_111_926 ();
 DECAPx1_ASAP7_75t_R FILLER_111_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_944 ();
 DECAPx6_ASAP7_75t_R FILLER_111_981 ();
 DECAPx1_ASAP7_75t_R FILLER_111_995 ();
 FILLER_ASAP7_75t_R FILLER_111_1011 ();
 DECAPx4_ASAP7_75t_R FILLER_111_1019 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1042 ();
 FILLER_ASAP7_75t_R FILLER_111_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1058 ();
 FILLER_ASAP7_75t_R FILLER_111_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1067 ();
 FILLER_ASAP7_75t_R FILLER_111_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1081 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1123 ();
 FILLER_ASAP7_75t_R FILLER_111_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1144 ();
 DECAPx4_ASAP7_75t_R FILLER_111_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1166 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_112_2 ();
 DECAPx10_ASAP7_75t_R FILLER_112_24 ();
 DECAPx10_ASAP7_75t_R FILLER_112_46 ();
 DECAPx10_ASAP7_75t_R FILLER_112_68 ();
 DECAPx2_ASAP7_75t_R FILLER_112_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_96 ();
 DECAPx1_ASAP7_75t_R FILLER_112_119 ();
 DECAPx10_ASAP7_75t_R FILLER_112_145 ();
 DECAPx6_ASAP7_75t_R FILLER_112_167 ();
 DECAPx2_ASAP7_75t_R FILLER_112_181 ();
 FILLER_ASAP7_75t_R FILLER_112_207 ();
 FILLER_ASAP7_75t_R FILLER_112_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_241 ();
 DECAPx4_ASAP7_75t_R FILLER_112_264 ();
 FILLER_ASAP7_75t_R FILLER_112_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_276 ();
 FILLER_ASAP7_75t_R FILLER_112_283 ();
 DECAPx1_ASAP7_75t_R FILLER_112_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_308 ();
 DECAPx2_ASAP7_75t_R FILLER_112_322 ();
 FILLER_ASAP7_75t_R FILLER_112_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_330 ();
 DECAPx1_ASAP7_75t_R FILLER_112_343 ();
 DECAPx6_ASAP7_75t_R FILLER_112_353 ();
 DECAPx2_ASAP7_75t_R FILLER_112_367 ();
 FILLER_ASAP7_75t_R FILLER_112_386 ();
 DECAPx4_ASAP7_75t_R FILLER_112_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_411 ();
 DECAPx10_ASAP7_75t_R FILLER_112_434 ();
 DECAPx10_ASAP7_75t_R FILLER_112_464 ();
 DECAPx2_ASAP7_75t_R FILLER_112_486 ();
 DECAPx6_ASAP7_75t_R FILLER_112_547 ();
 FILLER_ASAP7_75t_R FILLER_112_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_563 ();
 DECAPx2_ASAP7_75t_R FILLER_112_573 ();
 FILLER_ASAP7_75t_R FILLER_112_579 ();
 FILLER_ASAP7_75t_R FILLER_112_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_599 ();
 DECAPx1_ASAP7_75t_R FILLER_112_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_617 ();
 DECAPx10_ASAP7_75t_R FILLER_112_646 ();
 DECAPx2_ASAP7_75t_R FILLER_112_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_674 ();
 DECAPx10_ASAP7_75t_R FILLER_112_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_742 ();
 FILLER_ASAP7_75t_R FILLER_112_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_755 ();
 DECAPx10_ASAP7_75t_R FILLER_112_780 ();
 DECAPx2_ASAP7_75t_R FILLER_112_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_808 ();
 DECAPx1_ASAP7_75t_R FILLER_112_821 ();
 DECAPx2_ASAP7_75t_R FILLER_112_833 ();
 DECAPx1_ASAP7_75t_R FILLER_112_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_866 ();
 DECAPx4_ASAP7_75t_R FILLER_112_889 ();
 DECAPx10_ASAP7_75t_R FILLER_112_921 ();
 DECAPx2_ASAP7_75t_R FILLER_112_943 ();
 FILLER_ASAP7_75t_R FILLER_112_949 ();
 DECAPx4_ASAP7_75t_R FILLER_112_979 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_112_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1167 ();
 FILLER_ASAP7_75t_R FILLER_112_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_113_2 ();
 DECAPx10_ASAP7_75t_R FILLER_113_24 ();
 DECAPx10_ASAP7_75t_R FILLER_113_46 ();
 DECAPx2_ASAP7_75t_R FILLER_113_68 ();
 FILLER_ASAP7_75t_R FILLER_113_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_102 ();
 DECAPx2_ASAP7_75t_R FILLER_113_109 ();
 FILLER_ASAP7_75t_R FILLER_113_115 ();
 DECAPx10_ASAP7_75t_R FILLER_113_154 ();
 DECAPx4_ASAP7_75t_R FILLER_113_176 ();
 DECAPx1_ASAP7_75t_R FILLER_113_192 ();
 DECAPx10_ASAP7_75t_R FILLER_113_206 ();
 DECAPx2_ASAP7_75t_R FILLER_113_228 ();
 FILLER_ASAP7_75t_R FILLER_113_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_236 ();
 DECAPx4_ASAP7_75t_R FILLER_113_259 ();
 DECAPx2_ASAP7_75t_R FILLER_113_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_308 ();
 DECAPx2_ASAP7_75t_R FILLER_113_322 ();
 DECAPx1_ASAP7_75t_R FILLER_113_336 ();
 DECAPx2_ASAP7_75t_R FILLER_113_359 ();
 DECAPx1_ASAP7_75t_R FILLER_113_375 ();
 FILLER_ASAP7_75t_R FILLER_113_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_387 ();
 FILLER_ASAP7_75t_R FILLER_113_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_447 ();
 FILLER_ASAP7_75t_R FILLER_113_454 ();
 FILLER_ASAP7_75t_R FILLER_113_464 ();
 DECAPx1_ASAP7_75t_R FILLER_113_506 ();
 DECAPx4_ASAP7_75t_R FILLER_113_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_565 ();
 FILLER_ASAP7_75t_R FILLER_113_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_574 ();
 DECAPx6_ASAP7_75t_R FILLER_113_581 ();
 FILLER_ASAP7_75t_R FILLER_113_595 ();
 DECAPx2_ASAP7_75t_R FILLER_113_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_624 ();
 DECAPx10_ASAP7_75t_R FILLER_113_695 ();
 DECAPx6_ASAP7_75t_R FILLER_113_717 ();
 DECAPx1_ASAP7_75t_R FILLER_113_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_735 ();
 DECAPx1_ASAP7_75t_R FILLER_113_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_752 ();
 FILLER_ASAP7_75t_R FILLER_113_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_761 ();
 DECAPx4_ASAP7_75t_R FILLER_113_780 ();
 DECAPx6_ASAP7_75t_R FILLER_113_796 ();
 FILLER_ASAP7_75t_R FILLER_113_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_812 ();
 FILLER_ASAP7_75t_R FILLER_113_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_823 ();
 FILLER_ASAP7_75t_R FILLER_113_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_839 ();
 DECAPx1_ASAP7_75t_R FILLER_113_852 ();
 DECAPx4_ASAP7_75t_R FILLER_113_862 ();
 FILLER_ASAP7_75t_R FILLER_113_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_874 ();
 DECAPx1_ASAP7_75t_R FILLER_113_899 ();
 DECAPx6_ASAP7_75t_R FILLER_113_907 ();
 FILLER_ASAP7_75t_R FILLER_113_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_923 ();
 DECAPx6_ASAP7_75t_R FILLER_113_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_940 ();
 DECAPx6_ASAP7_75t_R FILLER_113_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_977 ();
 DECAPx10_ASAP7_75t_R FILLER_113_998 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1064 ();
 FILLER_ASAP7_75t_R FILLER_113_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1084 ();
 FILLER_ASAP7_75t_R FILLER_113_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1132 ();
 FILLER_ASAP7_75t_R FILLER_113_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1186 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1204 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_114_2 ();
 DECAPx10_ASAP7_75t_R FILLER_114_24 ();
 DECAPx10_ASAP7_75t_R FILLER_114_46 ();
 DECAPx6_ASAP7_75t_R FILLER_114_68 ();
 DECAPx2_ASAP7_75t_R FILLER_114_82 ();
 FILLER_ASAP7_75t_R FILLER_114_100 ();
 FILLER_ASAP7_75t_R FILLER_114_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_111 ();
 DECAPx1_ASAP7_75t_R FILLER_114_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_133 ();
 DECAPx2_ASAP7_75t_R FILLER_114_140 ();
 FILLER_ASAP7_75t_R FILLER_114_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_148 ();
 DECAPx2_ASAP7_75t_R FILLER_114_171 ();
 DECAPx6_ASAP7_75t_R FILLER_114_188 ();
 DECAPx2_ASAP7_75t_R FILLER_114_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_208 ();
 DECAPx6_ASAP7_75t_R FILLER_114_237 ();
 FILLER_ASAP7_75t_R FILLER_114_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_308 ();
 FILLER_ASAP7_75t_R FILLER_114_312 ();
 DECAPx2_ASAP7_75t_R FILLER_114_321 ();
 DECAPx4_ASAP7_75t_R FILLER_114_333 ();
 FILLER_ASAP7_75t_R FILLER_114_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_352 ();
 DECAPx10_ASAP7_75t_R FILLER_114_360 ();
 DECAPx2_ASAP7_75t_R FILLER_114_394 ();
 FILLER_ASAP7_75t_R FILLER_114_400 ();
 DECAPx6_ASAP7_75t_R FILLER_114_424 ();
 FILLER_ASAP7_75t_R FILLER_114_438 ();
 FILLER_ASAP7_75t_R FILLER_114_454 ();
 DECAPx6_ASAP7_75t_R FILLER_114_464 ();
 FILLER_ASAP7_75t_R FILLER_114_500 ();
 DECAPx10_ASAP7_75t_R FILLER_114_524 ();
 FILLER_ASAP7_75t_R FILLER_114_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_574 ();
 FILLER_ASAP7_75t_R FILLER_114_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_605 ();
 FILLER_ASAP7_75t_R FILLER_114_612 ();
 DECAPx10_ASAP7_75t_R FILLER_114_644 ();
 DECAPx10_ASAP7_75t_R FILLER_114_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_688 ();
 DECAPx6_ASAP7_75t_R FILLER_114_699 ();
 FILLER_ASAP7_75t_R FILLER_114_713 ();
 DECAPx2_ASAP7_75t_R FILLER_114_725 ();
 FILLER_ASAP7_75t_R FILLER_114_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_748 ();
 FILLER_ASAP7_75t_R FILLER_114_789 ();
 FILLER_ASAP7_75t_R FILLER_114_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_811 ();
 DECAPx2_ASAP7_75t_R FILLER_114_818 ();
 FILLER_ASAP7_75t_R FILLER_114_824 ();
 DECAPx1_ASAP7_75t_R FILLER_114_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_844 ();
 FILLER_ASAP7_75t_R FILLER_114_853 ();
 FILLER_ASAP7_75t_R FILLER_114_861 ();
 DECAPx10_ASAP7_75t_R FILLER_114_887 ();
 DECAPx6_ASAP7_75t_R FILLER_114_909 ();
 DECAPx1_ASAP7_75t_R FILLER_114_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_927 ();
 FILLER_ASAP7_75t_R FILLER_114_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_959 ();
 DECAPx4_ASAP7_75t_R FILLER_114_966 ();
 FILLER_ASAP7_75t_R FILLER_114_976 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1037 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1079 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1125 ();
 FILLER_ASAP7_75t_R FILLER_114_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_115_2 ();
 DECAPx10_ASAP7_75t_R FILLER_115_24 ();
 DECAPx10_ASAP7_75t_R FILLER_115_46 ();
 DECAPx4_ASAP7_75t_R FILLER_115_68 ();
 FILLER_ASAP7_75t_R FILLER_115_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_91 ();
 FILLER_ASAP7_75t_R FILLER_115_95 ();
 DECAPx1_ASAP7_75t_R FILLER_115_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_122 ();
 DECAPx1_ASAP7_75t_R FILLER_115_145 ();
 DECAPx10_ASAP7_75t_R FILLER_115_205 ();
 DECAPx10_ASAP7_75t_R FILLER_115_227 ();
 DECAPx1_ASAP7_75t_R FILLER_115_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_253 ();
 DECAPx6_ASAP7_75t_R FILLER_115_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_281 ();
 DECAPx6_ASAP7_75t_R FILLER_115_288 ();
 DECAPx2_ASAP7_75t_R FILLER_115_302 ();
 DECAPx2_ASAP7_75t_R FILLER_115_311 ();
 DECAPx10_ASAP7_75t_R FILLER_115_351 ();
 DECAPx10_ASAP7_75t_R FILLER_115_390 ();
 DECAPx2_ASAP7_75t_R FILLER_115_412 ();
 FILLER_ASAP7_75t_R FILLER_115_418 ();
 DECAPx4_ASAP7_75t_R FILLER_115_444 ();
 DECAPx6_ASAP7_75t_R FILLER_115_464 ();
 DECAPx1_ASAP7_75t_R FILLER_115_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_482 ();
 DECAPx2_ASAP7_75t_R FILLER_115_489 ();
 FILLER_ASAP7_75t_R FILLER_115_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_533 ();
 FILLER_ASAP7_75t_R FILLER_115_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_554 ();
 FILLER_ASAP7_75t_R FILLER_115_565 ();
 FILLER_ASAP7_75t_R FILLER_115_573 ();
 FILLER_ASAP7_75t_R FILLER_115_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_583 ();
 DECAPx1_ASAP7_75t_R FILLER_115_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_602 ();
 FILLER_ASAP7_75t_R FILLER_115_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_622 ();
 DECAPx6_ASAP7_75t_R FILLER_115_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_644 ();
 DECAPx10_ASAP7_75t_R FILLER_115_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_687 ();
 DECAPx4_ASAP7_75t_R FILLER_115_698 ();
 DECAPx2_ASAP7_75t_R FILLER_115_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_736 ();
 DECAPx2_ASAP7_75t_R FILLER_115_743 ();
 DECAPx1_ASAP7_75t_R FILLER_115_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_761 ();
 DECAPx4_ASAP7_75t_R FILLER_115_769 ();
 FILLER_ASAP7_75t_R FILLER_115_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_781 ();
 FILLER_ASAP7_75t_R FILLER_115_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_791 ();
 DECAPx2_ASAP7_75t_R FILLER_115_798 ();
 DECAPx2_ASAP7_75t_R FILLER_115_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_833 ();
 DECAPx4_ASAP7_75t_R FILLER_115_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_850 ();
 DECAPx6_ASAP7_75t_R FILLER_115_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_879 ();
 FILLER_ASAP7_75t_R FILLER_115_902 ();
 DECAPx6_ASAP7_75t_R FILLER_115_926 ();
 DECAPx1_ASAP7_75t_R FILLER_115_940 ();
 DECAPx10_ASAP7_75t_R FILLER_115_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_988 ();
 DECAPx4_ASAP7_75t_R FILLER_115_995 ();
 FILLER_ASAP7_75t_R FILLER_115_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_115_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1099 ();
 FILLER_ASAP7_75t_R FILLER_115_1106 ();
 FILLER_ASAP7_75t_R FILLER_115_1117 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1125 ();
 FILLER_ASAP7_75t_R FILLER_115_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1149 ();
 FILLER_ASAP7_75t_R FILLER_115_1159 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1167 ();
 FILLER_ASAP7_75t_R FILLER_115_1179 ();
 FILLER_ASAP7_75t_R FILLER_115_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1210 ();
 FILLER_ASAP7_75t_R FILLER_115_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_116_2 ();
 DECAPx10_ASAP7_75t_R FILLER_116_24 ();
 DECAPx10_ASAP7_75t_R FILLER_116_46 ();
 FILLER_ASAP7_75t_R FILLER_116_68 ();
 DECAPx2_ASAP7_75t_R FILLER_116_126 ();
 FILLER_ASAP7_75t_R FILLER_116_132 ();
 DECAPx4_ASAP7_75t_R FILLER_116_147 ();
 FILLER_ASAP7_75t_R FILLER_116_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_159 ();
 FILLER_ASAP7_75t_R FILLER_116_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_179 ();
 DECAPx10_ASAP7_75t_R FILLER_116_197 ();
 FILLER_ASAP7_75t_R FILLER_116_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_282 ();
 FILLER_ASAP7_75t_R FILLER_116_291 ();
 FILLER_ASAP7_75t_R FILLER_116_305 ();
 DECAPx1_ASAP7_75t_R FILLER_116_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_314 ();
 DECAPx2_ASAP7_75t_R FILLER_116_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_356 ();
 DECAPx2_ASAP7_75t_R FILLER_116_363 ();
 FILLER_ASAP7_75t_R FILLER_116_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_371 ();
 FILLER_ASAP7_75t_R FILLER_116_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_420 ();
 DECAPx4_ASAP7_75t_R FILLER_116_427 ();
 FILLER_ASAP7_75t_R FILLER_116_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_439 ();
 DECAPx2_ASAP7_75t_R FILLER_116_454 ();
 FILLER_ASAP7_75t_R FILLER_116_460 ();
 FILLER_ASAP7_75t_R FILLER_116_464 ();
 FILLER_ASAP7_75t_R FILLER_116_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_476 ();
 DECAPx10_ASAP7_75t_R FILLER_116_495 ();
 DECAPx2_ASAP7_75t_R FILLER_116_517 ();
 FILLER_ASAP7_75t_R FILLER_116_545 ();
 DECAPx4_ASAP7_75t_R FILLER_116_555 ();
 FILLER_ASAP7_75t_R FILLER_116_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_567 ();
 DECAPx1_ASAP7_75t_R FILLER_116_582 ();
 FILLER_ASAP7_75t_R FILLER_116_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_594 ();
 DECAPx4_ASAP7_75t_R FILLER_116_605 ();
 DECAPx1_ASAP7_75t_R FILLER_116_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_632 ();
 FILLER_ASAP7_75t_R FILLER_116_643 ();
 DECAPx10_ASAP7_75t_R FILLER_116_687 ();
 DECAPx2_ASAP7_75t_R FILLER_116_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_715 ();
 DECAPx4_ASAP7_75t_R FILLER_116_742 ();
 FILLER_ASAP7_75t_R FILLER_116_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_754 ();
 DECAPx4_ASAP7_75t_R FILLER_116_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_788 ();
 DECAPx6_ASAP7_75t_R FILLER_116_800 ();
 DECAPx1_ASAP7_75t_R FILLER_116_826 ();
 DECAPx6_ASAP7_75t_R FILLER_116_844 ();
 DECAPx2_ASAP7_75t_R FILLER_116_880 ();
 FILLER_ASAP7_75t_R FILLER_116_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_894 ();
 DECAPx2_ASAP7_75t_R FILLER_116_901 ();
 FILLER_ASAP7_75t_R FILLER_116_925 ();
 DECAPx2_ASAP7_75t_R FILLER_116_933 ();
 DECAPx2_ASAP7_75t_R FILLER_116_946 ();
 FILLER_ASAP7_75t_R FILLER_116_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_954 ();
 DECAPx10_ASAP7_75t_R FILLER_116_977 ();
 DECAPx2_ASAP7_75t_R FILLER_116_999 ();
 FILLER_ASAP7_75t_R FILLER_116_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1007 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1014 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1069 ();
 FILLER_ASAP7_75t_R FILLER_116_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1095 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1171 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_117_2 ();
 DECAPx10_ASAP7_75t_R FILLER_117_24 ();
 DECAPx10_ASAP7_75t_R FILLER_117_46 ();
 DECAPx6_ASAP7_75t_R FILLER_117_68 ();
 DECAPx6_ASAP7_75t_R FILLER_117_99 ();
 FILLER_ASAP7_75t_R FILLER_117_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_115 ();
 DECAPx4_ASAP7_75t_R FILLER_117_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_146 ();
 DECAPx6_ASAP7_75t_R FILLER_117_159 ();
 FILLER_ASAP7_75t_R FILLER_117_173 ();
 DECAPx10_ASAP7_75t_R FILLER_117_196 ();
 DECAPx10_ASAP7_75t_R FILLER_117_218 ();
 DECAPx2_ASAP7_75t_R FILLER_117_240 ();
 DECAPx6_ASAP7_75t_R FILLER_117_268 ();
 DECAPx10_ASAP7_75t_R FILLER_117_288 ();
 DECAPx1_ASAP7_75t_R FILLER_117_310 ();
 DECAPx6_ASAP7_75t_R FILLER_117_320 ();
 FILLER_ASAP7_75t_R FILLER_117_334 ();
 DECAPx4_ASAP7_75t_R FILLER_117_342 ();
 FILLER_ASAP7_75t_R FILLER_117_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_354 ();
 DECAPx10_ASAP7_75t_R FILLER_117_375 ();
 DECAPx2_ASAP7_75t_R FILLER_117_403 ();
 DECAPx1_ASAP7_75t_R FILLER_117_417 ();
 DECAPx2_ASAP7_75t_R FILLER_117_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_443 ();
 DECAPx1_ASAP7_75t_R FILLER_117_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_474 ();
 FILLER_ASAP7_75t_R FILLER_117_485 ();
 FILLER_ASAP7_75t_R FILLER_117_510 ();
 DECAPx6_ASAP7_75t_R FILLER_117_534 ();
 DECAPx1_ASAP7_75t_R FILLER_117_548 ();
 DECAPx6_ASAP7_75t_R FILLER_117_580 ();
 FILLER_ASAP7_75t_R FILLER_117_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_596 ();
 DECAPx2_ASAP7_75t_R FILLER_117_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_624 ();
 DECAPx6_ASAP7_75t_R FILLER_117_645 ();
 DECAPx2_ASAP7_75t_R FILLER_117_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_665 ();
 DECAPx2_ASAP7_75t_R FILLER_117_688 ();
 FILLER_ASAP7_75t_R FILLER_117_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_714 ();
 DECAPx4_ASAP7_75t_R FILLER_117_721 ();
 FILLER_ASAP7_75t_R FILLER_117_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_737 ();
 FILLER_ASAP7_75t_R FILLER_117_748 ();
 FILLER_ASAP7_75t_R FILLER_117_758 ();
 FILLER_ASAP7_75t_R FILLER_117_768 ();
 DECAPx4_ASAP7_75t_R FILLER_117_780 ();
 FILLER_ASAP7_75t_R FILLER_117_790 ();
 DECAPx10_ASAP7_75t_R FILLER_117_798 ();
 DECAPx6_ASAP7_75t_R FILLER_117_820 ();
 DECAPx1_ASAP7_75t_R FILLER_117_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_844 ();
 DECAPx10_ASAP7_75t_R FILLER_117_851 ();
 DECAPx4_ASAP7_75t_R FILLER_117_873 ();
 FILLER_ASAP7_75t_R FILLER_117_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_907 ();
 FILLER_ASAP7_75t_R FILLER_117_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_934 ();
 DECAPx6_ASAP7_75t_R FILLER_117_943 ();
 DECAPx2_ASAP7_75t_R FILLER_117_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_963 ();
 DECAPx4_ASAP7_75t_R FILLER_117_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_980 ();
 DECAPx10_ASAP7_75t_R FILLER_117_987 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1009 ();
 FILLER_ASAP7_75t_R FILLER_117_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1049 ();
 FILLER_ASAP7_75t_R FILLER_117_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1073 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1139 ();
 FILLER_ASAP7_75t_R FILLER_117_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1187 ();
 FILLER_ASAP7_75t_R FILLER_117_1203 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_118_2 ();
 DECAPx10_ASAP7_75t_R FILLER_118_24 ();
 DECAPx10_ASAP7_75t_R FILLER_118_46 ();
 DECAPx6_ASAP7_75t_R FILLER_118_68 ();
 FILLER_ASAP7_75t_R FILLER_118_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_84 ();
 DECAPx2_ASAP7_75t_R FILLER_118_107 ();
 FILLER_ASAP7_75t_R FILLER_118_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_148 ();
 DECAPx10_ASAP7_75t_R FILLER_118_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_177 ();
 FILLER_ASAP7_75t_R FILLER_118_186 ();
 DECAPx10_ASAP7_75t_R FILLER_118_194 ();
 DECAPx10_ASAP7_75t_R FILLER_118_216 ();
 DECAPx10_ASAP7_75t_R FILLER_118_238 ();
 DECAPx10_ASAP7_75t_R FILLER_118_260 ();
 DECAPx2_ASAP7_75t_R FILLER_118_282 ();
 DECAPx2_ASAP7_75t_R FILLER_118_330 ();
 FILLER_ASAP7_75t_R FILLER_118_336 ();
 DECAPx2_ASAP7_75t_R FILLER_118_346 ();
 FILLER_ASAP7_75t_R FILLER_118_374 ();
 DECAPx2_ASAP7_75t_R FILLER_118_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_427 ();
 DECAPx1_ASAP7_75t_R FILLER_118_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_444 ();
 FILLER_ASAP7_75t_R FILLER_118_448 ();
 FILLER_ASAP7_75t_R FILLER_118_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_464 ();
 DECAPx10_ASAP7_75t_R FILLER_118_471 ();
 DECAPx4_ASAP7_75t_R FILLER_118_493 ();
 DECAPx10_ASAP7_75t_R FILLER_118_513 ();
 DECAPx6_ASAP7_75t_R FILLER_118_535 ();
 FILLER_ASAP7_75t_R FILLER_118_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_551 ();
 DECAPx2_ASAP7_75t_R FILLER_118_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_568 ();
 DECAPx6_ASAP7_75t_R FILLER_118_589 ();
 FILLER_ASAP7_75t_R FILLER_118_603 ();
 DECAPx2_ASAP7_75t_R FILLER_118_611 ();
 DECAPx4_ASAP7_75t_R FILLER_118_627 ();
 FILLER_ASAP7_75t_R FILLER_118_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_639 ();
 DECAPx2_ASAP7_75t_R FILLER_118_660 ();
 DECAPx10_ASAP7_75t_R FILLER_118_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_738 ();
 FILLER_ASAP7_75t_R FILLER_118_749 ();
 FILLER_ASAP7_75t_R FILLER_118_757 ();
 FILLER_ASAP7_75t_R FILLER_118_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_769 ();
 DECAPx6_ASAP7_75t_R FILLER_118_776 ();
 FILLER_ASAP7_75t_R FILLER_118_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_801 ();
 FILLER_ASAP7_75t_R FILLER_118_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_814 ();
 FILLER_ASAP7_75t_R FILLER_118_829 ();
 FILLER_ASAP7_75t_R FILLER_118_843 ();
 DECAPx10_ASAP7_75t_R FILLER_118_851 ();
 DECAPx2_ASAP7_75t_R FILLER_118_873 ();
 DECAPx4_ASAP7_75t_R FILLER_118_897 ();
 FILLER_ASAP7_75t_R FILLER_118_913 ();
 FILLER_ASAP7_75t_R FILLER_118_921 ();
 FILLER_ASAP7_75t_R FILLER_118_937 ();
 DECAPx10_ASAP7_75t_R FILLER_118_947 ();
 DECAPx4_ASAP7_75t_R FILLER_118_969 ();
 FILLER_ASAP7_75t_R FILLER_118_979 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1052 ();
 FILLER_ASAP7_75t_R FILLER_118_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1112 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1134 ();
 FILLER_ASAP7_75t_R FILLER_118_1148 ();
 FILLER_ASAP7_75t_R FILLER_118_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1167 ();
 FILLER_ASAP7_75t_R FILLER_118_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1208 ();
 FILLER_ASAP7_75t_R FILLER_118_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_119_2 ();
 DECAPx10_ASAP7_75t_R FILLER_119_24 ();
 DECAPx10_ASAP7_75t_R FILLER_119_46 ();
 DECAPx6_ASAP7_75t_R FILLER_119_68 ();
 DECAPx2_ASAP7_75t_R FILLER_119_82 ();
 DECAPx10_ASAP7_75t_R FILLER_119_94 ();
 DECAPx10_ASAP7_75t_R FILLER_119_116 ();
 DECAPx2_ASAP7_75t_R FILLER_119_138 ();
 FILLER_ASAP7_75t_R FILLER_119_144 ();
 DECAPx6_ASAP7_75t_R FILLER_119_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_177 ();
 DECAPx10_ASAP7_75t_R FILLER_119_193 ();
 DECAPx10_ASAP7_75t_R FILLER_119_215 ();
 DECAPx6_ASAP7_75t_R FILLER_119_237 ();
 FILLER_ASAP7_75t_R FILLER_119_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_253 ();
 DECAPx6_ASAP7_75t_R FILLER_119_282 ();
 DECAPx2_ASAP7_75t_R FILLER_119_296 ();
 DECAPx10_ASAP7_75t_R FILLER_119_324 ();
 DECAPx1_ASAP7_75t_R FILLER_119_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_350 ();
 DECAPx10_ASAP7_75t_R FILLER_119_373 ();
 FILLER_ASAP7_75t_R FILLER_119_405 ();
 DECAPx2_ASAP7_75t_R FILLER_119_410 ();
 FILLER_ASAP7_75t_R FILLER_119_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_418 ();
 DECAPx4_ASAP7_75t_R FILLER_119_429 ();
 DECAPx1_ASAP7_75t_R FILLER_119_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_453 ();
 FILLER_ASAP7_75t_R FILLER_119_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_464 ();
 FILLER_ASAP7_75t_R FILLER_119_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_487 ();
 DECAPx2_ASAP7_75t_R FILLER_119_494 ();
 DECAPx4_ASAP7_75t_R FILLER_119_513 ();
 FILLER_ASAP7_75t_R FILLER_119_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_525 ();
 DECAPx2_ASAP7_75t_R FILLER_119_557 ();
 FILLER_ASAP7_75t_R FILLER_119_563 ();
 DECAPx6_ASAP7_75t_R FILLER_119_583 ();
 DECAPx1_ASAP7_75t_R FILLER_119_597 ();
 DECAPx10_ASAP7_75t_R FILLER_119_611 ();
 DECAPx10_ASAP7_75t_R FILLER_119_633 ();
 DECAPx6_ASAP7_75t_R FILLER_119_655 ();
 DECAPx6_ASAP7_75t_R FILLER_119_691 ();
 DECAPx1_ASAP7_75t_R FILLER_119_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_709 ();
 DECAPx4_ASAP7_75t_R FILLER_119_728 ();
 FILLER_ASAP7_75t_R FILLER_119_738 ();
 FILLER_ASAP7_75t_R FILLER_119_746 ();
 FILLER_ASAP7_75t_R FILLER_119_752 ();
 FILLER_ASAP7_75t_R FILLER_119_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_766 ();
 FILLER_ASAP7_75t_R FILLER_119_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_789 ();
 FILLER_ASAP7_75t_R FILLER_119_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_798 ();
 FILLER_ASAP7_75t_R FILLER_119_811 ();
 DECAPx2_ASAP7_75t_R FILLER_119_823 ();
 FILLER_ASAP7_75t_R FILLER_119_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_831 ();
 DECAPx4_ASAP7_75t_R FILLER_119_842 ();
 FILLER_ASAP7_75t_R FILLER_119_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_854 ();
 FILLER_ASAP7_75t_R FILLER_119_891 ();
 FILLER_ASAP7_75t_R FILLER_119_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_907 ();
 FILLER_ASAP7_75t_R FILLER_119_922 ();
 FILLER_ASAP7_75t_R FILLER_119_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_931 ();
 FILLER_ASAP7_75t_R FILLER_119_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_977 ();
 DECAPx2_ASAP7_75t_R FILLER_119_984 ();
 FILLER_ASAP7_75t_R FILLER_119_990 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1090 ();
 DECAPx6_ASAP7_75t_R FILLER_119_1112 ();
 FILLER_ASAP7_75t_R FILLER_119_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1150 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1182 ();
 FILLER_ASAP7_75t_R FILLER_119_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1190 ();
 FILLER_ASAP7_75t_R FILLER_119_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_120_2 ();
 DECAPx10_ASAP7_75t_R FILLER_120_24 ();
 DECAPx10_ASAP7_75t_R FILLER_120_46 ();
 DECAPx10_ASAP7_75t_R FILLER_120_68 ();
 DECAPx6_ASAP7_75t_R FILLER_120_90 ();
 DECAPx2_ASAP7_75t_R FILLER_120_110 ();
 DECAPx1_ASAP7_75t_R FILLER_120_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_137 ();
 DECAPx2_ASAP7_75t_R FILLER_120_146 ();
 DECAPx10_ASAP7_75t_R FILLER_120_217 ();
 DECAPx6_ASAP7_75t_R FILLER_120_239 ();
 DECAPx1_ASAP7_75t_R FILLER_120_253 ();
 DECAPx10_ASAP7_75t_R FILLER_120_283 ();
 DECAPx10_ASAP7_75t_R FILLER_120_325 ();
 DECAPx10_ASAP7_75t_R FILLER_120_347 ();
 DECAPx1_ASAP7_75t_R FILLER_120_369 ();
 FILLER_ASAP7_75t_R FILLER_120_405 ();
 DECAPx4_ASAP7_75t_R FILLER_120_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_461 ();
 DECAPx6_ASAP7_75t_R FILLER_120_464 ();
 DECAPx2_ASAP7_75t_R FILLER_120_502 ();
 FILLER_ASAP7_75t_R FILLER_120_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_518 ();
 DECAPx4_ASAP7_75t_R FILLER_120_539 ();
 FILLER_ASAP7_75t_R FILLER_120_555 ();
 DECAPx4_ASAP7_75t_R FILLER_120_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_571 ();
 FILLER_ASAP7_75t_R FILLER_120_602 ();
 DECAPx1_ASAP7_75t_R FILLER_120_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_618 ();
 DECAPx1_ASAP7_75t_R FILLER_120_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_643 ();
 DECAPx10_ASAP7_75t_R FILLER_120_666 ();
 DECAPx10_ASAP7_75t_R FILLER_120_688 ();
 FILLER_ASAP7_75t_R FILLER_120_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_712 ();
 DECAPx1_ASAP7_75t_R FILLER_120_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_727 ();
 DECAPx1_ASAP7_75t_R FILLER_120_753 ();
 DECAPx2_ASAP7_75t_R FILLER_120_782 ();
 DECAPx2_ASAP7_75t_R FILLER_120_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_806 ();
 DECAPx10_ASAP7_75t_R FILLER_120_813 ();
 DECAPx1_ASAP7_75t_R FILLER_120_867 ();
 FILLER_ASAP7_75t_R FILLER_120_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_909 ();
 DECAPx1_ASAP7_75t_R FILLER_120_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_936 ();
 DECAPx1_ASAP7_75t_R FILLER_120_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_948 ();
 DECAPx1_ASAP7_75t_R FILLER_120_971 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1014 ();
 FILLER_ASAP7_75t_R FILLER_120_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_120_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_120_1111 ();
 FILLER_ASAP7_75t_R FILLER_120_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_120_1152 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1185 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1200 ();
 FILLER_ASAP7_75t_R FILLER_120_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_121_2 ();
 DECAPx10_ASAP7_75t_R FILLER_121_24 ();
 DECAPx10_ASAP7_75t_R FILLER_121_46 ();
 DECAPx6_ASAP7_75t_R FILLER_121_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_82 ();
 DECAPx2_ASAP7_75t_R FILLER_121_94 ();
 FILLER_ASAP7_75t_R FILLER_121_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_124 ();
 DECAPx2_ASAP7_75t_R FILLER_121_145 ();
 FILLER_ASAP7_75t_R FILLER_121_151 ();
 DECAPx6_ASAP7_75t_R FILLER_121_166 ();
 DECAPx1_ASAP7_75t_R FILLER_121_180 ();
 FILLER_ASAP7_75t_R FILLER_121_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_208 ();
 DECAPx1_ASAP7_75t_R FILLER_121_233 ();
 FILLER_ASAP7_75t_R FILLER_121_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_259 ();
 DECAPx10_ASAP7_75t_R FILLER_121_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_304 ();
 DECAPx4_ASAP7_75t_R FILLER_121_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_322 ();
 DECAPx1_ASAP7_75t_R FILLER_121_329 ();
 DECAPx6_ASAP7_75t_R FILLER_121_377 ();
 DECAPx2_ASAP7_75t_R FILLER_121_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_406 ();
 FILLER_ASAP7_75t_R FILLER_121_416 ();
 DECAPx10_ASAP7_75t_R FILLER_121_424 ();
 DECAPx2_ASAP7_75t_R FILLER_121_446 ();
 FILLER_ASAP7_75t_R FILLER_121_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_454 ();
 DECAPx2_ASAP7_75t_R FILLER_121_461 ();
 DECAPx1_ASAP7_75t_R FILLER_121_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_479 ();
 DECAPx1_ASAP7_75t_R FILLER_121_486 ();
 FILLER_ASAP7_75t_R FILLER_121_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_513 ();
 DECAPx4_ASAP7_75t_R FILLER_121_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_546 ();
 DECAPx10_ASAP7_75t_R FILLER_121_561 ();
 DECAPx6_ASAP7_75t_R FILLER_121_583 ();
 DECAPx2_ASAP7_75t_R FILLER_121_608 ();
 FILLER_ASAP7_75t_R FILLER_121_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_616 ();
 DECAPx4_ASAP7_75t_R FILLER_121_661 ();
 DECAPx4_ASAP7_75t_R FILLER_121_681 ();
 FILLER_ASAP7_75t_R FILLER_121_691 ();
 DECAPx4_ASAP7_75t_R FILLER_121_716 ();
 DECAPx1_ASAP7_75t_R FILLER_121_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_737 ();
 DECAPx6_ASAP7_75t_R FILLER_121_748 ();
 DECAPx1_ASAP7_75t_R FILLER_121_762 ();
 DECAPx6_ASAP7_75t_R FILLER_121_772 ();
 FILLER_ASAP7_75t_R FILLER_121_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_788 ();
 DECAPx4_ASAP7_75t_R FILLER_121_795 ();
 FILLER_ASAP7_75t_R FILLER_121_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_807 ();
 FILLER_ASAP7_75t_R FILLER_121_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_832 ();
 DECAPx6_ASAP7_75t_R FILLER_121_840 ();
 FILLER_ASAP7_75t_R FILLER_121_854 ();
 DECAPx2_ASAP7_75t_R FILLER_121_862 ();
 DECAPx2_ASAP7_75t_R FILLER_121_918 ();
 DECAPx6_ASAP7_75t_R FILLER_121_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_940 ();
 DECAPx1_ASAP7_75t_R FILLER_121_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_953 ();
 DECAPx4_ASAP7_75t_R FILLER_121_976 ();
 FILLER_ASAP7_75t_R FILLER_121_986 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_121_1072 ();
 FILLER_ASAP7_75t_R FILLER_121_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1088 ();
 FILLER_ASAP7_75t_R FILLER_121_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1144 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1161 ();
 FILLER_ASAP7_75t_R FILLER_121_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_122_2 ();
 DECAPx10_ASAP7_75t_R FILLER_122_24 ();
 DECAPx10_ASAP7_75t_R FILLER_122_46 ();
 DECAPx2_ASAP7_75t_R FILLER_122_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_74 ();
 FILLER_ASAP7_75t_R FILLER_122_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_114 ();
 DECAPx10_ASAP7_75t_R FILLER_122_122 ();
 DECAPx2_ASAP7_75t_R FILLER_122_144 ();
 FILLER_ASAP7_75t_R FILLER_122_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_152 ();
 DECAPx1_ASAP7_75t_R FILLER_122_168 ();
 DECAPx6_ASAP7_75t_R FILLER_122_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_203 ();
 DECAPx1_ASAP7_75t_R FILLER_122_224 ();
 FILLER_ASAP7_75t_R FILLER_122_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_233 ();
 DECAPx2_ASAP7_75t_R FILLER_122_246 ();
 DECAPx4_ASAP7_75t_R FILLER_122_264 ();
 FILLER_ASAP7_75t_R FILLER_122_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_276 ();
 DECAPx4_ASAP7_75t_R FILLER_122_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_309 ();
 DECAPx2_ASAP7_75t_R FILLER_122_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_329 ();
 DECAPx6_ASAP7_75t_R FILLER_122_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_388 ();
 DECAPx1_ASAP7_75t_R FILLER_122_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_409 ();
 FILLER_ASAP7_75t_R FILLER_122_418 ();
 DECAPx1_ASAP7_75t_R FILLER_122_428 ();
 DECAPx2_ASAP7_75t_R FILLER_122_438 ();
 FILLER_ASAP7_75t_R FILLER_122_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_446 ();
 DECAPx2_ASAP7_75t_R FILLER_122_453 ();
 FILLER_ASAP7_75t_R FILLER_122_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_461 ();
 DECAPx2_ASAP7_75t_R FILLER_122_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_470 ();
 DECAPx2_ASAP7_75t_R FILLER_122_477 ();
 DECAPx2_ASAP7_75t_R FILLER_122_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_506 ();
 DECAPx1_ASAP7_75t_R FILLER_122_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_518 ();
 DECAPx2_ASAP7_75t_R FILLER_122_541 ();
 DECAPx4_ASAP7_75t_R FILLER_122_553 ();
 DECAPx4_ASAP7_75t_R FILLER_122_579 ();
 FILLER_ASAP7_75t_R FILLER_122_599 ();
 DECAPx4_ASAP7_75t_R FILLER_122_633 ();
 FILLER_ASAP7_75t_R FILLER_122_643 ();
 DECAPx10_ASAP7_75t_R FILLER_122_667 ();
 DECAPx10_ASAP7_75t_R FILLER_122_689 ();
 DECAPx4_ASAP7_75t_R FILLER_122_711 ();
 DECAPx6_ASAP7_75t_R FILLER_122_741 ();
 DECAPx2_ASAP7_75t_R FILLER_122_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_761 ();
 DECAPx2_ASAP7_75t_R FILLER_122_782 ();
 FILLER_ASAP7_75t_R FILLER_122_788 ();
 DECAPx4_ASAP7_75t_R FILLER_122_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_832 ();
 DECAPx2_ASAP7_75t_R FILLER_122_863 ();
 FILLER_ASAP7_75t_R FILLER_122_869 ();
 DECAPx10_ASAP7_75t_R FILLER_122_877 ();
 DECAPx10_ASAP7_75t_R FILLER_122_899 ();
 DECAPx2_ASAP7_75t_R FILLER_122_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_927 ();
 DECAPx2_ASAP7_75t_R FILLER_122_934 ();
 DECAPx6_ASAP7_75t_R FILLER_122_975 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1046 ();
 DECAPx4_ASAP7_75t_R FILLER_122_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1102 ();
 FILLER_ASAP7_75t_R FILLER_122_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1155 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1197 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1208 ();
 FILLER_ASAP7_75t_R FILLER_122_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_123_2 ();
 DECAPx10_ASAP7_75t_R FILLER_123_24 ();
 DECAPx10_ASAP7_75t_R FILLER_123_46 ();
 DECAPx4_ASAP7_75t_R FILLER_123_68 ();
 FILLER_ASAP7_75t_R FILLER_123_78 ();
 DECAPx6_ASAP7_75t_R FILLER_123_86 ();
 FILLER_ASAP7_75t_R FILLER_123_100 ();
 DECAPx4_ASAP7_75t_R FILLER_123_108 ();
 FILLER_ASAP7_75t_R FILLER_123_118 ();
 DECAPx2_ASAP7_75t_R FILLER_123_127 ();
 FILLER_ASAP7_75t_R FILLER_123_133 ();
 DECAPx6_ASAP7_75t_R FILLER_123_141 ();
 FILLER_ASAP7_75t_R FILLER_123_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_157 ();
 DECAPx4_ASAP7_75t_R FILLER_123_164 ();
 FILLER_ASAP7_75t_R FILLER_123_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_176 ();
 FILLER_ASAP7_75t_R FILLER_123_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_187 ();
 DECAPx6_ASAP7_75t_R FILLER_123_194 ();
 DECAPx2_ASAP7_75t_R FILLER_123_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_214 ();
 DECAPx6_ASAP7_75t_R FILLER_123_221 ();
 DECAPx1_ASAP7_75t_R FILLER_123_235 ();
 DECAPx2_ASAP7_75t_R FILLER_123_245 ();
 FILLER_ASAP7_75t_R FILLER_123_251 ();
 FILLER_ASAP7_75t_R FILLER_123_273 ();
 DECAPx2_ASAP7_75t_R FILLER_123_281 ();
 FILLER_ASAP7_75t_R FILLER_123_287 ();
 DECAPx6_ASAP7_75t_R FILLER_123_309 ();
 FILLER_ASAP7_75t_R FILLER_123_323 ();
 DECAPx10_ASAP7_75t_R FILLER_123_347 ();
 DECAPx1_ASAP7_75t_R FILLER_123_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_373 ();
 DECAPx1_ASAP7_75t_R FILLER_123_377 ();
 DECAPx1_ASAP7_75t_R FILLER_123_403 ();
 DECAPx2_ASAP7_75t_R FILLER_123_410 ();
 DECAPx4_ASAP7_75t_R FILLER_123_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_452 ();
 FILLER_ASAP7_75t_R FILLER_123_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_465 ();
 DECAPx4_ASAP7_75t_R FILLER_123_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_482 ();
 DECAPx10_ASAP7_75t_R FILLER_123_497 ();
 DECAPx10_ASAP7_75t_R FILLER_123_519 ();
 DECAPx1_ASAP7_75t_R FILLER_123_541 ();
 DECAPx2_ASAP7_75t_R FILLER_123_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_587 ();
 FILLER_ASAP7_75t_R FILLER_123_596 ();
 DECAPx2_ASAP7_75t_R FILLER_123_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_618 ();
 DECAPx2_ASAP7_75t_R FILLER_123_629 ();
 FILLER_ASAP7_75t_R FILLER_123_635 ();
 DECAPx4_ASAP7_75t_R FILLER_123_643 ();
 DECAPx1_ASAP7_75t_R FILLER_123_659 ();
 DECAPx10_ASAP7_75t_R FILLER_123_687 ();
 DECAPx10_ASAP7_75t_R FILLER_123_729 ();
 DECAPx2_ASAP7_75t_R FILLER_123_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_757 ();
 DECAPx10_ASAP7_75t_R FILLER_123_768 ();
 FILLER_ASAP7_75t_R FILLER_123_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_792 ();
 DECAPx10_ASAP7_75t_R FILLER_123_799 ();
 DECAPx2_ASAP7_75t_R FILLER_123_821 ();
 FILLER_ASAP7_75t_R FILLER_123_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_829 ();
 DECAPx10_ASAP7_75t_R FILLER_123_850 ();
 DECAPx6_ASAP7_75t_R FILLER_123_872 ();
 DECAPx2_ASAP7_75t_R FILLER_123_886 ();
 DECAPx6_ASAP7_75t_R FILLER_123_908 ();
 FILLER_ASAP7_75t_R FILLER_123_922 ();
 FILLER_ASAP7_75t_R FILLER_123_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_941 ();
 DECAPx6_ASAP7_75t_R FILLER_123_971 ();
 DECAPx1_ASAP7_75t_R FILLER_123_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_989 ();
 DECAPx10_ASAP7_75t_R FILLER_123_996 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1032 ();
 FILLER_ASAP7_75t_R FILLER_123_1044 ();
 FILLER_ASAP7_75t_R FILLER_123_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_123_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1160 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1217 ();
 DECAPx4_ASAP7_75t_R FILLER_124_2 ();
 FILLER_ASAP7_75t_R FILLER_124_12 ();
 DECAPx10_ASAP7_75t_R FILLER_124_20 ();
 DECAPx10_ASAP7_75t_R FILLER_124_42 ();
 DECAPx10_ASAP7_75t_R FILLER_124_64 ();
 DECAPx4_ASAP7_75t_R FILLER_124_86 ();
 DECAPx4_ASAP7_75t_R FILLER_124_119 ();
 FILLER_ASAP7_75t_R FILLER_124_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_131 ();
 DECAPx1_ASAP7_75t_R FILLER_124_154 ();
 DECAPx2_ASAP7_75t_R FILLER_124_180 ();
 FILLER_ASAP7_75t_R FILLER_124_186 ();
 FILLER_ASAP7_75t_R FILLER_124_210 ();
 FILLER_ASAP7_75t_R FILLER_124_234 ();
 DECAPx4_ASAP7_75t_R FILLER_124_242 ();
 FILLER_ASAP7_75t_R FILLER_124_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_254 ();
 DECAPx6_ASAP7_75t_R FILLER_124_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_275 ();
 FILLER_ASAP7_75t_R FILLER_124_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_303 ();
 DECAPx4_ASAP7_75t_R FILLER_124_312 ();
 DECAPx6_ASAP7_75t_R FILLER_124_342 ();
 DECAPx2_ASAP7_75t_R FILLER_124_356 ();
 DECAPx6_ASAP7_75t_R FILLER_124_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_396 ();
 DECAPx2_ASAP7_75t_R FILLER_124_405 ();
 FILLER_ASAP7_75t_R FILLER_124_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_413 ();
 DECAPx2_ASAP7_75t_R FILLER_124_428 ();
 FILLER_ASAP7_75t_R FILLER_124_434 ();
 DECAPx1_ASAP7_75t_R FILLER_124_458 ();
 FILLER_ASAP7_75t_R FILLER_124_464 ();
 DECAPx2_ASAP7_75t_R FILLER_124_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_478 ();
 DECAPx1_ASAP7_75t_R FILLER_124_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_487 ();
 FILLER_ASAP7_75t_R FILLER_124_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_493 ();
 DECAPx10_ASAP7_75t_R FILLER_124_516 ();
 DECAPx6_ASAP7_75t_R FILLER_124_538 ();
 DECAPx2_ASAP7_75t_R FILLER_124_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_558 ();
 DECAPx4_ASAP7_75t_R FILLER_124_572 ();
 FILLER_ASAP7_75t_R FILLER_124_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_595 ();
 DECAPx10_ASAP7_75t_R FILLER_124_609 ();
 DECAPx4_ASAP7_75t_R FILLER_124_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_656 ();
 FILLER_ASAP7_75t_R FILLER_124_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_665 ();
 FILLER_ASAP7_75t_R FILLER_124_686 ();
 DECAPx10_ASAP7_75t_R FILLER_124_694 ();
 DECAPx1_ASAP7_75t_R FILLER_124_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_720 ();
 DECAPx2_ASAP7_75t_R FILLER_124_761 ();
 FILLER_ASAP7_75t_R FILLER_124_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_769 ();
 DECAPx2_ASAP7_75t_R FILLER_124_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_818 ();
 DECAPx6_ASAP7_75t_R FILLER_124_863 ();
 DECAPx1_ASAP7_75t_R FILLER_124_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_887 ();
 DECAPx1_ASAP7_75t_R FILLER_124_902 ();
 FILLER_ASAP7_75t_R FILLER_124_914 ();
 DECAPx1_ASAP7_75t_R FILLER_124_922 ();
 DECAPx10_ASAP7_75t_R FILLER_124_941 ();
 DECAPx10_ASAP7_75t_R FILLER_124_963 ();
 DECAPx2_ASAP7_75t_R FILLER_124_985 ();
 FILLER_ASAP7_75t_R FILLER_124_991 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1005 ();
 FILLER_ASAP7_75t_R FILLER_124_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1034 ();
 FILLER_ASAP7_75t_R FILLER_124_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1067 ();
 FILLER_ASAP7_75t_R FILLER_124_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1167 ();
 FILLER_ASAP7_75t_R FILLER_124_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1184 ();
 FILLER_ASAP7_75t_R FILLER_124_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_2 ();
 DECAPx10_ASAP7_75t_R FILLER_125_9 ();
 DECAPx10_ASAP7_75t_R FILLER_125_31 ();
 DECAPx10_ASAP7_75t_R FILLER_125_53 ();
 DECAPx1_ASAP7_75t_R FILLER_125_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_79 ();
 DECAPx6_ASAP7_75t_R FILLER_125_146 ();
 DECAPx2_ASAP7_75t_R FILLER_125_182 ();
 FILLER_ASAP7_75t_R FILLER_125_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_233 ();
 DECAPx10_ASAP7_75t_R FILLER_125_260 ();
 DECAPx4_ASAP7_75t_R FILLER_125_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_292 ();
 DECAPx2_ASAP7_75t_R FILLER_125_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_303 ();
 DECAPx6_ASAP7_75t_R FILLER_125_310 ();
 DECAPx6_ASAP7_75t_R FILLER_125_331 ();
 DECAPx2_ASAP7_75t_R FILLER_125_345 ();
 DECAPx6_ASAP7_75t_R FILLER_125_371 ();
 DECAPx1_ASAP7_75t_R FILLER_125_385 ();
 DECAPx1_ASAP7_75t_R FILLER_125_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_409 ();
 DECAPx2_ASAP7_75t_R FILLER_125_426 ();
 FILLER_ASAP7_75t_R FILLER_125_432 ();
 DECAPx2_ASAP7_75t_R FILLER_125_450 ();
 FILLER_ASAP7_75t_R FILLER_125_456 ();
 DECAPx2_ASAP7_75t_R FILLER_125_468 ();
 DECAPx6_ASAP7_75t_R FILLER_125_508 ();
 DECAPx1_ASAP7_75t_R FILLER_125_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_526 ();
 FILLER_ASAP7_75t_R FILLER_125_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_584 ();
 FILLER_ASAP7_75t_R FILLER_125_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_600 ();
 DECAPx10_ASAP7_75t_R FILLER_125_607 ();
 DECAPx4_ASAP7_75t_R FILLER_125_629 ();
 FILLER_ASAP7_75t_R FILLER_125_639 ();
 DECAPx2_ASAP7_75t_R FILLER_125_647 ();
 FILLER_ASAP7_75t_R FILLER_125_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_655 ();
 DECAPx2_ASAP7_75t_R FILLER_125_664 ();
 DECAPx10_ASAP7_75t_R FILLER_125_684 ();
 FILLER_ASAP7_75t_R FILLER_125_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_708 ();
 DECAPx10_ASAP7_75t_R FILLER_125_729 ();
 DECAPx10_ASAP7_75t_R FILLER_125_751 ();
 DECAPx1_ASAP7_75t_R FILLER_125_773 ();
 DECAPx10_ASAP7_75t_R FILLER_125_797 ();
 DECAPx6_ASAP7_75t_R FILLER_125_819 ();
 DECAPx2_ASAP7_75t_R FILLER_125_833 ();
 FILLER_ASAP7_75t_R FILLER_125_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_869 ();
 DECAPx2_ASAP7_75t_R FILLER_125_884 ();
 FILLER_ASAP7_75t_R FILLER_125_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_904 ();
 FILLER_ASAP7_75t_R FILLER_125_911 ();
 FILLER_ASAP7_75t_R FILLER_125_919 ();
 FILLER_ASAP7_75t_R FILLER_125_926 ();
 FILLER_ASAP7_75t_R FILLER_125_939 ();
 DECAPx6_ASAP7_75t_R FILLER_125_949 ();
 FILLER_ASAP7_75t_R FILLER_125_963 ();
 FILLER_ASAP7_75t_R FILLER_125_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_973 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1031 ();
 FILLER_ASAP7_75t_R FILLER_125_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1090 ();
 FILLER_ASAP7_75t_R FILLER_125_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1098 ();
 FILLER_ASAP7_75t_R FILLER_125_1102 ();
 FILLER_ASAP7_75t_R FILLER_125_1110 ();
 FILLER_ASAP7_75t_R FILLER_125_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1149 ();
 FILLER_ASAP7_75t_R FILLER_125_1163 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_126_2 ();
 DECAPx10_ASAP7_75t_R FILLER_126_24 ();
 DECAPx10_ASAP7_75t_R FILLER_126_46 ();
 FILLER_ASAP7_75t_R FILLER_126_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_70 ();
 DECAPx2_ASAP7_75t_R FILLER_126_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_99 ();
 DECAPx4_ASAP7_75t_R FILLER_126_106 ();
 FILLER_ASAP7_75t_R FILLER_126_116 ();
 DECAPx1_ASAP7_75t_R FILLER_126_125 ();
 FILLER_ASAP7_75t_R FILLER_126_136 ();
 DECAPx6_ASAP7_75t_R FILLER_126_168 ();
 DECAPx1_ASAP7_75t_R FILLER_126_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_186 ();
 DECAPx2_ASAP7_75t_R FILLER_126_200 ();
 FILLER_ASAP7_75t_R FILLER_126_206 ();
 DECAPx6_ASAP7_75t_R FILLER_126_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_239 ();
 DECAPx2_ASAP7_75t_R FILLER_126_246 ();
 FILLER_ASAP7_75t_R FILLER_126_252 ();
 DECAPx2_ASAP7_75t_R FILLER_126_276 ();
 FILLER_ASAP7_75t_R FILLER_126_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_284 ();
 DECAPx1_ASAP7_75t_R FILLER_126_288 ();
 DECAPx2_ASAP7_75t_R FILLER_126_306 ();
 FILLER_ASAP7_75t_R FILLER_126_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_325 ();
 DECAPx4_ASAP7_75t_R FILLER_126_332 ();
 FILLER_ASAP7_75t_R FILLER_126_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_344 ();
 DECAPx2_ASAP7_75t_R FILLER_126_386 ();
 FILLER_ASAP7_75t_R FILLER_126_392 ();
 FILLER_ASAP7_75t_R FILLER_126_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_408 ();
 DECAPx6_ASAP7_75t_R FILLER_126_415 ();
 DECAPx1_ASAP7_75t_R FILLER_126_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_433 ();
 DECAPx2_ASAP7_75t_R FILLER_126_464 ();
 FILLER_ASAP7_75t_R FILLER_126_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_497 ();
 DECAPx10_ASAP7_75t_R FILLER_126_504 ();
 DECAPx6_ASAP7_75t_R FILLER_126_526 ();
 DECAPx2_ASAP7_75t_R FILLER_126_540 ();
 DECAPx4_ASAP7_75t_R FILLER_126_585 ();
 FILLER_ASAP7_75t_R FILLER_126_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_597 ();
 DECAPx4_ASAP7_75t_R FILLER_126_604 ();
 FILLER_ASAP7_75t_R FILLER_126_614 ();
 DECAPx4_ASAP7_75t_R FILLER_126_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_644 ();
 DECAPx2_ASAP7_75t_R FILLER_126_651 ();
 FILLER_ASAP7_75t_R FILLER_126_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_678 ();
 DECAPx6_ASAP7_75t_R FILLER_126_685 ();
 DECAPx2_ASAP7_75t_R FILLER_126_699 ();
 DECAPx4_ASAP7_75t_R FILLER_126_725 ();
 FILLER_ASAP7_75t_R FILLER_126_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_737 ();
 DECAPx6_ASAP7_75t_R FILLER_126_782 ();
 FILLER_ASAP7_75t_R FILLER_126_816 ();
 DECAPx10_ASAP7_75t_R FILLER_126_838 ();
 DECAPx2_ASAP7_75t_R FILLER_126_882 ();
 FILLER_ASAP7_75t_R FILLER_126_888 ();
 DECAPx4_ASAP7_75t_R FILLER_126_896 ();
 DECAPx6_ASAP7_75t_R FILLER_126_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_946 ();
 DECAPx1_ASAP7_75t_R FILLER_126_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_959 ();
 FILLER_ASAP7_75t_R FILLER_126_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_990 ();
 DECAPx6_ASAP7_75t_R FILLER_126_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1017 ();
 FILLER_ASAP7_75t_R FILLER_126_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_126_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1059 ();
 DECAPx6_ASAP7_75t_R FILLER_126_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1136 ();
 DECAPx6_ASAP7_75t_R FILLER_126_1158 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1179 ();
 FILLER_ASAP7_75t_R FILLER_126_1189 ();
 FILLER_ASAP7_75t_R FILLER_126_1197 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1212 ();
 FILLER_ASAP7_75t_R FILLER_126_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_127_2 ();
 DECAPx10_ASAP7_75t_R FILLER_127_24 ();
 DECAPx10_ASAP7_75t_R FILLER_127_46 ();
 DECAPx4_ASAP7_75t_R FILLER_127_68 ();
 FILLER_ASAP7_75t_R FILLER_127_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_80 ();
 DECAPx2_ASAP7_75t_R FILLER_127_87 ();
 FILLER_ASAP7_75t_R FILLER_127_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_101 ();
 DECAPx6_ASAP7_75t_R FILLER_127_110 ();
 DECAPx2_ASAP7_75t_R FILLER_127_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_130 ();
 DECAPx4_ASAP7_75t_R FILLER_127_143 ();
 FILLER_ASAP7_75t_R FILLER_127_153 ();
 DECAPx4_ASAP7_75t_R FILLER_127_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_180 ();
 DECAPx2_ASAP7_75t_R FILLER_127_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_207 ();
 DECAPx6_ASAP7_75t_R FILLER_127_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_232 ();
 DECAPx2_ASAP7_75t_R FILLER_127_239 ();
 DECAPx10_ASAP7_75t_R FILLER_127_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_273 ();
 DECAPx10_ASAP7_75t_R FILLER_127_286 ();
 FILLER_ASAP7_75t_R FILLER_127_308 ();
 FILLER_ASAP7_75t_R FILLER_127_316 ();
 FILLER_ASAP7_75t_R FILLER_127_344 ();
 FILLER_ASAP7_75t_R FILLER_127_352 ();
 DECAPx2_ASAP7_75t_R FILLER_127_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_399 ();
 DECAPx10_ASAP7_75t_R FILLER_127_406 ();
 DECAPx2_ASAP7_75t_R FILLER_127_428 ();
 FILLER_ASAP7_75t_R FILLER_127_434 ();
 DECAPx2_ASAP7_75t_R FILLER_127_442 ();
 DECAPx2_ASAP7_75t_R FILLER_127_454 ();
 FILLER_ASAP7_75t_R FILLER_127_460 ();
 DECAPx6_ASAP7_75t_R FILLER_127_474 ();
 FILLER_ASAP7_75t_R FILLER_127_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_507 ();
 DECAPx10_ASAP7_75t_R FILLER_127_515 ();
 DECAPx2_ASAP7_75t_R FILLER_127_537 ();
 FILLER_ASAP7_75t_R FILLER_127_553 ();
 DECAPx2_ASAP7_75t_R FILLER_127_563 ();
 DECAPx6_ASAP7_75t_R FILLER_127_578 ();
 DECAPx1_ASAP7_75t_R FILLER_127_605 ();
 FILLER_ASAP7_75t_R FILLER_127_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_623 ();
 DECAPx4_ASAP7_75t_R FILLER_127_644 ();
 DECAPx2_ASAP7_75t_R FILLER_127_660 ();
 DECAPx1_ASAP7_75t_R FILLER_127_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_676 ();
 FILLER_ASAP7_75t_R FILLER_127_685 ();
 DECAPx2_ASAP7_75t_R FILLER_127_737 ();
 FILLER_ASAP7_75t_R FILLER_127_743 ();
 DECAPx10_ASAP7_75t_R FILLER_127_789 ();
 DECAPx10_ASAP7_75t_R FILLER_127_811 ();
 DECAPx6_ASAP7_75t_R FILLER_127_833 ();
 DECAPx1_ASAP7_75t_R FILLER_127_847 ();
 DECAPx2_ASAP7_75t_R FILLER_127_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_908 ();
 DECAPx2_ASAP7_75t_R FILLER_127_915 ();
 FILLER_ASAP7_75t_R FILLER_127_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_923 ();
 DECAPx4_ASAP7_75t_R FILLER_127_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_936 ();
 DECAPx10_ASAP7_75t_R FILLER_127_959 ();
 DECAPx2_ASAP7_75t_R FILLER_127_981 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1015 ();
 FILLER_ASAP7_75t_R FILLER_127_1021 ();
 FILLER_ASAP7_75t_R FILLER_127_1029 ();
 FILLER_ASAP7_75t_R FILLER_127_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1042 ();
 FILLER_ASAP7_75t_R FILLER_127_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1066 ();
 DECAPx6_ASAP7_75t_R FILLER_127_1090 ();
 FILLER_ASAP7_75t_R FILLER_127_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_127_1135 ();
 FILLER_ASAP7_75t_R FILLER_127_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1157 ();
 FILLER_ASAP7_75t_R FILLER_127_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1189 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1210 ();
 FILLER_ASAP7_75t_R FILLER_127_1216 ();
 DECAPx4_ASAP7_75t_R FILLER_128_2 ();
 DECAPx10_ASAP7_75t_R FILLER_128_24 ();
 DECAPx10_ASAP7_75t_R FILLER_128_46 ();
 DECAPx4_ASAP7_75t_R FILLER_128_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_78 ();
 DECAPx1_ASAP7_75t_R FILLER_128_85 ();
 DECAPx1_ASAP7_75t_R FILLER_128_100 ();
 DECAPx6_ASAP7_75t_R FILLER_128_115 ();
 FILLER_ASAP7_75t_R FILLER_128_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_131 ();
 DECAPx2_ASAP7_75t_R FILLER_128_140 ();
 FILLER_ASAP7_75t_R FILLER_128_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_171 ();
 DECAPx10_ASAP7_75t_R FILLER_128_194 ();
 DECAPx6_ASAP7_75t_R FILLER_128_216 ();
 FILLER_ASAP7_75t_R FILLER_128_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_232 ();
 DECAPx4_ASAP7_75t_R FILLER_128_292 ();
 FILLER_ASAP7_75t_R FILLER_128_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_304 ();
 DECAPx1_ASAP7_75t_R FILLER_128_317 ();
 DECAPx6_ASAP7_75t_R FILLER_128_334 ();
 DECAPx1_ASAP7_75t_R FILLER_128_348 ();
 DECAPx6_ASAP7_75t_R FILLER_128_358 ();
 FILLER_ASAP7_75t_R FILLER_128_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_410 ();
 FILLER_ASAP7_75t_R FILLER_128_417 ();
 DECAPx2_ASAP7_75t_R FILLER_128_425 ();
 FILLER_ASAP7_75t_R FILLER_128_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_433 ();
 FILLER_ASAP7_75t_R FILLER_128_440 ();
 DECAPx2_ASAP7_75t_R FILLER_128_456 ();
 DECAPx2_ASAP7_75t_R FILLER_128_475 ();
 FILLER_ASAP7_75t_R FILLER_128_481 ();
 DECAPx2_ASAP7_75t_R FILLER_128_503 ();
 FILLER_ASAP7_75t_R FILLER_128_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_511 ();
 FILLER_ASAP7_75t_R FILLER_128_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_521 ();
 FILLER_ASAP7_75t_R FILLER_128_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_549 ();
 FILLER_ASAP7_75t_R FILLER_128_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_590 ();
 DECAPx10_ASAP7_75t_R FILLER_128_599 ();
 DECAPx2_ASAP7_75t_R FILLER_128_621 ();
 DECAPx1_ASAP7_75t_R FILLER_128_641 ();
 DECAPx2_ASAP7_75t_R FILLER_128_651 ();
 FILLER_ASAP7_75t_R FILLER_128_657 ();
 FILLER_ASAP7_75t_R FILLER_128_671 ();
 DECAPx1_ASAP7_75t_R FILLER_128_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_683 ();
 DECAPx10_ASAP7_75t_R FILLER_128_692 ();
 DECAPx10_ASAP7_75t_R FILLER_128_714 ();
 DECAPx6_ASAP7_75t_R FILLER_128_736 ();
 FILLER_ASAP7_75t_R FILLER_128_750 ();
 FILLER_ASAP7_75t_R FILLER_128_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_796 ();
 DECAPx10_ASAP7_75t_R FILLER_128_839 ();
 FILLER_ASAP7_75t_R FILLER_128_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_886 ();
 DECAPx2_ASAP7_75t_R FILLER_128_899 ();
 FILLER_ASAP7_75t_R FILLER_128_905 ();
 DECAPx10_ASAP7_75t_R FILLER_128_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_937 ();
 FILLER_ASAP7_75t_R FILLER_128_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_948 ();
 DECAPx6_ASAP7_75t_R FILLER_128_967 ();
 DECAPx4_ASAP7_75t_R FILLER_128_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1013 ();
 FILLER_ASAP7_75t_R FILLER_128_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1025 ();
 FILLER_ASAP7_75t_R FILLER_128_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1049 ();
 FILLER_ASAP7_75t_R FILLER_128_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1076 ();
 FILLER_ASAP7_75t_R FILLER_128_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1110 ();
 FILLER_ASAP7_75t_R FILLER_128_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1170 ();
 FILLER_ASAP7_75t_R FILLER_128_1178 ();
 FILLER_ASAP7_75t_R FILLER_128_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1215 ();
 FILLER_ASAP7_75t_R FILLER_128_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_129_2 ();
 DECAPx10_ASAP7_75t_R FILLER_129_24 ();
 DECAPx10_ASAP7_75t_R FILLER_129_46 ();
 DECAPx2_ASAP7_75t_R FILLER_129_68 ();
 FILLER_ASAP7_75t_R FILLER_129_74 ();
 DECAPx2_ASAP7_75t_R FILLER_129_98 ();
 FILLER_ASAP7_75t_R FILLER_129_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_150 ();
 DECAPx10_ASAP7_75t_R FILLER_129_159 ();
 DECAPx4_ASAP7_75t_R FILLER_129_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_191 ();
 DECAPx10_ASAP7_75t_R FILLER_129_195 ();
 DECAPx10_ASAP7_75t_R FILLER_129_217 ();
 DECAPx4_ASAP7_75t_R FILLER_129_239 ();
 FILLER_ASAP7_75t_R FILLER_129_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_277 ();
 FILLER_ASAP7_75t_R FILLER_129_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_298 ();
 FILLER_ASAP7_75t_R FILLER_129_305 ();
 DECAPx1_ASAP7_75t_R FILLER_129_318 ();
 DECAPx2_ASAP7_75t_R FILLER_129_336 ();
 DECAPx10_ASAP7_75t_R FILLER_129_348 ();
 DECAPx10_ASAP7_75t_R FILLER_129_370 ();
 DECAPx1_ASAP7_75t_R FILLER_129_392 ();
 FILLER_ASAP7_75t_R FILLER_129_402 ();
 DECAPx1_ASAP7_75t_R FILLER_129_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_414 ();
 DECAPx4_ASAP7_75t_R FILLER_129_423 ();
 FILLER_ASAP7_75t_R FILLER_129_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_435 ();
 DECAPx10_ASAP7_75t_R FILLER_129_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_466 ();
 DECAPx1_ASAP7_75t_R FILLER_129_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_477 ();
 DECAPx2_ASAP7_75t_R FILLER_129_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_506 ();
 DECAPx6_ASAP7_75t_R FILLER_129_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_529 ();
 DECAPx4_ASAP7_75t_R FILLER_129_536 ();
 FILLER_ASAP7_75t_R FILLER_129_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_554 ();
 FILLER_ASAP7_75t_R FILLER_129_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_569 ();
 DECAPx4_ASAP7_75t_R FILLER_129_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_586 ();
 DECAPx6_ASAP7_75t_R FILLER_129_595 ();
 DECAPx2_ASAP7_75t_R FILLER_129_609 ();
 DECAPx6_ASAP7_75t_R FILLER_129_625 ();
 DECAPx2_ASAP7_75t_R FILLER_129_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_657 ();
 FILLER_ASAP7_75t_R FILLER_129_666 ();
 DECAPx10_ASAP7_75t_R FILLER_129_676 ();
 DECAPx6_ASAP7_75t_R FILLER_129_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_712 ();
 DECAPx2_ASAP7_75t_R FILLER_129_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_741 ();
 DECAPx4_ASAP7_75t_R FILLER_129_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_758 ();
 DECAPx2_ASAP7_75t_R FILLER_129_792 ();
 FILLER_ASAP7_75t_R FILLER_129_798 ();
 DECAPx1_ASAP7_75t_R FILLER_129_813 ();
 FILLER_ASAP7_75t_R FILLER_129_837 ();
 DECAPx10_ASAP7_75t_R FILLER_129_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_864 ();
 DECAPx6_ASAP7_75t_R FILLER_129_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_901 ();
 DECAPx2_ASAP7_75t_R FILLER_129_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_942 ();
 DECAPx10_ASAP7_75t_R FILLER_129_953 ();
 DECAPx10_ASAP7_75t_R FILLER_129_975 ();
 DECAPx4_ASAP7_75t_R FILLER_129_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1007 ();
 FILLER_ASAP7_75t_R FILLER_129_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1031 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_129_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1111 ();
 FILLER_ASAP7_75t_R FILLER_129_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1134 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1141 ();
 FILLER_ASAP7_75t_R FILLER_129_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1153 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1175 ();
 FILLER_ASAP7_75t_R FILLER_129_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_130_2 ();
 DECAPx10_ASAP7_75t_R FILLER_130_24 ();
 DECAPx10_ASAP7_75t_R FILLER_130_46 ();
 DECAPx6_ASAP7_75t_R FILLER_130_68 ();
 FILLER_ASAP7_75t_R FILLER_130_82 ();
 DECAPx2_ASAP7_75t_R FILLER_130_101 ();
 FILLER_ASAP7_75t_R FILLER_130_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_109 ();
 DECAPx6_ASAP7_75t_R FILLER_130_116 ();
 DECAPx2_ASAP7_75t_R FILLER_130_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_136 ();
 DECAPx2_ASAP7_75t_R FILLER_130_148 ();
 DECAPx6_ASAP7_75t_R FILLER_130_171 ();
 DECAPx1_ASAP7_75t_R FILLER_130_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_212 ();
 DECAPx10_ASAP7_75t_R FILLER_130_216 ();
 DECAPx10_ASAP7_75t_R FILLER_130_238 ();
 DECAPx4_ASAP7_75t_R FILLER_130_260 ();
 FILLER_ASAP7_75t_R FILLER_130_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_293 ();
 FILLER_ASAP7_75t_R FILLER_130_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_318 ();
 DECAPx10_ASAP7_75t_R FILLER_130_334 ();
 DECAPx10_ASAP7_75t_R FILLER_130_356 ();
 DECAPx6_ASAP7_75t_R FILLER_130_378 ();
 DECAPx2_ASAP7_75t_R FILLER_130_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_398 ();
 DECAPx4_ASAP7_75t_R FILLER_130_407 ();
 FILLER_ASAP7_75t_R FILLER_130_417 ();
 DECAPx4_ASAP7_75t_R FILLER_130_425 ();
 FILLER_ASAP7_75t_R FILLER_130_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_443 ();
 DECAPx4_ASAP7_75t_R FILLER_130_464 ();
 FILLER_ASAP7_75t_R FILLER_130_488 ();
 DECAPx4_ASAP7_75t_R FILLER_130_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_507 ();
 DECAPx4_ASAP7_75t_R FILLER_130_518 ();
 FILLER_ASAP7_75t_R FILLER_130_528 ();
 FILLER_ASAP7_75t_R FILLER_130_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_562 ();
 FILLER_ASAP7_75t_R FILLER_130_579 ();
 DECAPx6_ASAP7_75t_R FILLER_130_598 ();
 FILLER_ASAP7_75t_R FILLER_130_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_624 ();
 DECAPx1_ASAP7_75t_R FILLER_130_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_641 ();
 DECAPx1_ASAP7_75t_R FILLER_130_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_660 ();
 FILLER_ASAP7_75t_R FILLER_130_673 ();
 DECAPx2_ASAP7_75t_R FILLER_130_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_736 ();
 DECAPx10_ASAP7_75t_R FILLER_130_750 ();
 DECAPx1_ASAP7_75t_R FILLER_130_772 ();
 DECAPx2_ASAP7_75t_R FILLER_130_788 ();
 FILLER_ASAP7_75t_R FILLER_130_794 ();
 FILLER_ASAP7_75t_R FILLER_130_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_817 ();
 FILLER_ASAP7_75t_R FILLER_130_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_840 ();
 FILLER_ASAP7_75t_R FILLER_130_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_863 ();
 DECAPx10_ASAP7_75t_R FILLER_130_870 ();
 DECAPx1_ASAP7_75t_R FILLER_130_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_916 ();
 DECAPx1_ASAP7_75t_R FILLER_130_936 ();
 DECAPx6_ASAP7_75t_R FILLER_130_950 ();
 DECAPx2_ASAP7_75t_R FILLER_130_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_993 ();
 DECAPx4_ASAP7_75t_R FILLER_130_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1102 ();
 DECAPx4_ASAP7_75t_R FILLER_130_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_130_1131 ();
 FILLER_ASAP7_75t_R FILLER_130_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1223 ();
 DECAPx1_ASAP7_75t_R FILLER_131_2 ();
 DECAPx10_ASAP7_75t_R FILLER_131_12 ();
 DECAPx10_ASAP7_75t_R FILLER_131_34 ();
 DECAPx10_ASAP7_75t_R FILLER_131_56 ();
 DECAPx6_ASAP7_75t_R FILLER_131_78 ();
 DECAPx1_ASAP7_75t_R FILLER_131_150 ();
 DECAPx2_ASAP7_75t_R FILLER_131_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_166 ();
 DECAPx6_ASAP7_75t_R FILLER_131_189 ();
 DECAPx1_ASAP7_75t_R FILLER_131_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_207 ();
 DECAPx4_ASAP7_75t_R FILLER_131_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_238 ();
 DECAPx6_ASAP7_75t_R FILLER_131_265 ();
 FILLER_ASAP7_75t_R FILLER_131_279 ();
 DECAPx2_ASAP7_75t_R FILLER_131_288 ();
 FILLER_ASAP7_75t_R FILLER_131_294 ();
 DECAPx1_ASAP7_75t_R FILLER_131_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_316 ();
 FILLER_ASAP7_75t_R FILLER_131_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_334 ();
 DECAPx10_ASAP7_75t_R FILLER_131_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_399 ();
 FILLER_ASAP7_75t_R FILLER_131_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_414 ();
 DECAPx2_ASAP7_75t_R FILLER_131_427 ();
 FILLER_ASAP7_75t_R FILLER_131_433 ();
 FILLER_ASAP7_75t_R FILLER_131_451 ();
 DECAPx4_ASAP7_75t_R FILLER_131_459 ();
 DECAPx4_ASAP7_75t_R FILLER_131_475 ();
 FILLER_ASAP7_75t_R FILLER_131_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_487 ();
 DECAPx1_ASAP7_75t_R FILLER_131_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_502 ();
 DECAPx6_ASAP7_75t_R FILLER_131_520 ();
 DECAPx2_ASAP7_75t_R FILLER_131_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_570 ();
 FILLER_ASAP7_75t_R FILLER_131_577 ();
 FILLER_ASAP7_75t_R FILLER_131_587 ();
 FILLER_ASAP7_75t_R FILLER_131_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_597 ();
 DECAPx2_ASAP7_75t_R FILLER_131_606 ();
 FILLER_ASAP7_75t_R FILLER_131_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_614 ();
 DECAPx4_ASAP7_75t_R FILLER_131_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_643 ();
 DECAPx2_ASAP7_75t_R FILLER_131_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_678 ();
 DECAPx6_ASAP7_75t_R FILLER_131_715 ();
 FILLER_ASAP7_75t_R FILLER_131_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_731 ();
 DECAPx1_ASAP7_75t_R FILLER_131_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_756 ();
 DECAPx1_ASAP7_75t_R FILLER_131_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_771 ();
 FILLER_ASAP7_75t_R FILLER_131_794 ();
 DECAPx10_ASAP7_75t_R FILLER_131_802 ();
 DECAPx6_ASAP7_75t_R FILLER_131_824 ();
 FILLER_ASAP7_75t_R FILLER_131_838 ();
 DECAPx10_ASAP7_75t_R FILLER_131_860 ();
 DECAPx6_ASAP7_75t_R FILLER_131_882 ();
 DECAPx6_ASAP7_75t_R FILLER_131_906 ();
 DECAPx1_ASAP7_75t_R FILLER_131_920 ();
 DECAPx6_ASAP7_75t_R FILLER_131_926 ();
 FILLER_ASAP7_75t_R FILLER_131_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_942 ();
 DECAPx4_ASAP7_75t_R FILLER_131_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_131_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1098 ();
 FILLER_ASAP7_75t_R FILLER_131_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1106 ();
 FILLER_ASAP7_75t_R FILLER_131_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_131_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1167 ();
 FILLER_ASAP7_75t_R FILLER_131_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_132_2 ();
 DECAPx10_ASAP7_75t_R FILLER_132_24 ();
 DECAPx10_ASAP7_75t_R FILLER_132_46 ();
 DECAPx10_ASAP7_75t_R FILLER_132_68 ();
 DECAPx10_ASAP7_75t_R FILLER_132_90 ();
 DECAPx10_ASAP7_75t_R FILLER_132_112 ();
 DECAPx6_ASAP7_75t_R FILLER_132_134 ();
 FILLER_ASAP7_75t_R FILLER_132_148 ();
 DECAPx4_ASAP7_75t_R FILLER_132_167 ();
 FILLER_ASAP7_75t_R FILLER_132_177 ();
 DECAPx10_ASAP7_75t_R FILLER_132_189 ();
 DECAPx6_ASAP7_75t_R FILLER_132_211 ();
 DECAPx1_ASAP7_75t_R FILLER_132_225 ();
 DECAPx4_ASAP7_75t_R FILLER_132_249 ();
 DECAPx6_ASAP7_75t_R FILLER_132_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_298 ();
 DECAPx6_ASAP7_75t_R FILLER_132_310 ();
 DECAPx4_ASAP7_75t_R FILLER_132_338 ();
 DECAPx10_ASAP7_75t_R FILLER_132_361 ();
 DECAPx6_ASAP7_75t_R FILLER_132_383 ();
 FILLER_ASAP7_75t_R FILLER_132_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_399 ();
 FILLER_ASAP7_75t_R FILLER_132_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_416 ();
 DECAPx2_ASAP7_75t_R FILLER_132_425 ();
 FILLER_ASAP7_75t_R FILLER_132_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_433 ();
 DECAPx4_ASAP7_75t_R FILLER_132_442 ();
 FILLER_ASAP7_75t_R FILLER_132_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_466 ();
 FILLER_ASAP7_75t_R FILLER_132_483 ();
 DECAPx1_ASAP7_75t_R FILLER_132_499 ();
 DECAPx10_ASAP7_75t_R FILLER_132_519 ();
 DECAPx10_ASAP7_75t_R FILLER_132_541 ();
 FILLER_ASAP7_75t_R FILLER_132_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_565 ();
 DECAPx1_ASAP7_75t_R FILLER_132_579 ();
 DECAPx6_ASAP7_75t_R FILLER_132_589 ();
 DECAPx2_ASAP7_75t_R FILLER_132_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_609 ();
 DECAPx10_ASAP7_75t_R FILLER_132_620 ();
 DECAPx6_ASAP7_75t_R FILLER_132_642 ();
 DECAPx1_ASAP7_75t_R FILLER_132_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_660 ();
 DECAPx10_ASAP7_75t_R FILLER_132_675 ();
 DECAPx10_ASAP7_75t_R FILLER_132_697 ();
 DECAPx2_ASAP7_75t_R FILLER_132_719 ();
 FILLER_ASAP7_75t_R FILLER_132_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_727 ();
 FILLER_ASAP7_75t_R FILLER_132_734 ();
 DECAPx4_ASAP7_75t_R FILLER_132_744 ();
 DECAPx1_ASAP7_75t_R FILLER_132_774 ();
 DECAPx2_ASAP7_75t_R FILLER_132_786 ();
 FILLER_ASAP7_75t_R FILLER_132_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_801 ();
 FILLER_ASAP7_75t_R FILLER_132_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_810 ();
 DECAPx6_ASAP7_75t_R FILLER_132_818 ();
 DECAPx1_ASAP7_75t_R FILLER_132_832 ();
 DECAPx1_ASAP7_75t_R FILLER_132_858 ();
 DECAPx2_ASAP7_75t_R FILLER_132_868 ();
 FILLER_ASAP7_75t_R FILLER_132_874 ();
 FILLER_ASAP7_75t_R FILLER_132_904 ();
 DECAPx1_ASAP7_75t_R FILLER_132_920 ();
 DECAPx2_ASAP7_75t_R FILLER_132_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_936 ();
 DECAPx4_ASAP7_75t_R FILLER_132_950 ();
 FILLER_ASAP7_75t_R FILLER_132_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_962 ();
 DECAPx1_ASAP7_75t_R FILLER_132_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_989 ();
 DECAPx4_ASAP7_75t_R FILLER_132_998 ();
 FILLER_ASAP7_75t_R FILLER_132_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1054 ();
 FILLER_ASAP7_75t_R FILLER_132_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1062 ();
 FILLER_ASAP7_75t_R FILLER_132_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1092 ();
 FILLER_ASAP7_75t_R FILLER_132_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1100 ();
 FILLER_ASAP7_75t_R FILLER_132_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1186 ();
 FILLER_ASAP7_75t_R FILLER_132_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1205 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_133_8 ();
 DECAPx10_ASAP7_75t_R FILLER_133_30 ();
 DECAPx10_ASAP7_75t_R FILLER_133_52 ();
 DECAPx10_ASAP7_75t_R FILLER_133_74 ();
 DECAPx10_ASAP7_75t_R FILLER_133_96 ();
 DECAPx10_ASAP7_75t_R FILLER_133_118 ();
 DECAPx6_ASAP7_75t_R FILLER_133_140 ();
 DECAPx2_ASAP7_75t_R FILLER_133_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_160 ();
 DECAPx10_ASAP7_75t_R FILLER_133_191 ();
 DECAPx10_ASAP7_75t_R FILLER_133_213 ();
 DECAPx2_ASAP7_75t_R FILLER_133_235 ();
 FILLER_ASAP7_75t_R FILLER_133_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_264 ();
 DECAPx2_ASAP7_75t_R FILLER_133_293 ();
 FILLER_ASAP7_75t_R FILLER_133_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_301 ();
 DECAPx2_ASAP7_75t_R FILLER_133_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_319 ();
 DECAPx1_ASAP7_75t_R FILLER_133_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_345 ();
 FILLER_ASAP7_75t_R FILLER_133_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_368 ();
 DECAPx4_ASAP7_75t_R FILLER_133_372 ();
 DECAPx6_ASAP7_75t_R FILLER_133_402 ();
 FILLER_ASAP7_75t_R FILLER_133_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_418 ();
 DECAPx2_ASAP7_75t_R FILLER_133_441 ();
 FILLER_ASAP7_75t_R FILLER_133_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_449 ();
 DECAPx1_ASAP7_75t_R FILLER_133_466 ();
 DECAPx2_ASAP7_75t_R FILLER_133_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_488 ();
 DECAPx10_ASAP7_75t_R FILLER_133_529 ();
 DECAPx10_ASAP7_75t_R FILLER_133_551 ();
 DECAPx4_ASAP7_75t_R FILLER_133_573 ();
 FILLER_ASAP7_75t_R FILLER_133_583 ();
 DECAPx2_ASAP7_75t_R FILLER_133_595 ();
 FILLER_ASAP7_75t_R FILLER_133_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_623 ();
 DECAPx2_ASAP7_75t_R FILLER_133_658 ();
 FILLER_ASAP7_75t_R FILLER_133_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_678 ();
 DECAPx10_ASAP7_75t_R FILLER_133_685 ();
 DECAPx6_ASAP7_75t_R FILLER_133_707 ();
 DECAPx2_ASAP7_75t_R FILLER_133_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_727 ();
 DECAPx2_ASAP7_75t_R FILLER_133_758 ();
 FILLER_ASAP7_75t_R FILLER_133_764 ();
 FILLER_ASAP7_75t_R FILLER_133_786 ();
 FILLER_ASAP7_75t_R FILLER_133_804 ();
 DECAPx10_ASAP7_75t_R FILLER_133_814 ();
 FILLER_ASAP7_75t_R FILLER_133_836 ();
 DECAPx2_ASAP7_75t_R FILLER_133_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_866 ();
 DECAPx1_ASAP7_75t_R FILLER_133_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_874 ();
 DECAPx2_ASAP7_75t_R FILLER_133_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_895 ();
 DECAPx2_ASAP7_75t_R FILLER_133_902 ();
 DECAPx4_ASAP7_75t_R FILLER_133_914 ();
 FILLER_ASAP7_75t_R FILLER_133_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_928 ();
 DECAPx2_ASAP7_75t_R FILLER_133_936 ();
 FILLER_ASAP7_75t_R FILLER_133_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_944 ();
 FILLER_ASAP7_75t_R FILLER_133_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_967 ();
 DECAPx2_ASAP7_75t_R FILLER_133_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_997 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1006 ();
 FILLER_ASAP7_75t_R FILLER_133_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_133_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1139 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1150 ();
 DECAPx6_ASAP7_75t_R FILLER_133_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1187 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_134_2 ();
 DECAPx10_ASAP7_75t_R FILLER_134_24 ();
 DECAPx10_ASAP7_75t_R FILLER_134_46 ();
 DECAPx4_ASAP7_75t_R FILLER_134_68 ();
 FILLER_ASAP7_75t_R FILLER_134_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_80 ();
 DECAPx6_ASAP7_75t_R FILLER_134_103 ();
 DECAPx1_ASAP7_75t_R FILLER_134_117 ();
 DECAPx4_ASAP7_75t_R FILLER_134_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_147 ();
 DECAPx10_ASAP7_75t_R FILLER_134_154 ();
 DECAPx10_ASAP7_75t_R FILLER_134_176 ();
 DECAPx10_ASAP7_75t_R FILLER_134_198 ();
 DECAPx10_ASAP7_75t_R FILLER_134_220 ();
 DECAPx4_ASAP7_75t_R FILLER_134_242 ();
 DECAPx2_ASAP7_75t_R FILLER_134_258 ();
 DECAPx4_ASAP7_75t_R FILLER_134_286 ();
 DECAPx4_ASAP7_75t_R FILLER_134_311 ();
 FILLER_ASAP7_75t_R FILLER_134_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_357 ();
 DECAPx6_ASAP7_75t_R FILLER_134_380 ();
 FILLER_ASAP7_75t_R FILLER_134_394 ();
 DECAPx6_ASAP7_75t_R FILLER_134_418 ();
 FILLER_ASAP7_75t_R FILLER_134_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_434 ();
 FILLER_ASAP7_75t_R FILLER_134_447 ();
 FILLER_ASAP7_75t_R FILLER_134_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_461 ();
 DECAPx4_ASAP7_75t_R FILLER_134_464 ();
 DECAPx1_ASAP7_75t_R FILLER_134_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_509 ();
 DECAPx10_ASAP7_75t_R FILLER_134_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_548 ();
 DECAPx10_ASAP7_75t_R FILLER_134_569 ();
 FILLER_ASAP7_75t_R FILLER_134_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_593 ();
 DECAPx1_ASAP7_75t_R FILLER_134_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_620 ();
 DECAPx1_ASAP7_75t_R FILLER_134_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_633 ();
 FILLER_ASAP7_75t_R FILLER_134_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_642 ();
 FILLER_ASAP7_75t_R FILLER_134_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_667 ();
 DECAPx1_ASAP7_75t_R FILLER_134_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_678 ();
 DECAPx4_ASAP7_75t_R FILLER_134_693 ();
 DECAPx6_ASAP7_75t_R FILLER_134_725 ();
 DECAPx1_ASAP7_75t_R FILLER_134_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_743 ();
 DECAPx6_ASAP7_75t_R FILLER_134_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_772 ();
 DECAPx2_ASAP7_75t_R FILLER_134_779 ();
 FILLER_ASAP7_75t_R FILLER_134_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_800 ();
 FILLER_ASAP7_75t_R FILLER_134_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_860 ();
 FILLER_ASAP7_75t_R FILLER_134_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_869 ();
 FILLER_ASAP7_75t_R FILLER_134_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_875 ();
 DECAPx2_ASAP7_75t_R FILLER_134_890 ();
 FILLER_ASAP7_75t_R FILLER_134_896 ();
 DECAPx2_ASAP7_75t_R FILLER_134_918 ();
 FILLER_ASAP7_75t_R FILLER_134_924 ();
 DECAPx1_ASAP7_75t_R FILLER_134_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_938 ();
 DECAPx2_ASAP7_75t_R FILLER_134_955 ();
 DECAPx6_ASAP7_75t_R FILLER_134_967 ();
 FILLER_ASAP7_75t_R FILLER_134_981 ();
 FILLER_ASAP7_75t_R FILLER_134_1015 ();
 FILLER_ASAP7_75t_R FILLER_134_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1045 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1060 ();
 FILLER_ASAP7_75t_R FILLER_134_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_134_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1100 ();
 FILLER_ASAP7_75t_R FILLER_134_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1193 ();
 DECAPx6_ASAP7_75t_R FILLER_135_2 ();
 DECAPx10_ASAP7_75t_R FILLER_135_22 ();
 DECAPx10_ASAP7_75t_R FILLER_135_44 ();
 DECAPx2_ASAP7_75t_R FILLER_135_66 ();
 FILLER_ASAP7_75t_R FILLER_135_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_74 ();
 DECAPx1_ASAP7_75t_R FILLER_135_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_85 ();
 DECAPx4_ASAP7_75t_R FILLER_135_92 ();
 DECAPx4_ASAP7_75t_R FILLER_135_108 ();
 DECAPx10_ASAP7_75t_R FILLER_135_140 ();
 DECAPx10_ASAP7_75t_R FILLER_135_162 ();
 DECAPx10_ASAP7_75t_R FILLER_135_184 ();
 DECAPx10_ASAP7_75t_R FILLER_135_206 ();
 DECAPx10_ASAP7_75t_R FILLER_135_228 ();
 DECAPx6_ASAP7_75t_R FILLER_135_250 ();
 FILLER_ASAP7_75t_R FILLER_135_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_266 ();
 FILLER_ASAP7_75t_R FILLER_135_327 ();
 FILLER_ASAP7_75t_R FILLER_135_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_337 ();
 DECAPx1_ASAP7_75t_R FILLER_135_344 ();
 DECAPx10_ASAP7_75t_R FILLER_135_361 ();
 DECAPx6_ASAP7_75t_R FILLER_135_383 ();
 DECAPx1_ASAP7_75t_R FILLER_135_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_401 ();
 DECAPx4_ASAP7_75t_R FILLER_135_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_434 ();
 FILLER_ASAP7_75t_R FILLER_135_441 ();
 DECAPx4_ASAP7_75t_R FILLER_135_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_504 ();
 FILLER_ASAP7_75t_R FILLER_135_511 ();
 DECAPx4_ASAP7_75t_R FILLER_135_523 ();
 FILLER_ASAP7_75t_R FILLER_135_533 ();
 DECAPx2_ASAP7_75t_R FILLER_135_553 ();
 FILLER_ASAP7_75t_R FILLER_135_559 ();
 DECAPx2_ASAP7_75t_R FILLER_135_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_611 ();
 FILLER_ASAP7_75t_R FILLER_135_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_640 ();
 FILLER_ASAP7_75t_R FILLER_135_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_649 ();
 DECAPx10_ASAP7_75t_R FILLER_135_656 ();
 DECAPx4_ASAP7_75t_R FILLER_135_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_688 ();
 DECAPx1_ASAP7_75t_R FILLER_135_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_721 ();
 DECAPx6_ASAP7_75t_R FILLER_135_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_742 ();
 DECAPx2_ASAP7_75t_R FILLER_135_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_765 ();
 DECAPx1_ASAP7_75t_R FILLER_135_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_789 ();
 FILLER_ASAP7_75t_R FILLER_135_796 ();
 FILLER_ASAP7_75t_R FILLER_135_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_806 ();
 DECAPx10_ASAP7_75t_R FILLER_135_813 ();
 DECAPx1_ASAP7_75t_R FILLER_135_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_839 ();
 DECAPx2_ASAP7_75t_R FILLER_135_862 ();
 FILLER_ASAP7_75t_R FILLER_135_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_870 ();
 DECAPx2_ASAP7_75t_R FILLER_135_885 ();
 FILLER_ASAP7_75t_R FILLER_135_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_900 ();
 DECAPx1_ASAP7_75t_R FILLER_135_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_923 ();
 FILLER_ASAP7_75t_R FILLER_135_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_936 ();
 DECAPx2_ASAP7_75t_R FILLER_135_943 ();
 FILLER_ASAP7_75t_R FILLER_135_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_951 ();
 DECAPx2_ASAP7_75t_R FILLER_135_974 ();
 DECAPx10_ASAP7_75t_R FILLER_135_986 ();
 DECAPx4_ASAP7_75t_R FILLER_135_1008 ();
 FILLER_ASAP7_75t_R FILLER_135_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1063 ();
 FILLER_ASAP7_75t_R FILLER_135_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1174 ();
 FILLER_ASAP7_75t_R FILLER_135_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_136_2 ();
 FILLER_ASAP7_75t_R FILLER_136_24 ();
 DECAPx10_ASAP7_75t_R FILLER_136_32 ();
 DECAPx4_ASAP7_75t_R FILLER_136_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_84 ();
 DECAPx2_ASAP7_75t_R FILLER_136_91 ();
 FILLER_ASAP7_75t_R FILLER_136_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_99 ();
 DECAPx10_ASAP7_75t_R FILLER_136_122 ();
 FILLER_ASAP7_75t_R FILLER_136_144 ();
 DECAPx6_ASAP7_75t_R FILLER_136_172 ();
 DECAPx1_ASAP7_75t_R FILLER_136_186 ();
 DECAPx10_ASAP7_75t_R FILLER_136_212 ();
 DECAPx4_ASAP7_75t_R FILLER_136_234 ();
 DECAPx2_ASAP7_75t_R FILLER_136_269 ();
 FILLER_ASAP7_75t_R FILLER_136_275 ();
 FILLER_ASAP7_75t_R FILLER_136_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_321 ();
 DECAPx10_ASAP7_75t_R FILLER_136_346 ();
 DECAPx10_ASAP7_75t_R FILLER_136_368 ();
 DECAPx10_ASAP7_75t_R FILLER_136_390 ();
 DECAPx1_ASAP7_75t_R FILLER_136_412 ();
 DECAPx4_ASAP7_75t_R FILLER_136_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_451 ();
 DECAPx1_ASAP7_75t_R FILLER_136_458 ();
 DECAPx4_ASAP7_75t_R FILLER_136_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_474 ();
 DECAPx2_ASAP7_75t_R FILLER_136_489 ();
 DECAPx1_ASAP7_75t_R FILLER_136_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_518 ();
 DECAPx10_ASAP7_75t_R FILLER_136_525 ();
 DECAPx4_ASAP7_75t_R FILLER_136_547 ();
 FILLER_ASAP7_75t_R FILLER_136_557 ();
 DECAPx2_ASAP7_75t_R FILLER_136_581 ();
 FILLER_ASAP7_75t_R FILLER_136_587 ();
 FILLER_ASAP7_75t_R FILLER_136_609 ();
 DECAPx1_ASAP7_75t_R FILLER_136_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_637 ();
 FILLER_ASAP7_75t_R FILLER_136_652 ();
 DECAPx6_ASAP7_75t_R FILLER_136_660 ();
 DECAPx2_ASAP7_75t_R FILLER_136_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_680 ();
 FILLER_ASAP7_75t_R FILLER_136_701 ();
 DECAPx6_ASAP7_75t_R FILLER_136_723 ();
 FILLER_ASAP7_75t_R FILLER_136_737 ();
 DECAPx4_ASAP7_75t_R FILLER_136_749 ();
 DECAPx2_ASAP7_75t_R FILLER_136_773 ();
 FILLER_ASAP7_75t_R FILLER_136_779 ();
 DECAPx2_ASAP7_75t_R FILLER_136_789 ();
 FILLER_ASAP7_75t_R FILLER_136_795 ();
 DECAPx2_ASAP7_75t_R FILLER_136_803 ();
 DECAPx10_ASAP7_75t_R FILLER_136_831 ();
 DECAPx6_ASAP7_75t_R FILLER_136_853 ();
 DECAPx6_ASAP7_75t_R FILLER_136_885 ();
 FILLER_ASAP7_75t_R FILLER_136_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_905 ();
 DECAPx1_ASAP7_75t_R FILLER_136_916 ();
 FILLER_ASAP7_75t_R FILLER_136_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_943 ();
 DECAPx10_ASAP7_75t_R FILLER_136_951 ();
 DECAPx1_ASAP7_75t_R FILLER_136_993 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1008 ();
 FILLER_ASAP7_75t_R FILLER_136_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1016 ();
 FILLER_ASAP7_75t_R FILLER_136_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1062 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1090 ();
 DECAPx6_ASAP7_75t_R FILLER_136_1094 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1176 ();
 FILLER_ASAP7_75t_R FILLER_136_1182 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1204 ();
 FILLER_ASAP7_75t_R FILLER_136_1214 ();
 FILLER_ASAP7_75t_R FILLER_136_1222 ();
 DECAPx4_ASAP7_75t_R FILLER_137_2 ();
 DECAPx10_ASAP7_75t_R FILLER_137_18 ();
 DECAPx10_ASAP7_75t_R FILLER_137_40 ();
 DECAPx4_ASAP7_75t_R FILLER_137_62 ();
 FILLER_ASAP7_75t_R FILLER_137_72 ();
 DECAPx6_ASAP7_75t_R FILLER_137_86 ();
 FILLER_ASAP7_75t_R FILLER_137_100 ();
 DECAPx1_ASAP7_75t_R FILLER_137_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_114 ();
 DECAPx6_ASAP7_75t_R FILLER_137_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_151 ();
 DECAPx2_ASAP7_75t_R FILLER_137_185 ();
 DECAPx2_ASAP7_75t_R FILLER_137_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_203 ();
 FILLER_ASAP7_75t_R FILLER_137_226 ();
 DECAPx2_ASAP7_75t_R FILLER_137_264 ();
 FILLER_ASAP7_75t_R FILLER_137_270 ();
 FILLER_ASAP7_75t_R FILLER_137_298 ();
 DECAPx6_ASAP7_75t_R FILLER_137_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_337 ();
 DECAPx10_ASAP7_75t_R FILLER_137_342 ();
 DECAPx10_ASAP7_75t_R FILLER_137_364 ();
 DECAPx6_ASAP7_75t_R FILLER_137_386 ();
 FILLER_ASAP7_75t_R FILLER_137_400 ();
 FILLER_ASAP7_75t_R FILLER_137_424 ();
 DECAPx2_ASAP7_75t_R FILLER_137_448 ();
 FILLER_ASAP7_75t_R FILLER_137_454 ();
 DECAPx10_ASAP7_75t_R FILLER_137_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_511 ();
 DECAPx10_ASAP7_75t_R FILLER_137_534 ();
 DECAPx10_ASAP7_75t_R FILLER_137_556 ();
 DECAPx10_ASAP7_75t_R FILLER_137_578 ();
 DECAPx2_ASAP7_75t_R FILLER_137_600 ();
 FILLER_ASAP7_75t_R FILLER_137_606 ();
 DECAPx10_ASAP7_75t_R FILLER_137_630 ();
 FILLER_ASAP7_75t_R FILLER_137_652 ();
 DECAPx6_ASAP7_75t_R FILLER_137_662 ();
 DECAPx1_ASAP7_75t_R FILLER_137_676 ();
 DECAPx4_ASAP7_75t_R FILLER_137_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_712 ();
 DECAPx6_ASAP7_75t_R FILLER_137_719 ();
 DECAPx2_ASAP7_75t_R FILLER_137_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_739 ();
 FILLER_ASAP7_75t_R FILLER_137_772 ();
 DECAPx6_ASAP7_75t_R FILLER_137_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_802 ();
 FILLER_ASAP7_75t_R FILLER_137_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_811 ();
 DECAPx1_ASAP7_75t_R FILLER_137_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_823 ();
 DECAPx6_ASAP7_75t_R FILLER_137_846 ();
 FILLER_ASAP7_75t_R FILLER_137_860 ();
 FILLER_ASAP7_75t_R FILLER_137_872 ();
 DECAPx10_ASAP7_75t_R FILLER_137_880 ();
 FILLER_ASAP7_75t_R FILLER_137_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_913 ();
 DECAPx1_ASAP7_75t_R FILLER_137_920 ();
 FILLER_ASAP7_75t_R FILLER_137_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_928 ();
 DECAPx4_ASAP7_75t_R FILLER_137_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_955 ();
 DECAPx6_ASAP7_75t_R FILLER_137_962 ();
 DECAPx1_ASAP7_75t_R FILLER_137_976 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1018 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1050 ();
 DECAPx6_ASAP7_75t_R FILLER_137_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1092 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1099 ();
 FILLER_ASAP7_75t_R FILLER_137_1109 ();
 DECAPx6_ASAP7_75t_R FILLER_137_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1190 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1212 ();
 FILLER_ASAP7_75t_R FILLER_137_1222 ();
 DECAPx4_ASAP7_75t_R FILLER_138_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_12 ();
 DECAPx10_ASAP7_75t_R FILLER_138_19 ();
 DECAPx10_ASAP7_75t_R FILLER_138_41 ();
 FILLER_ASAP7_75t_R FILLER_138_63 ();
 DECAPx1_ASAP7_75t_R FILLER_138_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_83 ();
 DECAPx1_ASAP7_75t_R FILLER_138_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_101 ();
 DECAPx2_ASAP7_75t_R FILLER_138_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_114 ();
 FILLER_ASAP7_75t_R FILLER_138_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_123 ();
 DECAPx1_ASAP7_75t_R FILLER_138_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_161 ();
 FILLER_ASAP7_75t_R FILLER_138_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_186 ();
 DECAPx2_ASAP7_75t_R FILLER_138_198 ();
 FILLER_ASAP7_75t_R FILLER_138_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_206 ();
 DECAPx10_ASAP7_75t_R FILLER_138_213 ();
 FILLER_ASAP7_75t_R FILLER_138_235 ();
 DECAPx4_ASAP7_75t_R FILLER_138_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_257 ();
 DECAPx1_ASAP7_75t_R FILLER_138_313 ();
 DECAPx4_ASAP7_75t_R FILLER_138_321 ();
 FILLER_ASAP7_75t_R FILLER_138_331 ();
 DECAPx6_ASAP7_75t_R FILLER_138_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_370 ();
 DECAPx1_ASAP7_75t_R FILLER_138_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_397 ();
 DECAPx2_ASAP7_75t_R FILLER_138_456 ();
 DECAPx4_ASAP7_75t_R FILLER_138_486 ();
 FILLER_ASAP7_75t_R FILLER_138_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_498 ();
 DECAPx10_ASAP7_75t_R FILLER_138_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_527 ();
 DECAPx6_ASAP7_75t_R FILLER_138_538 ();
 DECAPx2_ASAP7_75t_R FILLER_138_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_558 ();
 DECAPx2_ASAP7_75t_R FILLER_138_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_593 ();
 FILLER_ASAP7_75t_R FILLER_138_600 ();
 FILLER_ASAP7_75t_R FILLER_138_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_611 ();
 FILLER_ASAP7_75t_R FILLER_138_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_632 ();
 DECAPx1_ASAP7_75t_R FILLER_138_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_645 ();
 FILLER_ASAP7_75t_R FILLER_138_666 ();
 DECAPx1_ASAP7_75t_R FILLER_138_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_682 ();
 DECAPx10_ASAP7_75t_R FILLER_138_689 ();
 DECAPx1_ASAP7_75t_R FILLER_138_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_715 ();
 DECAPx2_ASAP7_75t_R FILLER_138_722 ();
 DECAPx4_ASAP7_75t_R FILLER_138_745 ();
 DECAPx2_ASAP7_75t_R FILLER_138_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_773 ();
 FILLER_ASAP7_75t_R FILLER_138_800 ();
 DECAPx2_ASAP7_75t_R FILLER_138_816 ();
 FILLER_ASAP7_75t_R FILLER_138_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_824 ();
 DECAPx10_ASAP7_75t_R FILLER_138_831 ();
 DECAPx2_ASAP7_75t_R FILLER_138_853 ();
 FILLER_ASAP7_75t_R FILLER_138_859 ();
 DECAPx4_ASAP7_75t_R FILLER_138_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_891 ();
 FILLER_ASAP7_75t_R FILLER_138_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_901 ();
 DECAPx4_ASAP7_75t_R FILLER_138_913 ();
 DECAPx2_ASAP7_75t_R FILLER_138_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_939 ();
 DECAPx2_ASAP7_75t_R FILLER_138_948 ();
 FILLER_ASAP7_75t_R FILLER_138_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_956 ();
 FILLER_ASAP7_75t_R FILLER_138_960 ();
 DECAPx2_ASAP7_75t_R FILLER_138_982 ();
 FILLER_ASAP7_75t_R FILLER_138_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_990 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1026 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1057 ();
 FILLER_ASAP7_75t_R FILLER_138_1071 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1079 ();
 FILLER_ASAP7_75t_R FILLER_138_1089 ();
 FILLER_ASAP7_75t_R FILLER_138_1113 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1131 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1152 ();
 FILLER_ASAP7_75t_R FILLER_138_1162 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1175 ();
 FILLER_ASAP7_75t_R FILLER_138_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1201 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1208 ();
 FILLER_ASAP7_75t_R FILLER_138_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_139_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_14 ();
 DECAPx4_ASAP7_75t_R FILLER_139_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_31 ();
 DECAPx6_ASAP7_75t_R FILLER_139_38 ();
 DECAPx1_ASAP7_75t_R FILLER_139_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_84 ();
 FILLER_ASAP7_75t_R FILLER_139_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_107 ();
 FILLER_ASAP7_75t_R FILLER_139_114 ();
 FILLER_ASAP7_75t_R FILLER_139_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_125 ();
 FILLER_ASAP7_75t_R FILLER_139_133 ();
 DECAPx1_ASAP7_75t_R FILLER_139_157 ();
 FILLER_ASAP7_75t_R FILLER_139_173 ();
 DECAPx10_ASAP7_75t_R FILLER_139_204 ();
 DECAPx2_ASAP7_75t_R FILLER_139_226 ();
 DECAPx6_ASAP7_75t_R FILLER_139_252 ();
 DECAPx1_ASAP7_75t_R FILLER_139_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_270 ();
 DECAPx2_ASAP7_75t_R FILLER_139_315 ();
 FILLER_ASAP7_75t_R FILLER_139_321 ();
 DECAPx10_ASAP7_75t_R FILLER_139_331 ();
 DECAPx6_ASAP7_75t_R FILLER_139_353 ();
 FILLER_ASAP7_75t_R FILLER_139_367 ();
 FILLER_ASAP7_75t_R FILLER_139_413 ();
 DECAPx2_ASAP7_75t_R FILLER_139_440 ();
 DECAPx6_ASAP7_75t_R FILLER_139_468 ();
 DECAPx1_ASAP7_75t_R FILLER_139_482 ();
 DECAPx10_ASAP7_75t_R FILLER_139_509 ();
 DECAPx10_ASAP7_75t_R FILLER_139_531 ();
 DECAPx1_ASAP7_75t_R FILLER_139_553 ();
 DECAPx2_ASAP7_75t_R FILLER_139_579 ();
 FILLER_ASAP7_75t_R FILLER_139_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_596 ();
 DECAPx6_ASAP7_75t_R FILLER_139_600 ();
 FILLER_ASAP7_75t_R FILLER_139_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_636 ();
 DECAPx2_ASAP7_75t_R FILLER_139_643 ();
 FILLER_ASAP7_75t_R FILLER_139_649 ();
 DECAPx10_ASAP7_75t_R FILLER_139_657 ();
 DECAPx10_ASAP7_75t_R FILLER_139_679 ();
 DECAPx2_ASAP7_75t_R FILLER_139_701 ();
 DECAPx2_ASAP7_75t_R FILLER_139_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_731 ();
 FILLER_ASAP7_75t_R FILLER_139_740 ();
 FILLER_ASAP7_75t_R FILLER_139_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_757 ();
 DECAPx2_ASAP7_75t_R FILLER_139_764 ();
 DECAPx6_ASAP7_75t_R FILLER_139_780 ();
 DECAPx2_ASAP7_75t_R FILLER_139_802 ();
 DECAPx4_ASAP7_75t_R FILLER_139_814 ();
 FILLER_ASAP7_75t_R FILLER_139_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_826 ();
 DECAPx6_ASAP7_75t_R FILLER_139_849 ();
 FILLER_ASAP7_75t_R FILLER_139_863 ();
 DECAPx2_ASAP7_75t_R FILLER_139_871 ();
 DECAPx2_ASAP7_75t_R FILLER_139_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_891 ();
 DECAPx2_ASAP7_75t_R FILLER_139_904 ();
 FILLER_ASAP7_75t_R FILLER_139_910 ();
 DECAPx4_ASAP7_75t_R FILLER_139_934 ();
 DECAPx1_ASAP7_75t_R FILLER_139_950 ();
 DECAPx6_ASAP7_75t_R FILLER_139_963 ();
 FILLER_ASAP7_75t_R FILLER_139_977 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1063 ();
 FILLER_ASAP7_75t_R FILLER_139_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1101 ();
 FILLER_ASAP7_75t_R FILLER_139_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_139_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_139_1220 ();
 FILLER_ASAP7_75t_R FILLER_140_8 ();
 DECAPx10_ASAP7_75t_R FILLER_140_16 ();
 DECAPx10_ASAP7_75t_R FILLER_140_38 ();
 FILLER_ASAP7_75t_R FILLER_140_60 ();
 FILLER_ASAP7_75t_R FILLER_140_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_76 ();
 FILLER_ASAP7_75t_R FILLER_140_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_96 ();
 DECAPx1_ASAP7_75t_R FILLER_140_126 ();
 FILLER_ASAP7_75t_R FILLER_140_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_139 ();
 DECAPx1_ASAP7_75t_R FILLER_140_158 ();
 DECAPx2_ASAP7_75t_R FILLER_140_170 ();
 FILLER_ASAP7_75t_R FILLER_140_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_178 ();
 DECAPx1_ASAP7_75t_R FILLER_140_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_201 ();
 DECAPx6_ASAP7_75t_R FILLER_140_211 ();
 DECAPx2_ASAP7_75t_R FILLER_140_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_231 ();
 DECAPx4_ASAP7_75t_R FILLER_140_238 ();
 FILLER_ASAP7_75t_R FILLER_140_248 ();
 DECAPx10_ASAP7_75t_R FILLER_140_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_285 ();
 DECAPx10_ASAP7_75t_R FILLER_140_346 ();
 DECAPx2_ASAP7_75t_R FILLER_140_368 ();
 FILLER_ASAP7_75t_R FILLER_140_374 ();
 DECAPx6_ASAP7_75t_R FILLER_140_398 ();
 DECAPx1_ASAP7_75t_R FILLER_140_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_468 ();
 DECAPx4_ASAP7_75t_R FILLER_140_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_501 ();
 DECAPx10_ASAP7_75t_R FILLER_140_522 ();
 DECAPx10_ASAP7_75t_R FILLER_140_544 ();
 DECAPx2_ASAP7_75t_R FILLER_140_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_572 ();
 DECAPx1_ASAP7_75t_R FILLER_140_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_622 ();
 FILLER_ASAP7_75t_R FILLER_140_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_643 ();
 DECAPx1_ASAP7_75t_R FILLER_140_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_656 ();
 DECAPx6_ASAP7_75t_R FILLER_140_679 ();
 FILLER_ASAP7_75t_R FILLER_140_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_709 ();
 FILLER_ASAP7_75t_R FILLER_140_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_732 ();
 FILLER_ASAP7_75t_R FILLER_140_739 ();
 DECAPx4_ASAP7_75t_R FILLER_140_749 ();
 FILLER_ASAP7_75t_R FILLER_140_759 ();
 DECAPx6_ASAP7_75t_R FILLER_140_780 ();
 FILLER_ASAP7_75t_R FILLER_140_800 ();
 DECAPx10_ASAP7_75t_R FILLER_140_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_838 ();
 FILLER_ASAP7_75t_R FILLER_140_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_882 ();
 DECAPx6_ASAP7_75t_R FILLER_140_889 ();
 DECAPx2_ASAP7_75t_R FILLER_140_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_925 ();
 DECAPx2_ASAP7_75t_R FILLER_140_942 ();
 FILLER_ASAP7_75t_R FILLER_140_948 ();
 DECAPx1_ASAP7_75t_R FILLER_140_953 ();
 FILLER_ASAP7_75t_R FILLER_140_971 ();
 DECAPx10_ASAP7_75t_R FILLER_140_995 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1046 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1093 ();
 DECAPx4_ASAP7_75t_R FILLER_140_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1147 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1160 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_141_2 ();
 DECAPx10_ASAP7_75t_R FILLER_141_24 ();
 DECAPx6_ASAP7_75t_R FILLER_141_46 ();
 DECAPx2_ASAP7_75t_R FILLER_141_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_66 ();
 DECAPx4_ASAP7_75t_R FILLER_141_89 ();
 FILLER_ASAP7_75t_R FILLER_141_105 ();
 DECAPx10_ASAP7_75t_R FILLER_141_129 ();
 DECAPx10_ASAP7_75t_R FILLER_141_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_232 ();
 DECAPx1_ASAP7_75t_R FILLER_141_244 ();
 DECAPx6_ASAP7_75t_R FILLER_141_258 ();
 FILLER_ASAP7_75t_R FILLER_141_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_274 ();
 DECAPx1_ASAP7_75t_R FILLER_141_279 ();
 DECAPx10_ASAP7_75t_R FILLER_141_307 ();
 DECAPx10_ASAP7_75t_R FILLER_141_329 ();
 DECAPx2_ASAP7_75t_R FILLER_141_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_357 ();
 DECAPx10_ASAP7_75t_R FILLER_141_386 ();
 DECAPx10_ASAP7_75t_R FILLER_141_408 ();
 DECAPx10_ASAP7_75t_R FILLER_141_430 ();
 DECAPx2_ASAP7_75t_R FILLER_141_452 ();
 DECAPx6_ASAP7_75t_R FILLER_141_480 ();
 FILLER_ASAP7_75t_R FILLER_141_494 ();
 DECAPx2_ASAP7_75t_R FILLER_141_518 ();
 FILLER_ASAP7_75t_R FILLER_141_524 ();
 DECAPx4_ASAP7_75t_R FILLER_141_544 ();
 FILLER_ASAP7_75t_R FILLER_141_574 ();
 DECAPx6_ASAP7_75t_R FILLER_141_596 ();
 DECAPx1_ASAP7_75t_R FILLER_141_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_614 ();
 DECAPx10_ASAP7_75t_R FILLER_141_649 ();
 FILLER_ASAP7_75t_R FILLER_141_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_701 ();
 DECAPx2_ASAP7_75t_R FILLER_141_708 ();
 FILLER_ASAP7_75t_R FILLER_141_714 ();
 DECAPx4_ASAP7_75t_R FILLER_141_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_740 ();
 DECAPx4_ASAP7_75t_R FILLER_141_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_766 ();
 DECAPx10_ASAP7_75t_R FILLER_141_775 ();
 DECAPx2_ASAP7_75t_R FILLER_141_803 ();
 FILLER_ASAP7_75t_R FILLER_141_809 ();
 DECAPx6_ASAP7_75t_R FILLER_141_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_864 ();
 FILLER_ASAP7_75t_R FILLER_141_873 ();
 FILLER_ASAP7_75t_R FILLER_141_883 ();
 DECAPx2_ASAP7_75t_R FILLER_141_908 ();
 DECAPx2_ASAP7_75t_R FILLER_141_926 ();
 FILLER_ASAP7_75t_R FILLER_141_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_958 ();
 DECAPx1_ASAP7_75t_R FILLER_141_991 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1039 ();
 FILLER_ASAP7_75t_R FILLER_141_1049 ();
 FILLER_ASAP7_75t_R FILLER_141_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1087 ();
 FILLER_ASAP7_75t_R FILLER_141_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1171 ();
 FILLER_ASAP7_75t_R FILLER_141_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1202 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1214 ();
 DECAPx4_ASAP7_75t_R FILLER_142_2 ();
 DECAPx10_ASAP7_75t_R FILLER_142_22 ();
 DECAPx10_ASAP7_75t_R FILLER_142_44 ();
 DECAPx10_ASAP7_75t_R FILLER_142_66 ();
 DECAPx10_ASAP7_75t_R FILLER_142_88 ();
 DECAPx1_ASAP7_75t_R FILLER_142_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_114 ();
 DECAPx2_ASAP7_75t_R FILLER_142_137 ();
 FILLER_ASAP7_75t_R FILLER_142_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_145 ();
 DECAPx2_ASAP7_75t_R FILLER_142_163 ();
 FILLER_ASAP7_75t_R FILLER_142_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_171 ();
 DECAPx2_ASAP7_75t_R FILLER_142_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_206 ();
 DECAPx6_ASAP7_75t_R FILLER_142_213 ();
 FILLER_ASAP7_75t_R FILLER_142_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_235 ();
 DECAPx4_ASAP7_75t_R FILLER_142_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_280 ();
 DECAPx4_ASAP7_75t_R FILLER_142_301 ();
 FILLER_ASAP7_75t_R FILLER_142_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_313 ();
 DECAPx6_ASAP7_75t_R FILLER_142_334 ();
 FILLER_ASAP7_75t_R FILLER_142_348 ();
 DECAPx2_ASAP7_75t_R FILLER_142_368 ();
 FILLER_ASAP7_75t_R FILLER_142_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_376 ();
 DECAPx6_ASAP7_75t_R FILLER_142_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_422 ();
 DECAPx4_ASAP7_75t_R FILLER_142_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_439 ();
 DECAPx10_ASAP7_75t_R FILLER_142_464 ();
 DECAPx2_ASAP7_75t_R FILLER_142_492 ();
 DECAPx10_ASAP7_75t_R FILLER_142_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_523 ();
 DECAPx10_ASAP7_75t_R FILLER_142_534 ();
 FILLER_ASAP7_75t_R FILLER_142_556 ();
 DECAPx4_ASAP7_75t_R FILLER_142_568 ();
 DECAPx10_ASAP7_75t_R FILLER_142_604 ();
 FILLER_ASAP7_75t_R FILLER_142_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_648 ();
 DECAPx10_ASAP7_75t_R FILLER_142_669 ();
 FILLER_ASAP7_75t_R FILLER_142_691 ();
 FILLER_ASAP7_75t_R FILLER_142_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_703 ();
 DECAPx2_ASAP7_75t_R FILLER_142_714 ();
 FILLER_ASAP7_75t_R FILLER_142_720 ();
 DECAPx4_ASAP7_75t_R FILLER_142_730 ();
 DECAPx4_ASAP7_75t_R FILLER_142_774 ();
 FILLER_ASAP7_75t_R FILLER_142_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_792 ();
 FILLER_ASAP7_75t_R FILLER_142_805 ();
 DECAPx10_ASAP7_75t_R FILLER_142_813 ();
 DECAPx2_ASAP7_75t_R FILLER_142_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_841 ();
 FILLER_ASAP7_75t_R FILLER_142_864 ();
 DECAPx1_ASAP7_75t_R FILLER_142_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_920 ();
 DECAPx4_ASAP7_75t_R FILLER_142_934 ();
 FILLER_ASAP7_75t_R FILLER_142_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_946 ();
 DECAPx10_ASAP7_75t_R FILLER_142_953 ();
 DECAPx1_ASAP7_75t_R FILLER_142_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_979 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1044 ();
 FILLER_ASAP7_75t_R FILLER_142_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1090 ();
 FILLER_ASAP7_75t_R FILLER_142_1100 ();
 FILLER_ASAP7_75t_R FILLER_142_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1136 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1165 ();
 FILLER_ASAP7_75t_R FILLER_142_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1205 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1218 ();
 DECAPx6_ASAP7_75t_R FILLER_143_2 ();
 DECAPx10_ASAP7_75t_R FILLER_143_26 ();
 DECAPx10_ASAP7_75t_R FILLER_143_48 ();
 DECAPx2_ASAP7_75t_R FILLER_143_70 ();
 FILLER_ASAP7_75t_R FILLER_143_76 ();
 DECAPx10_ASAP7_75t_R FILLER_143_106 ();
 DECAPx2_ASAP7_75t_R FILLER_143_145 ();
 FILLER_ASAP7_75t_R FILLER_143_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_153 ();
 DECAPx1_ASAP7_75t_R FILLER_143_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_180 ();
 FILLER_ASAP7_75t_R FILLER_143_191 ();
 DECAPx6_ASAP7_75t_R FILLER_143_206 ();
 DECAPx2_ASAP7_75t_R FILLER_143_220 ();
 FILLER_ASAP7_75t_R FILLER_143_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_240 ();
 FILLER_ASAP7_75t_R FILLER_143_249 ();
 DECAPx10_ASAP7_75t_R FILLER_143_257 ();
 DECAPx2_ASAP7_75t_R FILLER_143_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_285 ();
 DECAPx10_ASAP7_75t_R FILLER_143_292 ();
 DECAPx10_ASAP7_75t_R FILLER_143_314 ();
 DECAPx10_ASAP7_75t_R FILLER_143_336 ();
 DECAPx4_ASAP7_75t_R FILLER_143_358 ();
 FILLER_ASAP7_75t_R FILLER_143_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_405 ();
 DECAPx1_ASAP7_75t_R FILLER_143_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_434 ();
 DECAPx2_ASAP7_75t_R FILLER_143_443 ();
 FILLER_ASAP7_75t_R FILLER_143_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_451 ();
 DECAPx10_ASAP7_75t_R FILLER_143_480 ();
 FILLER_ASAP7_75t_R FILLER_143_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_514 ();
 DECAPx10_ASAP7_75t_R FILLER_143_535 ();
 DECAPx4_ASAP7_75t_R FILLER_143_557 ();
 FILLER_ASAP7_75t_R FILLER_143_567 ();
 FILLER_ASAP7_75t_R FILLER_143_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_595 ();
 DECAPx6_ASAP7_75t_R FILLER_143_606 ();
 DECAPx2_ASAP7_75t_R FILLER_143_620 ();
 DECAPx2_ASAP7_75t_R FILLER_143_632 ();
 FILLER_ASAP7_75t_R FILLER_143_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_647 ();
 DECAPx1_ASAP7_75t_R FILLER_143_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_660 ();
 FILLER_ASAP7_75t_R FILLER_143_683 ();
 DECAPx1_ASAP7_75t_R FILLER_143_694 ();
 FILLER_ASAP7_75t_R FILLER_143_718 ();
 DECAPx4_ASAP7_75t_R FILLER_143_736 ();
 FILLER_ASAP7_75t_R FILLER_143_746 ();
 DECAPx2_ASAP7_75t_R FILLER_143_754 ();
 FILLER_ASAP7_75t_R FILLER_143_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_762 ();
 DECAPx2_ASAP7_75t_R FILLER_143_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_775 ();
 DECAPx4_ASAP7_75t_R FILLER_143_782 ();
 DECAPx4_ASAP7_75t_R FILLER_143_808 ();
 FILLER_ASAP7_75t_R FILLER_143_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_820 ();
 DECAPx4_ASAP7_75t_R FILLER_143_841 ();
 FILLER_ASAP7_75t_R FILLER_143_851 ();
 FILLER_ASAP7_75t_R FILLER_143_882 ();
 DECAPx6_ASAP7_75t_R FILLER_143_898 ();
 DECAPx1_ASAP7_75t_R FILLER_143_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_916 ();
 DECAPx2_ASAP7_75t_R FILLER_143_941 ();
 DECAPx10_ASAP7_75t_R FILLER_143_969 ();
 DECAPx2_ASAP7_75t_R FILLER_143_991 ();
 FILLER_ASAP7_75t_R FILLER_143_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_999 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1081 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1118 ();
 FILLER_ASAP7_75t_R FILLER_143_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1126 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_144_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_8 ();
 FILLER_ASAP7_75t_R FILLER_144_15 ();
 DECAPx10_ASAP7_75t_R FILLER_144_43 ();
 DECAPx10_ASAP7_75t_R FILLER_144_65 ();
 DECAPx2_ASAP7_75t_R FILLER_144_87 ();
 FILLER_ASAP7_75t_R FILLER_144_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_95 ();
 DECAPx4_ASAP7_75t_R FILLER_144_107 ();
 FILLER_ASAP7_75t_R FILLER_144_117 ();
 DECAPx4_ASAP7_75t_R FILLER_144_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_137 ();
 DECAPx10_ASAP7_75t_R FILLER_144_164 ();
 DECAPx2_ASAP7_75t_R FILLER_144_186 ();
 FILLER_ASAP7_75t_R FILLER_144_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_194 ();
 DECAPx10_ASAP7_75t_R FILLER_144_201 ();
 DECAPx10_ASAP7_75t_R FILLER_144_223 ();
 DECAPx2_ASAP7_75t_R FILLER_144_245 ();
 FILLER_ASAP7_75t_R FILLER_144_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_253 ();
 DECAPx4_ASAP7_75t_R FILLER_144_271 ();
 FILLER_ASAP7_75t_R FILLER_144_281 ();
 DECAPx6_ASAP7_75t_R FILLER_144_287 ();
 DECAPx1_ASAP7_75t_R FILLER_144_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_305 ();
 DECAPx10_ASAP7_75t_R FILLER_144_330 ();
 DECAPx6_ASAP7_75t_R FILLER_144_352 ();
 DECAPx2_ASAP7_75t_R FILLER_144_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_378 ();
 DECAPx4_ASAP7_75t_R FILLER_144_385 ();
 FILLER_ASAP7_75t_R FILLER_144_401 ();
 DECAPx6_ASAP7_75t_R FILLER_144_415 ();
 DECAPx1_ASAP7_75t_R FILLER_144_429 ();
 FILLER_ASAP7_75t_R FILLER_144_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_447 ();
 DECAPx1_ASAP7_75t_R FILLER_144_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_468 ();
 DECAPx2_ASAP7_75t_R FILLER_144_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_497 ();
 DECAPx2_ASAP7_75t_R FILLER_144_506 ();
 FILLER_ASAP7_75t_R FILLER_144_512 ();
 DECAPx10_ASAP7_75t_R FILLER_144_521 ();
 DECAPx10_ASAP7_75t_R FILLER_144_543 ();
 DECAPx6_ASAP7_75t_R FILLER_144_565 ();
 DECAPx2_ASAP7_75t_R FILLER_144_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_585 ();
 DECAPx1_ASAP7_75t_R FILLER_144_622 ();
 DECAPx10_ASAP7_75t_R FILLER_144_654 ();
 DECAPx1_ASAP7_75t_R FILLER_144_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_715 ();
 DECAPx6_ASAP7_75t_R FILLER_144_728 ();
 FILLER_ASAP7_75t_R FILLER_144_742 ();
 FILLER_ASAP7_75t_R FILLER_144_752 ();
 FILLER_ASAP7_75t_R FILLER_144_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_762 ();
 DECAPx1_ASAP7_75t_R FILLER_144_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_775 ();
 FILLER_ASAP7_75t_R FILLER_144_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_800 ();
 DECAPx10_ASAP7_75t_R FILLER_144_815 ();
 DECAPx10_ASAP7_75t_R FILLER_144_837 ();
 DECAPx2_ASAP7_75t_R FILLER_144_859 ();
 DECAPx1_ASAP7_75t_R FILLER_144_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_879 ();
 DECAPx1_ASAP7_75t_R FILLER_144_908 ();
 FILLER_ASAP7_75t_R FILLER_144_916 ();
 FILLER_ASAP7_75t_R FILLER_144_932 ();
 DECAPx6_ASAP7_75t_R FILLER_144_948 ();
 DECAPx2_ASAP7_75t_R FILLER_144_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_968 ();
 DECAPx4_ASAP7_75t_R FILLER_144_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_997 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1004 ();
 FILLER_ASAP7_75t_R FILLER_144_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1054 ();
 FILLER_ASAP7_75t_R FILLER_144_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1062 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1078 ();
 FILLER_ASAP7_75t_R FILLER_144_1084 ();
 FILLER_ASAP7_75t_R FILLER_144_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1197 ();
 FILLER_ASAP7_75t_R FILLER_144_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_145_2 ();
 DECAPx10_ASAP7_75t_R FILLER_145_24 ();
 DECAPx10_ASAP7_75t_R FILLER_145_46 ();
 DECAPx4_ASAP7_75t_R FILLER_145_68 ();
 FILLER_ASAP7_75t_R FILLER_145_78 ();
 DECAPx4_ASAP7_75t_R FILLER_145_122 ();
 FILLER_ASAP7_75t_R FILLER_145_132 ();
 DECAPx10_ASAP7_75t_R FILLER_145_142 ();
 DECAPx6_ASAP7_75t_R FILLER_145_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_178 ();
 FILLER_ASAP7_75t_R FILLER_145_201 ();
 FILLER_ASAP7_75t_R FILLER_145_237 ();
 FILLER_ASAP7_75t_R FILLER_145_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_262 ();
 DECAPx10_ASAP7_75t_R FILLER_145_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_352 ();
 FILLER_ASAP7_75t_R FILLER_145_375 ();
 FILLER_ASAP7_75t_R FILLER_145_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_394 ();
 DECAPx4_ASAP7_75t_R FILLER_145_401 ();
 FILLER_ASAP7_75t_R FILLER_145_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_413 ();
 FILLER_ASAP7_75t_R FILLER_145_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_429 ();
 DECAPx1_ASAP7_75t_R FILLER_145_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_444 ();
 FILLER_ASAP7_75t_R FILLER_145_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_468 ();
 DECAPx2_ASAP7_75t_R FILLER_145_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_483 ();
 DECAPx2_ASAP7_75t_R FILLER_145_490 ();
 DECAPx10_ASAP7_75t_R FILLER_145_506 ();
 DECAPx2_ASAP7_75t_R FILLER_145_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_573 ();
 DECAPx1_ASAP7_75t_R FILLER_145_581 ();
 FILLER_ASAP7_75t_R FILLER_145_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_603 ();
 DECAPx6_ASAP7_75t_R FILLER_145_620 ();
 DECAPx2_ASAP7_75t_R FILLER_145_634 ();
 DECAPx10_ASAP7_75t_R FILLER_145_646 ();
 DECAPx2_ASAP7_75t_R FILLER_145_668 ();
 FILLER_ASAP7_75t_R FILLER_145_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_676 ();
 DECAPx2_ASAP7_75t_R FILLER_145_694 ();
 FILLER_ASAP7_75t_R FILLER_145_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_709 ();
 FILLER_ASAP7_75t_R FILLER_145_717 ();
 DECAPx4_ASAP7_75t_R FILLER_145_729 ();
 FILLER_ASAP7_75t_R FILLER_145_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_741 ();
 DECAPx1_ASAP7_75t_R FILLER_145_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_773 ();
 FILLER_ASAP7_75t_R FILLER_145_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_782 ();
 FILLER_ASAP7_75t_R FILLER_145_789 ();
 DECAPx10_ASAP7_75t_R FILLER_145_811 ();
 DECAPx10_ASAP7_75t_R FILLER_145_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_855 ();
 DECAPx6_ASAP7_75t_R FILLER_145_873 ();
 DECAPx2_ASAP7_75t_R FILLER_145_893 ();
 DECAPx6_ASAP7_75t_R FILLER_145_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_935 ();
 DECAPx4_ASAP7_75t_R FILLER_145_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_954 ();
 DECAPx10_ASAP7_75t_R FILLER_145_983 ();
 FILLER_ASAP7_75t_R FILLER_145_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1056 ();
 FILLER_ASAP7_75t_R FILLER_145_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1071 ();
 FILLER_ASAP7_75t_R FILLER_145_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1080 ();
 FILLER_ASAP7_75t_R FILLER_145_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1156 ();
 FILLER_ASAP7_75t_R FILLER_145_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1217 ();
 FILLER_ASAP7_75t_R FILLER_146_2 ();
 DECAPx4_ASAP7_75t_R FILLER_146_14 ();
 FILLER_ASAP7_75t_R FILLER_146_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_26 ();
 DECAPx6_ASAP7_75t_R FILLER_146_37 ();
 DECAPx1_ASAP7_75t_R FILLER_146_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_55 ();
 DECAPx1_ASAP7_75t_R FILLER_146_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_82 ();
 DECAPx6_ASAP7_75t_R FILLER_146_89 ();
 FILLER_ASAP7_75t_R FILLER_146_109 ();
 FILLER_ASAP7_75t_R FILLER_146_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_133 ();
 DECAPx2_ASAP7_75t_R FILLER_146_156 ();
 FILLER_ASAP7_75t_R FILLER_146_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_164 ();
 DECAPx1_ASAP7_75t_R FILLER_146_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_175 ();
 DECAPx1_ASAP7_75t_R FILLER_146_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_190 ();
 DECAPx2_ASAP7_75t_R FILLER_146_197 ();
 DECAPx2_ASAP7_75t_R FILLER_146_217 ();
 FILLER_ASAP7_75t_R FILLER_146_223 ();
 FILLER_ASAP7_75t_R FILLER_146_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_234 ();
 DECAPx10_ASAP7_75t_R FILLER_146_247 ();
 DECAPx10_ASAP7_75t_R FILLER_146_269 ();
 DECAPx10_ASAP7_75t_R FILLER_146_291 ();
 DECAPx6_ASAP7_75t_R FILLER_146_313 ();
 DECAPx1_ASAP7_75t_R FILLER_146_327 ();
 DECAPx6_ASAP7_75t_R FILLER_146_337 ();
 FILLER_ASAP7_75t_R FILLER_146_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_381 ();
 DECAPx4_ASAP7_75t_R FILLER_146_394 ();
 FILLER_ASAP7_75t_R FILLER_146_404 ();
 DECAPx2_ASAP7_75t_R FILLER_146_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_418 ();
 DECAPx2_ASAP7_75t_R FILLER_146_425 ();
 FILLER_ASAP7_75t_R FILLER_146_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_433 ();
 FILLER_ASAP7_75t_R FILLER_146_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_446 ();
 FILLER_ASAP7_75t_R FILLER_146_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_461 ();
 FILLER_ASAP7_75t_R FILLER_146_464 ();
 DECAPx10_ASAP7_75t_R FILLER_146_474 ();
 DECAPx10_ASAP7_75t_R FILLER_146_508 ();
 DECAPx2_ASAP7_75t_R FILLER_146_530 ();
 DECAPx2_ASAP7_75t_R FILLER_146_542 ();
 FILLER_ASAP7_75t_R FILLER_146_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_580 ();
 DECAPx6_ASAP7_75t_R FILLER_146_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_598 ();
 DECAPx6_ASAP7_75t_R FILLER_146_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_628 ();
 FILLER_ASAP7_75t_R FILLER_146_679 ();
 DECAPx4_ASAP7_75t_R FILLER_146_694 ();
 DECAPx10_ASAP7_75t_R FILLER_146_711 ();
 FILLER_ASAP7_75t_R FILLER_146_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_745 ();
 DECAPx10_ASAP7_75t_R FILLER_146_762 ();
 DECAPx6_ASAP7_75t_R FILLER_146_784 ();
 DECAPx2_ASAP7_75t_R FILLER_146_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_810 ();
 DECAPx2_ASAP7_75t_R FILLER_146_834 ();
 FILLER_ASAP7_75t_R FILLER_146_840 ();
 FILLER_ASAP7_75t_R FILLER_146_862 ();
 DECAPx2_ASAP7_75t_R FILLER_146_874 ();
 DECAPx1_ASAP7_75t_R FILLER_146_892 ();
 DECAPx10_ASAP7_75t_R FILLER_146_953 ();
 DECAPx10_ASAP7_75t_R FILLER_146_975 ();
 DECAPx10_ASAP7_75t_R FILLER_146_997 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1043 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1052 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1088 ();
 FILLER_ASAP7_75t_R FILLER_146_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1107 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1134 ();
 DECAPx4_ASAP7_75t_R FILLER_146_1174 ();
 FILLER_ASAP7_75t_R FILLER_146_1184 ();
 FILLER_ASAP7_75t_R FILLER_146_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_147_2 ();
 DECAPx10_ASAP7_75t_R FILLER_147_24 ();
 DECAPx6_ASAP7_75t_R FILLER_147_46 ();
 FILLER_ASAP7_75t_R FILLER_147_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_80 ();
 DECAPx2_ASAP7_75t_R FILLER_147_92 ();
 FILLER_ASAP7_75t_R FILLER_147_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_100 ();
 DECAPx1_ASAP7_75t_R FILLER_147_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_127 ();
 DECAPx2_ASAP7_75t_R FILLER_147_140 ();
 FILLER_ASAP7_75t_R FILLER_147_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_148 ();
 FILLER_ASAP7_75t_R FILLER_147_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_196 ();
 DECAPx10_ASAP7_75t_R FILLER_147_274 ();
 DECAPx10_ASAP7_75t_R FILLER_147_296 ();
 DECAPx1_ASAP7_75t_R FILLER_147_318 ();
 FILLER_ASAP7_75t_R FILLER_147_344 ();
 DECAPx6_ASAP7_75t_R FILLER_147_366 ();
 DECAPx1_ASAP7_75t_R FILLER_147_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_384 ();
 DECAPx2_ASAP7_75t_R FILLER_147_391 ();
 FILLER_ASAP7_75t_R FILLER_147_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_407 ();
 DECAPx1_ASAP7_75t_R FILLER_147_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_427 ();
 DECAPx4_ASAP7_75t_R FILLER_147_436 ();
 FILLER_ASAP7_75t_R FILLER_147_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_460 ();
 DECAPx6_ASAP7_75t_R FILLER_147_479 ();
 FILLER_ASAP7_75t_R FILLER_147_493 ();
 DECAPx2_ASAP7_75t_R FILLER_147_509 ();
 FILLER_ASAP7_75t_R FILLER_147_515 ();
 DECAPx10_ASAP7_75t_R FILLER_147_537 ();
 DECAPx6_ASAP7_75t_R FILLER_147_559 ();
 DECAPx2_ASAP7_75t_R FILLER_147_573 ();
 DECAPx4_ASAP7_75t_R FILLER_147_593 ();
 DECAPx2_ASAP7_75t_R FILLER_147_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_621 ();
 DECAPx6_ASAP7_75t_R FILLER_147_658 ();
 DECAPx1_ASAP7_75t_R FILLER_147_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_676 ();
 DECAPx2_ASAP7_75t_R FILLER_147_699 ();
 FILLER_ASAP7_75t_R FILLER_147_726 ();
 DECAPx2_ASAP7_75t_R FILLER_147_746 ();
 FILLER_ASAP7_75t_R FILLER_147_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_754 ();
 DECAPx2_ASAP7_75t_R FILLER_147_765 ();
 FILLER_ASAP7_75t_R FILLER_147_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_795 ();
 DECAPx2_ASAP7_75t_R FILLER_147_818 ();
 DECAPx6_ASAP7_75t_R FILLER_147_827 ();
 DECAPx2_ASAP7_75t_R FILLER_147_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_847 ();
 DECAPx2_ASAP7_75t_R FILLER_147_870 ();
 DECAPx4_ASAP7_75t_R FILLER_147_903 ();
 FILLER_ASAP7_75t_R FILLER_147_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_915 ();
 DECAPx1_ASAP7_75t_R FILLER_147_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_934 ();
 DECAPx10_ASAP7_75t_R FILLER_147_946 ();
 DECAPx1_ASAP7_75t_R FILLER_147_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_975 ();
 DECAPx10_ASAP7_75t_R FILLER_147_999 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_147_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1097 ();
 FILLER_ASAP7_75t_R FILLER_147_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1139 ();
 DECAPx1_ASAP7_75t_R FILLER_147_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1161 ();
 FILLER_ASAP7_75t_R FILLER_147_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1196 ();
 DECAPx6_ASAP7_75t_R FILLER_147_1208 ();
 FILLER_ASAP7_75t_R FILLER_147_1222 ();
 DECAPx6_ASAP7_75t_R FILLER_148_2 ();
 DECAPx1_ASAP7_75t_R FILLER_148_16 ();
 DECAPx10_ASAP7_75t_R FILLER_148_26 ();
 DECAPx10_ASAP7_75t_R FILLER_148_48 ();
 DECAPx4_ASAP7_75t_R FILLER_148_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_80 ();
 DECAPx1_ASAP7_75t_R FILLER_148_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_99 ();
 DECAPx10_ASAP7_75t_R FILLER_148_106 ();
 DECAPx10_ASAP7_75t_R FILLER_148_128 ();
 DECAPx10_ASAP7_75t_R FILLER_148_150 ();
 DECAPx6_ASAP7_75t_R FILLER_148_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_186 ();
 DECAPx1_ASAP7_75t_R FILLER_148_209 ();
 DECAPx6_ASAP7_75t_R FILLER_148_225 ();
 DECAPx1_ASAP7_75t_R FILLER_148_239 ();
 DECAPx6_ASAP7_75t_R FILLER_148_249 ();
 DECAPx1_ASAP7_75t_R FILLER_148_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_267 ();
 DECAPx10_ASAP7_75t_R FILLER_148_298 ();
 DECAPx6_ASAP7_75t_R FILLER_148_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_334 ();
 DECAPx4_ASAP7_75t_R FILLER_148_363 ();
 FILLER_ASAP7_75t_R FILLER_148_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_398 ();
 FILLER_ASAP7_75t_R FILLER_148_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_433 ();
 FILLER_ASAP7_75t_R FILLER_148_454 ();
 FILLER_ASAP7_75t_R FILLER_148_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_466 ();
 DECAPx6_ASAP7_75t_R FILLER_148_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_510 ();
 FILLER_ASAP7_75t_R FILLER_148_524 ();
 DECAPx6_ASAP7_75t_R FILLER_148_538 ();
 FILLER_ASAP7_75t_R FILLER_148_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_554 ();
 FILLER_ASAP7_75t_R FILLER_148_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_599 ();
 FILLER_ASAP7_75t_R FILLER_148_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_620 ();
 FILLER_ASAP7_75t_R FILLER_148_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_633 ();
 DECAPx4_ASAP7_75t_R FILLER_148_648 ();
 FILLER_ASAP7_75t_R FILLER_148_658 ();
 DECAPx10_ASAP7_75t_R FILLER_148_663 ();
 DECAPx2_ASAP7_75t_R FILLER_148_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_699 ();
 DECAPx2_ASAP7_75t_R FILLER_148_727 ();
 FILLER_ASAP7_75t_R FILLER_148_733 ();
 DECAPx2_ASAP7_75t_R FILLER_148_751 ();
 FILLER_ASAP7_75t_R FILLER_148_779 ();
 DECAPx4_ASAP7_75t_R FILLER_148_803 ();
 FILLER_ASAP7_75t_R FILLER_148_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_895 ();
 DECAPx10_ASAP7_75t_R FILLER_148_917 ();
 DECAPx10_ASAP7_75t_R FILLER_148_939 ();
 DECAPx1_ASAP7_75t_R FILLER_148_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_965 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1032 ();
 FILLER_ASAP7_75t_R FILLER_148_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1069 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1091 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1151 ();
 FILLER_ASAP7_75t_R FILLER_148_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1162 ();
 DECAPx1_ASAP7_75t_R FILLER_148_1183 ();
 FILLER_ASAP7_75t_R FILLER_148_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_148_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1213 ();
 DECAPx1_ASAP7_75t_R FILLER_148_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_149_2 ();
 DECAPx10_ASAP7_75t_R FILLER_149_24 ();
 DECAPx10_ASAP7_75t_R FILLER_149_46 ();
 DECAPx4_ASAP7_75t_R FILLER_149_85 ();
 DECAPx1_ASAP7_75t_R FILLER_149_109 ();
 DECAPx4_ASAP7_75t_R FILLER_149_120 ();
 FILLER_ASAP7_75t_R FILLER_149_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_132 ();
 DECAPx2_ASAP7_75t_R FILLER_149_141 ();
 FILLER_ASAP7_75t_R FILLER_149_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_149 ();
 DECAPx10_ASAP7_75t_R FILLER_149_178 ();
 DECAPx2_ASAP7_75t_R FILLER_149_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_206 ();
 DECAPx4_ASAP7_75t_R FILLER_149_229 ();
 FILLER_ASAP7_75t_R FILLER_149_239 ();
 DECAPx10_ASAP7_75t_R FILLER_149_263 ();
 DECAPx10_ASAP7_75t_R FILLER_149_285 ();
 DECAPx2_ASAP7_75t_R FILLER_149_307 ();
 FILLER_ASAP7_75t_R FILLER_149_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_315 ();
 DECAPx2_ASAP7_75t_R FILLER_149_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_366 ();
 DECAPx6_ASAP7_75t_R FILLER_149_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_410 ();
 DECAPx2_ASAP7_75t_R FILLER_149_420 ();
 FILLER_ASAP7_75t_R FILLER_149_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_428 ();
 DECAPx2_ASAP7_75t_R FILLER_149_439 ();
 FILLER_ASAP7_75t_R FILLER_149_445 ();
 DECAPx10_ASAP7_75t_R FILLER_149_466 ();
 FILLER_ASAP7_75t_R FILLER_149_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_521 ();
 DECAPx10_ASAP7_75t_R FILLER_149_530 ();
 DECAPx4_ASAP7_75t_R FILLER_149_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_562 ();
 FILLER_ASAP7_75t_R FILLER_149_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_575 ();
 DECAPx4_ASAP7_75t_R FILLER_149_588 ();
 FILLER_ASAP7_75t_R FILLER_149_601 ();
 DECAPx4_ASAP7_75t_R FILLER_149_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_621 ();
 DECAPx1_ASAP7_75t_R FILLER_149_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_641 ();
 DECAPx10_ASAP7_75t_R FILLER_149_662 ();
 FILLER_ASAP7_75t_R FILLER_149_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_692 ();
 FILLER_ASAP7_75t_R FILLER_149_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_702 ();
 DECAPx10_ASAP7_75t_R FILLER_149_731 ();
 DECAPx2_ASAP7_75t_R FILLER_149_753 ();
 DECAPx6_ASAP7_75t_R FILLER_149_781 ();
 DECAPx1_ASAP7_75t_R FILLER_149_795 ();
 FILLER_ASAP7_75t_R FILLER_149_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_823 ();
 DECAPx10_ASAP7_75t_R FILLER_149_827 ();
 DECAPx6_ASAP7_75t_R FILLER_149_849 ();
 FILLER_ASAP7_75t_R FILLER_149_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_865 ();
 DECAPx2_ASAP7_75t_R FILLER_149_908 ();
 DECAPx4_ASAP7_75t_R FILLER_149_926 ();
 DECAPx1_ASAP7_75t_R FILLER_149_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1020 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1048 ();
 DECAPx4_ASAP7_75t_R FILLER_149_1082 ();
 FILLER_ASAP7_75t_R FILLER_149_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_149_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1162 ();
 FILLER_ASAP7_75t_R FILLER_149_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1186 ();
 DECAPx4_ASAP7_75t_R FILLER_149_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_150_2 ();
 DECAPx10_ASAP7_75t_R FILLER_150_24 ();
 DECAPx4_ASAP7_75t_R FILLER_150_46 ();
 FILLER_ASAP7_75t_R FILLER_150_56 ();
 DECAPx1_ASAP7_75t_R FILLER_150_80 ();
 DECAPx10_ASAP7_75t_R FILLER_150_92 ();
 DECAPx4_ASAP7_75t_R FILLER_150_114 ();
 FILLER_ASAP7_75t_R FILLER_150_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_126 ();
 FILLER_ASAP7_75t_R FILLER_150_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_151 ();
 DECAPx10_ASAP7_75t_R FILLER_150_177 ();
 DECAPx10_ASAP7_75t_R FILLER_150_199 ();
 DECAPx1_ASAP7_75t_R FILLER_150_221 ();
 DECAPx1_ASAP7_75t_R FILLER_150_233 ();
 DECAPx2_ASAP7_75t_R FILLER_150_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_254 ();
 DECAPx6_ASAP7_75t_R FILLER_150_278 ();
 DECAPx2_ASAP7_75t_R FILLER_150_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_298 ();
 DECAPx6_ASAP7_75t_R FILLER_150_319 ();
 FILLER_ASAP7_75t_R FILLER_150_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_335 ();
 DECAPx1_ASAP7_75t_R FILLER_150_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_368 ();
 DECAPx2_ASAP7_75t_R FILLER_150_375 ();
 DECAPx6_ASAP7_75t_R FILLER_150_396 ();
 DECAPx1_ASAP7_75t_R FILLER_150_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_423 ();
 DECAPx2_ASAP7_75t_R FILLER_150_442 ();
 DECAPx6_ASAP7_75t_R FILLER_150_464 ();
 DECAPx6_ASAP7_75t_R FILLER_150_500 ();
 DECAPx4_ASAP7_75t_R FILLER_150_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_546 ();
 FILLER_ASAP7_75t_R FILLER_150_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_604 ();
 FILLER_ASAP7_75t_R FILLER_150_615 ();
 FILLER_ASAP7_75t_R FILLER_150_629 ();
 DECAPx1_ASAP7_75t_R FILLER_150_646 ();
 FILLER_ASAP7_75t_R FILLER_150_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_674 ();
 FILLER_ASAP7_75t_R FILLER_150_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_688 ();
 FILLER_ASAP7_75t_R FILLER_150_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_698 ();
 FILLER_ASAP7_75t_R FILLER_150_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_707 ();
 DECAPx6_ASAP7_75t_R FILLER_150_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_736 ();
 DECAPx10_ASAP7_75t_R FILLER_150_757 ();
 DECAPx10_ASAP7_75t_R FILLER_150_779 ();
 DECAPx2_ASAP7_75t_R FILLER_150_801 ();
 DECAPx10_ASAP7_75t_R FILLER_150_827 ();
 DECAPx6_ASAP7_75t_R FILLER_150_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_863 ();
 DECAPx10_ASAP7_75t_R FILLER_150_898 ();
 DECAPx10_ASAP7_75t_R FILLER_150_920 ();
 DECAPx4_ASAP7_75t_R FILLER_150_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_952 ();
 DECAPx1_ASAP7_75t_R FILLER_150_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1010 ();
 DECAPx4_ASAP7_75t_R FILLER_150_1021 ();
 FILLER_ASAP7_75t_R FILLER_150_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1033 ();
 FILLER_ASAP7_75t_R FILLER_150_1040 ();
 FILLER_ASAP7_75t_R FILLER_150_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1072 ();
 DECAPx6_ASAP7_75t_R FILLER_150_1103 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1117 ();
 FILLER_ASAP7_75t_R FILLER_150_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1142 ();
 DECAPx4_ASAP7_75t_R FILLER_150_1164 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1186 ();
 DECAPx4_ASAP7_75t_R FILLER_150_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_151_2 ();
 DECAPx10_ASAP7_75t_R FILLER_151_24 ();
 DECAPx10_ASAP7_75t_R FILLER_151_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_68 ();
 FILLER_ASAP7_75t_R FILLER_151_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_77 ();
 FILLER_ASAP7_75t_R FILLER_151_90 ();
 DECAPx2_ASAP7_75t_R FILLER_151_100 ();
 DECAPx1_ASAP7_75t_R FILLER_151_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_163 ();
 FILLER_ASAP7_75t_R FILLER_151_186 ();
 FILLER_ASAP7_75t_R FILLER_151_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_241 ();
 DECAPx6_ASAP7_75t_R FILLER_151_249 ();
 DECAPx2_ASAP7_75t_R FILLER_151_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_269 ();
 DECAPx4_ASAP7_75t_R FILLER_151_316 ();
 FILLER_ASAP7_75t_R FILLER_151_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_328 ();
 FILLER_ASAP7_75t_R FILLER_151_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_335 ();
 DECAPx1_ASAP7_75t_R FILLER_151_364 ();
 DECAPx1_ASAP7_75t_R FILLER_151_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_380 ();
 DECAPx1_ASAP7_75t_R FILLER_151_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_388 ();
 DECAPx1_ASAP7_75t_R FILLER_151_421 ();
 DECAPx6_ASAP7_75t_R FILLER_151_432 ();
 FILLER_ASAP7_75t_R FILLER_151_446 ();
 DECAPx10_ASAP7_75t_R FILLER_151_458 ();
 DECAPx1_ASAP7_75t_R FILLER_151_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_484 ();
 DECAPx1_ASAP7_75t_R FILLER_151_495 ();
 DECAPx2_ASAP7_75t_R FILLER_151_505 ();
 DECAPx10_ASAP7_75t_R FILLER_151_540 ();
 DECAPx4_ASAP7_75t_R FILLER_151_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_572 ();
 FILLER_ASAP7_75t_R FILLER_151_576 ();
 DECAPx1_ASAP7_75t_R FILLER_151_596 ();
 DECAPx2_ASAP7_75t_R FILLER_151_607 ();
 FILLER_ASAP7_75t_R FILLER_151_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_615 ();
 DECAPx2_ASAP7_75t_R FILLER_151_630 ();
 DECAPx10_ASAP7_75t_R FILLER_151_642 ();
 DECAPx2_ASAP7_75t_R FILLER_151_664 ();
 DECAPx2_ASAP7_75t_R FILLER_151_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_697 ();
 DECAPx1_ASAP7_75t_R FILLER_151_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_714 ();
 DECAPx6_ASAP7_75t_R FILLER_151_722 ();
 DECAPx6_ASAP7_75t_R FILLER_151_756 ();
 FILLER_ASAP7_75t_R FILLER_151_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_772 ();
 DECAPx4_ASAP7_75t_R FILLER_151_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_786 ();
 FILLER_ASAP7_75t_R FILLER_151_809 ();
 DECAPx6_ASAP7_75t_R FILLER_151_814 ();
 FILLER_ASAP7_75t_R FILLER_151_828 ();
 DECAPx10_ASAP7_75t_R FILLER_151_880 ();
 DECAPx4_ASAP7_75t_R FILLER_151_902 ();
 FILLER_ASAP7_75t_R FILLER_151_912 ();
 DECAPx1_ASAP7_75t_R FILLER_151_926 ();
 DECAPx1_ASAP7_75t_R FILLER_151_948 ();
 DECAPx1_ASAP7_75t_R FILLER_151_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_960 ();
 FILLER_ASAP7_75t_R FILLER_151_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_969 ();
 DECAPx2_ASAP7_75t_R FILLER_151_985 ();
 FILLER_ASAP7_75t_R FILLER_151_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_151_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1054 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_151_1132 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_151_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_151_1209 ();
 FILLER_ASAP7_75t_R FILLER_151_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_152_2 ();
 DECAPx10_ASAP7_75t_R FILLER_152_24 ();
 DECAPx10_ASAP7_75t_R FILLER_152_46 ();
 DECAPx6_ASAP7_75t_R FILLER_152_68 ();
 FILLER_ASAP7_75t_R FILLER_152_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_106 ();
 DECAPx2_ASAP7_75t_R FILLER_152_128 ();
 FILLER_ASAP7_75t_R FILLER_152_141 ();
 DECAPx10_ASAP7_75t_R FILLER_152_154 ();
 DECAPx1_ASAP7_75t_R FILLER_152_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_180 ();
 DECAPx6_ASAP7_75t_R FILLER_152_198 ();
 DECAPx2_ASAP7_75t_R FILLER_152_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_218 ();
 DECAPx4_ASAP7_75t_R FILLER_152_231 ();
 FILLER_ASAP7_75t_R FILLER_152_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_243 ();
 DECAPx1_ASAP7_75t_R FILLER_152_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_282 ();
 DECAPx10_ASAP7_75t_R FILLER_152_306 ();
 FILLER_ASAP7_75t_R FILLER_152_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_330 ();
 DECAPx6_ASAP7_75t_R FILLER_152_353 ();
 DECAPx1_ASAP7_75t_R FILLER_152_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_371 ();
 DECAPx2_ASAP7_75t_R FILLER_152_400 ();
 FILLER_ASAP7_75t_R FILLER_152_406 ();
 DECAPx4_ASAP7_75t_R FILLER_152_422 ();
 FILLER_ASAP7_75t_R FILLER_152_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_434 ();
 FILLER_ASAP7_75t_R FILLER_152_445 ();
 DECAPx6_ASAP7_75t_R FILLER_152_464 ();
 DECAPx2_ASAP7_75t_R FILLER_152_478 ();
 FILLER_ASAP7_75t_R FILLER_152_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_494 ();
 FILLER_ASAP7_75t_R FILLER_152_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_518 ();
 DECAPx2_ASAP7_75t_R FILLER_152_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_534 ();
 DECAPx10_ASAP7_75t_R FILLER_152_541 ();
 FILLER_ASAP7_75t_R FILLER_152_563 ();
 FILLER_ASAP7_75t_R FILLER_152_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_589 ();
 DECAPx4_ASAP7_75t_R FILLER_152_608 ();
 FILLER_ASAP7_75t_R FILLER_152_618 ();
 DECAPx1_ASAP7_75t_R FILLER_152_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_636 ();
 DECAPx2_ASAP7_75t_R FILLER_152_659 ();
 FILLER_ASAP7_75t_R FILLER_152_665 ();
 DECAPx2_ASAP7_75t_R FILLER_152_670 ();
 FILLER_ASAP7_75t_R FILLER_152_681 ();
 FILLER_ASAP7_75t_R FILLER_152_689 ();
 FILLER_ASAP7_75t_R FILLER_152_707 ();
 DECAPx2_ASAP7_75t_R FILLER_152_731 ();
 FILLER_ASAP7_75t_R FILLER_152_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_775 ();
 DECAPx10_ASAP7_75t_R FILLER_152_798 ();
 DECAPx10_ASAP7_75t_R FILLER_152_820 ();
 DECAPx10_ASAP7_75t_R FILLER_152_842 ();
 DECAPx6_ASAP7_75t_R FILLER_152_864 ();
 DECAPx4_ASAP7_75t_R FILLER_152_920 ();
 DECAPx4_ASAP7_75t_R FILLER_152_940 ();
 FILLER_ASAP7_75t_R FILLER_152_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_952 ();
 FILLER_ASAP7_75t_R FILLER_152_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_970 ();
 DECAPx1_ASAP7_75t_R FILLER_152_998 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1071 ();
 FILLER_ASAP7_75t_R FILLER_152_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1153 ();
 FILLER_ASAP7_75t_R FILLER_152_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1185 ();
 FILLER_ASAP7_75t_R FILLER_152_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_153_2 ();
 DECAPx10_ASAP7_75t_R FILLER_153_24 ();
 DECAPx6_ASAP7_75t_R FILLER_153_46 ();
 DECAPx1_ASAP7_75t_R FILLER_153_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_64 ();
 DECAPx2_ASAP7_75t_R FILLER_153_95 ();
 DECAPx2_ASAP7_75t_R FILLER_153_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_114 ();
 DECAPx6_ASAP7_75t_R FILLER_153_129 ();
 DECAPx2_ASAP7_75t_R FILLER_153_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_149 ();
 DECAPx6_ASAP7_75t_R FILLER_153_172 ();
 DECAPx2_ASAP7_75t_R FILLER_153_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_192 ();
 DECAPx10_ASAP7_75t_R FILLER_153_199 ();
 DECAPx6_ASAP7_75t_R FILLER_153_221 ();
 DECAPx1_ASAP7_75t_R FILLER_153_235 ();
 DECAPx6_ASAP7_75t_R FILLER_153_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_268 ();
 DECAPx10_ASAP7_75t_R FILLER_153_291 ();
 DECAPx10_ASAP7_75t_R FILLER_153_313 ();
 DECAPx2_ASAP7_75t_R FILLER_153_335 ();
 FILLER_ASAP7_75t_R FILLER_153_341 ();
 DECAPx2_ASAP7_75t_R FILLER_153_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_392 ();
 DECAPx10_ASAP7_75t_R FILLER_153_399 ();
 DECAPx4_ASAP7_75t_R FILLER_153_421 ();
 FILLER_ASAP7_75t_R FILLER_153_431 ();
 DECAPx2_ASAP7_75t_R FILLER_153_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_461 ();
 DECAPx1_ASAP7_75t_R FILLER_153_480 ();
 DECAPx1_ASAP7_75t_R FILLER_153_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_508 ();
 DECAPx1_ASAP7_75t_R FILLER_153_515 ();
 DECAPx2_ASAP7_75t_R FILLER_153_554 ();
 FILLER_ASAP7_75t_R FILLER_153_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_596 ();
 FILLER_ASAP7_75t_R FILLER_153_607 ();
 FILLER_ASAP7_75t_R FILLER_153_616 ();
 FILLER_ASAP7_75t_R FILLER_153_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_626 ();
 DECAPx6_ASAP7_75t_R FILLER_153_633 ();
 DECAPx1_ASAP7_75t_R FILLER_153_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_651 ();
 DECAPx2_ASAP7_75t_R FILLER_153_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_705 ();
 DECAPx10_ASAP7_75t_R FILLER_153_710 ();
 DECAPx6_ASAP7_75t_R FILLER_153_732 ();
 FILLER_ASAP7_75t_R FILLER_153_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_748 ();
 DECAPx2_ASAP7_75t_R FILLER_153_752 ();
 FILLER_ASAP7_75t_R FILLER_153_758 ();
 FILLER_ASAP7_75t_R FILLER_153_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_782 ();
 DECAPx4_ASAP7_75t_R FILLER_153_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_819 ();
 DECAPx4_ASAP7_75t_R FILLER_153_841 ();
 DECAPx10_ASAP7_75t_R FILLER_153_871 ();
 DECAPx2_ASAP7_75t_R FILLER_153_893 ();
 FILLER_ASAP7_75t_R FILLER_153_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_933 ();
 DECAPx6_ASAP7_75t_R FILLER_153_940 ();
 FILLER_ASAP7_75t_R FILLER_153_972 ();
 FILLER_ASAP7_75t_R FILLER_153_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_983 ();
 DECAPx2_ASAP7_75t_R FILLER_153_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_996 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1019 ();
 FILLER_ASAP7_75t_R FILLER_153_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_153_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1132 ();
 FILLER_ASAP7_75t_R FILLER_153_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_153_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1223 ();
 DECAPx6_ASAP7_75t_R FILLER_154_2 ();
 FILLER_ASAP7_75t_R FILLER_154_16 ();
 DECAPx10_ASAP7_75t_R FILLER_154_24 ();
 DECAPx6_ASAP7_75t_R FILLER_154_46 ();
 DECAPx10_ASAP7_75t_R FILLER_154_82 ();
 DECAPx10_ASAP7_75t_R FILLER_154_104 ();
 DECAPx4_ASAP7_75t_R FILLER_154_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_150 ();
 DECAPx6_ASAP7_75t_R FILLER_154_157 ();
 DECAPx2_ASAP7_75t_R FILLER_154_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_177 ();
 DECAPx2_ASAP7_75t_R FILLER_154_184 ();
 FILLER_ASAP7_75t_R FILLER_154_190 ();
 FILLER_ASAP7_75t_R FILLER_154_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_236 ();
 FILLER_ASAP7_75t_R FILLER_154_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_284 ();
 DECAPx10_ASAP7_75t_R FILLER_154_288 ();
 DECAPx6_ASAP7_75t_R FILLER_154_310 ();
 DECAPx1_ASAP7_75t_R FILLER_154_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_351 ();
 FILLER_ASAP7_75t_R FILLER_154_362 ();
 DECAPx2_ASAP7_75t_R FILLER_154_384 ();
 FILLER_ASAP7_75t_R FILLER_154_390 ();
 DECAPx1_ASAP7_75t_R FILLER_154_400 ();
 FILLER_ASAP7_75t_R FILLER_154_412 ();
 DECAPx2_ASAP7_75t_R FILLER_154_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_426 ();
 DECAPx2_ASAP7_75t_R FILLER_154_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_453 ();
 DECAPx4_ASAP7_75t_R FILLER_154_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_493 ();
 DECAPx4_ASAP7_75t_R FILLER_154_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_510 ();
 DECAPx1_ASAP7_75t_R FILLER_154_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_525 ();
 DECAPx10_ASAP7_75t_R FILLER_154_538 ();
 DECAPx4_ASAP7_75t_R FILLER_154_560 ();
 FILLER_ASAP7_75t_R FILLER_154_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_572 ();
 DECAPx1_ASAP7_75t_R FILLER_154_593 ();
 DECAPx4_ASAP7_75t_R FILLER_154_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_614 ();
 DECAPx4_ASAP7_75t_R FILLER_154_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_643 ();
 DECAPx4_ASAP7_75t_R FILLER_154_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_674 ();
 FILLER_ASAP7_75t_R FILLER_154_686 ();
 DECAPx10_ASAP7_75t_R FILLER_154_691 ();
 DECAPx4_ASAP7_75t_R FILLER_154_713 ();
 DECAPx2_ASAP7_75t_R FILLER_154_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_733 ();
 DECAPx6_ASAP7_75t_R FILLER_154_756 ();
 DECAPx1_ASAP7_75t_R FILLER_154_770 ();
 DECAPx10_ASAP7_75t_R FILLER_154_797 ();
 DECAPx10_ASAP7_75t_R FILLER_154_819 ();
 DECAPx10_ASAP7_75t_R FILLER_154_841 ();
 DECAPx2_ASAP7_75t_R FILLER_154_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_891 ();
 DECAPx10_ASAP7_75t_R FILLER_154_914 ();
 DECAPx2_ASAP7_75t_R FILLER_154_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_956 ();
 DECAPx10_ASAP7_75t_R FILLER_154_987 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1019 ();
 FILLER_ASAP7_75t_R FILLER_154_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1052 ();
 FILLER_ASAP7_75t_R FILLER_154_1066 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1090 ();
 FILLER_ASAP7_75t_R FILLER_154_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1148 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1170 ();
 FILLER_ASAP7_75t_R FILLER_154_1180 ();
 FILLER_ASAP7_75t_R FILLER_154_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1218 ();
 DECAPx4_ASAP7_75t_R FILLER_155_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_12 ();
 DECAPx2_ASAP7_75t_R FILLER_155_19 ();
 DECAPx10_ASAP7_75t_R FILLER_155_31 ();
 DECAPx10_ASAP7_75t_R FILLER_155_53 ();
 DECAPx2_ASAP7_75t_R FILLER_155_75 ();
 FILLER_ASAP7_75t_R FILLER_155_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_83 ();
 DECAPx1_ASAP7_75t_R FILLER_155_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_129 ();
 DECAPx2_ASAP7_75t_R FILLER_155_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_186 ();
 DECAPx6_ASAP7_75t_R FILLER_155_198 ();
 FILLER_ASAP7_75t_R FILLER_155_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_236 ();
 FILLER_ASAP7_75t_R FILLER_155_243 ();
 DECAPx6_ASAP7_75t_R FILLER_155_267 ();
 FILLER_ASAP7_75t_R FILLER_155_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_304 ();
 FILLER_ASAP7_75t_R FILLER_155_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_313 ();
 DECAPx4_ASAP7_75t_R FILLER_155_336 ();
 FILLER_ASAP7_75t_R FILLER_155_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_348 ();
 DECAPx10_ASAP7_75t_R FILLER_155_355 ();
 FILLER_ASAP7_75t_R FILLER_155_377 ();
 FILLER_ASAP7_75t_R FILLER_155_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_403 ();
 DECAPx1_ASAP7_75t_R FILLER_155_423 ();
 DECAPx6_ASAP7_75t_R FILLER_155_430 ();
 DECAPx4_ASAP7_75t_R FILLER_155_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_461 ();
 DECAPx2_ASAP7_75t_R FILLER_155_476 ();
 FILLER_ASAP7_75t_R FILLER_155_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_484 ();
 DECAPx1_ASAP7_75t_R FILLER_155_488 ();
 FILLER_ASAP7_75t_R FILLER_155_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_504 ();
 DECAPx10_ASAP7_75t_R FILLER_155_533 ();
 DECAPx10_ASAP7_75t_R FILLER_155_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_577 ();
 DECAPx4_ASAP7_75t_R FILLER_155_584 ();
 FILLER_ASAP7_75t_R FILLER_155_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_596 ();
 DECAPx10_ASAP7_75t_R FILLER_155_613 ();
 DECAPx4_ASAP7_75t_R FILLER_155_635 ();
 DECAPx1_ASAP7_75t_R FILLER_155_651 ();
 DECAPx10_ASAP7_75t_R FILLER_155_675 ();
 DECAPx1_ASAP7_75t_R FILLER_155_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_723 ();
 DECAPx1_ASAP7_75t_R FILLER_155_749 ();
 DECAPx6_ASAP7_75t_R FILLER_155_775 ();
 DECAPx1_ASAP7_75t_R FILLER_155_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_793 ();
 DECAPx10_ASAP7_75t_R FILLER_155_834 ();
 DECAPx2_ASAP7_75t_R FILLER_155_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_862 ();
 DECAPx6_ASAP7_75t_R FILLER_155_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_889 ();
 DECAPx10_ASAP7_75t_R FILLER_155_902 ();
 DECAPx6_ASAP7_75t_R FILLER_155_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_940 ();
 FILLER_ASAP7_75t_R FILLER_155_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_964 ();
 DECAPx4_ASAP7_75t_R FILLER_155_971 ();
 FILLER_ASAP7_75t_R FILLER_155_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_983 ();
 FILLER_ASAP7_75t_R FILLER_155_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_994 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1072 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1102 ();
 DECAPx4_ASAP7_75t_R FILLER_155_1106 ();
 FILLER_ASAP7_75t_R FILLER_155_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1138 ();
 FILLER_ASAP7_75t_R FILLER_155_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1172 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1208 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1218 ();
 FILLER_ASAP7_75t_R FILLER_156_2 ();
 DECAPx10_ASAP7_75t_R FILLER_156_10 ();
 DECAPx10_ASAP7_75t_R FILLER_156_32 ();
 DECAPx10_ASAP7_75t_R FILLER_156_54 ();
 DECAPx2_ASAP7_75t_R FILLER_156_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_93 ();
 DECAPx1_ASAP7_75t_R FILLER_156_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_104 ();
 DECAPx4_ASAP7_75t_R FILLER_156_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_121 ();
 FILLER_ASAP7_75t_R FILLER_156_128 ();
 DECAPx6_ASAP7_75t_R FILLER_156_147 ();
 DECAPx2_ASAP7_75t_R FILLER_156_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_167 ();
 FILLER_ASAP7_75t_R FILLER_156_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_189 ();
 DECAPx6_ASAP7_75t_R FILLER_156_197 ();
 FILLER_ASAP7_75t_R FILLER_156_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_219 ();
 DECAPx10_ASAP7_75t_R FILLER_156_235 ();
 DECAPx10_ASAP7_75t_R FILLER_156_257 ();
 DECAPx1_ASAP7_75t_R FILLER_156_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_283 ();
 DECAPx10_ASAP7_75t_R FILLER_156_296 ();
 DECAPx10_ASAP7_75t_R FILLER_156_318 ();
 DECAPx4_ASAP7_75t_R FILLER_156_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_350 ();
 FILLER_ASAP7_75t_R FILLER_156_373 ();
 DECAPx2_ASAP7_75t_R FILLER_156_389 ();
 FILLER_ASAP7_75t_R FILLER_156_395 ();
 DECAPx1_ASAP7_75t_R FILLER_156_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_410 ();
 FILLER_ASAP7_75t_R FILLER_156_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_419 ();
 DECAPx6_ASAP7_75t_R FILLER_156_434 ();
 DECAPx2_ASAP7_75t_R FILLER_156_448 ();
 DECAPx6_ASAP7_75t_R FILLER_156_464 ();
 DECAPx2_ASAP7_75t_R FILLER_156_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_484 ();
 DECAPx6_ASAP7_75t_R FILLER_156_488 ();
 DECAPx6_ASAP7_75t_R FILLER_156_528 ();
 DECAPx1_ASAP7_75t_R FILLER_156_542 ();
 DECAPx6_ASAP7_75t_R FILLER_156_552 ();
 DECAPx1_ASAP7_75t_R FILLER_156_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_570 ();
 DECAPx10_ASAP7_75t_R FILLER_156_599 ();
 DECAPx10_ASAP7_75t_R FILLER_156_621 ();
 DECAPx2_ASAP7_75t_R FILLER_156_643 ();
 FILLER_ASAP7_75t_R FILLER_156_649 ();
 DECAPx4_ASAP7_75t_R FILLER_156_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_681 ();
 DECAPx10_ASAP7_75t_R FILLER_156_724 ();
 DECAPx2_ASAP7_75t_R FILLER_156_746 ();
 DECAPx1_ASAP7_75t_R FILLER_156_759 ();
 DECAPx2_ASAP7_75t_R FILLER_156_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_789 ();
 DECAPx1_ASAP7_75t_R FILLER_156_810 ();
 DECAPx10_ASAP7_75t_R FILLER_156_821 ();
 FILLER_ASAP7_75t_R FILLER_156_843 ();
 DECAPx6_ASAP7_75t_R FILLER_156_867 ();
 FILLER_ASAP7_75t_R FILLER_156_881 ();
 DECAPx4_ASAP7_75t_R FILLER_156_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_915 ();
 DECAPx4_ASAP7_75t_R FILLER_156_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_948 ();
 DECAPx2_ASAP7_75t_R FILLER_156_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_969 ();
 FILLER_ASAP7_75t_R FILLER_156_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_991 ();
 FILLER_ASAP7_75t_R FILLER_156_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1025 ();
 DECAPx4_ASAP7_75t_R FILLER_156_1086 ();
 DECAPx4_ASAP7_75t_R FILLER_156_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_156_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1165 ();
 DECAPx4_ASAP7_75t_R FILLER_156_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_156_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_157_2 ();
 DECAPx10_ASAP7_75t_R FILLER_157_24 ();
 DECAPx10_ASAP7_75t_R FILLER_157_46 ();
 DECAPx10_ASAP7_75t_R FILLER_157_68 ();
 DECAPx4_ASAP7_75t_R FILLER_157_90 ();
 FILLER_ASAP7_75t_R FILLER_157_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_102 ();
 DECAPx6_ASAP7_75t_R FILLER_157_125 ();
 FILLER_ASAP7_75t_R FILLER_157_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_141 ();
 DECAPx6_ASAP7_75t_R FILLER_157_164 ();
 DECAPx2_ASAP7_75t_R FILLER_157_199 ();
 DECAPx1_ASAP7_75t_R FILLER_157_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_225 ();
 DECAPx1_ASAP7_75t_R FILLER_157_233 ();
 DECAPx4_ASAP7_75t_R FILLER_157_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_259 ();
 DECAPx1_ASAP7_75t_R FILLER_157_286 ();
 DECAPx10_ASAP7_75t_R FILLER_157_316 ();
 DECAPx6_ASAP7_75t_R FILLER_157_338 ();
 FILLER_ASAP7_75t_R FILLER_157_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_354 ();
 DECAPx6_ASAP7_75t_R FILLER_157_375 ();
 DECAPx1_ASAP7_75t_R FILLER_157_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_393 ();
 DECAPx6_ASAP7_75t_R FILLER_157_408 ();
 DECAPx1_ASAP7_75t_R FILLER_157_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_426 ();
 DECAPx4_ASAP7_75t_R FILLER_157_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_459 ();
 FILLER_ASAP7_75t_R FILLER_157_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_482 ();
 DECAPx1_ASAP7_75t_R FILLER_157_493 ();
 DECAPx2_ASAP7_75t_R FILLER_157_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_513 ();
 DECAPx4_ASAP7_75t_R FILLER_157_526 ();
 FILLER_ASAP7_75t_R FILLER_157_536 ();
 DECAPx1_ASAP7_75t_R FILLER_157_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_592 ();
 DECAPx10_ASAP7_75t_R FILLER_157_615 ();
 DECAPx6_ASAP7_75t_R FILLER_157_663 ();
 DECAPx1_ASAP7_75t_R FILLER_157_677 ();
 DECAPx10_ASAP7_75t_R FILLER_157_703 ();
 FILLER_ASAP7_75t_R FILLER_157_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_727 ();
 DECAPx2_ASAP7_75t_R FILLER_157_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_754 ();
 DECAPx1_ASAP7_75t_R FILLER_157_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_771 ();
 FILLER_ASAP7_75t_R FILLER_157_785 ();
 DECAPx6_ASAP7_75t_R FILLER_157_823 ();
 DECAPx2_ASAP7_75t_R FILLER_157_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_843 ();
 DECAPx4_ASAP7_75t_R FILLER_157_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_881 ();
 FILLER_ASAP7_75t_R FILLER_157_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_902 ();
 DECAPx4_ASAP7_75t_R FILLER_157_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_923 ();
 FILLER_ASAP7_75t_R FILLER_157_926 ();
 DECAPx4_ASAP7_75t_R FILLER_157_940 ();
 FILLER_ASAP7_75t_R FILLER_157_950 ();
 DECAPx2_ASAP7_75t_R FILLER_157_972 ();
 FILLER_ASAP7_75t_R FILLER_157_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_992 ();
 DECAPx1_ASAP7_75t_R FILLER_157_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1067 ();
 FILLER_ASAP7_75t_R FILLER_157_1073 ();
 FILLER_ASAP7_75t_R FILLER_157_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1105 ();
 FILLER_ASAP7_75t_R FILLER_157_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_157_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_157_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1198 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1208 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_158_2 ();
 DECAPx10_ASAP7_75t_R FILLER_158_24 ();
 DECAPx10_ASAP7_75t_R FILLER_158_46 ();
 DECAPx10_ASAP7_75t_R FILLER_158_68 ();
 DECAPx10_ASAP7_75t_R FILLER_158_90 ();
 DECAPx1_ASAP7_75t_R FILLER_158_112 ();
 DECAPx10_ASAP7_75t_R FILLER_158_127 ();
 DECAPx6_ASAP7_75t_R FILLER_158_149 ();
 FILLER_ASAP7_75t_R FILLER_158_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_165 ();
 DECAPx2_ASAP7_75t_R FILLER_158_183 ();
 FILLER_ASAP7_75t_R FILLER_158_189 ();
 FILLER_ASAP7_75t_R FILLER_158_231 ();
 FILLER_ASAP7_75t_R FILLER_158_240 ();
 DECAPx4_ASAP7_75t_R FILLER_158_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_260 ();
 DECAPx4_ASAP7_75t_R FILLER_158_267 ();
 FILLER_ASAP7_75t_R FILLER_158_277 ();
 DECAPx6_ASAP7_75t_R FILLER_158_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_313 ();
 FILLER_ASAP7_75t_R FILLER_158_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_338 ();
 FILLER_ASAP7_75t_R FILLER_158_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_347 ();
 FILLER_ASAP7_75t_R FILLER_158_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_360 ();
 DECAPx1_ASAP7_75t_R FILLER_158_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_371 ();
 DECAPx1_ASAP7_75t_R FILLER_158_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_382 ();
 FILLER_ASAP7_75t_R FILLER_158_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_392 ();
 FILLER_ASAP7_75t_R FILLER_158_415 ();
 DECAPx4_ASAP7_75t_R FILLER_158_430 ();
 FILLER_ASAP7_75t_R FILLER_158_440 ();
 DECAPx2_ASAP7_75t_R FILLER_158_464 ();
 DECAPx6_ASAP7_75t_R FILLER_158_476 ();
 DECAPx1_ASAP7_75t_R FILLER_158_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_494 ();
 DECAPx1_ASAP7_75t_R FILLER_158_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_509 ();
 DECAPx10_ASAP7_75t_R FILLER_158_516 ();
 DECAPx2_ASAP7_75t_R FILLER_158_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_544 ();
 DECAPx2_ASAP7_75t_R FILLER_158_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_568 ();
 DECAPx2_ASAP7_75t_R FILLER_158_575 ();
 FILLER_ASAP7_75t_R FILLER_158_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_583 ();
 DECAPx6_ASAP7_75t_R FILLER_158_595 ();
 DECAPx10_ASAP7_75t_R FILLER_158_631 ();
 DECAPx10_ASAP7_75t_R FILLER_158_653 ();
 DECAPx4_ASAP7_75t_R FILLER_158_675 ();
 FILLER_ASAP7_75t_R FILLER_158_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_687 ();
 DECAPx4_ASAP7_75t_R FILLER_158_691 ();
 DECAPx2_ASAP7_75t_R FILLER_158_711 ();
 FILLER_ASAP7_75t_R FILLER_158_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_719 ();
 DECAPx1_ASAP7_75t_R FILLER_158_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_742 ();
 DECAPx1_ASAP7_75t_R FILLER_158_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_754 ();
 DECAPx4_ASAP7_75t_R FILLER_158_761 ();
 FILLER_ASAP7_75t_R FILLER_158_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_773 ();
 DECAPx10_ASAP7_75t_R FILLER_158_784 ();
 FILLER_ASAP7_75t_R FILLER_158_806 ();
 DECAPx1_ASAP7_75t_R FILLER_158_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_825 ();
 FILLER_ASAP7_75t_R FILLER_158_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_844 ();
 FILLER_ASAP7_75t_R FILLER_158_865 ();
 DECAPx1_ASAP7_75t_R FILLER_158_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_875 ();
 FILLER_ASAP7_75t_R FILLER_158_937 ();
 DECAPx4_ASAP7_75t_R FILLER_158_947 ();
 FILLER_ASAP7_75t_R FILLER_158_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_966 ();
 DECAPx1_ASAP7_75t_R FILLER_158_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_993 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1007 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_158_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1054 ();
 FILLER_ASAP7_75t_R FILLER_158_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1092 ();
 FILLER_ASAP7_75t_R FILLER_158_1132 ();
 FILLER_ASAP7_75t_R FILLER_158_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_159_2 ();
 DECAPx10_ASAP7_75t_R FILLER_159_24 ();
 DECAPx10_ASAP7_75t_R FILLER_159_46 ();
 DECAPx10_ASAP7_75t_R FILLER_159_68 ();
 DECAPx10_ASAP7_75t_R FILLER_159_90 ();
 DECAPx2_ASAP7_75t_R FILLER_159_112 ();
 DECAPx6_ASAP7_75t_R FILLER_159_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_154 ();
 DECAPx1_ASAP7_75t_R FILLER_159_183 ();
 DECAPx10_ASAP7_75t_R FILLER_159_198 ();
 DECAPx4_ASAP7_75t_R FILLER_159_220 ();
 FILLER_ASAP7_75t_R FILLER_159_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_239 ();
 DECAPx6_ASAP7_75t_R FILLER_159_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_276 ();
 DECAPx4_ASAP7_75t_R FILLER_159_303 ();
 FILLER_ASAP7_75t_R FILLER_159_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_315 ();
 DECAPx1_ASAP7_75t_R FILLER_159_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_340 ();
 FILLER_ASAP7_75t_R FILLER_159_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_351 ();
 DECAPx1_ASAP7_75t_R FILLER_159_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_364 ();
 DECAPx1_ASAP7_75t_R FILLER_159_394 ();
 DECAPx6_ASAP7_75t_R FILLER_159_424 ();
 DECAPx2_ASAP7_75t_R FILLER_159_438 ();
 DECAPx2_ASAP7_75t_R FILLER_159_464 ();
 FILLER_ASAP7_75t_R FILLER_159_470 ();
 DECAPx6_ASAP7_75t_R FILLER_159_514 ();
 FILLER_ASAP7_75t_R FILLER_159_528 ();
 DECAPx10_ASAP7_75t_R FILLER_159_556 ();
 DECAPx2_ASAP7_75t_R FILLER_159_578 ();
 DECAPx2_ASAP7_75t_R FILLER_159_590 ();
 FILLER_ASAP7_75t_R FILLER_159_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_598 ();
 DECAPx10_ASAP7_75t_R FILLER_159_616 ();
 DECAPx6_ASAP7_75t_R FILLER_159_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_652 ();
 DECAPx6_ASAP7_75t_R FILLER_159_689 ();
 FILLER_ASAP7_75t_R FILLER_159_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_705 ();
 FILLER_ASAP7_75t_R FILLER_159_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_715 ();
 DECAPx2_ASAP7_75t_R FILLER_159_726 ();
 FILLER_ASAP7_75t_R FILLER_159_732 ();
 DECAPx1_ASAP7_75t_R FILLER_159_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_745 ();
 DECAPx2_ASAP7_75t_R FILLER_159_764 ();
 FILLER_ASAP7_75t_R FILLER_159_770 ();
 DECAPx4_ASAP7_75t_R FILLER_159_780 ();
 DECAPx1_ASAP7_75t_R FILLER_159_803 ();
 DECAPx2_ASAP7_75t_R FILLER_159_819 ();
 FILLER_ASAP7_75t_R FILLER_159_825 ();
 DECAPx4_ASAP7_75t_R FILLER_159_833 ();
 FILLER_ASAP7_75t_R FILLER_159_843 ();
 DECAPx2_ASAP7_75t_R FILLER_159_853 ();
 FILLER_ASAP7_75t_R FILLER_159_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_861 ();
 DECAPx6_ASAP7_75t_R FILLER_159_896 ();
 FILLER_ASAP7_75t_R FILLER_159_910 ();
 FILLER_ASAP7_75t_R FILLER_159_922 ();
 FILLER_ASAP7_75t_R FILLER_159_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_928 ();
 DECAPx6_ASAP7_75t_R FILLER_159_939 ();
 DECAPx1_ASAP7_75t_R FILLER_159_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_957 ();
 DECAPx1_ASAP7_75t_R FILLER_159_974 ();
 FILLER_ASAP7_75t_R FILLER_159_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_983 ();
 DECAPx1_ASAP7_75t_R FILLER_159_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1029 ();
 FILLER_ASAP7_75t_R FILLER_159_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_159_1059 ();
 FILLER_ASAP7_75t_R FILLER_159_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1086 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1100 ();
 FILLER_ASAP7_75t_R FILLER_159_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1178 ();
 FILLER_ASAP7_75t_R FILLER_159_1184 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1216 ();
 FILLER_ASAP7_75t_R FILLER_159_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_160_2 ();
 DECAPx10_ASAP7_75t_R FILLER_160_24 ();
 DECAPx10_ASAP7_75t_R FILLER_160_46 ();
 DECAPx10_ASAP7_75t_R FILLER_160_68 ();
 DECAPx10_ASAP7_75t_R FILLER_160_90 ();
 DECAPx4_ASAP7_75t_R FILLER_160_112 ();
 DECAPx10_ASAP7_75t_R FILLER_160_128 ();
 DECAPx10_ASAP7_75t_R FILLER_160_150 ();
 DECAPx4_ASAP7_75t_R FILLER_160_172 ();
 FILLER_ASAP7_75t_R FILLER_160_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_184 ();
 DECAPx2_ASAP7_75t_R FILLER_160_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_230 ();
 DECAPx10_ASAP7_75t_R FILLER_160_248 ();
 DECAPx4_ASAP7_75t_R FILLER_160_270 ();
 DECAPx6_ASAP7_75t_R FILLER_160_286 ();
 FILLER_ASAP7_75t_R FILLER_160_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_302 ();
 DECAPx2_ASAP7_75t_R FILLER_160_328 ();
 FILLER_ASAP7_75t_R FILLER_160_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_336 ();
 FILLER_ASAP7_75t_R FILLER_160_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_355 ();
 DECAPx6_ASAP7_75t_R FILLER_160_364 ();
 DECAPx6_ASAP7_75t_R FILLER_160_406 ();
 FILLER_ASAP7_75t_R FILLER_160_420 ();
 DECAPx4_ASAP7_75t_R FILLER_160_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_461 ();
 DECAPx4_ASAP7_75t_R FILLER_160_464 ();
 FILLER_ASAP7_75t_R FILLER_160_474 ();
 DECAPx10_ASAP7_75t_R FILLER_160_482 ();
 FILLER_ASAP7_75t_R FILLER_160_504 ();
 DECAPx2_ASAP7_75t_R FILLER_160_536 ();
 DECAPx4_ASAP7_75t_R FILLER_160_551 ();
 FILLER_ASAP7_75t_R FILLER_160_561 ();
 DECAPx1_ASAP7_75t_R FILLER_160_569 ();
 DECAPx1_ASAP7_75t_R FILLER_160_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_595 ();
 DECAPx1_ASAP7_75t_R FILLER_160_604 ();
 DECAPx1_ASAP7_75t_R FILLER_160_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_634 ();
 DECAPx10_ASAP7_75t_R FILLER_160_641 ();
 DECAPx1_ASAP7_75t_R FILLER_160_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_667 ();
 DECAPx6_ASAP7_75t_R FILLER_160_686 ();
 DECAPx1_ASAP7_75t_R FILLER_160_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_704 ();
 FILLER_ASAP7_75t_R FILLER_160_723 ();
 DECAPx2_ASAP7_75t_R FILLER_160_734 ();
 FILLER_ASAP7_75t_R FILLER_160_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_758 ();
 FILLER_ASAP7_75t_R FILLER_160_765 ();
 FILLER_ASAP7_75t_R FILLER_160_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_778 ();
 DECAPx6_ASAP7_75t_R FILLER_160_789 ();
 DECAPx2_ASAP7_75t_R FILLER_160_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_809 ();
 DECAPx2_ASAP7_75t_R FILLER_160_817 ();
 DECAPx2_ASAP7_75t_R FILLER_160_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_845 ();
 DECAPx6_ASAP7_75t_R FILLER_160_854 ();
 DECAPx2_ASAP7_75t_R FILLER_160_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_887 ();
 DECAPx6_ASAP7_75t_R FILLER_160_910 ();
 DECAPx1_ASAP7_75t_R FILLER_160_924 ();
 DECAPx2_ASAP7_75t_R FILLER_160_934 ();
 DECAPx10_ASAP7_75t_R FILLER_160_946 ();
 DECAPx1_ASAP7_75t_R FILLER_160_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_972 ();
 DECAPx2_ASAP7_75t_R FILLER_160_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_983 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1000 ();
 FILLER_ASAP7_75t_R FILLER_160_1010 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1111 ();
 FILLER_ASAP7_75t_R FILLER_160_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1131 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1144 ();
 FILLER_ASAP7_75t_R FILLER_160_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1180 ();
 FILLER_ASAP7_75t_R FILLER_160_1213 ();
 FILLER_ASAP7_75t_R FILLER_160_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_161_2 ();
 DECAPx10_ASAP7_75t_R FILLER_161_24 ();
 DECAPx10_ASAP7_75t_R FILLER_161_46 ();
 DECAPx10_ASAP7_75t_R FILLER_161_68 ();
 DECAPx10_ASAP7_75t_R FILLER_161_90 ();
 DECAPx10_ASAP7_75t_R FILLER_161_112 ();
 DECAPx10_ASAP7_75t_R FILLER_161_134 ();
 DECAPx4_ASAP7_75t_R FILLER_161_156 ();
 FILLER_ASAP7_75t_R FILLER_161_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_168 ();
 DECAPx10_ASAP7_75t_R FILLER_161_183 ();
 DECAPx4_ASAP7_75t_R FILLER_161_205 ();
 FILLER_ASAP7_75t_R FILLER_161_215 ();
 DECAPx1_ASAP7_75t_R FILLER_161_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_243 ();
 DECAPx1_ASAP7_75t_R FILLER_161_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_270 ();
 DECAPx1_ASAP7_75t_R FILLER_161_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_297 ();
 DECAPx1_ASAP7_75t_R FILLER_161_318 ();
 DECAPx6_ASAP7_75t_R FILLER_161_326 ();
 DECAPx6_ASAP7_75t_R FILLER_161_354 ();
 DECAPx1_ASAP7_75t_R FILLER_161_368 ();
 DECAPx1_ASAP7_75t_R FILLER_161_398 ();
 DECAPx2_ASAP7_75t_R FILLER_161_446 ();
 FILLER_ASAP7_75t_R FILLER_161_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_454 ();
 FILLER_ASAP7_75t_R FILLER_161_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_477 ();
 DECAPx10_ASAP7_75t_R FILLER_161_504 ();
 DECAPx6_ASAP7_75t_R FILLER_161_526 ();
 DECAPx1_ASAP7_75t_R FILLER_161_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_544 ();
 DECAPx2_ASAP7_75t_R FILLER_161_551 ();
 FILLER_ASAP7_75t_R FILLER_161_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_559 ();
 DECAPx4_ASAP7_75t_R FILLER_161_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_607 ();
 DECAPx1_ASAP7_75t_R FILLER_161_620 ();
 FILLER_ASAP7_75t_R FILLER_161_635 ();
 DECAPx4_ASAP7_75t_R FILLER_161_659 ();
 DECAPx6_ASAP7_75t_R FILLER_161_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_712 ();
 DECAPx2_ASAP7_75t_R FILLER_161_733 ();
 FILLER_ASAP7_75t_R FILLER_161_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_741 ();
 DECAPx2_ASAP7_75t_R FILLER_161_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_760 ();
 DECAPx1_ASAP7_75t_R FILLER_161_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_771 ();
 DECAPx4_ASAP7_75t_R FILLER_161_782 ();
 DECAPx1_ASAP7_75t_R FILLER_161_804 ();
 DECAPx2_ASAP7_75t_R FILLER_161_820 ();
 DECAPx2_ASAP7_75t_R FILLER_161_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_842 ();
 DECAPx10_ASAP7_75t_R FILLER_161_856 ();
 DECAPx10_ASAP7_75t_R FILLER_161_878 ();
 DECAPx10_ASAP7_75t_R FILLER_161_900 ();
 FILLER_ASAP7_75t_R FILLER_161_922 ();
 DECAPx1_ASAP7_75t_R FILLER_161_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_946 ();
 DECAPx1_ASAP7_75t_R FILLER_161_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_968 ();
 DECAPx1_ASAP7_75t_R FILLER_161_985 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1004 ();
 FILLER_ASAP7_75t_R FILLER_161_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1026 ();
 FILLER_ASAP7_75t_R FILLER_161_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1083 ();
 FILLER_ASAP7_75t_R FILLER_161_1093 ();
 FILLER_ASAP7_75t_R FILLER_161_1107 ();
 FILLER_ASAP7_75t_R FILLER_161_1117 ();
 FILLER_ASAP7_75t_R FILLER_161_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1154 ();
 FILLER_ASAP7_75t_R FILLER_161_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1205 ();
 FILLER_ASAP7_75t_R FILLER_161_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_162_2 ();
 DECAPx10_ASAP7_75t_R FILLER_162_24 ();
 DECAPx10_ASAP7_75t_R FILLER_162_46 ();
 DECAPx10_ASAP7_75t_R FILLER_162_68 ();
 DECAPx10_ASAP7_75t_R FILLER_162_90 ();
 DECAPx10_ASAP7_75t_R FILLER_162_112 ();
 DECAPx4_ASAP7_75t_R FILLER_162_134 ();
 FILLER_ASAP7_75t_R FILLER_162_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_146 ();
 DECAPx1_ASAP7_75t_R FILLER_162_169 ();
 DECAPx2_ASAP7_75t_R FILLER_162_212 ();
 FILLER_ASAP7_75t_R FILLER_162_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_220 ();
 FILLER_ASAP7_75t_R FILLER_162_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_229 ();
 DECAPx1_ASAP7_75t_R FILLER_162_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_245 ();
 DECAPx2_ASAP7_75t_R FILLER_162_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_258 ();
 DECAPx4_ASAP7_75t_R FILLER_162_265 ();
 DECAPx6_ASAP7_75t_R FILLER_162_281 ();
 DECAPx2_ASAP7_75t_R FILLER_162_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_301 ();
 DECAPx10_ASAP7_75t_R FILLER_162_305 ();
 DECAPx4_ASAP7_75t_R FILLER_162_327 ();
 FILLER_ASAP7_75t_R FILLER_162_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_339 ();
 FILLER_ASAP7_75t_R FILLER_162_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_350 ();
 DECAPx2_ASAP7_75t_R FILLER_162_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_367 ();
 DECAPx10_ASAP7_75t_R FILLER_162_375 ();
 DECAPx10_ASAP7_75t_R FILLER_162_397 ();
 DECAPx4_ASAP7_75t_R FILLER_162_432 ();
 DECAPx2_ASAP7_75t_R FILLER_162_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_470 ();
 FILLER_ASAP7_75t_R FILLER_162_491 ();
 FILLER_ASAP7_75t_R FILLER_162_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_503 ();
 DECAPx10_ASAP7_75t_R FILLER_162_510 ();
 DECAPx1_ASAP7_75t_R FILLER_162_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_536 ();
 DECAPx2_ASAP7_75t_R FILLER_162_570 ();
 FILLER_ASAP7_75t_R FILLER_162_576 ();
 DECAPx2_ASAP7_75t_R FILLER_162_614 ();
 DECAPx10_ASAP7_75t_R FILLER_162_626 ();
 DECAPx6_ASAP7_75t_R FILLER_162_648 ();
 DECAPx1_ASAP7_75t_R FILLER_162_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_689 ();
 DECAPx1_ASAP7_75t_R FILLER_162_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_716 ();
 DECAPx2_ASAP7_75t_R FILLER_162_737 ();
 DECAPx1_ASAP7_75t_R FILLER_162_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_774 ();
 FILLER_ASAP7_75t_R FILLER_162_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_784 ();
 DECAPx2_ASAP7_75t_R FILLER_162_791 ();
 DECAPx4_ASAP7_75t_R FILLER_162_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_813 ();
 DECAPx4_ASAP7_75t_R FILLER_162_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_841 ();
 DECAPx4_ASAP7_75t_R FILLER_162_876 ();
 FILLER_ASAP7_75t_R FILLER_162_886 ();
 DECAPx4_ASAP7_75t_R FILLER_162_910 ();
 FILLER_ASAP7_75t_R FILLER_162_920 ();
 FILLER_ASAP7_75t_R FILLER_162_942 ();
 DECAPx2_ASAP7_75t_R FILLER_162_951 ();
 FILLER_ASAP7_75t_R FILLER_162_957 ();
 DECAPx6_ASAP7_75t_R FILLER_162_969 ();
 DECAPx2_ASAP7_75t_R FILLER_162_983 ();
 FILLER_ASAP7_75t_R FILLER_162_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1092 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1099 ();
 FILLER_ASAP7_75t_R FILLER_162_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1115 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1125 ();
 FILLER_ASAP7_75t_R FILLER_162_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1148 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1175 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1199 ();
 FILLER_ASAP7_75t_R FILLER_162_1209 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_163_2 ();
 DECAPx10_ASAP7_75t_R FILLER_163_24 ();
 DECAPx10_ASAP7_75t_R FILLER_163_46 ();
 DECAPx10_ASAP7_75t_R FILLER_163_68 ();
 DECAPx10_ASAP7_75t_R FILLER_163_90 ();
 DECAPx6_ASAP7_75t_R FILLER_163_112 ();
 DECAPx1_ASAP7_75t_R FILLER_163_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_148 ();
 DECAPx4_ASAP7_75t_R FILLER_163_191 ();
 FILLER_ASAP7_75t_R FILLER_163_201 ();
 DECAPx10_ASAP7_75t_R FILLER_163_225 ();
 DECAPx2_ASAP7_75t_R FILLER_163_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_253 ();
 DECAPx6_ASAP7_75t_R FILLER_163_274 ();
 FILLER_ASAP7_75t_R FILLER_163_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_290 ();
 DECAPx2_ASAP7_75t_R FILLER_163_301 ();
 FILLER_ASAP7_75t_R FILLER_163_316 ();
 FILLER_ASAP7_75t_R FILLER_163_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_378 ();
 DECAPx10_ASAP7_75t_R FILLER_163_423 ();
 DECAPx6_ASAP7_75t_R FILLER_163_445 ();
 DECAPx2_ASAP7_75t_R FILLER_163_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_465 ();
 DECAPx1_ASAP7_75t_R FILLER_163_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_494 ();
 DECAPx6_ASAP7_75t_R FILLER_163_517 ();
 DECAPx2_ASAP7_75t_R FILLER_163_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_537 ();
 DECAPx10_ASAP7_75t_R FILLER_163_555 ();
 DECAPx1_ASAP7_75t_R FILLER_163_577 ();
 DECAPx6_ASAP7_75t_R FILLER_163_596 ();
 DECAPx10_ASAP7_75t_R FILLER_163_618 ();
 DECAPx10_ASAP7_75t_R FILLER_163_640 ();
 DECAPx6_ASAP7_75t_R FILLER_163_662 ();
 FILLER_ASAP7_75t_R FILLER_163_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_691 ();
 FILLER_ASAP7_75t_R FILLER_163_700 ();
 FILLER_ASAP7_75t_R FILLER_163_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_719 ();
 FILLER_ASAP7_75t_R FILLER_163_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_738 ();
 DECAPx1_ASAP7_75t_R FILLER_163_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_770 ();
 DECAPx2_ASAP7_75t_R FILLER_163_820 ();
 DECAPx2_ASAP7_75t_R FILLER_163_839 ();
 DECAPx4_ASAP7_75t_R FILLER_163_851 ();
 FILLER_ASAP7_75t_R FILLER_163_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_863 ();
 DECAPx1_ASAP7_75t_R FILLER_163_867 ();
 DECAPx10_ASAP7_75t_R FILLER_163_893 ();
 DECAPx2_ASAP7_75t_R FILLER_163_915 ();
 FILLER_ASAP7_75t_R FILLER_163_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_923 ();
 FILLER_ASAP7_75t_R FILLER_163_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_928 ();
 DECAPx1_ASAP7_75t_R FILLER_163_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_959 ();
 DECAPx2_ASAP7_75t_R FILLER_163_966 ();
 DECAPx1_ASAP7_75t_R FILLER_163_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_996 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1001 ();
 FILLER_ASAP7_75t_R FILLER_163_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1092 ();
 FILLER_ASAP7_75t_R FILLER_163_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1171 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1193 ();
 FILLER_ASAP7_75t_R FILLER_163_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1215 ();
 FILLER_ASAP7_75t_R FILLER_163_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_164_2 ();
 DECAPx10_ASAP7_75t_R FILLER_164_24 ();
 DECAPx10_ASAP7_75t_R FILLER_164_46 ();
 DECAPx10_ASAP7_75t_R FILLER_164_68 ();
 DECAPx10_ASAP7_75t_R FILLER_164_90 ();
 DECAPx6_ASAP7_75t_R FILLER_164_112 ();
 FILLER_ASAP7_75t_R FILLER_164_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_150 ();
 DECAPx4_ASAP7_75t_R FILLER_164_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_176 ();
 FILLER_ASAP7_75t_R FILLER_164_183 ();
 DECAPx10_ASAP7_75t_R FILLER_164_191 ();
 DECAPx2_ASAP7_75t_R FILLER_164_213 ();
 FILLER_ASAP7_75t_R FILLER_164_219 ();
 DECAPx6_ASAP7_75t_R FILLER_164_249 ();
 FILLER_ASAP7_75t_R FILLER_164_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_265 ();
 DECAPx4_ASAP7_75t_R FILLER_164_278 ();
 FILLER_ASAP7_75t_R FILLER_164_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_310 ();
 FILLER_ASAP7_75t_R FILLER_164_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_335 ();
 FILLER_ASAP7_75t_R FILLER_164_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_349 ();
 FILLER_ASAP7_75t_R FILLER_164_370 ();
 FILLER_ASAP7_75t_R FILLER_164_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_414 ();
 DECAPx10_ASAP7_75t_R FILLER_164_440 ();
 FILLER_ASAP7_75t_R FILLER_164_464 ();
 DECAPx10_ASAP7_75t_R FILLER_164_486 ();
 DECAPx6_ASAP7_75t_R FILLER_164_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_522 ();
 DECAPx10_ASAP7_75t_R FILLER_164_551 ();
 DECAPx1_ASAP7_75t_R FILLER_164_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_577 ();
 DECAPx4_ASAP7_75t_R FILLER_164_600 ();
 FILLER_ASAP7_75t_R FILLER_164_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_626 ();
 FILLER_ASAP7_75t_R FILLER_164_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_635 ();
 DECAPx10_ASAP7_75t_R FILLER_164_642 ();
 DECAPx6_ASAP7_75t_R FILLER_164_664 ();
 FILLER_ASAP7_75t_R FILLER_164_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_680 ();
 DECAPx2_ASAP7_75t_R FILLER_164_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_718 ();
 DECAPx6_ASAP7_75t_R FILLER_164_736 ();
 DECAPx1_ASAP7_75t_R FILLER_164_750 ();
 FILLER_ASAP7_75t_R FILLER_164_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_777 ();
 DECAPx1_ASAP7_75t_R FILLER_164_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_788 ();
 DECAPx4_ASAP7_75t_R FILLER_164_799 ();
 FILLER_ASAP7_75t_R FILLER_164_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_811 ();
 DECAPx1_ASAP7_75t_R FILLER_164_821 ();
 DECAPx1_ASAP7_75t_R FILLER_164_843 ();
 DECAPx4_ASAP7_75t_R FILLER_164_853 ();
 FILLER_ASAP7_75t_R FILLER_164_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_865 ();
 FILLER_ASAP7_75t_R FILLER_164_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_888 ();
 DECAPx2_ASAP7_75t_R FILLER_164_893 ();
 FILLER_ASAP7_75t_R FILLER_164_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_901 ();
 DECAPx4_ASAP7_75t_R FILLER_164_922 ();
 FILLER_ASAP7_75t_R FILLER_164_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_944 ();
 DECAPx4_ASAP7_75t_R FILLER_164_948 ();
 DECAPx1_ASAP7_75t_R FILLER_164_965 ();
 DECAPx10_ASAP7_75t_R FILLER_164_978 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1000 ();
 FILLER_ASAP7_75t_R FILLER_164_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_164_1029 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1122 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1152 ();
 DECAPx6_ASAP7_75t_R FILLER_164_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1182 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1211 ();
 FILLER_ASAP7_75t_R FILLER_164_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_165_2 ();
 DECAPx10_ASAP7_75t_R FILLER_165_24 ();
 DECAPx10_ASAP7_75t_R FILLER_165_46 ();
 DECAPx10_ASAP7_75t_R FILLER_165_68 ();
 DECAPx10_ASAP7_75t_R FILLER_165_90 ();
 DECAPx10_ASAP7_75t_R FILLER_165_112 ();
 DECAPx6_ASAP7_75t_R FILLER_165_134 ();
 DECAPx10_ASAP7_75t_R FILLER_165_203 ();
 DECAPx6_ASAP7_75t_R FILLER_165_225 ();
 DECAPx1_ASAP7_75t_R FILLER_165_239 ();
 DECAPx4_ASAP7_75t_R FILLER_165_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_259 ();
 FILLER_ASAP7_75t_R FILLER_165_266 ();
 DECAPx2_ASAP7_75t_R FILLER_165_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_294 ();
 DECAPx6_ASAP7_75t_R FILLER_165_317 ();
 FILLER_ASAP7_75t_R FILLER_165_342 ();
 DECAPx10_ASAP7_75t_R FILLER_165_365 ();
 DECAPx6_ASAP7_75t_R FILLER_165_387 ();
 DECAPx1_ASAP7_75t_R FILLER_165_401 ();
 DECAPx10_ASAP7_75t_R FILLER_165_411 ();
 DECAPx10_ASAP7_75t_R FILLER_165_433 ();
 DECAPx6_ASAP7_75t_R FILLER_165_455 ();
 DECAPx6_ASAP7_75t_R FILLER_165_475 ();
 DECAPx2_ASAP7_75t_R FILLER_165_489 ();
 DECAPx10_ASAP7_75t_R FILLER_165_517 ();
 DECAPx1_ASAP7_75t_R FILLER_165_539 ();
 DECAPx1_ASAP7_75t_R FILLER_165_550 ();
 DECAPx6_ASAP7_75t_R FILLER_165_582 ();
 DECAPx1_ASAP7_75t_R FILLER_165_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_634 ();
 DECAPx6_ASAP7_75t_R FILLER_165_657 ();
 DECAPx1_ASAP7_75t_R FILLER_165_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_690 ();
 DECAPx1_ASAP7_75t_R FILLER_165_697 ();
 DECAPx2_ASAP7_75t_R FILLER_165_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_722 ();
 FILLER_ASAP7_75t_R FILLER_165_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_738 ();
 DECAPx6_ASAP7_75t_R FILLER_165_742 ();
 DECAPx4_ASAP7_75t_R FILLER_165_759 ();
 FILLER_ASAP7_75t_R FILLER_165_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_771 ();
 DECAPx10_ASAP7_75t_R FILLER_165_775 ();
 DECAPx4_ASAP7_75t_R FILLER_165_797 ();
 FILLER_ASAP7_75t_R FILLER_165_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_809 ();
 DECAPx2_ASAP7_75t_R FILLER_165_822 ();
 FILLER_ASAP7_75t_R FILLER_165_828 ();
 DECAPx1_ASAP7_75t_R FILLER_165_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_847 ();
 DECAPx1_ASAP7_75t_R FILLER_165_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_860 ();
 DECAPx6_ASAP7_75t_R FILLER_165_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_895 ();
 FILLER_ASAP7_75t_R FILLER_165_922 ();
 DECAPx4_ASAP7_75t_R FILLER_165_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_936 ();
 FILLER_ASAP7_75t_R FILLER_165_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_953 ();
 FILLER_ASAP7_75t_R FILLER_165_970 ();
 FILLER_ASAP7_75t_R FILLER_165_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_988 ();
 FILLER_ASAP7_75t_R FILLER_165_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_994 ();
 FILLER_ASAP7_75t_R FILLER_165_1001 ();
 FILLER_ASAP7_75t_R FILLER_165_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1011 ();
 FILLER_ASAP7_75t_R FILLER_165_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1024 ();
 FILLER_ASAP7_75t_R FILLER_165_1045 ();
 DECAPx1_ASAP7_75t_R FILLER_165_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1081 ();
 DECAPx4_ASAP7_75t_R FILLER_165_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_165_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1153 ();
 FILLER_ASAP7_75t_R FILLER_165_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1164 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1186 ();
 DECAPx4_ASAP7_75t_R FILLER_165_1206 ();
 FILLER_ASAP7_75t_R FILLER_165_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_166_2 ();
 DECAPx10_ASAP7_75t_R FILLER_166_24 ();
 DECAPx10_ASAP7_75t_R FILLER_166_46 ();
 DECAPx10_ASAP7_75t_R FILLER_166_68 ();
 DECAPx10_ASAP7_75t_R FILLER_166_90 ();
 DECAPx10_ASAP7_75t_R FILLER_166_112 ();
 DECAPx2_ASAP7_75t_R FILLER_166_144 ();
 DECAPx6_ASAP7_75t_R FILLER_166_173 ();
 FILLER_ASAP7_75t_R FILLER_166_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_200 ();
 DECAPx4_ASAP7_75t_R FILLER_166_229 ();
 FILLER_ASAP7_75t_R FILLER_166_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_241 ();
 DECAPx10_ASAP7_75t_R FILLER_166_264 ();
 DECAPx4_ASAP7_75t_R FILLER_166_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_302 ();
 DECAPx2_ASAP7_75t_R FILLER_166_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_338 ();
 DECAPx6_ASAP7_75t_R FILLER_166_378 ();
 FILLER_ASAP7_75t_R FILLER_166_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_394 ();
 DECAPx6_ASAP7_75t_R FILLER_166_421 ();
 DECAPx1_ASAP7_75t_R FILLER_166_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_461 ();
 FILLER_ASAP7_75t_R FILLER_166_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_466 ();
 DECAPx2_ASAP7_75t_R FILLER_166_475 ();
 FILLER_ASAP7_75t_R FILLER_166_481 ();
 DECAPx2_ASAP7_75t_R FILLER_166_499 ();
 FILLER_ASAP7_75t_R FILLER_166_505 ();
 DECAPx4_ASAP7_75t_R FILLER_166_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_545 ();
 FILLER_ASAP7_75t_R FILLER_166_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_561 ();
 FILLER_ASAP7_75t_R FILLER_166_568 ();
 DECAPx6_ASAP7_75t_R FILLER_166_582 ();
 FILLER_ASAP7_75t_R FILLER_166_596 ();
 DECAPx2_ASAP7_75t_R FILLER_166_620 ();
 FILLER_ASAP7_75t_R FILLER_166_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_628 ();
 DECAPx10_ASAP7_75t_R FILLER_166_640 ();
 DECAPx6_ASAP7_75t_R FILLER_166_662 ();
 DECAPx2_ASAP7_75t_R FILLER_166_676 ();
 DECAPx4_ASAP7_75t_R FILLER_166_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_704 ();
 DECAPx2_ASAP7_75t_R FILLER_166_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_717 ();
 DECAPx1_ASAP7_75t_R FILLER_166_725 ();
 DECAPx1_ASAP7_75t_R FILLER_166_735 ();
 DECAPx4_ASAP7_75t_R FILLER_166_749 ();
 FILLER_ASAP7_75t_R FILLER_166_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_761 ();
 DECAPx1_ASAP7_75t_R FILLER_166_786 ();
 DECAPx2_ASAP7_75t_R FILLER_166_802 ();
 DECAPx10_ASAP7_75t_R FILLER_166_820 ();
 DECAPx2_ASAP7_75t_R FILLER_166_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_848 ();
 DECAPx10_ASAP7_75t_R FILLER_166_856 ();
 FILLER_ASAP7_75t_R FILLER_166_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_880 ();
 FILLER_ASAP7_75t_R FILLER_166_925 ();
 FILLER_ASAP7_75t_R FILLER_166_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_945 ();
 FILLER_ASAP7_75t_R FILLER_166_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_992 ();
 DECAPx2_ASAP7_75t_R FILLER_166_996 ();
 FILLER_ASAP7_75t_R FILLER_166_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_166_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1118 ();
 FILLER_ASAP7_75t_R FILLER_166_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1185 ();
 FILLER_ASAP7_75t_R FILLER_166_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_167_2 ();
 DECAPx10_ASAP7_75t_R FILLER_167_24 ();
 DECAPx10_ASAP7_75t_R FILLER_167_46 ();
 DECAPx10_ASAP7_75t_R FILLER_167_68 ();
 DECAPx10_ASAP7_75t_R FILLER_167_90 ();
 DECAPx6_ASAP7_75t_R FILLER_167_112 ();
 FILLER_ASAP7_75t_R FILLER_167_126 ();
 DECAPx2_ASAP7_75t_R FILLER_167_138 ();
 DECAPx2_ASAP7_75t_R FILLER_167_150 ();
 DECAPx6_ASAP7_75t_R FILLER_167_170 ();
 DECAPx2_ASAP7_75t_R FILLER_167_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_190 ();
 FILLER_ASAP7_75t_R FILLER_167_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_199 ();
 DECAPx1_ASAP7_75t_R FILLER_167_231 ();
 DECAPx4_ASAP7_75t_R FILLER_167_245 ();
 FILLER_ASAP7_75t_R FILLER_167_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_257 ();
 DECAPx6_ASAP7_75t_R FILLER_167_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_278 ();
 DECAPx6_ASAP7_75t_R FILLER_167_285 ();
 FILLER_ASAP7_75t_R FILLER_167_299 ();
 FILLER_ASAP7_75t_R FILLER_167_313 ();
 FILLER_ASAP7_75t_R FILLER_167_332 ();
 FILLER_ASAP7_75t_R FILLER_167_347 ();
 DECAPx6_ASAP7_75t_R FILLER_167_356 ();
 DECAPx1_ASAP7_75t_R FILLER_167_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_396 ();
 DECAPx6_ASAP7_75t_R FILLER_167_431 ();
 DECAPx1_ASAP7_75t_R FILLER_167_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_470 ();
 DECAPx1_ASAP7_75t_R FILLER_167_491 ();
 DECAPx2_ASAP7_75t_R FILLER_167_515 ();
 FILLER_ASAP7_75t_R FILLER_167_521 ();
 FILLER_ASAP7_75t_R FILLER_167_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_547 ();
 DECAPx2_ASAP7_75t_R FILLER_167_554 ();
 DECAPx4_ASAP7_75t_R FILLER_167_568 ();
 DECAPx10_ASAP7_75t_R FILLER_167_595 ();
 FILLER_ASAP7_75t_R FILLER_167_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_619 ();
 DECAPx6_ASAP7_75t_R FILLER_167_684 ();
 FILLER_ASAP7_75t_R FILLER_167_698 ();
 DECAPx4_ASAP7_75t_R FILLER_167_710 ();
 DECAPx1_ASAP7_75t_R FILLER_167_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_753 ();
 DECAPx1_ASAP7_75t_R FILLER_167_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_764 ();
 DECAPx1_ASAP7_75t_R FILLER_167_771 ();
 DECAPx4_ASAP7_75t_R FILLER_167_781 ();
 FILLER_ASAP7_75t_R FILLER_167_791 ();
 DECAPx4_ASAP7_75t_R FILLER_167_799 ();
 DECAPx1_ASAP7_75t_R FILLER_167_821 ();
 DECAPx2_ASAP7_75t_R FILLER_167_838 ();
 DECAPx10_ASAP7_75t_R FILLER_167_856 ();
 DECAPx10_ASAP7_75t_R FILLER_167_878 ();
 DECAPx10_ASAP7_75t_R FILLER_167_900 ();
 FILLER_ASAP7_75t_R FILLER_167_922 ();
 DECAPx10_ASAP7_75t_R FILLER_167_940 ();
 DECAPx10_ASAP7_75t_R FILLER_167_962 ();
 DECAPx6_ASAP7_75t_R FILLER_167_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1014 ();
 FILLER_ASAP7_75t_R FILLER_167_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_167_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1091 ();
 FILLER_ASAP7_75t_R FILLER_167_1098 ();
 FILLER_ASAP7_75t_R FILLER_167_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_167_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1201 ();
 FILLER_ASAP7_75t_R FILLER_167_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1216 ();
 FILLER_ASAP7_75t_R FILLER_167_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_168_2 ();
 DECAPx10_ASAP7_75t_R FILLER_168_24 ();
 DECAPx10_ASAP7_75t_R FILLER_168_46 ();
 DECAPx10_ASAP7_75t_R FILLER_168_68 ();
 DECAPx10_ASAP7_75t_R FILLER_168_90 ();
 DECAPx2_ASAP7_75t_R FILLER_168_112 ();
 FILLER_ASAP7_75t_R FILLER_168_118 ();
 DECAPx1_ASAP7_75t_R FILLER_168_130 ();
 DECAPx6_ASAP7_75t_R FILLER_168_163 ();
 DECAPx4_ASAP7_75t_R FILLER_168_185 ();
 FILLER_ASAP7_75t_R FILLER_168_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_197 ();
 DECAPx1_ASAP7_75t_R FILLER_168_218 ();
 DECAPx10_ASAP7_75t_R FILLER_168_248 ();
 DECAPx6_ASAP7_75t_R FILLER_168_292 ();
 FILLER_ASAP7_75t_R FILLER_168_306 ();
 DECAPx1_ASAP7_75t_R FILLER_168_314 ();
 FILLER_ASAP7_75t_R FILLER_168_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_333 ();
 DECAPx1_ASAP7_75t_R FILLER_168_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_347 ();
 DECAPx10_ASAP7_75t_R FILLER_168_356 ();
 DECAPx4_ASAP7_75t_R FILLER_168_378 ();
 FILLER_ASAP7_75t_R FILLER_168_388 ();
 DECAPx1_ASAP7_75t_R FILLER_168_412 ();
 DECAPx2_ASAP7_75t_R FILLER_168_436 ();
 FILLER_ASAP7_75t_R FILLER_168_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_466 ();
 DECAPx6_ASAP7_75t_R FILLER_168_481 ();
 DECAPx2_ASAP7_75t_R FILLER_168_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_501 ();
 FILLER_ASAP7_75t_R FILLER_168_510 ();
 DECAPx2_ASAP7_75t_R FILLER_168_522 ();
 FILLER_ASAP7_75t_R FILLER_168_556 ();
 DECAPx1_ASAP7_75t_R FILLER_168_572 ();
 DECAPx10_ASAP7_75t_R FILLER_168_584 ();
 DECAPx4_ASAP7_75t_R FILLER_168_606 ();
 FILLER_ASAP7_75t_R FILLER_168_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_618 ();
 DECAPx10_ASAP7_75t_R FILLER_168_631 ();
 DECAPx6_ASAP7_75t_R FILLER_168_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_667 ();
 DECAPx4_ASAP7_75t_R FILLER_168_690 ();
 FILLER_ASAP7_75t_R FILLER_168_700 ();
 DECAPx10_ASAP7_75t_R FILLER_168_714 ();
 DECAPx1_ASAP7_75t_R FILLER_168_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_740 ();
 FILLER_ASAP7_75t_R FILLER_168_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_757 ();
 FILLER_ASAP7_75t_R FILLER_168_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_784 ();
 DECAPx1_ASAP7_75t_R FILLER_168_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_802 ();
 DECAPx1_ASAP7_75t_R FILLER_168_816 ();
 FILLER_ASAP7_75t_R FILLER_168_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_847 ();
 FILLER_ASAP7_75t_R FILLER_168_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_857 ();
 DECAPx10_ASAP7_75t_R FILLER_168_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_925 ();
 DECAPx6_ASAP7_75t_R FILLER_168_950 ();
 DECAPx1_ASAP7_75t_R FILLER_168_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_968 ();
 DECAPx1_ASAP7_75t_R FILLER_168_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_976 ();
 DECAPx4_ASAP7_75t_R FILLER_168_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_168_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1107 ();
 FILLER_ASAP7_75t_R FILLER_168_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1123 ();
 FILLER_ASAP7_75t_R FILLER_168_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_168_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_168_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_169_2 ();
 DECAPx10_ASAP7_75t_R FILLER_169_24 ();
 DECAPx10_ASAP7_75t_R FILLER_169_46 ();
 DECAPx10_ASAP7_75t_R FILLER_169_68 ();
 DECAPx10_ASAP7_75t_R FILLER_169_90 ();
 DECAPx10_ASAP7_75t_R FILLER_169_112 ();
 DECAPx1_ASAP7_75t_R FILLER_169_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_138 ();
 DECAPx4_ASAP7_75t_R FILLER_169_150 ();
 DECAPx1_ASAP7_75t_R FILLER_169_182 ();
 DECAPx6_ASAP7_75t_R FILLER_169_210 ();
 FILLER_ASAP7_75t_R FILLER_169_224 ();
 DECAPx6_ASAP7_75t_R FILLER_169_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_250 ();
 DECAPx1_ASAP7_75t_R FILLER_169_277 ();
 DECAPx6_ASAP7_75t_R FILLER_169_309 ();
 DECAPx2_ASAP7_75t_R FILLER_169_323 ();
 FILLER_ASAP7_75t_R FILLER_169_349 ();
 DECAPx10_ASAP7_75t_R FILLER_169_362 ();
 FILLER_ASAP7_75t_R FILLER_169_384 ();
 DECAPx10_ASAP7_75t_R FILLER_169_406 ();
 DECAPx6_ASAP7_75t_R FILLER_169_450 ();
 FILLER_ASAP7_75t_R FILLER_169_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_466 ();
 DECAPx10_ASAP7_75t_R FILLER_169_489 ();
 DECAPx2_ASAP7_75t_R FILLER_169_511 ();
 FILLER_ASAP7_75t_R FILLER_169_517 ();
 DECAPx2_ASAP7_75t_R FILLER_169_552 ();
 FILLER_ASAP7_75t_R FILLER_169_606 ();
 FILLER_ASAP7_75t_R FILLER_169_624 ();
 DECAPx6_ASAP7_75t_R FILLER_169_643 ();
 DECAPx1_ASAP7_75t_R FILLER_169_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_738 ();
 FILLER_ASAP7_75t_R FILLER_169_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_760 ();
 DECAPx2_ASAP7_75t_R FILLER_169_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_773 ();
 FILLER_ASAP7_75t_R FILLER_169_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_788 ();
 DECAPx1_ASAP7_75t_R FILLER_169_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_805 ();
 DECAPx4_ASAP7_75t_R FILLER_169_818 ();
 FILLER_ASAP7_75t_R FILLER_169_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_830 ();
 DECAPx4_ASAP7_75t_R FILLER_169_837 ();
 FILLER_ASAP7_75t_R FILLER_169_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_849 ();
 DECAPx4_ASAP7_75t_R FILLER_169_879 ();
 FILLER_ASAP7_75t_R FILLER_169_889 ();
 DECAPx4_ASAP7_75t_R FILLER_169_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_923 ();
 DECAPx2_ASAP7_75t_R FILLER_169_926 ();
 FILLER_ASAP7_75t_R FILLER_169_932 ();
 FILLER_ASAP7_75t_R FILLER_169_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_952 ();
 DECAPx4_ASAP7_75t_R FILLER_169_975 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1013 ();
 FILLER_ASAP7_75t_R FILLER_169_1038 ();
 DECAPx6_ASAP7_75t_R FILLER_169_1046 ();
 FILLER_ASAP7_75t_R FILLER_169_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_170_2 ();
 DECAPx10_ASAP7_75t_R FILLER_170_24 ();
 DECAPx10_ASAP7_75t_R FILLER_170_46 ();
 DECAPx10_ASAP7_75t_R FILLER_170_68 ();
 DECAPx10_ASAP7_75t_R FILLER_170_90 ();
 DECAPx1_ASAP7_75t_R FILLER_170_112 ();
 DECAPx10_ASAP7_75t_R FILLER_170_122 ();
 FILLER_ASAP7_75t_R FILLER_170_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_146 ();
 FILLER_ASAP7_75t_R FILLER_170_153 ();
 DECAPx1_ASAP7_75t_R FILLER_170_171 ();
 DECAPx10_ASAP7_75t_R FILLER_170_192 ();
 DECAPx10_ASAP7_75t_R FILLER_170_214 ();
 FILLER_ASAP7_75t_R FILLER_170_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_238 ();
 DECAPx1_ASAP7_75t_R FILLER_170_259 ();
 FILLER_ASAP7_75t_R FILLER_170_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_311 ();
 DECAPx1_ASAP7_75t_R FILLER_170_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_334 ();
 DECAPx2_ASAP7_75t_R FILLER_170_343 ();
 FILLER_ASAP7_75t_R FILLER_170_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_351 ();
 DECAPx10_ASAP7_75t_R FILLER_170_355 ();
 DECAPx10_ASAP7_75t_R FILLER_170_377 ();
 DECAPx6_ASAP7_75t_R FILLER_170_399 ();
 FILLER_ASAP7_75t_R FILLER_170_413 ();
 DECAPx1_ASAP7_75t_R FILLER_170_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_441 ();
 DECAPx1_ASAP7_75t_R FILLER_170_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_468 ();
 DECAPx1_ASAP7_75t_R FILLER_170_475 ();
 DECAPx4_ASAP7_75t_R FILLER_170_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_493 ();
 FILLER_ASAP7_75t_R FILLER_170_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_511 ();
 DECAPx2_ASAP7_75t_R FILLER_170_532 ();
 DECAPx1_ASAP7_75t_R FILLER_170_548 ();
 DECAPx6_ASAP7_75t_R FILLER_170_573 ();
 DECAPx1_ASAP7_75t_R FILLER_170_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_591 ();
 FILLER_ASAP7_75t_R FILLER_170_605 ();
 DECAPx1_ASAP7_75t_R FILLER_170_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_617 ();
 FILLER_ASAP7_75t_R FILLER_170_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_634 ();
 DECAPx10_ASAP7_75t_R FILLER_170_657 ();
 DECAPx10_ASAP7_75t_R FILLER_170_679 ();
 DECAPx4_ASAP7_75t_R FILLER_170_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_737 ();
 DECAPx4_ASAP7_75t_R FILLER_170_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_792 ();
 DECAPx2_ASAP7_75t_R FILLER_170_800 ();
 FILLER_ASAP7_75t_R FILLER_170_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_808 ();
 DECAPx4_ASAP7_75t_R FILLER_170_822 ();
 FILLER_ASAP7_75t_R FILLER_170_832 ();
 DECAPx1_ASAP7_75t_R FILLER_170_841 ();
 DECAPx10_ASAP7_75t_R FILLER_170_857 ();
 DECAPx10_ASAP7_75t_R FILLER_170_879 ();
 DECAPx10_ASAP7_75t_R FILLER_170_901 ();
 DECAPx2_ASAP7_75t_R FILLER_170_923 ();
 FILLER_ASAP7_75t_R FILLER_170_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_931 ();
 DECAPx2_ASAP7_75t_R FILLER_170_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_952 ();
 DECAPx1_ASAP7_75t_R FILLER_170_960 ();
 DECAPx6_ASAP7_75t_R FILLER_170_984 ();
 DECAPx1_ASAP7_75t_R FILLER_170_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1064 ();
 FILLER_ASAP7_75t_R FILLER_170_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1072 ();
 FILLER_ASAP7_75t_R FILLER_170_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1103 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1148 ();
 FILLER_ASAP7_75t_R FILLER_170_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1160 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1195 ();
 FILLER_ASAP7_75t_R FILLER_170_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1203 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1212 ();
 FILLER_ASAP7_75t_R FILLER_170_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_171_2 ();
 DECAPx10_ASAP7_75t_R FILLER_171_24 ();
 DECAPx10_ASAP7_75t_R FILLER_171_46 ();
 DECAPx10_ASAP7_75t_R FILLER_171_68 ();
 DECAPx10_ASAP7_75t_R FILLER_171_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_112 ();
 DECAPx1_ASAP7_75t_R FILLER_171_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_137 ();
 DECAPx2_ASAP7_75t_R FILLER_171_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_175 ();
 DECAPx2_ASAP7_75t_R FILLER_171_198 ();
 FILLER_ASAP7_75t_R FILLER_171_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_206 ();
 FILLER_ASAP7_75t_R FILLER_171_215 ();
 DECAPx10_ASAP7_75t_R FILLER_171_223 ();
 DECAPx4_ASAP7_75t_R FILLER_171_245 ();
 DECAPx1_ASAP7_75t_R FILLER_171_261 ();
 DECAPx4_ASAP7_75t_R FILLER_171_287 ();
 DECAPx2_ASAP7_75t_R FILLER_171_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_331 ();
 FILLER_ASAP7_75t_R FILLER_171_340 ();
 FILLER_ASAP7_75t_R FILLER_171_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_359 ();
 DECAPx2_ASAP7_75t_R FILLER_171_402 ();
 DECAPx6_ASAP7_75t_R FILLER_171_414 ();
 DECAPx4_ASAP7_75t_R FILLER_171_434 ();
 FILLER_ASAP7_75t_R FILLER_171_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_446 ();
 DECAPx4_ASAP7_75t_R FILLER_171_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_460 ();
 DECAPx1_ASAP7_75t_R FILLER_171_467 ();
 DECAPx2_ASAP7_75t_R FILLER_171_477 ();
 FILLER_ASAP7_75t_R FILLER_171_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_485 ();
 FILLER_ASAP7_75t_R FILLER_171_500 ();
 DECAPx10_ASAP7_75t_R FILLER_171_508 ();
 DECAPx10_ASAP7_75t_R FILLER_171_530 ();
 DECAPx1_ASAP7_75t_R FILLER_171_552 ();
 DECAPx2_ASAP7_75t_R FILLER_171_562 ();
 DECAPx2_ASAP7_75t_R FILLER_171_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_580 ();
 DECAPx10_ASAP7_75t_R FILLER_171_613 ();
 DECAPx10_ASAP7_75t_R FILLER_171_635 ();
 DECAPx4_ASAP7_75t_R FILLER_171_657 ();
 FILLER_ASAP7_75t_R FILLER_171_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_669 ();
 DECAPx10_ASAP7_75t_R FILLER_171_710 ();
 FILLER_ASAP7_75t_R FILLER_171_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_734 ();
 DECAPx1_ASAP7_75t_R FILLER_171_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_761 ();
 DECAPx10_ASAP7_75t_R FILLER_171_783 ();
 FILLER_ASAP7_75t_R FILLER_171_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_807 ();
 DECAPx1_ASAP7_75t_R FILLER_171_826 ();
 DECAPx2_ASAP7_75t_R FILLER_171_842 ();
 FILLER_ASAP7_75t_R FILLER_171_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_857 ();
 DECAPx4_ASAP7_75t_R FILLER_171_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_888 ();
 DECAPx4_ASAP7_75t_R FILLER_171_911 ();
 FILLER_ASAP7_75t_R FILLER_171_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_923 ();
 DECAPx2_ASAP7_75t_R FILLER_171_926 ();
 FILLER_ASAP7_75t_R FILLER_171_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_934 ();
 DECAPx2_ASAP7_75t_R FILLER_171_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_950 ();
 DECAPx1_ASAP7_75t_R FILLER_171_968 ();
 DECAPx2_ASAP7_75t_R FILLER_171_975 ();
 FILLER_ASAP7_75t_R FILLER_171_981 ();
 FILLER_ASAP7_75t_R FILLER_171_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1126 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1183 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_172_2 ();
 DECAPx10_ASAP7_75t_R FILLER_172_24 ();
 DECAPx10_ASAP7_75t_R FILLER_172_46 ();
 DECAPx10_ASAP7_75t_R FILLER_172_68 ();
 DECAPx10_ASAP7_75t_R FILLER_172_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_112 ();
 FILLER_ASAP7_75t_R FILLER_172_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_130 ();
 DECAPx10_ASAP7_75t_R FILLER_172_137 ();
 FILLER_ASAP7_75t_R FILLER_172_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_167 ();
 DECAPx10_ASAP7_75t_R FILLER_172_180 ();
 FILLER_ASAP7_75t_R FILLER_172_220 ();
 DECAPx2_ASAP7_75t_R FILLER_172_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_256 ();
 DECAPx1_ASAP7_75t_R FILLER_172_277 ();
 FILLER_ASAP7_75t_R FILLER_172_303 ();
 FILLER_ASAP7_75t_R FILLER_172_324 ();
 DECAPx1_ASAP7_75t_R FILLER_172_336 ();
 DECAPx10_ASAP7_75t_R FILLER_172_350 ();
 DECAPx2_ASAP7_75t_R FILLER_172_372 ();
 FILLER_ASAP7_75t_R FILLER_172_378 ();
 FILLER_ASAP7_75t_R FILLER_172_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_427 ();
 DECAPx4_ASAP7_75t_R FILLER_172_450 ();
 FILLER_ASAP7_75t_R FILLER_172_460 ();
 DECAPx10_ASAP7_75t_R FILLER_172_464 ();
 FILLER_ASAP7_75t_R FILLER_172_498 ();
 FILLER_ASAP7_75t_R FILLER_172_511 ();
 DECAPx1_ASAP7_75t_R FILLER_172_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_543 ();
 DECAPx4_ASAP7_75t_R FILLER_172_555 ();
 FILLER_ASAP7_75t_R FILLER_172_565 ();
 DECAPx6_ASAP7_75t_R FILLER_172_577 ();
 DECAPx1_ASAP7_75t_R FILLER_172_591 ();
 DECAPx2_ASAP7_75t_R FILLER_172_610 ();
 FILLER_ASAP7_75t_R FILLER_172_616 ();
 DECAPx10_ASAP7_75t_R FILLER_172_629 ();
 DECAPx4_ASAP7_75t_R FILLER_172_651 ();
 FILLER_ASAP7_75t_R FILLER_172_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_663 ();
 DECAPx10_ASAP7_75t_R FILLER_172_667 ();
 DECAPx1_ASAP7_75t_R FILLER_172_689 ();
 DECAPx2_ASAP7_75t_R FILLER_172_699 ();
 FILLER_ASAP7_75t_R FILLER_172_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_707 ();
 FILLER_ASAP7_75t_R FILLER_172_734 ();
 DECAPx4_ASAP7_75t_R FILLER_172_748 ();
 FILLER_ASAP7_75t_R FILLER_172_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_760 ();
 DECAPx2_ASAP7_75t_R FILLER_172_767 ();
 FILLER_ASAP7_75t_R FILLER_172_773 ();
 DECAPx1_ASAP7_75t_R FILLER_172_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_799 ();
 FILLER_ASAP7_75t_R FILLER_172_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_809 ();
 DECAPx4_ASAP7_75t_R FILLER_172_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_834 ();
 DECAPx2_ASAP7_75t_R FILLER_172_842 ();
 DECAPx2_ASAP7_75t_R FILLER_172_855 ();
 FILLER_ASAP7_75t_R FILLER_172_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_863 ();
 DECAPx1_ASAP7_75t_R FILLER_172_884 ();
 DECAPx1_ASAP7_75t_R FILLER_172_930 ();
 DECAPx2_ASAP7_75t_R FILLER_172_948 ();
 FILLER_ASAP7_75t_R FILLER_172_954 ();
 FILLER_ASAP7_75t_R FILLER_172_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_970 ();
 DECAPx6_ASAP7_75t_R FILLER_172_997 ();
 FILLER_ASAP7_75t_R FILLER_172_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1051 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1073 ();
 FILLER_ASAP7_75t_R FILLER_172_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1215 ();
 FILLER_ASAP7_75t_R FILLER_172_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_173_2 ();
 DECAPx10_ASAP7_75t_R FILLER_173_24 ();
 DECAPx10_ASAP7_75t_R FILLER_173_46 ();
 DECAPx10_ASAP7_75t_R FILLER_173_68 ();
 DECAPx6_ASAP7_75t_R FILLER_173_90 ();
 DECAPx1_ASAP7_75t_R FILLER_173_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_108 ();
 FILLER_ASAP7_75t_R FILLER_173_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_128 ();
 DECAPx4_ASAP7_75t_R FILLER_173_151 ();
 FILLER_ASAP7_75t_R FILLER_173_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_172 ();
 DECAPx1_ASAP7_75t_R FILLER_173_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_190 ();
 FILLER_ASAP7_75t_R FILLER_173_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_215 ();
 DECAPx10_ASAP7_75t_R FILLER_173_223 ();
 DECAPx10_ASAP7_75t_R FILLER_173_245 ();
 DECAPx4_ASAP7_75t_R FILLER_173_267 ();
 FILLER_ASAP7_75t_R FILLER_173_277 ();
 DECAPx6_ASAP7_75t_R FILLER_173_285 ();
 DECAPx1_ASAP7_75t_R FILLER_173_299 ();
 DECAPx1_ASAP7_75t_R FILLER_173_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_342 ();
 DECAPx10_ASAP7_75t_R FILLER_173_346 ();
 DECAPx10_ASAP7_75t_R FILLER_173_368 ();
 DECAPx4_ASAP7_75t_R FILLER_173_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_400 ();
 DECAPx1_ASAP7_75t_R FILLER_173_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_431 ();
 DECAPx1_ASAP7_75t_R FILLER_173_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_487 ();
 DECAPx2_ASAP7_75t_R FILLER_173_491 ();
 DECAPx2_ASAP7_75t_R FILLER_173_524 ();
 FILLER_ASAP7_75t_R FILLER_173_530 ();
 DECAPx4_ASAP7_75t_R FILLER_173_538 ();
 FILLER_ASAP7_75t_R FILLER_173_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_550 ();
 DECAPx1_ASAP7_75t_R FILLER_173_571 ();
 DECAPx10_ASAP7_75t_R FILLER_173_629 ();
 DECAPx6_ASAP7_75t_R FILLER_173_651 ();
 DECAPx1_ASAP7_75t_R FILLER_173_665 ();
 DECAPx2_ASAP7_75t_R FILLER_173_679 ();
 FILLER_ASAP7_75t_R FILLER_173_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_687 ();
 DECAPx2_ASAP7_75t_R FILLER_173_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_710 ();
 DECAPx2_ASAP7_75t_R FILLER_173_733 ();
 FILLER_ASAP7_75t_R FILLER_173_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_741 ();
 DECAPx6_ASAP7_75t_R FILLER_173_767 ();
 FILLER_ASAP7_75t_R FILLER_173_781 ();
 FILLER_ASAP7_75t_R FILLER_173_805 ();
 DECAPx2_ASAP7_75t_R FILLER_173_826 ();
 DECAPx2_ASAP7_75t_R FILLER_173_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_864 ();
 DECAPx6_ASAP7_75t_R FILLER_173_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_923 ();
 DECAPx2_ASAP7_75t_R FILLER_173_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_932 ();
 DECAPx2_ASAP7_75t_R FILLER_173_940 ();
 FILLER_ASAP7_75t_R FILLER_173_946 ();
 DECAPx1_ASAP7_75t_R FILLER_173_955 ();
 FILLER_ASAP7_75t_R FILLER_173_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_968 ();
 FILLER_ASAP7_75t_R FILLER_173_975 ();
 DECAPx10_ASAP7_75t_R FILLER_173_991 ();
 DECAPx6_ASAP7_75t_R FILLER_173_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1033 ();
 DECAPx6_ASAP7_75t_R FILLER_173_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_173_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1147 ();
 DECAPx4_ASAP7_75t_R FILLER_173_1199 ();
 FILLER_ASAP7_75t_R FILLER_173_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1214 ();
 DECAPx1_ASAP7_75t_R FILLER_173_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_174_2 ();
 DECAPx10_ASAP7_75t_R FILLER_174_24 ();
 DECAPx10_ASAP7_75t_R FILLER_174_46 ();
 DECAPx10_ASAP7_75t_R FILLER_174_68 ();
 DECAPx2_ASAP7_75t_R FILLER_174_90 ();
 FILLER_ASAP7_75t_R FILLER_174_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_98 ();
 DECAPx1_ASAP7_75t_R FILLER_174_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_125 ();
 DECAPx4_ASAP7_75t_R FILLER_174_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_145 ();
 DECAPx6_ASAP7_75t_R FILLER_174_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_223 ();
 DECAPx10_ASAP7_75t_R FILLER_174_258 ();
 DECAPx10_ASAP7_75t_R FILLER_174_280 ();
 DECAPx4_ASAP7_75t_R FILLER_174_302 ();
 DECAPx10_ASAP7_75t_R FILLER_174_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_337 ();
 DECAPx10_ASAP7_75t_R FILLER_174_382 ();
 FILLER_ASAP7_75t_R FILLER_174_404 ();
 DECAPx2_ASAP7_75t_R FILLER_174_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_479 ();
 DECAPx1_ASAP7_75t_R FILLER_174_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_490 ();
 DECAPx6_ASAP7_75t_R FILLER_174_512 ();
 FILLER_ASAP7_75t_R FILLER_174_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_528 ();
 FILLER_ASAP7_75t_R FILLER_174_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_551 ();
 DECAPx6_ASAP7_75t_R FILLER_174_558 ();
 FILLER_ASAP7_75t_R FILLER_174_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_574 ();
 DECAPx2_ASAP7_75t_R FILLER_174_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_589 ();
 DECAPx10_ASAP7_75t_R FILLER_174_618 ();
 FILLER_ASAP7_75t_R FILLER_174_640 ();
 DECAPx2_ASAP7_75t_R FILLER_174_672 ();
 FILLER_ASAP7_75t_R FILLER_174_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_680 ();
 FILLER_ASAP7_75t_R FILLER_174_689 ();
 DECAPx10_ASAP7_75t_R FILLER_174_714 ();
 DECAPx10_ASAP7_75t_R FILLER_174_736 ();
 DECAPx6_ASAP7_75t_R FILLER_174_765 ();
 DECAPx2_ASAP7_75t_R FILLER_174_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_799 ();
 FILLER_ASAP7_75t_R FILLER_174_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_821 ();
 FILLER_ASAP7_75t_R FILLER_174_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_842 ();
 DECAPx10_ASAP7_75t_R FILLER_174_862 ();
 DECAPx6_ASAP7_75t_R FILLER_174_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_908 ();
 FILLER_ASAP7_75t_R FILLER_174_931 ();
 DECAPx1_ASAP7_75t_R FILLER_174_943 ();
 FILLER_ASAP7_75t_R FILLER_174_960 ();
 DECAPx10_ASAP7_75t_R FILLER_174_972 ();
 DECAPx6_ASAP7_75t_R FILLER_174_994 ();
 FILLER_ASAP7_75t_R FILLER_174_1008 ();
 FILLER_ASAP7_75t_R FILLER_174_1034 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1072 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1096 ();
 FILLER_ASAP7_75t_R FILLER_174_1122 ();
 DECAPx4_ASAP7_75t_R FILLER_174_1130 ();
 FILLER_ASAP7_75t_R FILLER_174_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1187 ();
 FILLER_ASAP7_75t_R FILLER_174_1211 ();
 FILLER_ASAP7_75t_R FILLER_174_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_175_2 ();
 DECAPx10_ASAP7_75t_R FILLER_175_24 ();
 DECAPx10_ASAP7_75t_R FILLER_175_46 ();
 DECAPx10_ASAP7_75t_R FILLER_175_68 ();
 DECAPx10_ASAP7_75t_R FILLER_175_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_112 ();
 DECAPx1_ASAP7_75t_R FILLER_175_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_123 ();
 DECAPx10_ASAP7_75t_R FILLER_175_131 ();
 DECAPx4_ASAP7_75t_R FILLER_175_176 ();
 DECAPx6_ASAP7_75t_R FILLER_175_208 ();
 FILLER_ASAP7_75t_R FILLER_175_222 ();
 DECAPx10_ASAP7_75t_R FILLER_175_232 ();
 DECAPx2_ASAP7_75t_R FILLER_175_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_260 ();
 FILLER_ASAP7_75t_R FILLER_175_309 ();
 DECAPx10_ASAP7_75t_R FILLER_175_314 ();
 DECAPx4_ASAP7_75t_R FILLER_175_336 ();
 FILLER_ASAP7_75t_R FILLER_175_346 ();
 DECAPx4_ASAP7_75t_R FILLER_175_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_406 ();
 DECAPx6_ASAP7_75t_R FILLER_175_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_427 ();
 FILLER_ASAP7_75t_R FILLER_175_434 ();
 DECAPx1_ASAP7_75t_R FILLER_175_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_466 ();
 DECAPx1_ASAP7_75t_R FILLER_175_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_509 ();
 DECAPx10_ASAP7_75t_R FILLER_175_516 ();
 DECAPx2_ASAP7_75t_R FILLER_175_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_544 ();
 DECAPx1_ASAP7_75t_R FILLER_175_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_555 ();
 DECAPx6_ASAP7_75t_R FILLER_175_567 ();
 FILLER_ASAP7_75t_R FILLER_175_581 ();
 DECAPx1_ASAP7_75t_R FILLER_175_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_599 ();
 DECAPx10_ASAP7_75t_R FILLER_175_622 ();
 FILLER_ASAP7_75t_R FILLER_175_644 ();
 DECAPx10_ASAP7_75t_R FILLER_175_673 ();
 DECAPx4_ASAP7_75t_R FILLER_175_695 ();
 DECAPx4_ASAP7_75t_R FILLER_175_718 ();
 FILLER_ASAP7_75t_R FILLER_175_728 ();
 DECAPx10_ASAP7_75t_R FILLER_175_752 ();
 DECAPx10_ASAP7_75t_R FILLER_175_778 ();
 DECAPx1_ASAP7_75t_R FILLER_175_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_811 ();
 FILLER_ASAP7_75t_R FILLER_175_818 ();
 DECAPx2_ASAP7_75t_R FILLER_175_839 ();
 FILLER_ASAP7_75t_R FILLER_175_845 ();
 DECAPx2_ASAP7_75t_R FILLER_175_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_860 ();
 DECAPx6_ASAP7_75t_R FILLER_175_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_895 ();
 DECAPx6_ASAP7_75t_R FILLER_175_904 ();
 DECAPx2_ASAP7_75t_R FILLER_175_918 ();
 DECAPx1_ASAP7_75t_R FILLER_175_926 ();
 DECAPx2_ASAP7_75t_R FILLER_175_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_962 ();
 FILLER_ASAP7_75t_R FILLER_175_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1058 ();
 FILLER_ASAP7_75t_R FILLER_175_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1074 ();
 FILLER_ASAP7_75t_R FILLER_175_1097 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1105 ();
 FILLER_ASAP7_75t_R FILLER_175_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1193 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1218 ();
 FILLER_ASAP7_75t_R FILLER_175_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_176_2 ();
 DECAPx10_ASAP7_75t_R FILLER_176_24 ();
 DECAPx10_ASAP7_75t_R FILLER_176_46 ();
 DECAPx10_ASAP7_75t_R FILLER_176_68 ();
 DECAPx10_ASAP7_75t_R FILLER_176_90 ();
 DECAPx2_ASAP7_75t_R FILLER_176_112 ();
 FILLER_ASAP7_75t_R FILLER_176_118 ();
 DECAPx2_ASAP7_75t_R FILLER_176_138 ();
 FILLER_ASAP7_75t_R FILLER_176_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_146 ();
 DECAPx1_ASAP7_75t_R FILLER_176_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_163 ();
 DECAPx6_ASAP7_75t_R FILLER_176_186 ();
 DECAPx10_ASAP7_75t_R FILLER_176_223 ();
 DECAPx10_ASAP7_75t_R FILLER_176_245 ();
 DECAPx2_ASAP7_75t_R FILLER_176_267 ();
 FILLER_ASAP7_75t_R FILLER_176_273 ();
 DECAPx1_ASAP7_75t_R FILLER_176_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_308 ();
 DECAPx10_ASAP7_75t_R FILLER_176_329 ();
 DECAPx6_ASAP7_75t_R FILLER_176_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_365 ();
 DECAPx1_ASAP7_75t_R FILLER_176_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_374 ();
 DECAPx6_ASAP7_75t_R FILLER_176_379 ();
 DECAPx2_ASAP7_75t_R FILLER_176_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_406 ();
 FILLER_ASAP7_75t_R FILLER_176_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_429 ();
 DECAPx2_ASAP7_75t_R FILLER_176_450 ();
 FILLER_ASAP7_75t_R FILLER_176_464 ();
 DECAPx2_ASAP7_75t_R FILLER_176_478 ();
 FILLER_ASAP7_75t_R FILLER_176_484 ();
 FILLER_ASAP7_75t_R FILLER_176_508 ();
 DECAPx4_ASAP7_75t_R FILLER_176_533 ();
 FILLER_ASAP7_75t_R FILLER_176_543 ();
 DECAPx10_ASAP7_75t_R FILLER_176_613 ();
 FILLER_ASAP7_75t_R FILLER_176_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_637 ();
 FILLER_ASAP7_75t_R FILLER_176_645 ();
 DECAPx1_ASAP7_75t_R FILLER_176_654 ();
 DECAPx4_ASAP7_75t_R FILLER_176_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_692 ();
 DECAPx2_ASAP7_75t_R FILLER_176_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_702 ();
 FILLER_ASAP7_75t_R FILLER_176_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_718 ();
 DECAPx4_ASAP7_75t_R FILLER_176_741 ();
 FILLER_ASAP7_75t_R FILLER_176_751 ();
 DECAPx2_ASAP7_75t_R FILLER_176_797 ();
 FILLER_ASAP7_75t_R FILLER_176_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_805 ();
 DECAPx6_ASAP7_75t_R FILLER_176_820 ();
 DECAPx2_ASAP7_75t_R FILLER_176_834 ();
 DECAPx1_ASAP7_75t_R FILLER_176_880 ();
 DECAPx6_ASAP7_75t_R FILLER_176_887 ();
 DECAPx2_ASAP7_75t_R FILLER_176_921 ();
 FILLER_ASAP7_75t_R FILLER_176_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_929 ();
 DECAPx6_ASAP7_75t_R FILLER_176_933 ();
 FILLER_ASAP7_75t_R FILLER_176_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_949 ();
 DECAPx2_ASAP7_75t_R FILLER_176_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_965 ();
 DECAPx10_ASAP7_75t_R FILLER_176_975 ();
 FILLER_ASAP7_75t_R FILLER_176_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1034 ();
 DECAPx6_ASAP7_75t_R FILLER_176_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1052 ();
 DECAPx4_ASAP7_75t_R FILLER_176_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1187 ();
 DECAPx4_ASAP7_75t_R FILLER_176_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_177_2 ();
 DECAPx10_ASAP7_75t_R FILLER_177_24 ();
 DECAPx10_ASAP7_75t_R FILLER_177_46 ();
 DECAPx10_ASAP7_75t_R FILLER_177_68 ();
 DECAPx6_ASAP7_75t_R FILLER_177_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_104 ();
 DECAPx4_ASAP7_75t_R FILLER_177_133 ();
 FILLER_ASAP7_75t_R FILLER_177_143 ();
 DECAPx2_ASAP7_75t_R FILLER_177_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_157 ();
 DECAPx10_ASAP7_75t_R FILLER_177_164 ();
 DECAPx10_ASAP7_75t_R FILLER_177_186 ();
 DECAPx2_ASAP7_75t_R FILLER_177_208 ();
 FILLER_ASAP7_75t_R FILLER_177_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_216 ();
 DECAPx6_ASAP7_75t_R FILLER_177_243 ();
 FILLER_ASAP7_75t_R FILLER_177_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_263 ();
 DECAPx4_ASAP7_75t_R FILLER_177_290 ();
 FILLER_ASAP7_75t_R FILLER_177_300 ();
 DECAPx2_ASAP7_75t_R FILLER_177_322 ();
 FILLER_ASAP7_75t_R FILLER_177_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_334 ();
 DECAPx4_ASAP7_75t_R FILLER_177_355 ();
 DECAPx4_ASAP7_75t_R FILLER_177_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_423 ();
 DECAPx2_ASAP7_75t_R FILLER_177_453 ();
 FILLER_ASAP7_75t_R FILLER_177_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_474 ();
 DECAPx2_ASAP7_75t_R FILLER_177_481 ();
 FILLER_ASAP7_75t_R FILLER_177_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_496 ();
 FILLER_ASAP7_75t_R FILLER_177_516 ();
 DECAPx1_ASAP7_75t_R FILLER_177_524 ();
 DECAPx10_ASAP7_75t_R FILLER_177_531 ();
 DECAPx10_ASAP7_75t_R FILLER_177_553 ();
 FILLER_ASAP7_75t_R FILLER_177_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_577 ();
 DECAPx4_ASAP7_75t_R FILLER_177_584 ();
 DECAPx10_ASAP7_75t_R FILLER_177_606 ();
 DECAPx4_ASAP7_75t_R FILLER_177_628 ();
 FILLER_ASAP7_75t_R FILLER_177_638 ();
 DECAPx6_ASAP7_75t_R FILLER_177_656 ();
 FILLER_ASAP7_75t_R FILLER_177_670 ();
 DECAPx1_ASAP7_75t_R FILLER_177_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_692 ();
 DECAPx6_ASAP7_75t_R FILLER_177_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_717 ();
 DECAPx4_ASAP7_75t_R FILLER_177_725 ();
 FILLER_ASAP7_75t_R FILLER_177_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_758 ();
 DECAPx2_ASAP7_75t_R FILLER_177_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_787 ();
 DECAPx10_ASAP7_75t_R FILLER_177_810 ();
 DECAPx10_ASAP7_75t_R FILLER_177_832 ();
 DECAPx6_ASAP7_75t_R FILLER_177_854 ();
 DECAPx2_ASAP7_75t_R FILLER_177_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_874 ();
 DECAPx2_ASAP7_75t_R FILLER_177_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_926 ();
 FILLER_ASAP7_75t_R FILLER_177_947 ();
 DECAPx1_ASAP7_75t_R FILLER_177_963 ();
 DECAPx2_ASAP7_75t_R FILLER_177_981 ();
 FILLER_ASAP7_75t_R FILLER_177_987 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_178_2 ();
 DECAPx10_ASAP7_75t_R FILLER_178_24 ();
 DECAPx10_ASAP7_75t_R FILLER_178_46 ();
 DECAPx10_ASAP7_75t_R FILLER_178_68 ();
 DECAPx10_ASAP7_75t_R FILLER_178_90 ();
 DECAPx1_ASAP7_75t_R FILLER_178_112 ();
 DECAPx2_ASAP7_75t_R FILLER_178_127 ();
 FILLER_ASAP7_75t_R FILLER_178_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_135 ();
 FILLER_ASAP7_75t_R FILLER_178_148 ();
 DECAPx6_ASAP7_75t_R FILLER_178_163 ();
 FILLER_ASAP7_75t_R FILLER_178_177 ();
 FILLER_ASAP7_75t_R FILLER_178_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_189 ();
 FILLER_ASAP7_75t_R FILLER_178_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_212 ();
 DECAPx10_ASAP7_75t_R FILLER_178_233 ();
 DECAPx2_ASAP7_75t_R FILLER_178_255 ();
 FILLER_ASAP7_75t_R FILLER_178_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_263 ();
 DECAPx10_ASAP7_75t_R FILLER_178_294 ();
 DECAPx10_ASAP7_75t_R FILLER_178_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_358 ();
 FILLER_ASAP7_75t_R FILLER_178_363 ();
 DECAPx4_ASAP7_75t_R FILLER_178_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_381 ();
 DECAPx6_ASAP7_75t_R FILLER_178_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_402 ();
 DECAPx1_ASAP7_75t_R FILLER_178_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_413 ();
 DECAPx6_ASAP7_75t_R FILLER_178_426 ();
 FILLER_ASAP7_75t_R FILLER_178_440 ();
 FILLER_ASAP7_75t_R FILLER_178_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_466 ();
 DECAPx4_ASAP7_75t_R FILLER_178_479 ();
 FILLER_ASAP7_75t_R FILLER_178_489 ();
 FILLER_ASAP7_75t_R FILLER_178_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_516 ();
 FILLER_ASAP7_75t_R FILLER_178_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_525 ();
 DECAPx10_ASAP7_75t_R FILLER_178_532 ();
 DECAPx10_ASAP7_75t_R FILLER_178_554 ();
 DECAPx2_ASAP7_75t_R FILLER_178_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_590 ();
 DECAPx10_ASAP7_75t_R FILLER_178_603 ();
 DECAPx2_ASAP7_75t_R FILLER_178_625 ();
 FILLER_ASAP7_75t_R FILLER_178_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_645 ();
 FILLER_ASAP7_75t_R FILLER_178_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_669 ();
 DECAPx2_ASAP7_75t_R FILLER_178_685 ();
 DECAPx6_ASAP7_75t_R FILLER_178_701 ();
 DECAPx1_ASAP7_75t_R FILLER_178_715 ();
 FILLER_ASAP7_75t_R FILLER_178_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_735 ();
 DECAPx2_ASAP7_75t_R FILLER_178_743 ();
 FILLER_ASAP7_75t_R FILLER_178_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_751 ();
 DECAPx6_ASAP7_75t_R FILLER_178_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_773 ();
 DECAPx10_ASAP7_75t_R FILLER_178_796 ();
 DECAPx10_ASAP7_75t_R FILLER_178_818 ();
 DECAPx2_ASAP7_75t_R FILLER_178_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_846 ();
 DECAPx6_ASAP7_75t_R FILLER_178_851 ();
 FILLER_ASAP7_75t_R FILLER_178_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_887 ();
 DECAPx10_ASAP7_75t_R FILLER_178_896 ();
 DECAPx10_ASAP7_75t_R FILLER_178_918 ();
 DECAPx4_ASAP7_75t_R FILLER_178_940 ();
 FILLER_ASAP7_75t_R FILLER_178_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_952 ();
 DECAPx4_ASAP7_75t_R FILLER_178_959 ();
 FILLER_ASAP7_75t_R FILLER_178_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_971 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1000 ();
 DECAPx1_ASAP7_75t_R FILLER_178_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1040 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1105 ();
 FILLER_ASAP7_75t_R FILLER_178_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_179_2 ();
 DECAPx10_ASAP7_75t_R FILLER_179_24 ();
 DECAPx10_ASAP7_75t_R FILLER_179_46 ();
 DECAPx10_ASAP7_75t_R FILLER_179_68 ();
 DECAPx6_ASAP7_75t_R FILLER_179_90 ();
 DECAPx1_ASAP7_75t_R FILLER_179_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_108 ();
 DECAPx2_ASAP7_75t_R FILLER_179_131 ();
 FILLER_ASAP7_75t_R FILLER_179_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_139 ();
 FILLER_ASAP7_75t_R FILLER_179_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_150 ();
 FILLER_ASAP7_75t_R FILLER_179_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_182 ();
 FILLER_ASAP7_75t_R FILLER_179_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_214 ();
 FILLER_ASAP7_75t_R FILLER_179_224 ();
 DECAPx4_ASAP7_75t_R FILLER_179_243 ();
 FILLER_ASAP7_75t_R FILLER_179_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_255 ();
 DECAPx1_ASAP7_75t_R FILLER_179_300 ();
 DECAPx10_ASAP7_75t_R FILLER_179_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_332 ();
 DECAPx4_ASAP7_75t_R FILLER_179_339 ();
 FILLER_ASAP7_75t_R FILLER_179_367 ();
 DECAPx6_ASAP7_75t_R FILLER_179_391 ();
 DECAPx2_ASAP7_75t_R FILLER_179_405 ();
 FILLER_ASAP7_75t_R FILLER_179_417 ();
 FILLER_ASAP7_75t_R FILLER_179_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_427 ();
 DECAPx1_ASAP7_75t_R FILLER_179_448 ();
 DECAPx2_ASAP7_75t_R FILLER_179_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_468 ();
 DECAPx6_ASAP7_75t_R FILLER_179_475 ();
 FILLER_ASAP7_75t_R FILLER_179_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_503 ();
 DECAPx10_ASAP7_75t_R FILLER_179_510 ();
 FILLER_ASAP7_75t_R FILLER_179_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_534 ();
 DECAPx1_ASAP7_75t_R FILLER_179_555 ();
 DECAPx4_ASAP7_75t_R FILLER_179_563 ();
 FILLER_ASAP7_75t_R FILLER_179_573 ();
 DECAPx1_ASAP7_75t_R FILLER_179_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_591 ();
 DECAPx10_ASAP7_75t_R FILLER_179_599 ();
 FILLER_ASAP7_75t_R FILLER_179_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_651 ();
 FILLER_ASAP7_75t_R FILLER_179_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_662 ();
 FILLER_ASAP7_75t_R FILLER_179_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_672 ();
 FILLER_ASAP7_75t_R FILLER_179_680 ();
 FILLER_ASAP7_75t_R FILLER_179_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_691 ();
 DECAPx1_ASAP7_75t_R FILLER_179_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_758 ();
 DECAPx4_ASAP7_75t_R FILLER_179_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_791 ();
 FILLER_ASAP7_75t_R FILLER_179_895 ();
 FILLER_ASAP7_75t_R FILLER_179_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_905 ();
 FILLER_ASAP7_75t_R FILLER_179_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_923 ();
 DECAPx6_ASAP7_75t_R FILLER_179_926 ();
 DECAPx6_ASAP7_75t_R FILLER_179_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_974 ();
 DECAPx2_ASAP7_75t_R FILLER_179_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1129 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1151 ();
 FILLER_ASAP7_75t_R FILLER_179_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1182 ();
 DECAPx6_ASAP7_75t_R FILLER_179_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_180_2 ();
 DECAPx10_ASAP7_75t_R FILLER_180_24 ();
 DECAPx10_ASAP7_75t_R FILLER_180_46 ();
 DECAPx10_ASAP7_75t_R FILLER_180_68 ();
 DECAPx10_ASAP7_75t_R FILLER_180_90 ();
 DECAPx2_ASAP7_75t_R FILLER_180_112 ();
 DECAPx4_ASAP7_75t_R FILLER_180_124 ();
 DECAPx6_ASAP7_75t_R FILLER_180_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_170 ();
 DECAPx6_ASAP7_75t_R FILLER_180_188 ();
 DECAPx4_ASAP7_75t_R FILLER_180_258 ();
 FILLER_ASAP7_75t_R FILLER_180_268 ();
 FILLER_ASAP7_75t_R FILLER_180_276 ();
 DECAPx10_ASAP7_75t_R FILLER_180_281 ();
 DECAPx2_ASAP7_75t_R FILLER_180_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_331 ();
 DECAPx1_ASAP7_75t_R FILLER_180_354 ();
 DECAPx6_ASAP7_75t_R FILLER_180_375 ();
 FILLER_ASAP7_75t_R FILLER_180_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_391 ();
 DECAPx2_ASAP7_75t_R FILLER_180_412 ();
 FILLER_ASAP7_75t_R FILLER_180_418 ();
 DECAPx1_ASAP7_75t_R FILLER_180_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_468 ();
 DECAPx1_ASAP7_75t_R FILLER_180_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_476 ();
 DECAPx2_ASAP7_75t_R FILLER_180_481 ();
 FILLER_ASAP7_75t_R FILLER_180_487 ();
 DECAPx10_ASAP7_75t_R FILLER_180_499 ();
 DECAPx2_ASAP7_75t_R FILLER_180_521 ();
 FILLER_ASAP7_75t_R FILLER_180_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_529 ();
 DECAPx4_ASAP7_75t_R FILLER_180_554 ();
 FILLER_ASAP7_75t_R FILLER_180_600 ();
 DECAPx6_ASAP7_75t_R FILLER_180_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_638 ();
 FILLER_ASAP7_75t_R FILLER_180_658 ();
 FILLER_ASAP7_75t_R FILLER_180_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_704 ();
 DECAPx6_ASAP7_75t_R FILLER_180_733 ();
 FILLER_ASAP7_75t_R FILLER_180_747 ();
 DECAPx6_ASAP7_75t_R FILLER_180_755 ();
 DECAPx1_ASAP7_75t_R FILLER_180_769 ();
 DECAPx10_ASAP7_75t_R FILLER_180_795 ();
 DECAPx10_ASAP7_75t_R FILLER_180_817 ();
 DECAPx10_ASAP7_75t_R FILLER_180_839 ();
 DECAPx2_ASAP7_75t_R FILLER_180_861 ();
 FILLER_ASAP7_75t_R FILLER_180_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_869 ();
 FILLER_ASAP7_75t_R FILLER_180_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_894 ();
 DECAPx1_ASAP7_75t_R FILLER_180_940 ();
 DECAPx4_ASAP7_75t_R FILLER_180_948 ();
 DECAPx6_ASAP7_75t_R FILLER_180_980 ();
 FILLER_ASAP7_75t_R FILLER_180_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_996 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1010 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1059 ();
 FILLER_ASAP7_75t_R FILLER_180_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1204 ();
 DECAPx6_ASAP7_75t_R FILLER_180_1208 ();
 FILLER_ASAP7_75t_R FILLER_180_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_181_2 ();
 DECAPx10_ASAP7_75t_R FILLER_181_24 ();
 DECAPx10_ASAP7_75t_R FILLER_181_46 ();
 DECAPx10_ASAP7_75t_R FILLER_181_68 ();
 DECAPx10_ASAP7_75t_R FILLER_181_90 ();
 DECAPx10_ASAP7_75t_R FILLER_181_112 ();
 DECAPx2_ASAP7_75t_R FILLER_181_134 ();
 FILLER_ASAP7_75t_R FILLER_181_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_142 ();
 DECAPx2_ASAP7_75t_R FILLER_181_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_166 ();
 DECAPx10_ASAP7_75t_R FILLER_181_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_209 ();
 DECAPx10_ASAP7_75t_R FILLER_181_232 ();
 DECAPx10_ASAP7_75t_R FILLER_181_254 ();
 DECAPx10_ASAP7_75t_R FILLER_181_276 ();
 DECAPx1_ASAP7_75t_R FILLER_181_298 ();
 DECAPx1_ASAP7_75t_R FILLER_181_322 ();
 DECAPx10_ASAP7_75t_R FILLER_181_337 ();
 FILLER_ASAP7_75t_R FILLER_181_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_361 ();
 DECAPx1_ASAP7_75t_R FILLER_181_368 ();
 DECAPx1_ASAP7_75t_R FILLER_181_406 ();
 DECAPx10_ASAP7_75t_R FILLER_181_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_438 ();
 DECAPx6_ASAP7_75t_R FILLER_181_445 ();
 FILLER_ASAP7_75t_R FILLER_181_459 ();
 DECAPx6_ASAP7_75t_R FILLER_181_512 ();
 DECAPx2_ASAP7_75t_R FILLER_181_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_532 ();
 DECAPx4_ASAP7_75t_R FILLER_181_557 ();
 FILLER_ASAP7_75t_R FILLER_181_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_575 ();
 DECAPx1_ASAP7_75t_R FILLER_181_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_591 ();
 DECAPx10_ASAP7_75t_R FILLER_181_609 ();
 DECAPx4_ASAP7_75t_R FILLER_181_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_641 ();
 DECAPx1_ASAP7_75t_R FILLER_181_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_668 ();
 DECAPx1_ASAP7_75t_R FILLER_181_686 ();
 DECAPx2_ASAP7_75t_R FILLER_181_703 ();
 FILLER_ASAP7_75t_R FILLER_181_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_711 ();
 DECAPx6_ASAP7_75t_R FILLER_181_718 ();
 DECAPx2_ASAP7_75t_R FILLER_181_740 ();
 FILLER_ASAP7_75t_R FILLER_181_746 ();
 DECAPx1_ASAP7_75t_R FILLER_181_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_765 ();
 DECAPx6_ASAP7_75t_R FILLER_181_779 ();
 DECAPx2_ASAP7_75t_R FILLER_181_837 ();
 FILLER_ASAP7_75t_R FILLER_181_843 ();
 FILLER_ASAP7_75t_R FILLER_181_867 ();
 DECAPx6_ASAP7_75t_R FILLER_181_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_886 ();
 DECAPx2_ASAP7_75t_R FILLER_181_894 ();
 FILLER_ASAP7_75t_R FILLER_181_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_902 ();
 DECAPx2_ASAP7_75t_R FILLER_181_915 ();
 FILLER_ASAP7_75t_R FILLER_181_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_923 ();
 DECAPx4_ASAP7_75t_R FILLER_181_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_936 ();
 DECAPx6_ASAP7_75t_R FILLER_181_967 ();
 DECAPx1_ASAP7_75t_R FILLER_181_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_985 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1008 ();
 FILLER_ASAP7_75t_R FILLER_181_1030 ();
 FILLER_ASAP7_75t_R FILLER_181_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1070 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1079 ();
 FILLER_ASAP7_75t_R FILLER_181_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1095 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1130 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1154 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1187 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1198 ();
 FILLER_ASAP7_75t_R FILLER_181_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_181_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_182_2 ();
 DECAPx10_ASAP7_75t_R FILLER_182_24 ();
 DECAPx10_ASAP7_75t_R FILLER_182_46 ();
 DECAPx10_ASAP7_75t_R FILLER_182_68 ();
 DECAPx10_ASAP7_75t_R FILLER_182_90 ();
 DECAPx6_ASAP7_75t_R FILLER_182_112 ();
 FILLER_ASAP7_75t_R FILLER_182_126 ();
 DECAPx6_ASAP7_75t_R FILLER_182_139 ();
 DECAPx1_ASAP7_75t_R FILLER_182_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_157 ();
 DECAPx6_ASAP7_75t_R FILLER_182_180 ();
 DECAPx1_ASAP7_75t_R FILLER_182_194 ();
 DECAPx10_ASAP7_75t_R FILLER_182_237 ();
 DECAPx10_ASAP7_75t_R FILLER_182_259 ();
 DECAPx6_ASAP7_75t_R FILLER_182_281 ();
 DECAPx2_ASAP7_75t_R FILLER_182_295 ();
 DECAPx10_ASAP7_75t_R FILLER_182_313 ();
 DECAPx10_ASAP7_75t_R FILLER_182_335 ();
 DECAPx4_ASAP7_75t_R FILLER_182_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_373 ();
 DECAPx10_ASAP7_75t_R FILLER_182_382 ();
 DECAPx2_ASAP7_75t_R FILLER_182_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_410 ();
 DECAPx2_ASAP7_75t_R FILLER_182_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_439 ();
 DECAPx4_ASAP7_75t_R FILLER_182_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_474 ();
 DECAPx2_ASAP7_75t_R FILLER_182_498 ();
 DECAPx1_ASAP7_75t_R FILLER_182_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_538 ();
 FILLER_ASAP7_75t_R FILLER_182_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_551 ();
 FILLER_ASAP7_75t_R FILLER_182_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_601 ();
 DECAPx10_ASAP7_75t_R FILLER_182_608 ();
 DECAPx6_ASAP7_75t_R FILLER_182_630 ();
 FILLER_ASAP7_75t_R FILLER_182_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_646 ();
 FILLER_ASAP7_75t_R FILLER_182_652 ();
 DECAPx6_ASAP7_75t_R FILLER_182_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_676 ();
 DECAPx1_ASAP7_75t_R FILLER_182_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_689 ();
 DECAPx6_ASAP7_75t_R FILLER_182_710 ();
 FILLER_ASAP7_75t_R FILLER_182_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_736 ();
 DECAPx6_ASAP7_75t_R FILLER_182_743 ();
 DECAPx1_ASAP7_75t_R FILLER_182_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_761 ();
 DECAPx4_ASAP7_75t_R FILLER_182_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_785 ();
 DECAPx6_ASAP7_75t_R FILLER_182_830 ();
 DECAPx1_ASAP7_75t_R FILLER_182_844 ();
 DECAPx6_ASAP7_75t_R FILLER_182_854 ();
 DECAPx2_ASAP7_75t_R FILLER_182_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_874 ();
 DECAPx6_ASAP7_75t_R FILLER_182_886 ();
 DECAPx2_ASAP7_75t_R FILLER_182_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_906 ();
 FILLER_ASAP7_75t_R FILLER_182_914 ();
 DECAPx10_ASAP7_75t_R FILLER_182_936 ();
 FILLER_ASAP7_75t_R FILLER_182_958 ();
 DECAPx10_ASAP7_75t_R FILLER_182_982 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1083 ();
 FILLER_ASAP7_75t_R FILLER_182_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1184 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1206 ();
 FILLER_ASAP7_75t_R FILLER_182_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_183_2 ();
 DECAPx10_ASAP7_75t_R FILLER_183_24 ();
 DECAPx10_ASAP7_75t_R FILLER_183_46 ();
 DECAPx10_ASAP7_75t_R FILLER_183_68 ();
 DECAPx10_ASAP7_75t_R FILLER_183_90 ();
 DECAPx6_ASAP7_75t_R FILLER_183_112 ();
 DECAPx2_ASAP7_75t_R FILLER_183_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_132 ();
 FILLER_ASAP7_75t_R FILLER_183_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_157 ();
 DECAPx10_ASAP7_75t_R FILLER_183_164 ();
 FILLER_ASAP7_75t_R FILLER_183_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_188 ();
 DECAPx10_ASAP7_75t_R FILLER_183_233 ();
 DECAPx10_ASAP7_75t_R FILLER_183_255 ();
 DECAPx4_ASAP7_75t_R FILLER_183_277 ();
 FILLER_ASAP7_75t_R FILLER_183_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_300 ();
 DECAPx10_ASAP7_75t_R FILLER_183_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_332 ();
 DECAPx1_ASAP7_75t_R FILLER_183_381 ();
 DECAPx10_ASAP7_75t_R FILLER_183_392 ();
 DECAPx1_ASAP7_75t_R FILLER_183_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_438 ();
 FILLER_ASAP7_75t_R FILLER_183_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_447 ();
 DECAPx1_ASAP7_75t_R FILLER_183_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_472 ();
 DECAPx10_ASAP7_75t_R FILLER_183_499 ();
 DECAPx1_ASAP7_75t_R FILLER_183_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_525 ();
 DECAPx1_ASAP7_75t_R FILLER_183_530 ();
 DECAPx6_ASAP7_75t_R FILLER_183_556 ();
 FILLER_ASAP7_75t_R FILLER_183_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_572 ();
 DECAPx2_ASAP7_75t_R FILLER_183_587 ();
 FILLER_ASAP7_75t_R FILLER_183_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_624 ();
 FILLER_ASAP7_75t_R FILLER_183_640 ();
 DECAPx1_ASAP7_75t_R FILLER_183_664 ();
 DECAPx2_ASAP7_75t_R FILLER_183_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_692 ();
 DECAPx2_ASAP7_75t_R FILLER_183_696 ();
 FILLER_ASAP7_75t_R FILLER_183_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_704 ();
 DECAPx6_ASAP7_75t_R FILLER_183_708 ();
 FILLER_ASAP7_75t_R FILLER_183_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_724 ();
 FILLER_ASAP7_75t_R FILLER_183_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_738 ();
 DECAPx6_ASAP7_75t_R FILLER_183_745 ();
 FILLER_ASAP7_75t_R FILLER_183_759 ();
 DECAPx2_ASAP7_75t_R FILLER_183_780 ();
 FILLER_ASAP7_75t_R FILLER_183_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_853 ();
 DECAPx1_ASAP7_75t_R FILLER_183_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_875 ();
 FILLER_ASAP7_75t_R FILLER_183_906 ();
 DECAPx1_ASAP7_75t_R FILLER_183_926 ();
 DECAPx4_ASAP7_75t_R FILLER_183_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_960 ();
 DECAPx10_ASAP7_75t_R FILLER_183_967 ();
 FILLER_ASAP7_75t_R FILLER_183_989 ();
 DECAPx4_ASAP7_75t_R FILLER_183_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1011 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_183_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1078 ();
 DECAPx4_ASAP7_75t_R FILLER_183_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1177 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_184_2 ();
 DECAPx10_ASAP7_75t_R FILLER_184_24 ();
 DECAPx10_ASAP7_75t_R FILLER_184_46 ();
 DECAPx10_ASAP7_75t_R FILLER_184_68 ();
 DECAPx10_ASAP7_75t_R FILLER_184_90 ();
 DECAPx10_ASAP7_75t_R FILLER_184_112 ();
 DECAPx10_ASAP7_75t_R FILLER_184_140 ();
 DECAPx10_ASAP7_75t_R FILLER_184_162 ();
 DECAPx6_ASAP7_75t_R FILLER_184_184 ();
 FILLER_ASAP7_75t_R FILLER_184_198 ();
 DECAPx2_ASAP7_75t_R FILLER_184_206 ();
 FILLER_ASAP7_75t_R FILLER_184_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_214 ();
 DECAPx10_ASAP7_75t_R FILLER_184_221 ();
 DECAPx10_ASAP7_75t_R FILLER_184_243 ();
 DECAPx6_ASAP7_75t_R FILLER_184_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_316 ();
 FILLER_ASAP7_75t_R FILLER_184_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_334 ();
 DECAPx2_ASAP7_75t_R FILLER_184_341 ();
 DECAPx1_ASAP7_75t_R FILLER_184_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_358 ();
 DECAPx1_ASAP7_75t_R FILLER_184_366 ();
 DECAPx6_ASAP7_75t_R FILLER_184_392 ();
 DECAPx1_ASAP7_75t_R FILLER_184_406 ();
 DECAPx1_ASAP7_75t_R FILLER_184_430 ();
 DECAPx10_ASAP7_75t_R FILLER_184_464 ();
 DECAPx10_ASAP7_75t_R FILLER_184_486 ();
 DECAPx1_ASAP7_75t_R FILLER_184_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_512 ();
 DECAPx2_ASAP7_75t_R FILLER_184_541 ();
 FILLER_ASAP7_75t_R FILLER_184_547 ();
 DECAPx2_ASAP7_75t_R FILLER_184_571 ();
 FILLER_ASAP7_75t_R FILLER_184_577 ();
 DECAPx10_ASAP7_75t_R FILLER_184_601 ();
 FILLER_ASAP7_75t_R FILLER_184_623 ();
 FILLER_ASAP7_75t_R FILLER_184_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_666 ();
 FILLER_ASAP7_75t_R FILLER_184_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_683 ();
 DECAPx2_ASAP7_75t_R FILLER_184_696 ();
 FILLER_ASAP7_75t_R FILLER_184_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_727 ();
 FILLER_ASAP7_75t_R FILLER_184_738 ();
 DECAPx2_ASAP7_75t_R FILLER_184_746 ();
 DECAPx1_ASAP7_75t_R FILLER_184_759 ();
 DECAPx4_ASAP7_75t_R FILLER_184_770 ();
 FILLER_ASAP7_75t_R FILLER_184_780 ();
 DECAPx10_ASAP7_75t_R FILLER_184_785 ();
 DECAPx10_ASAP7_75t_R FILLER_184_807 ();
 DECAPx10_ASAP7_75t_R FILLER_184_829 ();
 FILLER_ASAP7_75t_R FILLER_184_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_880 ();
 FILLER_ASAP7_75t_R FILLER_184_887 ();
 DECAPx6_ASAP7_75t_R FILLER_184_918 ();
 FILLER_ASAP7_75t_R FILLER_184_932 ();
 DECAPx6_ASAP7_75t_R FILLER_184_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_978 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1001 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1014 ();
 FILLER_ASAP7_75t_R FILLER_184_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1060 ();
 FILLER_ASAP7_75t_R FILLER_184_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1071 ();
 DECAPx4_ASAP7_75t_R FILLER_184_1078 ();
 DECAPx4_ASAP7_75t_R FILLER_184_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1166 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1188 ();
 FILLER_ASAP7_75t_R FILLER_184_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_185_2 ();
 DECAPx10_ASAP7_75t_R FILLER_185_24 ();
 DECAPx10_ASAP7_75t_R FILLER_185_46 ();
 DECAPx10_ASAP7_75t_R FILLER_185_68 ();
 DECAPx10_ASAP7_75t_R FILLER_185_90 ();
 DECAPx10_ASAP7_75t_R FILLER_185_112 ();
 DECAPx10_ASAP7_75t_R FILLER_185_134 ();
 DECAPx10_ASAP7_75t_R FILLER_185_156 ();
 DECAPx10_ASAP7_75t_R FILLER_185_178 ();
 DECAPx10_ASAP7_75t_R FILLER_185_200 ();
 DECAPx10_ASAP7_75t_R FILLER_185_222 ();
 DECAPx10_ASAP7_75t_R FILLER_185_244 ();
 DECAPx10_ASAP7_75t_R FILLER_185_266 ();
 FILLER_ASAP7_75t_R FILLER_185_288 ();
 DECAPx4_ASAP7_75t_R FILLER_185_296 ();
 DECAPx1_ASAP7_75t_R FILLER_185_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_342 ();
 FILLER_ASAP7_75t_R FILLER_185_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_366 ();
 DECAPx4_ASAP7_75t_R FILLER_185_379 ();
 FILLER_ASAP7_75t_R FILLER_185_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_413 ();
 FILLER_ASAP7_75t_R FILLER_185_434 ();
 DECAPx2_ASAP7_75t_R FILLER_185_469 ();
 FILLER_ASAP7_75t_R FILLER_185_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_480 ();
 FILLER_ASAP7_75t_R FILLER_185_484 ();
 DECAPx1_ASAP7_75t_R FILLER_185_506 ();
 DECAPx6_ASAP7_75t_R FILLER_185_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_550 ();
 FILLER_ASAP7_75t_R FILLER_185_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_559 ();
 DECAPx10_ASAP7_75t_R FILLER_185_571 ();
 DECAPx10_ASAP7_75t_R FILLER_185_593 ();
 DECAPx6_ASAP7_75t_R FILLER_185_615 ();
 DECAPx1_ASAP7_75t_R FILLER_185_629 ();
 DECAPx2_ASAP7_75t_R FILLER_185_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_649 ();
 DECAPx4_ASAP7_75t_R FILLER_185_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_697 ();
 DECAPx1_ASAP7_75t_R FILLER_185_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_708 ();
 DECAPx4_ASAP7_75t_R FILLER_185_716 ();
 DECAPx6_ASAP7_75t_R FILLER_185_755 ();
 DECAPx1_ASAP7_75t_R FILLER_185_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_773 ();
 DECAPx10_ASAP7_75t_R FILLER_185_808 ();
 DECAPx10_ASAP7_75t_R FILLER_185_830 ();
 DECAPx1_ASAP7_75t_R FILLER_185_858 ();
 DECAPx2_ASAP7_75t_R FILLER_185_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_888 ();
 FILLER_ASAP7_75t_R FILLER_185_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_899 ();
 FILLER_ASAP7_75t_R FILLER_185_908 ();
 DECAPx2_ASAP7_75t_R FILLER_185_916 ();
 FILLER_ASAP7_75t_R FILLER_185_922 ();
 DECAPx2_ASAP7_75t_R FILLER_185_932 ();
 FILLER_ASAP7_75t_R FILLER_185_938 ();
 DECAPx4_ASAP7_75t_R FILLER_185_962 ();
 FILLER_ASAP7_75t_R FILLER_185_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_974 ();
 DECAPx2_ASAP7_75t_R FILLER_185_988 ();
 FILLER_ASAP7_75t_R FILLER_185_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_996 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1020 ();
 FILLER_ASAP7_75t_R FILLER_185_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1077 ();
 FILLER_ASAP7_75t_R FILLER_185_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1085 ();
 DECAPx6_ASAP7_75t_R FILLER_185_1112 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1195 ();
 FILLER_ASAP7_75t_R FILLER_185_1212 ();
 FILLER_ASAP7_75t_R FILLER_185_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_186_2 ();
 DECAPx10_ASAP7_75t_R FILLER_186_24 ();
 DECAPx10_ASAP7_75t_R FILLER_186_46 ();
 DECAPx10_ASAP7_75t_R FILLER_186_68 ();
 DECAPx10_ASAP7_75t_R FILLER_186_90 ();
 DECAPx10_ASAP7_75t_R FILLER_186_112 ();
 DECAPx10_ASAP7_75t_R FILLER_186_134 ();
 DECAPx10_ASAP7_75t_R FILLER_186_156 ();
 DECAPx10_ASAP7_75t_R FILLER_186_178 ();
 DECAPx10_ASAP7_75t_R FILLER_186_200 ();
 DECAPx10_ASAP7_75t_R FILLER_186_222 ();
 DECAPx10_ASAP7_75t_R FILLER_186_244 ();
 DECAPx10_ASAP7_75t_R FILLER_186_266 ();
 DECAPx1_ASAP7_75t_R FILLER_186_288 ();
 FILLER_ASAP7_75t_R FILLER_186_309 ();
 DECAPx6_ASAP7_75t_R FILLER_186_317 ();
 DECAPx4_ASAP7_75t_R FILLER_186_337 ();
 FILLER_ASAP7_75t_R FILLER_186_347 ();
 DECAPx10_ASAP7_75t_R FILLER_186_355 ();
 DECAPx2_ASAP7_75t_R FILLER_186_377 ();
 FILLER_ASAP7_75t_R FILLER_186_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_385 ();
 DECAPx10_ASAP7_75t_R FILLER_186_398 ();
 DECAPx2_ASAP7_75t_R FILLER_186_420 ();
 FILLER_ASAP7_75t_R FILLER_186_426 ();
 FILLER_ASAP7_75t_R FILLER_186_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_461 ();
 DECAPx2_ASAP7_75t_R FILLER_186_464 ();
 FILLER_ASAP7_75t_R FILLER_186_470 ();
 DECAPx2_ASAP7_75t_R FILLER_186_494 ();
 FILLER_ASAP7_75t_R FILLER_186_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_502 ();
 FILLER_ASAP7_75t_R FILLER_186_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_521 ();
 DECAPx10_ASAP7_75t_R FILLER_186_528 ();
 DECAPx10_ASAP7_75t_R FILLER_186_550 ();
 DECAPx10_ASAP7_75t_R FILLER_186_572 ();
 DECAPx1_ASAP7_75t_R FILLER_186_594 ();
 DECAPx2_ASAP7_75t_R FILLER_186_618 ();
 FILLER_ASAP7_75t_R FILLER_186_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_633 ();
 DECAPx6_ASAP7_75t_R FILLER_186_640 ();
 FILLER_ASAP7_75t_R FILLER_186_654 ();
 DECAPx2_ASAP7_75t_R FILLER_186_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_669 ();
 DECAPx6_ASAP7_75t_R FILLER_186_682 ();
 FILLER_ASAP7_75t_R FILLER_186_696 ();
 DECAPx10_ASAP7_75t_R FILLER_186_710 ();
 FILLER_ASAP7_75t_R FILLER_186_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_734 ();
 DECAPx4_ASAP7_75t_R FILLER_186_738 ();
 DECAPx2_ASAP7_75t_R FILLER_186_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_760 ();
 DECAPx1_ASAP7_75t_R FILLER_186_771 ();
 DECAPx6_ASAP7_75t_R FILLER_186_781 ();
 FILLER_ASAP7_75t_R FILLER_186_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_850 ();
 DECAPx1_ASAP7_75t_R FILLER_186_871 ();
 DECAPx2_ASAP7_75t_R FILLER_186_878 ();
 FILLER_ASAP7_75t_R FILLER_186_912 ();
 FILLER_ASAP7_75t_R FILLER_186_922 ();
 DECAPx4_ASAP7_75t_R FILLER_186_946 ();
 FILLER_ASAP7_75t_R FILLER_186_956 ();
 DECAPx6_ASAP7_75t_R FILLER_186_980 ();
 FILLER_ASAP7_75t_R FILLER_186_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1017 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1024 ();
 FILLER_ASAP7_75t_R FILLER_186_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1047 ();
 FILLER_ASAP7_75t_R FILLER_186_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1083 ();
 FILLER_ASAP7_75t_R FILLER_186_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_186_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_187_2 ();
 DECAPx10_ASAP7_75t_R FILLER_187_24 ();
 DECAPx10_ASAP7_75t_R FILLER_187_46 ();
 DECAPx10_ASAP7_75t_R FILLER_187_68 ();
 DECAPx10_ASAP7_75t_R FILLER_187_90 ();
 DECAPx10_ASAP7_75t_R FILLER_187_112 ();
 DECAPx10_ASAP7_75t_R FILLER_187_134 ();
 DECAPx10_ASAP7_75t_R FILLER_187_156 ();
 DECAPx10_ASAP7_75t_R FILLER_187_178 ();
 DECAPx10_ASAP7_75t_R FILLER_187_200 ();
 DECAPx10_ASAP7_75t_R FILLER_187_222 ();
 DECAPx10_ASAP7_75t_R FILLER_187_244 ();
 DECAPx6_ASAP7_75t_R FILLER_187_266 ();
 DECAPx1_ASAP7_75t_R FILLER_187_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_284 ();
 DECAPx2_ASAP7_75t_R FILLER_187_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_346 ();
 DECAPx2_ASAP7_75t_R FILLER_187_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_375 ();
 DECAPx4_ASAP7_75t_R FILLER_187_382 ();
 FILLER_ASAP7_75t_R FILLER_187_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_402 ();
 DECAPx2_ASAP7_75t_R FILLER_187_420 ();
 FILLER_ASAP7_75t_R FILLER_187_426 ();
 DECAPx10_ASAP7_75t_R FILLER_187_452 ();
 FILLER_ASAP7_75t_R FILLER_187_474 ();
 DECAPx1_ASAP7_75t_R FILLER_187_479 ();
 FILLER_ASAP7_75t_R FILLER_187_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_505 ();
 DECAPx2_ASAP7_75t_R FILLER_187_510 ();
 FILLER_ASAP7_75t_R FILLER_187_516 ();
 DECAPx2_ASAP7_75t_R FILLER_187_540 ();
 FILLER_ASAP7_75t_R FILLER_187_546 ();
 FILLER_ASAP7_75t_R FILLER_187_559 ();
 FILLER_ASAP7_75t_R FILLER_187_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_570 ();
 DECAPx6_ASAP7_75t_R FILLER_187_593 ();
 DECAPx1_ASAP7_75t_R FILLER_187_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_633 ();
 DECAPx2_ASAP7_75t_R FILLER_187_650 ();
 DECAPx10_ASAP7_75t_R FILLER_187_668 ();
 DECAPx10_ASAP7_75t_R FILLER_187_690 ();
 FILLER_ASAP7_75t_R FILLER_187_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_714 ();
 DECAPx2_ASAP7_75t_R FILLER_187_721 ();
 FILLER_ASAP7_75t_R FILLER_187_727 ();
 FILLER_ASAP7_75t_R FILLER_187_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_737 ();
 FILLER_ASAP7_75t_R FILLER_187_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_748 ();
 DECAPx6_ASAP7_75t_R FILLER_187_759 ();
 DECAPx6_ASAP7_75t_R FILLER_187_779 ();
 DECAPx1_ASAP7_75t_R FILLER_187_793 ();
 DECAPx10_ASAP7_75t_R FILLER_187_817 ();
 FILLER_ASAP7_75t_R FILLER_187_839 ();
 DECAPx2_ASAP7_75t_R FILLER_187_863 ();
 DECAPx6_ASAP7_75t_R FILLER_187_875 ();
 DECAPx1_ASAP7_75t_R FILLER_187_889 ();
 DECAPx2_ASAP7_75t_R FILLER_187_906 ();
 FILLER_ASAP7_75t_R FILLER_187_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_914 ();
 FILLER_ASAP7_75t_R FILLER_187_922 ();
 DECAPx2_ASAP7_75t_R FILLER_187_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_965 ();
 FILLER_ASAP7_75t_R FILLER_187_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_995 ();
 FILLER_ASAP7_75t_R FILLER_187_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_187_1062 ();
 FILLER_ASAP7_75t_R FILLER_187_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_187_1192 ();
 DECAPx1_ASAP7_75t_R FILLER_187_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_188_2 ();
 DECAPx10_ASAP7_75t_R FILLER_188_24 ();
 DECAPx10_ASAP7_75t_R FILLER_188_46 ();
 DECAPx10_ASAP7_75t_R FILLER_188_68 ();
 DECAPx10_ASAP7_75t_R FILLER_188_90 ();
 DECAPx10_ASAP7_75t_R FILLER_188_112 ();
 DECAPx10_ASAP7_75t_R FILLER_188_134 ();
 DECAPx10_ASAP7_75t_R FILLER_188_156 ();
 DECAPx10_ASAP7_75t_R FILLER_188_178 ();
 DECAPx10_ASAP7_75t_R FILLER_188_200 ();
 DECAPx10_ASAP7_75t_R FILLER_188_222 ();
 DECAPx10_ASAP7_75t_R FILLER_188_244 ();
 DECAPx10_ASAP7_75t_R FILLER_188_266 ();
 DECAPx10_ASAP7_75t_R FILLER_188_288 ();
 DECAPx6_ASAP7_75t_R FILLER_188_310 ();
 DECAPx2_ASAP7_75t_R FILLER_188_324 ();
 DECAPx10_ASAP7_75t_R FILLER_188_336 ();
 DECAPx6_ASAP7_75t_R FILLER_188_358 ();
 FILLER_ASAP7_75t_R FILLER_188_372 ();
 DECAPx4_ASAP7_75t_R FILLER_188_404 ();
 DECAPx2_ASAP7_75t_R FILLER_188_436 ();
 DECAPx4_ASAP7_75t_R FILLER_188_452 ();
 DECAPx10_ASAP7_75t_R FILLER_188_464 ();
 DECAPx6_ASAP7_75t_R FILLER_188_486 ();
 FILLER_ASAP7_75t_R FILLER_188_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_502 ();
 FILLER_ASAP7_75t_R FILLER_188_509 ();
 DECAPx1_ASAP7_75t_R FILLER_188_517 ();
 DECAPx6_ASAP7_75t_R FILLER_188_527 ();
 FILLER_ASAP7_75t_R FILLER_188_541 ();
 FILLER_ASAP7_75t_R FILLER_188_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_565 ();
 DECAPx1_ASAP7_75t_R FILLER_188_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_584 ();
 DECAPx4_ASAP7_75t_R FILLER_188_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_615 ();
 DECAPx4_ASAP7_75t_R FILLER_188_626 ();
 DECAPx4_ASAP7_75t_R FILLER_188_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_652 ();
 DECAPx2_ASAP7_75t_R FILLER_188_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_681 ();
 DECAPx2_ASAP7_75t_R FILLER_188_692 ();
 FILLER_ASAP7_75t_R FILLER_188_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_700 ();
 DECAPx1_ASAP7_75t_R FILLER_188_719 ();
 DECAPx1_ASAP7_75t_R FILLER_188_761 ();
 DECAPx1_ASAP7_75t_R FILLER_188_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_809 ();
 DECAPx1_ASAP7_75t_R FILLER_188_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_824 ();
 DECAPx6_ASAP7_75t_R FILLER_188_828 ();
 DECAPx1_ASAP7_75t_R FILLER_188_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_846 ();
 DECAPx6_ASAP7_75t_R FILLER_188_853 ();
 DECAPx10_ASAP7_75t_R FILLER_188_887 ();
 DECAPx2_ASAP7_75t_R FILLER_188_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_915 ();
 DECAPx10_ASAP7_75t_R FILLER_188_922 ();
 DECAPx6_ASAP7_75t_R FILLER_188_944 ();
 FILLER_ASAP7_75t_R FILLER_188_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_982 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1025 ();
 FILLER_ASAP7_75t_R FILLER_188_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1050 ();
 FILLER_ASAP7_75t_R FILLER_188_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1098 ();
 FILLER_ASAP7_75t_R FILLER_188_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1121 ();
 FILLER_ASAP7_75t_R FILLER_188_1125 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1134 ();
 FILLER_ASAP7_75t_R FILLER_188_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_189_2 ();
 DECAPx10_ASAP7_75t_R FILLER_189_24 ();
 DECAPx10_ASAP7_75t_R FILLER_189_46 ();
 DECAPx10_ASAP7_75t_R FILLER_189_68 ();
 DECAPx10_ASAP7_75t_R FILLER_189_90 ();
 DECAPx10_ASAP7_75t_R FILLER_189_112 ();
 DECAPx10_ASAP7_75t_R FILLER_189_134 ();
 DECAPx10_ASAP7_75t_R FILLER_189_156 ();
 DECAPx10_ASAP7_75t_R FILLER_189_178 ();
 DECAPx10_ASAP7_75t_R FILLER_189_200 ();
 DECAPx10_ASAP7_75t_R FILLER_189_222 ();
 DECAPx10_ASAP7_75t_R FILLER_189_244 ();
 DECAPx10_ASAP7_75t_R FILLER_189_266 ();
 DECAPx6_ASAP7_75t_R FILLER_189_288 ();
 DECAPx1_ASAP7_75t_R FILLER_189_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_306 ();
 DECAPx6_ASAP7_75t_R FILLER_189_318 ();
 DECAPx1_ASAP7_75t_R FILLER_189_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_358 ();
 FILLER_ASAP7_75t_R FILLER_189_369 ();
 DECAPx4_ASAP7_75t_R FILLER_189_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_387 ();
 DECAPx10_ASAP7_75t_R FILLER_189_402 ();
 DECAPx10_ASAP7_75t_R FILLER_189_424 ();
 DECAPx10_ASAP7_75t_R FILLER_189_446 ();
 DECAPx2_ASAP7_75t_R FILLER_189_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_529 ();
 DECAPx2_ASAP7_75t_R FILLER_189_537 ();
 FILLER_ASAP7_75t_R FILLER_189_543 ();
 FILLER_ASAP7_75t_R FILLER_189_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_575 ();
 DECAPx2_ASAP7_75t_R FILLER_189_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_599 ();
 DECAPx2_ASAP7_75t_R FILLER_189_622 ();
 FILLER_ASAP7_75t_R FILLER_189_628 ();
 DECAPx4_ASAP7_75t_R FILLER_189_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_678 ();
 DECAPx1_ASAP7_75t_R FILLER_189_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_703 ();
 FILLER_ASAP7_75t_R FILLER_189_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_724 ();
 FILLER_ASAP7_75t_R FILLER_189_732 ();
 DECAPx1_ASAP7_75t_R FILLER_189_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_760 ();
 DECAPx2_ASAP7_75t_R FILLER_189_767 ();
 FILLER_ASAP7_75t_R FILLER_189_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_775 ();
 DECAPx4_ASAP7_75t_R FILLER_189_782 ();
 FILLER_ASAP7_75t_R FILLER_189_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_794 ();
 DECAPx10_ASAP7_75t_R FILLER_189_839 ();
 DECAPx10_ASAP7_75t_R FILLER_189_861 ();
 DECAPx1_ASAP7_75t_R FILLER_189_883 ();
 FILLER_ASAP7_75t_R FILLER_189_905 ();
 DECAPx4_ASAP7_75t_R FILLER_189_911 ();
 FILLER_ASAP7_75t_R FILLER_189_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_923 ();
 DECAPx6_ASAP7_75t_R FILLER_189_926 ();
 FILLER_ASAP7_75t_R FILLER_189_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_964 ();
 DECAPx4_ASAP7_75t_R FILLER_189_971 ();
 FILLER_ASAP7_75t_R FILLER_189_981 ();
 DECAPx2_ASAP7_75t_R FILLER_189_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_995 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1002 ();
 DECAPx4_ASAP7_75t_R FILLER_189_1024 ();
 FILLER_ASAP7_75t_R FILLER_189_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1036 ();
 FILLER_ASAP7_75t_R FILLER_189_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1175 ();
 FILLER_ASAP7_75t_R FILLER_189_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1192 ();
 FILLER_ASAP7_75t_R FILLER_189_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_190_2 ();
 DECAPx10_ASAP7_75t_R FILLER_190_24 ();
 DECAPx10_ASAP7_75t_R FILLER_190_46 ();
 DECAPx10_ASAP7_75t_R FILLER_190_68 ();
 DECAPx10_ASAP7_75t_R FILLER_190_90 ();
 DECAPx10_ASAP7_75t_R FILLER_190_112 ();
 DECAPx10_ASAP7_75t_R FILLER_190_134 ();
 DECAPx10_ASAP7_75t_R FILLER_190_156 ();
 DECAPx10_ASAP7_75t_R FILLER_190_178 ();
 DECAPx10_ASAP7_75t_R FILLER_190_200 ();
 DECAPx10_ASAP7_75t_R FILLER_190_222 ();
 DECAPx10_ASAP7_75t_R FILLER_190_244 ();
 DECAPx10_ASAP7_75t_R FILLER_190_266 ();
 FILLER_ASAP7_75t_R FILLER_190_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_290 ();
 DECAPx6_ASAP7_75t_R FILLER_190_297 ();
 FILLER_ASAP7_75t_R FILLER_190_331 ();
 DECAPx10_ASAP7_75t_R FILLER_190_341 ();
 DECAPx10_ASAP7_75t_R FILLER_190_363 ();
 DECAPx2_ASAP7_75t_R FILLER_190_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_405 ();
 DECAPx4_ASAP7_75t_R FILLER_190_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_433 ();
 DECAPx2_ASAP7_75t_R FILLER_190_454 ();
 FILLER_ASAP7_75t_R FILLER_190_460 ();
 DECAPx2_ASAP7_75t_R FILLER_190_464 ();
 DECAPx2_ASAP7_75t_R FILLER_190_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_499 ();
 DECAPx10_ASAP7_75t_R FILLER_190_530 ();
 DECAPx4_ASAP7_75t_R FILLER_190_552 ();
 FILLER_ASAP7_75t_R FILLER_190_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_564 ();
 FILLER_ASAP7_75t_R FILLER_190_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_573 ();
 DECAPx1_ASAP7_75t_R FILLER_190_596 ();
 DECAPx2_ASAP7_75t_R FILLER_190_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_616 ();
 DECAPx1_ASAP7_75t_R FILLER_190_642 ();
 DECAPx1_ASAP7_75t_R FILLER_190_668 ();
 DECAPx1_ASAP7_75t_R FILLER_190_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_682 ();
 FILLER_ASAP7_75t_R FILLER_190_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_695 ();
 DECAPx2_ASAP7_75t_R FILLER_190_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_726 ();
 DECAPx10_ASAP7_75t_R FILLER_190_733 ();
 DECAPx10_ASAP7_75t_R FILLER_190_755 ();
 FILLER_ASAP7_75t_R FILLER_190_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_806 ();
 DECAPx6_ASAP7_75t_R FILLER_190_817 ();
 FILLER_ASAP7_75t_R FILLER_190_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_843 ();
 DECAPx10_ASAP7_75t_R FILLER_190_870 ();
 FILLER_ASAP7_75t_R FILLER_190_899 ();
 DECAPx10_ASAP7_75t_R FILLER_190_921 ();
 DECAPx10_ASAP7_75t_R FILLER_190_943 ();
 DECAPx10_ASAP7_75t_R FILLER_190_965 ();
 FILLER_ASAP7_75t_R FILLER_190_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_996 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1045 ();
 FILLER_ASAP7_75t_R FILLER_190_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1176 ();
 FILLER_ASAP7_75t_R FILLER_190_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1187 ();
 DECAPx4_ASAP7_75t_R FILLER_190_1193 ();
 FILLER_ASAP7_75t_R FILLER_190_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1205 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_191_2 ();
 DECAPx10_ASAP7_75t_R FILLER_191_24 ();
 DECAPx10_ASAP7_75t_R FILLER_191_46 ();
 DECAPx10_ASAP7_75t_R FILLER_191_68 ();
 DECAPx10_ASAP7_75t_R FILLER_191_90 ();
 DECAPx10_ASAP7_75t_R FILLER_191_112 ();
 DECAPx10_ASAP7_75t_R FILLER_191_134 ();
 DECAPx10_ASAP7_75t_R FILLER_191_156 ();
 DECAPx10_ASAP7_75t_R FILLER_191_178 ();
 DECAPx10_ASAP7_75t_R FILLER_191_200 ();
 DECAPx10_ASAP7_75t_R FILLER_191_222 ();
 DECAPx10_ASAP7_75t_R FILLER_191_244 ();
 DECAPx6_ASAP7_75t_R FILLER_191_266 ();
 DECAPx2_ASAP7_75t_R FILLER_191_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_286 ();
 DECAPx1_ASAP7_75t_R FILLER_191_309 ();
 DECAPx6_ASAP7_75t_R FILLER_191_319 ();
 DECAPx2_ASAP7_75t_R FILLER_191_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_367 ();
 DECAPx1_ASAP7_75t_R FILLER_191_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_388 ();
 FILLER_ASAP7_75t_R FILLER_191_419 ();
 DECAPx4_ASAP7_75t_R FILLER_191_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_437 ();
 DECAPx4_ASAP7_75t_R FILLER_191_441 ();
 FILLER_ASAP7_75t_R FILLER_191_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_476 ();
 DECAPx10_ASAP7_75t_R FILLER_191_481 ();
 FILLER_ASAP7_75t_R FILLER_191_507 ();
 FILLER_ASAP7_75t_R FILLER_191_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_517 ();
 DECAPx6_ASAP7_75t_R FILLER_191_536 ();
 DECAPx1_ASAP7_75t_R FILLER_191_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_574 ();
 DECAPx10_ASAP7_75t_R FILLER_191_592 ();
 FILLER_ASAP7_75t_R FILLER_191_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_616 ();
 FILLER_ASAP7_75t_R FILLER_191_645 ();
 DECAPx6_ASAP7_75t_R FILLER_191_653 ();
 DECAPx1_ASAP7_75t_R FILLER_191_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_699 ();
 DECAPx6_ASAP7_75t_R FILLER_191_706 ();
 FILLER_ASAP7_75t_R FILLER_191_720 ();
 DECAPx2_ASAP7_75t_R FILLER_191_736 ();
 FILLER_ASAP7_75t_R FILLER_191_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_744 ();
 DECAPx2_ASAP7_75t_R FILLER_191_757 ();
 FILLER_ASAP7_75t_R FILLER_191_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_765 ();
 DECAPx6_ASAP7_75t_R FILLER_191_786 ();
 FILLER_ASAP7_75t_R FILLER_191_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_802 ();
 DECAPx6_ASAP7_75t_R FILLER_191_815 ();
 DECAPx2_ASAP7_75t_R FILLER_191_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_835 ();
 FILLER_ASAP7_75t_R FILLER_191_856 ();
 FILLER_ASAP7_75t_R FILLER_191_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_926 ();
 DECAPx10_ASAP7_75t_R FILLER_191_931 ();
 DECAPx10_ASAP7_75t_R FILLER_191_953 ();
 DECAPx1_ASAP7_75t_R FILLER_191_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_979 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1022 ();
 FILLER_ASAP7_75t_R FILLER_191_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1079 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1159 ();
 FILLER_ASAP7_75t_R FILLER_191_1181 ();
 FILLER_ASAP7_75t_R FILLER_191_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1209 ();
 FILLER_ASAP7_75t_R FILLER_191_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_192_2 ();
 DECAPx10_ASAP7_75t_R FILLER_192_24 ();
 DECAPx10_ASAP7_75t_R FILLER_192_46 ();
 DECAPx10_ASAP7_75t_R FILLER_192_68 ();
 DECAPx10_ASAP7_75t_R FILLER_192_90 ();
 DECAPx10_ASAP7_75t_R FILLER_192_112 ();
 DECAPx10_ASAP7_75t_R FILLER_192_134 ();
 DECAPx10_ASAP7_75t_R FILLER_192_156 ();
 DECAPx10_ASAP7_75t_R FILLER_192_178 ();
 DECAPx10_ASAP7_75t_R FILLER_192_200 ();
 DECAPx10_ASAP7_75t_R FILLER_192_222 ();
 DECAPx10_ASAP7_75t_R FILLER_192_244 ();
 DECAPx10_ASAP7_75t_R FILLER_192_266 ();
 DECAPx2_ASAP7_75t_R FILLER_192_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_294 ();
 DECAPx6_ASAP7_75t_R FILLER_192_306 ();
 FILLER_ASAP7_75t_R FILLER_192_320 ();
 DECAPx2_ASAP7_75t_R FILLER_192_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_334 ();
 DECAPx2_ASAP7_75t_R FILLER_192_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_361 ();
 FILLER_ASAP7_75t_R FILLER_192_377 ();
 DECAPx2_ASAP7_75t_R FILLER_192_385 ();
 FILLER_ASAP7_75t_R FILLER_192_399 ();
 DECAPx4_ASAP7_75t_R FILLER_192_411 ();
 DECAPx6_ASAP7_75t_R FILLER_192_443 ();
 DECAPx1_ASAP7_75t_R FILLER_192_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_461 ();
 DECAPx10_ASAP7_75t_R FILLER_192_464 ();
 DECAPx2_ASAP7_75t_R FILLER_192_486 ();
 FILLER_ASAP7_75t_R FILLER_192_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_514 ();
 DECAPx6_ASAP7_75t_R FILLER_192_528 ();
 DECAPx10_ASAP7_75t_R FILLER_192_584 ();
 DECAPx4_ASAP7_75t_R FILLER_192_606 ();
 FILLER_ASAP7_75t_R FILLER_192_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_640 ();
 DECAPx2_ASAP7_75t_R FILLER_192_669 ();
 FILLER_ASAP7_75t_R FILLER_192_675 ();
 DECAPx2_ASAP7_75t_R FILLER_192_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_691 ();
 DECAPx4_ASAP7_75t_R FILLER_192_706 ();
 FILLER_ASAP7_75t_R FILLER_192_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_718 ();
 FILLER_ASAP7_75t_R FILLER_192_725 ();
 DECAPx2_ASAP7_75t_R FILLER_192_739 ();
 FILLER_ASAP7_75t_R FILLER_192_745 ();
 DECAPx1_ASAP7_75t_R FILLER_192_774 ();
 FILLER_ASAP7_75t_R FILLER_192_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_800 ();
 DECAPx1_ASAP7_75t_R FILLER_192_807 ();
 DECAPx6_ASAP7_75t_R FILLER_192_844 ();
 DECAPx2_ASAP7_75t_R FILLER_192_858 ();
 FILLER_ASAP7_75t_R FILLER_192_870 ();
 DECAPx2_ASAP7_75t_R FILLER_192_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_906 ();
 DECAPx2_ASAP7_75t_R FILLER_192_917 ();
 FILLER_ASAP7_75t_R FILLER_192_923 ();
 DECAPx10_ASAP7_75t_R FILLER_192_931 ();
 DECAPx1_ASAP7_75t_R FILLER_192_953 ();
 DECAPx6_ASAP7_75t_R FILLER_192_961 ();
 DECAPx1_ASAP7_75t_R FILLER_192_975 ();
 DECAPx2_ASAP7_75t_R FILLER_192_985 ();
 FILLER_ASAP7_75t_R FILLER_192_991 ();
 DECAPx1_ASAP7_75t_R FILLER_192_999 ();
 DECAPx2_ASAP7_75t_R FILLER_192_1023 ();
 FILLER_ASAP7_75t_R FILLER_192_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1085 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1107 ();
 FILLER_ASAP7_75t_R FILLER_192_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1193 ();
 FILLER_ASAP7_75t_R FILLER_192_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_193_2 ();
 DECAPx10_ASAP7_75t_R FILLER_193_24 ();
 DECAPx10_ASAP7_75t_R FILLER_193_46 ();
 DECAPx10_ASAP7_75t_R FILLER_193_68 ();
 DECAPx10_ASAP7_75t_R FILLER_193_90 ();
 DECAPx10_ASAP7_75t_R FILLER_193_112 ();
 DECAPx10_ASAP7_75t_R FILLER_193_134 ();
 DECAPx10_ASAP7_75t_R FILLER_193_156 ();
 DECAPx10_ASAP7_75t_R FILLER_193_178 ();
 DECAPx10_ASAP7_75t_R FILLER_193_200 ();
 DECAPx10_ASAP7_75t_R FILLER_193_222 ();
 DECAPx10_ASAP7_75t_R FILLER_193_244 ();
 DECAPx10_ASAP7_75t_R FILLER_193_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_288 ();
 FILLER_ASAP7_75t_R FILLER_193_300 ();
 DECAPx2_ASAP7_75t_R FILLER_193_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_321 ();
 DECAPx2_ASAP7_75t_R FILLER_193_358 ();
 DECAPx10_ASAP7_75t_R FILLER_193_386 ();
 DECAPx10_ASAP7_75t_R FILLER_193_408 ();
 DECAPx10_ASAP7_75t_R FILLER_193_430 ();
 DECAPx2_ASAP7_75t_R FILLER_193_452 ();
 DECAPx4_ASAP7_75t_R FILLER_193_469 ();
 FILLER_ASAP7_75t_R FILLER_193_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_501 ();
 FILLER_ASAP7_75t_R FILLER_193_523 ();
 DECAPx1_ASAP7_75t_R FILLER_193_547 ();
 DECAPx1_ASAP7_75t_R FILLER_193_557 ();
 FILLER_ASAP7_75t_R FILLER_193_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_570 ();
 DECAPx10_ASAP7_75t_R FILLER_193_579 ();
 DECAPx6_ASAP7_75t_R FILLER_193_601 ();
 DECAPx1_ASAP7_75t_R FILLER_193_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_619 ();
 DECAPx10_ASAP7_75t_R FILLER_193_642 ();
 DECAPx2_ASAP7_75t_R FILLER_193_680 ();
 FILLER_ASAP7_75t_R FILLER_193_686 ();
 DECAPx2_ASAP7_75t_R FILLER_193_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_729 ();
 FILLER_ASAP7_75t_R FILLER_193_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_752 ();
 FILLER_ASAP7_75t_R FILLER_193_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_768 ();
 DECAPx2_ASAP7_75t_R FILLER_193_775 ();
 FILLER_ASAP7_75t_R FILLER_193_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_783 ();
 DECAPx6_ASAP7_75t_R FILLER_193_836 ();
 FILLER_ASAP7_75t_R FILLER_193_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_874 ();
 DECAPx1_ASAP7_75t_R FILLER_193_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_896 ();
 DECAPx2_ASAP7_75t_R FILLER_193_915 ();
 FILLER_ASAP7_75t_R FILLER_193_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_923 ();
 FILLER_ASAP7_75t_R FILLER_193_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_954 ();
 DECAPx6_ASAP7_75t_R FILLER_193_969 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1009 ();
 FILLER_ASAP7_75t_R FILLER_193_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_193_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1077 ();
 FILLER_ASAP7_75t_R FILLER_193_1083 ();
 FILLER_ASAP7_75t_R FILLER_193_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_193_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1146 ();
 DECAPx6_ASAP7_75t_R FILLER_193_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1181 ();
 FILLER_ASAP7_75t_R FILLER_193_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1211 ();
 FILLER_ASAP7_75t_R FILLER_193_1217 ();
 FILLER_ASAP7_75t_R FILLER_193_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_194_2 ();
 DECAPx10_ASAP7_75t_R FILLER_194_24 ();
 DECAPx10_ASAP7_75t_R FILLER_194_46 ();
 DECAPx10_ASAP7_75t_R FILLER_194_68 ();
 DECAPx10_ASAP7_75t_R FILLER_194_90 ();
 DECAPx10_ASAP7_75t_R FILLER_194_112 ();
 DECAPx10_ASAP7_75t_R FILLER_194_134 ();
 DECAPx10_ASAP7_75t_R FILLER_194_156 ();
 DECAPx10_ASAP7_75t_R FILLER_194_178 ();
 DECAPx10_ASAP7_75t_R FILLER_194_200 ();
 DECAPx10_ASAP7_75t_R FILLER_194_222 ();
 DECAPx10_ASAP7_75t_R FILLER_194_244 ();
 DECAPx4_ASAP7_75t_R FILLER_194_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_276 ();
 DECAPx1_ASAP7_75t_R FILLER_194_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_303 ();
 DECAPx10_ASAP7_75t_R FILLER_194_312 ();
 DECAPx2_ASAP7_75t_R FILLER_194_334 ();
 FILLER_ASAP7_75t_R FILLER_194_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_342 ();
 DECAPx6_ASAP7_75t_R FILLER_194_355 ();
 DECAPx2_ASAP7_75t_R FILLER_194_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_375 ();
 DECAPx10_ASAP7_75t_R FILLER_194_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_415 ();
 FILLER_ASAP7_75t_R FILLER_194_460 ();
 FILLER_ASAP7_75t_R FILLER_194_464 ();
 DECAPx2_ASAP7_75t_R FILLER_194_488 ();
 FILLER_ASAP7_75t_R FILLER_194_494 ();
 DECAPx4_ASAP7_75t_R FILLER_194_508 ();
 DECAPx10_ASAP7_75t_R FILLER_194_530 ();
 DECAPx2_ASAP7_75t_R FILLER_194_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_558 ();
 DECAPx1_ASAP7_75t_R FILLER_194_567 ();
 DECAPx10_ASAP7_75t_R FILLER_194_588 ();
 DECAPx6_ASAP7_75t_R FILLER_194_610 ();
 FILLER_ASAP7_75t_R FILLER_194_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_626 ();
 DECAPx10_ASAP7_75t_R FILLER_194_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_671 ();
 DECAPx10_ASAP7_75t_R FILLER_194_678 ();
 DECAPx4_ASAP7_75t_R FILLER_194_700 ();
 FILLER_ASAP7_75t_R FILLER_194_724 ();
 DECAPx6_ASAP7_75t_R FILLER_194_738 ();
 FILLER_ASAP7_75t_R FILLER_194_752 ();
 DECAPx4_ASAP7_75t_R FILLER_194_766 ();
 DECAPx6_ASAP7_75t_R FILLER_194_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_818 ();
 DECAPx10_ASAP7_75t_R FILLER_194_825 ();
 DECAPx2_ASAP7_75t_R FILLER_194_847 ();
 DECAPx10_ASAP7_75t_R FILLER_194_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_881 ();
 DECAPx10_ASAP7_75t_R FILLER_194_888 ();
 FILLER_ASAP7_75t_R FILLER_194_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_912 ();
 DECAPx6_ASAP7_75t_R FILLER_194_922 ();
 FILLER_ASAP7_75t_R FILLER_194_936 ();
 DECAPx6_ASAP7_75t_R FILLER_194_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1002 ();
 FILLER_ASAP7_75t_R FILLER_194_1023 ();
 FILLER_ASAP7_75t_R FILLER_194_1031 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_194_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1106 ();
 FILLER_ASAP7_75t_R FILLER_194_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1132 ();
 FILLER_ASAP7_75t_R FILLER_194_1154 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1172 ();
 FILLER_ASAP7_75t_R FILLER_194_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_195_2 ();
 DECAPx10_ASAP7_75t_R FILLER_195_24 ();
 DECAPx10_ASAP7_75t_R FILLER_195_46 ();
 DECAPx10_ASAP7_75t_R FILLER_195_68 ();
 DECAPx10_ASAP7_75t_R FILLER_195_90 ();
 DECAPx10_ASAP7_75t_R FILLER_195_112 ();
 DECAPx10_ASAP7_75t_R FILLER_195_134 ();
 DECAPx10_ASAP7_75t_R FILLER_195_156 ();
 DECAPx10_ASAP7_75t_R FILLER_195_178 ();
 DECAPx10_ASAP7_75t_R FILLER_195_200 ();
 DECAPx10_ASAP7_75t_R FILLER_195_222 ();
 DECAPx10_ASAP7_75t_R FILLER_195_244 ();
 DECAPx10_ASAP7_75t_R FILLER_195_266 ();
 FILLER_ASAP7_75t_R FILLER_195_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_290 ();
 DECAPx1_ASAP7_75t_R FILLER_195_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_301 ();
 DECAPx4_ASAP7_75t_R FILLER_195_309 ();
 DECAPx4_ASAP7_75t_R FILLER_195_330 ();
 FILLER_ASAP7_75t_R FILLER_195_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_342 ();
 DECAPx2_ASAP7_75t_R FILLER_195_357 ();
 FILLER_ASAP7_75t_R FILLER_195_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_365 ();
 DECAPx2_ASAP7_75t_R FILLER_195_377 ();
 FILLER_ASAP7_75t_R FILLER_195_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_385 ();
 DECAPx4_ASAP7_75t_R FILLER_195_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_429 ();
 DECAPx6_ASAP7_75t_R FILLER_195_436 ();
 DECAPx4_ASAP7_75t_R FILLER_195_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_466 ();
 DECAPx10_ASAP7_75t_R FILLER_195_473 ();
 DECAPx1_ASAP7_75t_R FILLER_195_495 ();
 DECAPx4_ASAP7_75t_R FILLER_195_510 ();
 DECAPx6_ASAP7_75t_R FILLER_195_532 ();
 DECAPx2_ASAP7_75t_R FILLER_195_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_552 ();
 DECAPx2_ASAP7_75t_R FILLER_195_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_581 ();
 DECAPx10_ASAP7_75t_R FILLER_195_604 ();
 DECAPx1_ASAP7_75t_R FILLER_195_626 ();
 FILLER_ASAP7_75t_R FILLER_195_637 ();
 DECAPx2_ASAP7_75t_R FILLER_195_667 ();
 DECAPx6_ASAP7_75t_R FILLER_195_681 ();
 DECAPx2_ASAP7_75t_R FILLER_195_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_727 ();
 DECAPx1_ASAP7_75t_R FILLER_195_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_739 ();
 DECAPx6_ASAP7_75t_R FILLER_195_764 ();
 DECAPx4_ASAP7_75t_R FILLER_195_808 ();
 DECAPx10_ASAP7_75t_R FILLER_195_826 ();
 DECAPx2_ASAP7_75t_R FILLER_195_848 ();
 FILLER_ASAP7_75t_R FILLER_195_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_856 ();
 FILLER_ASAP7_75t_R FILLER_195_863 ();
 DECAPx2_ASAP7_75t_R FILLER_195_887 ();
 FILLER_ASAP7_75t_R FILLER_195_893 ();
 DECAPx2_ASAP7_75t_R FILLER_195_918 ();
 DECAPx4_ASAP7_75t_R FILLER_195_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_956 ();
 DECAPx2_ASAP7_75t_R FILLER_195_961 ();
 DECAPx1_ASAP7_75t_R FILLER_195_991 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_196_2 ();
 DECAPx10_ASAP7_75t_R FILLER_196_24 ();
 DECAPx10_ASAP7_75t_R FILLER_196_46 ();
 DECAPx10_ASAP7_75t_R FILLER_196_68 ();
 DECAPx10_ASAP7_75t_R FILLER_196_90 ();
 DECAPx10_ASAP7_75t_R FILLER_196_112 ();
 DECAPx10_ASAP7_75t_R FILLER_196_134 ();
 DECAPx10_ASAP7_75t_R FILLER_196_156 ();
 DECAPx10_ASAP7_75t_R FILLER_196_178 ();
 DECAPx10_ASAP7_75t_R FILLER_196_200 ();
 DECAPx10_ASAP7_75t_R FILLER_196_222 ();
 DECAPx10_ASAP7_75t_R FILLER_196_244 ();
 DECAPx10_ASAP7_75t_R FILLER_196_266 ();
 DECAPx6_ASAP7_75t_R FILLER_196_288 ();
 FILLER_ASAP7_75t_R FILLER_196_302 ();
 DECAPx1_ASAP7_75t_R FILLER_196_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_342 ();
 DECAPx4_ASAP7_75t_R FILLER_196_365 ();
 DECAPx6_ASAP7_75t_R FILLER_196_381 ();
 DECAPx2_ASAP7_75t_R FILLER_196_395 ();
 DECAPx4_ASAP7_75t_R FILLER_196_431 ();
 FILLER_ASAP7_75t_R FILLER_196_441 ();
 FILLER_ASAP7_75t_R FILLER_196_454 ();
 DECAPx6_ASAP7_75t_R FILLER_196_486 ();
 DECAPx1_ASAP7_75t_R FILLER_196_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_504 ();
 DECAPx2_ASAP7_75t_R FILLER_196_527 ();
 FILLER_ASAP7_75t_R FILLER_196_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_535 ();
 FILLER_ASAP7_75t_R FILLER_196_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_566 ();
 DECAPx6_ASAP7_75t_R FILLER_196_600 ();
 DECAPx2_ASAP7_75t_R FILLER_196_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_620 ();
 DECAPx6_ASAP7_75t_R FILLER_196_626 ();
 DECAPx2_ASAP7_75t_R FILLER_196_662 ();
 FILLER_ASAP7_75t_R FILLER_196_668 ();
 FILLER_ASAP7_75t_R FILLER_196_708 ();
 DECAPx10_ASAP7_75t_R FILLER_196_720 ();
 DECAPx2_ASAP7_75t_R FILLER_196_742 ();
 FILLER_ASAP7_75t_R FILLER_196_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_750 ();
 DECAPx10_ASAP7_75t_R FILLER_196_758 ();
 DECAPx6_ASAP7_75t_R FILLER_196_780 ();
 FILLER_ASAP7_75t_R FILLER_196_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_796 ();
 DECAPx4_ASAP7_75t_R FILLER_196_805 ();
 DECAPx6_ASAP7_75t_R FILLER_196_825 ();
 DECAPx2_ASAP7_75t_R FILLER_196_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_871 ();
 FILLER_ASAP7_75t_R FILLER_196_878 ();
 DECAPx10_ASAP7_75t_R FILLER_196_906 ();
 DECAPx1_ASAP7_75t_R FILLER_196_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_932 ();
 DECAPx6_ASAP7_75t_R FILLER_196_937 ();
 DECAPx10_ASAP7_75t_R FILLER_196_954 ();
 DECAPx4_ASAP7_75t_R FILLER_196_976 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1006 ();
 FILLER_ASAP7_75t_R FILLER_196_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1137 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1159 ();
 FILLER_ASAP7_75t_R FILLER_196_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1182 ();
 FILLER_ASAP7_75t_R FILLER_196_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1196 ();
 FILLER_ASAP7_75t_R FILLER_196_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1212 ();
 FILLER_ASAP7_75t_R FILLER_196_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_197_2 ();
 DECAPx10_ASAP7_75t_R FILLER_197_24 ();
 DECAPx10_ASAP7_75t_R FILLER_197_46 ();
 DECAPx10_ASAP7_75t_R FILLER_197_68 ();
 DECAPx10_ASAP7_75t_R FILLER_197_90 ();
 DECAPx10_ASAP7_75t_R FILLER_197_112 ();
 DECAPx10_ASAP7_75t_R FILLER_197_134 ();
 DECAPx10_ASAP7_75t_R FILLER_197_156 ();
 DECAPx10_ASAP7_75t_R FILLER_197_178 ();
 DECAPx10_ASAP7_75t_R FILLER_197_200 ();
 DECAPx10_ASAP7_75t_R FILLER_197_222 ();
 DECAPx10_ASAP7_75t_R FILLER_197_244 ();
 DECAPx10_ASAP7_75t_R FILLER_197_266 ();
 FILLER_ASAP7_75t_R FILLER_197_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_318 ();
 DECAPx6_ASAP7_75t_R FILLER_197_326 ();
 FILLER_ASAP7_75t_R FILLER_197_340 ();
 FILLER_ASAP7_75t_R FILLER_197_348 ();
 DECAPx6_ASAP7_75t_R FILLER_197_356 ();
 DECAPx1_ASAP7_75t_R FILLER_197_392 ();
 FILLER_ASAP7_75t_R FILLER_197_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_415 ();
 DECAPx4_ASAP7_75t_R FILLER_197_438 ();
 FILLER_ASAP7_75t_R FILLER_197_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_450 ();
 DECAPx2_ASAP7_75t_R FILLER_197_468 ();
 FILLER_ASAP7_75t_R FILLER_197_474 ();
 DECAPx1_ASAP7_75t_R FILLER_197_504 ();
 DECAPx2_ASAP7_75t_R FILLER_197_514 ();
 FILLER_ASAP7_75t_R FILLER_197_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_522 ();
 DECAPx4_ASAP7_75t_R FILLER_197_546 ();
 FILLER_ASAP7_75t_R FILLER_197_556 ();
 DECAPx1_ASAP7_75t_R FILLER_197_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_568 ();
 DECAPx2_ASAP7_75t_R FILLER_197_576 ();
 FILLER_ASAP7_75t_R FILLER_197_582 ();
 FILLER_ASAP7_75t_R FILLER_197_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_603 ();
 DECAPx1_ASAP7_75t_R FILLER_197_632 ();
 DECAPx2_ASAP7_75t_R FILLER_197_642 ();
 DECAPx1_ASAP7_75t_R FILLER_197_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_668 ();
 FILLER_ASAP7_75t_R FILLER_197_689 ();
 FILLER_ASAP7_75t_R FILLER_197_697 ();
 FILLER_ASAP7_75t_R FILLER_197_713 ();
 DECAPx6_ASAP7_75t_R FILLER_197_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_735 ();
 DECAPx1_ASAP7_75t_R FILLER_197_749 ();
 DECAPx2_ASAP7_75t_R FILLER_197_760 ();
 DECAPx6_ASAP7_75t_R FILLER_197_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_822 ();
 DECAPx6_ASAP7_75t_R FILLER_197_833 ();
 DECAPx2_ASAP7_75t_R FILLER_197_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_853 ();
 DECAPx4_ASAP7_75t_R FILLER_197_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_870 ();
 FILLER_ASAP7_75t_R FILLER_197_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_893 ();
 DECAPx1_ASAP7_75t_R FILLER_197_914 ();
 DECAPx6_ASAP7_75t_R FILLER_197_926 ();
 FILLER_ASAP7_75t_R FILLER_197_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_948 ();
 DECAPx10_ASAP7_75t_R FILLER_197_969 ();
 DECAPx10_ASAP7_75t_R FILLER_197_991 ();
 FILLER_ASAP7_75t_R FILLER_197_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1041 ();
 FILLER_ASAP7_75t_R FILLER_197_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1050 ();
 FILLER_ASAP7_75t_R FILLER_197_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1073 ();
 DECAPx6_ASAP7_75t_R FILLER_197_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1120 ();
 DECAPx6_ASAP7_75t_R FILLER_197_1142 ();
 FILLER_ASAP7_75t_R FILLER_197_1156 ();
 DECAPx6_ASAP7_75t_R FILLER_197_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1208 ();
 FILLER_ASAP7_75t_R FILLER_197_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_198_2 ();
 DECAPx10_ASAP7_75t_R FILLER_198_24 ();
 DECAPx10_ASAP7_75t_R FILLER_198_46 ();
 DECAPx10_ASAP7_75t_R FILLER_198_68 ();
 DECAPx10_ASAP7_75t_R FILLER_198_90 ();
 DECAPx10_ASAP7_75t_R FILLER_198_112 ();
 DECAPx10_ASAP7_75t_R FILLER_198_134 ();
 DECAPx10_ASAP7_75t_R FILLER_198_156 ();
 DECAPx10_ASAP7_75t_R FILLER_198_178 ();
 DECAPx10_ASAP7_75t_R FILLER_198_200 ();
 DECAPx10_ASAP7_75t_R FILLER_198_222 ();
 DECAPx10_ASAP7_75t_R FILLER_198_244 ();
 DECAPx10_ASAP7_75t_R FILLER_198_266 ();
 DECAPx6_ASAP7_75t_R FILLER_198_288 ();
 FILLER_ASAP7_75t_R FILLER_198_302 ();
 DECAPx10_ASAP7_75t_R FILLER_198_343 ();
 DECAPx10_ASAP7_75t_R FILLER_198_365 ();
 DECAPx6_ASAP7_75t_R FILLER_198_387 ();
 FILLER_ASAP7_75t_R FILLER_198_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_403 ();
 DECAPx6_ASAP7_75t_R FILLER_198_443 ();
 DECAPx1_ASAP7_75t_R FILLER_198_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_461 ();
 DECAPx4_ASAP7_75t_R FILLER_198_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_474 ();
 DECAPx6_ASAP7_75t_R FILLER_198_486 ();
 FILLER_ASAP7_75t_R FILLER_198_500 ();
 DECAPx10_ASAP7_75t_R FILLER_198_508 ();
 DECAPx10_ASAP7_75t_R FILLER_198_530 ();
 DECAPx2_ASAP7_75t_R FILLER_198_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_558 ();
 DECAPx6_ASAP7_75t_R FILLER_198_578 ();
 FILLER_ASAP7_75t_R FILLER_198_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_594 ();
 DECAPx4_ASAP7_75t_R FILLER_198_623 ();
 FILLER_ASAP7_75t_R FILLER_198_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_635 ();
 FILLER_ASAP7_75t_R FILLER_198_658 ();
 FILLER_ASAP7_75t_R FILLER_198_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_684 ();
 DECAPx2_ASAP7_75t_R FILLER_198_688 ();
 FILLER_ASAP7_75t_R FILLER_198_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_696 ();
 DECAPx1_ASAP7_75t_R FILLER_198_705 ();
 DECAPx1_ASAP7_75t_R FILLER_198_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_740 ();
 FILLER_ASAP7_75t_R FILLER_198_747 ();
 DECAPx1_ASAP7_75t_R FILLER_198_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_759 ();
 DECAPx4_ASAP7_75t_R FILLER_198_772 ();
 FILLER_ASAP7_75t_R FILLER_198_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_803 ();
 FILLER_ASAP7_75t_R FILLER_198_812 ();
 DECAPx6_ASAP7_75t_R FILLER_198_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_846 ();
 DECAPx10_ASAP7_75t_R FILLER_198_867 ();
 FILLER_ASAP7_75t_R FILLER_198_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_891 ();
 DECAPx4_ASAP7_75t_R FILLER_198_898 ();
 FILLER_ASAP7_75t_R FILLER_198_908 ();
 DECAPx2_ASAP7_75t_R FILLER_198_930 ();
 FILLER_ASAP7_75t_R FILLER_198_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_938 ();
 DECAPx10_ASAP7_75t_R FILLER_198_961 ();
 DECAPx2_ASAP7_75t_R FILLER_198_983 ();
 FILLER_ASAP7_75t_R FILLER_198_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_991 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1016 ();
 FILLER_ASAP7_75t_R FILLER_198_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1047 ();
 FILLER_ASAP7_75t_R FILLER_198_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_198_1140 ();
 FILLER_ASAP7_75t_R FILLER_198_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1160 ();
 FILLER_ASAP7_75t_R FILLER_198_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1185 ();
 FILLER_ASAP7_75t_R FILLER_198_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_199_2 ();
 DECAPx10_ASAP7_75t_R FILLER_199_24 ();
 DECAPx10_ASAP7_75t_R FILLER_199_46 ();
 DECAPx10_ASAP7_75t_R FILLER_199_68 ();
 DECAPx10_ASAP7_75t_R FILLER_199_90 ();
 DECAPx10_ASAP7_75t_R FILLER_199_112 ();
 DECAPx10_ASAP7_75t_R FILLER_199_134 ();
 DECAPx10_ASAP7_75t_R FILLER_199_156 ();
 DECAPx10_ASAP7_75t_R FILLER_199_178 ();
 DECAPx10_ASAP7_75t_R FILLER_199_200 ();
 DECAPx10_ASAP7_75t_R FILLER_199_222 ();
 DECAPx10_ASAP7_75t_R FILLER_199_244 ();
 DECAPx10_ASAP7_75t_R FILLER_199_266 ();
 DECAPx10_ASAP7_75t_R FILLER_199_288 ();
 DECAPx4_ASAP7_75t_R FILLER_199_310 ();
 FILLER_ASAP7_75t_R FILLER_199_320 ();
 FILLER_ASAP7_75t_R FILLER_199_336 ();
 DECAPx4_ASAP7_75t_R FILLER_199_344 ();
 FILLER_ASAP7_75t_R FILLER_199_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_356 ();
 DECAPx1_ASAP7_75t_R FILLER_199_367 ();
 DECAPx2_ASAP7_75t_R FILLER_199_403 ();
 DECAPx1_ASAP7_75t_R FILLER_199_426 ();
 DECAPx6_ASAP7_75t_R FILLER_199_438 ();
 DECAPx2_ASAP7_75t_R FILLER_199_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_458 ();
 FILLER_ASAP7_75t_R FILLER_199_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_474 ();
 DECAPx6_ASAP7_75t_R FILLER_199_481 ();
 FILLER_ASAP7_75t_R FILLER_199_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_520 ();
 FILLER_ASAP7_75t_R FILLER_199_549 ();
 FILLER_ASAP7_75t_R FILLER_199_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_583 ();
 DECAPx10_ASAP7_75t_R FILLER_199_590 ();
 DECAPx1_ASAP7_75t_R FILLER_199_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_616 ();
 DECAPx10_ASAP7_75t_R FILLER_199_624 ();
 DECAPx10_ASAP7_75t_R FILLER_199_646 ();
 DECAPx4_ASAP7_75t_R FILLER_199_668 ();
 FILLER_ASAP7_75t_R FILLER_199_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_680 ();
 DECAPx6_ASAP7_75t_R FILLER_199_703 ();
 DECAPx1_ASAP7_75t_R FILLER_199_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_728 ();
 FILLER_ASAP7_75t_R FILLER_199_743 ();
 DECAPx2_ASAP7_75t_R FILLER_199_767 ();
 FILLER_ASAP7_75t_R FILLER_199_783 ();
 DECAPx1_ASAP7_75t_R FILLER_199_792 ();
 DECAPx1_ASAP7_75t_R FILLER_199_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_834 ();
 DECAPx4_ASAP7_75t_R FILLER_199_855 ();
 DECAPx6_ASAP7_75t_R FILLER_199_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_885 ();
 FILLER_ASAP7_75t_R FILLER_199_922 ();
 DECAPx10_ASAP7_75t_R FILLER_199_946 ();
 FILLER_ASAP7_75t_R FILLER_199_971 ();
 FILLER_ASAP7_75t_R FILLER_199_993 ();
 FILLER_ASAP7_75t_R FILLER_199_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1013 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1052 ();
 FILLER_ASAP7_75t_R FILLER_199_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_199_1171 ();
 FILLER_ASAP7_75t_R FILLER_199_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1191 ();
 FILLER_ASAP7_75t_R FILLER_199_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_200_2 ();
 DECAPx10_ASAP7_75t_R FILLER_200_24 ();
 DECAPx10_ASAP7_75t_R FILLER_200_46 ();
 DECAPx10_ASAP7_75t_R FILLER_200_68 ();
 DECAPx10_ASAP7_75t_R FILLER_200_90 ();
 DECAPx10_ASAP7_75t_R FILLER_200_112 ();
 DECAPx10_ASAP7_75t_R FILLER_200_134 ();
 DECAPx10_ASAP7_75t_R FILLER_200_156 ();
 DECAPx10_ASAP7_75t_R FILLER_200_178 ();
 DECAPx10_ASAP7_75t_R FILLER_200_200 ();
 DECAPx10_ASAP7_75t_R FILLER_200_222 ();
 DECAPx10_ASAP7_75t_R FILLER_200_244 ();
 DECAPx10_ASAP7_75t_R FILLER_200_266 ();
 DECAPx4_ASAP7_75t_R FILLER_200_288 ();
 FILLER_ASAP7_75t_R FILLER_200_298 ();
 DECAPx1_ASAP7_75t_R FILLER_200_311 ();
 FILLER_ASAP7_75t_R FILLER_200_327 ();
 DECAPx6_ASAP7_75t_R FILLER_200_357 ();
 FILLER_ASAP7_75t_R FILLER_200_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_373 ();
 DECAPx4_ASAP7_75t_R FILLER_200_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_390 ();
 DECAPx4_ASAP7_75t_R FILLER_200_403 ();
 DECAPx2_ASAP7_75t_R FILLER_200_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_432 ();
 DECAPx2_ASAP7_75t_R FILLER_200_456 ();
 FILLER_ASAP7_75t_R FILLER_200_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_466 ();
 DECAPx10_ASAP7_75t_R FILLER_200_484 ();
 DECAPx6_ASAP7_75t_R FILLER_200_506 ();
 FILLER_ASAP7_75t_R FILLER_200_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_529 ();
 DECAPx10_ASAP7_75t_R FILLER_200_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_565 ();
 DECAPx6_ASAP7_75t_R FILLER_200_601 ();
 FILLER_ASAP7_75t_R FILLER_200_615 ();
 DECAPx2_ASAP7_75t_R FILLER_200_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_635 ();
 FILLER_ASAP7_75t_R FILLER_200_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_651 ();
 DECAPx6_ASAP7_75t_R FILLER_200_656 ();
 FILLER_ASAP7_75t_R FILLER_200_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_672 ();
 DECAPx4_ASAP7_75t_R FILLER_200_717 ();
 FILLER_ASAP7_75t_R FILLER_200_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_743 ();
 DECAPx2_ASAP7_75t_R FILLER_200_750 ();
 FILLER_ASAP7_75t_R FILLER_200_756 ();
 DECAPx6_ASAP7_75t_R FILLER_200_764 ();
 DECAPx2_ASAP7_75t_R FILLER_200_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_784 ();
 FILLER_ASAP7_75t_R FILLER_200_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_814 ();
 FILLER_ASAP7_75t_R FILLER_200_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_829 ();
 DECAPx2_ASAP7_75t_R FILLER_200_837 ();
 FILLER_ASAP7_75t_R FILLER_200_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_845 ();
 DECAPx1_ASAP7_75t_R FILLER_200_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_890 ();
 DECAPx10_ASAP7_75t_R FILLER_200_894 ();
 DECAPx10_ASAP7_75t_R FILLER_200_916 ();
 DECAPx10_ASAP7_75t_R FILLER_200_938 ();
 DECAPx10_ASAP7_75t_R FILLER_200_960 ();
 DECAPx6_ASAP7_75t_R FILLER_200_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_996 ();
 FILLER_ASAP7_75t_R FILLER_200_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1173 ();
 FILLER_ASAP7_75t_R FILLER_200_1179 ();
 FILLER_ASAP7_75t_R FILLER_200_1184 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_201_2 ();
 DECAPx10_ASAP7_75t_R FILLER_201_24 ();
 DECAPx10_ASAP7_75t_R FILLER_201_46 ();
 DECAPx10_ASAP7_75t_R FILLER_201_68 ();
 DECAPx10_ASAP7_75t_R FILLER_201_90 ();
 DECAPx10_ASAP7_75t_R FILLER_201_112 ();
 DECAPx10_ASAP7_75t_R FILLER_201_134 ();
 DECAPx10_ASAP7_75t_R FILLER_201_156 ();
 DECAPx10_ASAP7_75t_R FILLER_201_178 ();
 DECAPx10_ASAP7_75t_R FILLER_201_200 ();
 DECAPx10_ASAP7_75t_R FILLER_201_222 ();
 DECAPx10_ASAP7_75t_R FILLER_201_244 ();
 DECAPx10_ASAP7_75t_R FILLER_201_266 ();
 DECAPx4_ASAP7_75t_R FILLER_201_288 ();
 DECAPx10_ASAP7_75t_R FILLER_201_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_398 ();
 DECAPx2_ASAP7_75t_R FILLER_201_406 ();
 DECAPx4_ASAP7_75t_R FILLER_201_418 ();
 FILLER_ASAP7_75t_R FILLER_201_428 ();
 DECAPx2_ASAP7_75t_R FILLER_201_438 ();
 DECAPx4_ASAP7_75t_R FILLER_201_464 ();
 DECAPx4_ASAP7_75t_R FILLER_201_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_523 ();
 DECAPx10_ASAP7_75t_R FILLER_201_533 ();
 FILLER_ASAP7_75t_R FILLER_201_555 ();
 DECAPx10_ASAP7_75t_R FILLER_201_573 ();
 DECAPx10_ASAP7_75t_R FILLER_201_595 ();
 DECAPx1_ASAP7_75t_R FILLER_201_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_659 ();
 DECAPx4_ASAP7_75t_R FILLER_201_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_680 ();
 DECAPx10_ASAP7_75t_R FILLER_201_687 ();
 DECAPx10_ASAP7_75t_R FILLER_201_709 ();
 FILLER_ASAP7_75t_R FILLER_201_731 ();
 DECAPx6_ASAP7_75t_R FILLER_201_739 ();
 FILLER_ASAP7_75t_R FILLER_201_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_755 ();
 DECAPx2_ASAP7_75t_R FILLER_201_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_782 ();
 FILLER_ASAP7_75t_R FILLER_201_795 ();
 FILLER_ASAP7_75t_R FILLER_201_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_805 ();
 DECAPx1_ASAP7_75t_R FILLER_201_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_816 ();
 DECAPx10_ASAP7_75t_R FILLER_201_836 ();
 DECAPx10_ASAP7_75t_R FILLER_201_858 ();
 DECAPx2_ASAP7_75t_R FILLER_201_880 ();
 FILLER_ASAP7_75t_R FILLER_201_886 ();
 DECAPx4_ASAP7_75t_R FILLER_201_912 ();
 FILLER_ASAP7_75t_R FILLER_201_922 ();
 DECAPx10_ASAP7_75t_R FILLER_201_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_952 ();
 DECAPx10_ASAP7_75t_R FILLER_201_975 ();
 FILLER_ASAP7_75t_R FILLER_201_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_999 ();
 FILLER_ASAP7_75t_R FILLER_201_1006 ();
 FILLER_ASAP7_75t_R FILLER_201_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1041 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1158 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1188 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_202_2 ();
 DECAPx10_ASAP7_75t_R FILLER_202_24 ();
 DECAPx10_ASAP7_75t_R FILLER_202_46 ();
 DECAPx10_ASAP7_75t_R FILLER_202_68 ();
 DECAPx10_ASAP7_75t_R FILLER_202_90 ();
 DECAPx10_ASAP7_75t_R FILLER_202_112 ();
 DECAPx10_ASAP7_75t_R FILLER_202_134 ();
 DECAPx10_ASAP7_75t_R FILLER_202_156 ();
 DECAPx10_ASAP7_75t_R FILLER_202_178 ();
 DECAPx10_ASAP7_75t_R FILLER_202_200 ();
 DECAPx10_ASAP7_75t_R FILLER_202_222 ();
 DECAPx10_ASAP7_75t_R FILLER_202_244 ();
 DECAPx10_ASAP7_75t_R FILLER_202_266 ();
 DECAPx6_ASAP7_75t_R FILLER_202_288 ();
 FILLER_ASAP7_75t_R FILLER_202_302 ();
 DECAPx4_ASAP7_75t_R FILLER_202_310 ();
 DECAPx10_ASAP7_75t_R FILLER_202_337 ();
 DECAPx6_ASAP7_75t_R FILLER_202_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_402 ();
 DECAPx1_ASAP7_75t_R FILLER_202_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_414 ();
 DECAPx6_ASAP7_75t_R FILLER_202_423 ();
 FILLER_ASAP7_75t_R FILLER_202_437 ();
 FILLER_ASAP7_75t_R FILLER_202_447 ();
 DECAPx1_ASAP7_75t_R FILLER_202_458 ();
 DECAPx2_ASAP7_75t_R FILLER_202_464 ();
 FILLER_ASAP7_75t_R FILLER_202_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_472 ();
 DECAPx2_ASAP7_75t_R FILLER_202_488 ();
 FILLER_ASAP7_75t_R FILLER_202_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_516 ();
 FILLER_ASAP7_75t_R FILLER_202_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_525 ();
 DECAPx6_ASAP7_75t_R FILLER_202_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_546 ();
 DECAPx1_ASAP7_75t_R FILLER_202_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_557 ();
 DECAPx4_ASAP7_75t_R FILLER_202_569 ();
 FILLER_ASAP7_75t_R FILLER_202_579 ();
 DECAPx4_ASAP7_75t_R FILLER_202_591 ();
 FILLER_ASAP7_75t_R FILLER_202_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_630 ();
 FILLER_ASAP7_75t_R FILLER_202_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_647 ();
 DECAPx2_ASAP7_75t_R FILLER_202_654 ();
 FILLER_ASAP7_75t_R FILLER_202_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_662 ();
 DECAPx2_ASAP7_75t_R FILLER_202_670 ();
 DECAPx6_ASAP7_75t_R FILLER_202_692 ();
 DECAPx1_ASAP7_75t_R FILLER_202_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_710 ();
 DECAPx2_ASAP7_75t_R FILLER_202_731 ();
 FILLER_ASAP7_75t_R FILLER_202_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_739 ();
 DECAPx4_ASAP7_75t_R FILLER_202_762 ();
 FILLER_ASAP7_75t_R FILLER_202_772 ();
 FILLER_ASAP7_75t_R FILLER_202_795 ();
 DECAPx4_ASAP7_75t_R FILLER_202_800 ();
 FILLER_ASAP7_75t_R FILLER_202_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_812 ();
 DECAPx10_ASAP7_75t_R FILLER_202_827 ();
 DECAPx10_ASAP7_75t_R FILLER_202_849 ();
 DECAPx6_ASAP7_75t_R FILLER_202_871 ();
 FILLER_ASAP7_75t_R FILLER_202_885 ();
 DECAPx4_ASAP7_75t_R FILLER_202_897 ();
 FILLER_ASAP7_75t_R FILLER_202_907 ();
 DECAPx4_ASAP7_75t_R FILLER_202_931 ();
 FILLER_ASAP7_75t_R FILLER_202_941 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_202_1023 ();
 FILLER_ASAP7_75t_R FILLER_202_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1035 ();
 FILLER_ASAP7_75t_R FILLER_202_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1126 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1148 ();
 FILLER_ASAP7_75t_R FILLER_202_1154 ();
 FILLER_ASAP7_75t_R FILLER_202_1164 ();
 FILLER_ASAP7_75t_R FILLER_202_1177 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1187 ();
 FILLER_ASAP7_75t_R FILLER_202_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_203_2 ();
 DECAPx10_ASAP7_75t_R FILLER_203_24 ();
 DECAPx10_ASAP7_75t_R FILLER_203_46 ();
 DECAPx10_ASAP7_75t_R FILLER_203_68 ();
 DECAPx10_ASAP7_75t_R FILLER_203_90 ();
 DECAPx10_ASAP7_75t_R FILLER_203_112 ();
 DECAPx10_ASAP7_75t_R FILLER_203_134 ();
 DECAPx10_ASAP7_75t_R FILLER_203_156 ();
 DECAPx10_ASAP7_75t_R FILLER_203_178 ();
 DECAPx10_ASAP7_75t_R FILLER_203_200 ();
 DECAPx10_ASAP7_75t_R FILLER_203_222 ();
 DECAPx10_ASAP7_75t_R FILLER_203_244 ();
 DECAPx10_ASAP7_75t_R FILLER_203_266 ();
 DECAPx10_ASAP7_75t_R FILLER_203_288 ();
 DECAPx10_ASAP7_75t_R FILLER_203_310 ();
 DECAPx6_ASAP7_75t_R FILLER_203_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_346 ();
 DECAPx6_ASAP7_75t_R FILLER_203_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_396 ();
 DECAPx4_ASAP7_75t_R FILLER_203_404 ();
 DECAPx10_ASAP7_75t_R FILLER_203_448 ();
 FILLER_ASAP7_75t_R FILLER_203_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_472 ();
 DECAPx10_ASAP7_75t_R FILLER_203_489 ();
 DECAPx4_ASAP7_75t_R FILLER_203_511 ();
 FILLER_ASAP7_75t_R FILLER_203_521 ();
 DECAPx2_ASAP7_75t_R FILLER_203_540 ();
 DECAPx4_ASAP7_75t_R FILLER_203_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_578 ();
 DECAPx6_ASAP7_75t_R FILLER_203_599 ();
 FILLER_ASAP7_75t_R FILLER_203_613 ();
 FILLER_ASAP7_75t_R FILLER_203_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_637 ();
 DECAPx2_ASAP7_75t_R FILLER_203_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_663 ();
 DECAPx6_ASAP7_75t_R FILLER_203_674 ();
 DECAPx1_ASAP7_75t_R FILLER_203_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_692 ();
 DECAPx4_ASAP7_75t_R FILLER_203_716 ();
 DECAPx2_ASAP7_75t_R FILLER_203_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_735 ();
 DECAPx10_ASAP7_75t_R FILLER_203_764 ();
 DECAPx4_ASAP7_75t_R FILLER_203_786 ();
 FILLER_ASAP7_75t_R FILLER_203_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_828 ();
 DECAPx1_ASAP7_75t_R FILLER_203_839 ();
 FILLER_ASAP7_75t_R FILLER_203_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_909 ();
 DECAPx2_ASAP7_75t_R FILLER_203_916 ();
 FILLER_ASAP7_75t_R FILLER_203_922 ();
 FILLER_ASAP7_75t_R FILLER_203_926 ();
 DECAPx2_ASAP7_75t_R FILLER_203_934 ();
 DECAPx2_ASAP7_75t_R FILLER_203_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_996 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1058 ();
 DECAPx6_ASAP7_75t_R FILLER_203_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1208 ();
 FILLER_ASAP7_75t_R FILLER_203_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_204_2 ();
 DECAPx10_ASAP7_75t_R FILLER_204_24 ();
 DECAPx10_ASAP7_75t_R FILLER_204_46 ();
 DECAPx10_ASAP7_75t_R FILLER_204_68 ();
 DECAPx10_ASAP7_75t_R FILLER_204_90 ();
 DECAPx10_ASAP7_75t_R FILLER_204_112 ();
 DECAPx10_ASAP7_75t_R FILLER_204_134 ();
 DECAPx10_ASAP7_75t_R FILLER_204_156 ();
 DECAPx10_ASAP7_75t_R FILLER_204_178 ();
 DECAPx10_ASAP7_75t_R FILLER_204_200 ();
 DECAPx10_ASAP7_75t_R FILLER_204_222 ();
 DECAPx10_ASAP7_75t_R FILLER_204_244 ();
 DECAPx10_ASAP7_75t_R FILLER_204_266 ();
 DECAPx10_ASAP7_75t_R FILLER_204_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_310 ();
 DECAPx6_ASAP7_75t_R FILLER_204_317 ();
 DECAPx2_ASAP7_75t_R FILLER_204_331 ();
 FILLER_ASAP7_75t_R FILLER_204_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_362 ();
 DECAPx10_ASAP7_75t_R FILLER_204_375 ();
 DECAPx6_ASAP7_75t_R FILLER_204_397 ();
 DECAPx1_ASAP7_75t_R FILLER_204_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_415 ();
 DECAPx6_ASAP7_75t_R FILLER_204_422 ();
 DECAPx1_ASAP7_75t_R FILLER_204_458 ();
 DECAPx6_ASAP7_75t_R FILLER_204_464 ();
 DECAPx1_ASAP7_75t_R FILLER_204_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_504 ();
 DECAPx1_ASAP7_75t_R FILLER_204_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_553 ();
 FILLER_ASAP7_75t_R FILLER_204_571 ();
 DECAPx4_ASAP7_75t_R FILLER_204_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_591 ();
 DECAPx4_ASAP7_75t_R FILLER_204_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_634 ();
 DECAPx1_ASAP7_75t_R FILLER_204_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_645 ();
 DECAPx6_ASAP7_75t_R FILLER_204_656 ();
 DECAPx2_ASAP7_75t_R FILLER_204_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_676 ();
 DECAPx10_ASAP7_75t_R FILLER_204_715 ();
 DECAPx10_ASAP7_75t_R FILLER_204_737 ();
 DECAPx6_ASAP7_75t_R FILLER_204_759 ();
 FILLER_ASAP7_75t_R FILLER_204_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_797 ();
 DECAPx2_ASAP7_75t_R FILLER_204_804 ();
 FILLER_ASAP7_75t_R FILLER_204_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_812 ();
 FILLER_ASAP7_75t_R FILLER_204_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_834 ();
 DECAPx2_ASAP7_75t_R FILLER_204_841 ();
 DECAPx2_ASAP7_75t_R FILLER_204_856 ();
 FILLER_ASAP7_75t_R FILLER_204_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_864 ();
 DECAPx4_ASAP7_75t_R FILLER_204_888 ();
 FILLER_ASAP7_75t_R FILLER_204_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_900 ();
 FILLER_ASAP7_75t_R FILLER_204_912 ();
 DECAPx1_ASAP7_75t_R FILLER_204_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_963 ();
 DECAPx2_ASAP7_75t_R FILLER_204_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_977 ();
 FILLER_ASAP7_75t_R FILLER_204_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1074 ();
 DECAPx6_ASAP7_75t_R FILLER_204_1096 ();
 FILLER_ASAP7_75t_R FILLER_204_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1182 ();
 FILLER_ASAP7_75t_R FILLER_204_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1208 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_205_2 ();
 DECAPx10_ASAP7_75t_R FILLER_205_24 ();
 DECAPx10_ASAP7_75t_R FILLER_205_46 ();
 DECAPx10_ASAP7_75t_R FILLER_205_68 ();
 DECAPx10_ASAP7_75t_R FILLER_205_90 ();
 DECAPx10_ASAP7_75t_R FILLER_205_112 ();
 DECAPx10_ASAP7_75t_R FILLER_205_134 ();
 DECAPx10_ASAP7_75t_R FILLER_205_156 ();
 DECAPx10_ASAP7_75t_R FILLER_205_178 ();
 DECAPx10_ASAP7_75t_R FILLER_205_200 ();
 DECAPx10_ASAP7_75t_R FILLER_205_222 ();
 DECAPx10_ASAP7_75t_R FILLER_205_244 ();
 DECAPx10_ASAP7_75t_R FILLER_205_266 ();
 DECAPx6_ASAP7_75t_R FILLER_205_288 ();
 DECAPx1_ASAP7_75t_R FILLER_205_302 ();
 DECAPx10_ASAP7_75t_R FILLER_205_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_348 ();
 FILLER_ASAP7_75t_R FILLER_205_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_400 ();
 DECAPx2_ASAP7_75t_R FILLER_205_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_416 ();
 DECAPx10_ASAP7_75t_R FILLER_205_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_461 ();
 DECAPx10_ASAP7_75t_R FILLER_205_472 ();
 DECAPx10_ASAP7_75t_R FILLER_205_494 ();
 DECAPx6_ASAP7_75t_R FILLER_205_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_550 ();
 DECAPx1_ASAP7_75t_R FILLER_205_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_568 ();
 DECAPx10_ASAP7_75t_R FILLER_205_581 ();
 DECAPx6_ASAP7_75t_R FILLER_205_603 ();
 DECAPx1_ASAP7_75t_R FILLER_205_617 ();
 DECAPx4_ASAP7_75t_R FILLER_205_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_651 ();
 DECAPx1_ASAP7_75t_R FILLER_205_672 ();
 FILLER_ASAP7_75t_R FILLER_205_682 ();
 DECAPx10_ASAP7_75t_R FILLER_205_712 ();
 DECAPx6_ASAP7_75t_R FILLER_205_756 ();
 DECAPx1_ASAP7_75t_R FILLER_205_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_774 ();
 DECAPx4_ASAP7_75t_R FILLER_205_801 ();
 FILLER_ASAP7_75t_R FILLER_205_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_827 ();
 DECAPx10_ASAP7_75t_R FILLER_205_834 ();
 DECAPx4_ASAP7_75t_R FILLER_205_856 ();
 FILLER_ASAP7_75t_R FILLER_205_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_868 ();
 DECAPx1_ASAP7_75t_R FILLER_205_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_879 ();
 FILLER_ASAP7_75t_R FILLER_205_895 ();
 DECAPx4_ASAP7_75t_R FILLER_205_912 ();
 FILLER_ASAP7_75t_R FILLER_205_922 ();
 DECAPx6_ASAP7_75t_R FILLER_205_926 ();
 FILLER_ASAP7_75t_R FILLER_205_940 ();
 DECAPx4_ASAP7_75t_R FILLER_205_948 ();
 FILLER_ASAP7_75t_R FILLER_205_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_960 ();
 DECAPx2_ASAP7_75t_R FILLER_205_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_981 ();
 FILLER_ASAP7_75t_R FILLER_205_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_992 ();
 DECAPx10_ASAP7_75t_R FILLER_205_999 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1043 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1090 ();
 FILLER_ASAP7_75t_R FILLER_205_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1114 ();
 DECAPx4_ASAP7_75t_R FILLER_205_1120 ();
 FILLER_ASAP7_75t_R FILLER_205_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1158 ();
 FILLER_ASAP7_75t_R FILLER_205_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1189 ();
 FILLER_ASAP7_75t_R FILLER_205_1193 ();
 DECAPx4_ASAP7_75t_R FILLER_205_1203 ();
 FILLER_ASAP7_75t_R FILLER_205_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_206_2 ();
 DECAPx10_ASAP7_75t_R FILLER_206_24 ();
 DECAPx10_ASAP7_75t_R FILLER_206_46 ();
 DECAPx10_ASAP7_75t_R FILLER_206_68 ();
 DECAPx10_ASAP7_75t_R FILLER_206_90 ();
 DECAPx10_ASAP7_75t_R FILLER_206_112 ();
 DECAPx10_ASAP7_75t_R FILLER_206_134 ();
 DECAPx10_ASAP7_75t_R FILLER_206_156 ();
 DECAPx10_ASAP7_75t_R FILLER_206_178 ();
 DECAPx10_ASAP7_75t_R FILLER_206_200 ();
 DECAPx10_ASAP7_75t_R FILLER_206_222 ();
 DECAPx10_ASAP7_75t_R FILLER_206_244 ();
 DECAPx10_ASAP7_75t_R FILLER_206_266 ();
 DECAPx10_ASAP7_75t_R FILLER_206_288 ();
 DECAPx10_ASAP7_75t_R FILLER_206_310 ();
 DECAPx6_ASAP7_75t_R FILLER_206_332 ();
 DECAPx1_ASAP7_75t_R FILLER_206_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_367 ();
 FILLER_ASAP7_75t_R FILLER_206_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_377 ();
 DECAPx2_ASAP7_75t_R FILLER_206_392 ();
 FILLER_ASAP7_75t_R FILLER_206_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_406 ();
 DECAPx6_ASAP7_75t_R FILLER_206_424 ();
 DECAPx1_ASAP7_75t_R FILLER_206_438 ();
 DECAPx10_ASAP7_75t_R FILLER_206_482 ();
 DECAPx2_ASAP7_75t_R FILLER_206_504 ();
 FILLER_ASAP7_75t_R FILLER_206_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_512 ();
 DECAPx6_ASAP7_75t_R FILLER_206_538 ();
 FILLER_ASAP7_75t_R FILLER_206_552 ();
 FILLER_ASAP7_75t_R FILLER_206_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_573 ();
 DECAPx4_ASAP7_75t_R FILLER_206_596 ();
 FILLER_ASAP7_75t_R FILLER_206_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_641 ();
 DECAPx4_ASAP7_75t_R FILLER_206_666 ();
 FILLER_ASAP7_75t_R FILLER_206_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_711 ();
 FILLER_ASAP7_75t_R FILLER_206_754 ();
 DECAPx2_ASAP7_75t_R FILLER_206_762 ();
 FILLER_ASAP7_75t_R FILLER_206_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_770 ();
 DECAPx6_ASAP7_75t_R FILLER_206_777 ();
 DECAPx6_ASAP7_75t_R FILLER_206_797 ();
 FILLER_ASAP7_75t_R FILLER_206_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_813 ();
 FILLER_ASAP7_75t_R FILLER_206_832 ();
 DECAPx10_ASAP7_75t_R FILLER_206_854 ();
 DECAPx1_ASAP7_75t_R FILLER_206_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_880 ();
 DECAPx2_ASAP7_75t_R FILLER_206_892 ();
 FILLER_ASAP7_75t_R FILLER_206_898 ();
 DECAPx4_ASAP7_75t_R FILLER_206_913 ();
 DECAPx4_ASAP7_75t_R FILLER_206_931 ();
 FILLER_ASAP7_75t_R FILLER_206_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_965 ();
 DECAPx1_ASAP7_75t_R FILLER_206_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_976 ();
 FILLER_ASAP7_75t_R FILLER_206_983 ();
 DECAPx1_ASAP7_75t_R FILLER_206_992 ();
 FILLER_ASAP7_75t_R FILLER_206_1003 ();
 FILLER_ASAP7_75t_R FILLER_206_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1143 ();
 DECAPx6_ASAP7_75t_R FILLER_206_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1179 ();
 FILLER_ASAP7_75t_R FILLER_206_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_207_2 ();
 DECAPx10_ASAP7_75t_R FILLER_207_24 ();
 DECAPx10_ASAP7_75t_R FILLER_207_46 ();
 DECAPx10_ASAP7_75t_R FILLER_207_68 ();
 DECAPx10_ASAP7_75t_R FILLER_207_90 ();
 DECAPx10_ASAP7_75t_R FILLER_207_112 ();
 DECAPx10_ASAP7_75t_R FILLER_207_134 ();
 DECAPx10_ASAP7_75t_R FILLER_207_156 ();
 DECAPx10_ASAP7_75t_R FILLER_207_178 ();
 DECAPx10_ASAP7_75t_R FILLER_207_200 ();
 DECAPx10_ASAP7_75t_R FILLER_207_222 ();
 DECAPx10_ASAP7_75t_R FILLER_207_244 ();
 DECAPx10_ASAP7_75t_R FILLER_207_266 ();
 DECAPx10_ASAP7_75t_R FILLER_207_288 ();
 DECAPx1_ASAP7_75t_R FILLER_207_310 ();
 DECAPx6_ASAP7_75t_R FILLER_207_326 ();
 DECAPx2_ASAP7_75t_R FILLER_207_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_346 ();
 DECAPx1_ASAP7_75t_R FILLER_207_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_379 ();
 DECAPx4_ASAP7_75t_R FILLER_207_392 ();
 DECAPx10_ASAP7_75t_R FILLER_207_409 ();
 FILLER_ASAP7_75t_R FILLER_207_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_433 ();
 DECAPx1_ASAP7_75t_R FILLER_207_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_474 ();
 DECAPx2_ASAP7_75t_R FILLER_207_503 ();
 FILLER_ASAP7_75t_R FILLER_207_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_511 ();
 FILLER_ASAP7_75t_R FILLER_207_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_530 ();
 DECAPx4_ASAP7_75t_R FILLER_207_553 ();
 FILLER_ASAP7_75t_R FILLER_207_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_565 ();
 DECAPx4_ASAP7_75t_R FILLER_207_596 ();
 FILLER_ASAP7_75t_R FILLER_207_606 ();
 DECAPx4_ASAP7_75t_R FILLER_207_614 ();
 FILLER_ASAP7_75t_R FILLER_207_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_626 ();
 FILLER_ASAP7_75t_R FILLER_207_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_635 ();
 DECAPx2_ASAP7_75t_R FILLER_207_642 ();
 DECAPx4_ASAP7_75t_R FILLER_207_668 ();
 FILLER_ASAP7_75t_R FILLER_207_678 ();
 DECAPx10_ASAP7_75t_R FILLER_207_686 ();
 DECAPx10_ASAP7_75t_R FILLER_207_708 ();
 DECAPx6_ASAP7_75t_R FILLER_207_730 ();
 FILLER_ASAP7_75t_R FILLER_207_744 ();
 FILLER_ASAP7_75t_R FILLER_207_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_754 ();
 DECAPx2_ASAP7_75t_R FILLER_207_781 ();
 FILLER_ASAP7_75t_R FILLER_207_787 ();
 DECAPx6_ASAP7_75t_R FILLER_207_811 ();
 FILLER_ASAP7_75t_R FILLER_207_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_827 ();
 DECAPx1_ASAP7_75t_R FILLER_207_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_844 ();
 DECAPx6_ASAP7_75t_R FILLER_207_851 ();
 DECAPx2_ASAP7_75t_R FILLER_207_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_871 ();
 FILLER_ASAP7_75t_R FILLER_207_894 ();
 DECAPx1_ASAP7_75t_R FILLER_207_932 ();
 DECAPx6_ASAP7_75t_R FILLER_207_942 ();
 DECAPx1_ASAP7_75t_R FILLER_207_956 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1061 ();
 DECAPx4_ASAP7_75t_R FILLER_207_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1201 ();
 FILLER_ASAP7_75t_R FILLER_207_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_208_2 ();
 DECAPx10_ASAP7_75t_R FILLER_208_24 ();
 DECAPx10_ASAP7_75t_R FILLER_208_46 ();
 DECAPx10_ASAP7_75t_R FILLER_208_68 ();
 DECAPx10_ASAP7_75t_R FILLER_208_90 ();
 DECAPx10_ASAP7_75t_R FILLER_208_112 ();
 DECAPx10_ASAP7_75t_R FILLER_208_134 ();
 DECAPx10_ASAP7_75t_R FILLER_208_156 ();
 DECAPx10_ASAP7_75t_R FILLER_208_178 ();
 DECAPx10_ASAP7_75t_R FILLER_208_200 ();
 DECAPx10_ASAP7_75t_R FILLER_208_222 ();
 DECAPx10_ASAP7_75t_R FILLER_208_244 ();
 DECAPx10_ASAP7_75t_R FILLER_208_266 ();
 DECAPx1_ASAP7_75t_R FILLER_208_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_292 ();
 FILLER_ASAP7_75t_R FILLER_208_315 ();
 DECAPx10_ASAP7_75t_R FILLER_208_320 ();
 FILLER_ASAP7_75t_R FILLER_208_342 ();
 DECAPx4_ASAP7_75t_R FILLER_208_388 ();
 FILLER_ASAP7_75t_R FILLER_208_398 ();
 FILLER_ASAP7_75t_R FILLER_208_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_470 ();
 DECAPx4_ASAP7_75t_R FILLER_208_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_503 ();
 FILLER_ASAP7_75t_R FILLER_208_521 ();
 DECAPx2_ASAP7_75t_R FILLER_208_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_542 ();
 FILLER_ASAP7_75t_R FILLER_208_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_556 ();
 DECAPx6_ASAP7_75t_R FILLER_208_568 ();
 FILLER_ASAP7_75t_R FILLER_208_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_584 ();
 DECAPx4_ASAP7_75t_R FILLER_208_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_625 ();
 DECAPx6_ASAP7_75t_R FILLER_208_632 ();
 DECAPx2_ASAP7_75t_R FILLER_208_646 ();
 DECAPx2_ASAP7_75t_R FILLER_208_673 ();
 DECAPx10_ASAP7_75t_R FILLER_208_691 ();
 DECAPx2_ASAP7_75t_R FILLER_208_713 ();
 FILLER_ASAP7_75t_R FILLER_208_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_721 ();
 DECAPx2_ASAP7_75t_R FILLER_208_744 ();
 FILLER_ASAP7_75t_R FILLER_208_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_773 ();
 DECAPx4_ASAP7_75t_R FILLER_208_780 ();
 FILLER_ASAP7_75t_R FILLER_208_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_815 ();
 DECAPx1_ASAP7_75t_R FILLER_208_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_827 ();
 DECAPx6_ASAP7_75t_R FILLER_208_850 ();
 FILLER_ASAP7_75t_R FILLER_208_864 ();
 DECAPx2_ASAP7_75t_R FILLER_208_892 ();
 FILLER_ASAP7_75t_R FILLER_208_898 ();
 FILLER_ASAP7_75t_R FILLER_208_918 ();
 DECAPx6_ASAP7_75t_R FILLER_208_942 ();
 DECAPx1_ASAP7_75t_R FILLER_208_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_960 ();
 DECAPx6_ASAP7_75t_R FILLER_208_968 ();
 DECAPx2_ASAP7_75t_R FILLER_208_982 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1162 ();
 DECAPx4_ASAP7_75t_R FILLER_208_1184 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1200 ();
 FILLER_ASAP7_75t_R FILLER_208_1214 ();
 FILLER_ASAP7_75t_R FILLER_208_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_209_2 ();
 DECAPx10_ASAP7_75t_R FILLER_209_24 ();
 DECAPx10_ASAP7_75t_R FILLER_209_46 ();
 DECAPx10_ASAP7_75t_R FILLER_209_68 ();
 DECAPx10_ASAP7_75t_R FILLER_209_90 ();
 DECAPx10_ASAP7_75t_R FILLER_209_112 ();
 DECAPx10_ASAP7_75t_R FILLER_209_134 ();
 DECAPx10_ASAP7_75t_R FILLER_209_156 ();
 DECAPx10_ASAP7_75t_R FILLER_209_178 ();
 DECAPx10_ASAP7_75t_R FILLER_209_200 ();
 DECAPx10_ASAP7_75t_R FILLER_209_222 ();
 DECAPx10_ASAP7_75t_R FILLER_209_244 ();
 DECAPx10_ASAP7_75t_R FILLER_209_266 ();
 DECAPx2_ASAP7_75t_R FILLER_209_288 ();
 FILLER_ASAP7_75t_R FILLER_209_294 ();
 DECAPx1_ASAP7_75t_R FILLER_209_302 ();
 DECAPx2_ASAP7_75t_R FILLER_209_323 ();
 FILLER_ASAP7_75t_R FILLER_209_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_331 ();
 DECAPx10_ASAP7_75t_R FILLER_209_338 ();
 DECAPx6_ASAP7_75t_R FILLER_209_377 ();
 DECAPx2_ASAP7_75t_R FILLER_209_391 ();
 FILLER_ASAP7_75t_R FILLER_209_408 ();
 DECAPx10_ASAP7_75t_R FILLER_209_416 ();
 DECAPx10_ASAP7_75t_R FILLER_209_438 ();
 DECAPx6_ASAP7_75t_R FILLER_209_477 ();
 DECAPx1_ASAP7_75t_R FILLER_209_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_495 ();
 DECAPx10_ASAP7_75t_R FILLER_209_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_540 ();
 DECAPx2_ASAP7_75t_R FILLER_209_591 ();
 FILLER_ASAP7_75t_R FILLER_209_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_641 ();
 DECAPx10_ASAP7_75t_R FILLER_209_654 ();
 FILLER_ASAP7_75t_R FILLER_209_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_678 ();
 DECAPx4_ASAP7_75t_R FILLER_209_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_701 ();
 DECAPx2_ASAP7_75t_R FILLER_209_735 ();
 FILLER_ASAP7_75t_R FILLER_209_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_743 ();
 DECAPx1_ASAP7_75t_R FILLER_209_750 ();
 DECAPx6_ASAP7_75t_R FILLER_209_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_774 ();
 DECAPx6_ASAP7_75t_R FILLER_209_795 ();
 FILLER_ASAP7_75t_R FILLER_209_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_824 ();
 FILLER_ASAP7_75t_R FILLER_209_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_876 ();
 DECAPx6_ASAP7_75t_R FILLER_209_904 ();
 DECAPx2_ASAP7_75t_R FILLER_209_918 ();
 DECAPx2_ASAP7_75t_R FILLER_209_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_943 ();
 DECAPx2_ASAP7_75t_R FILLER_209_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_968 ();
 DECAPx4_ASAP7_75t_R FILLER_209_975 ();
 FILLER_ASAP7_75t_R FILLER_209_985 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_209_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1121 ();
 DECAPx4_ASAP7_75t_R FILLER_209_1143 ();
 FILLER_ASAP7_75t_R FILLER_209_1153 ();
 FILLER_ASAP7_75t_R FILLER_209_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1165 ();
 FILLER_ASAP7_75t_R FILLER_209_1187 ();
 FILLER_ASAP7_75t_R FILLER_209_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1199 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_209_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_210_2 ();
 DECAPx10_ASAP7_75t_R FILLER_210_24 ();
 DECAPx10_ASAP7_75t_R FILLER_210_46 ();
 DECAPx10_ASAP7_75t_R FILLER_210_68 ();
 DECAPx10_ASAP7_75t_R FILLER_210_90 ();
 DECAPx10_ASAP7_75t_R FILLER_210_112 ();
 DECAPx10_ASAP7_75t_R FILLER_210_134 ();
 DECAPx10_ASAP7_75t_R FILLER_210_156 ();
 DECAPx10_ASAP7_75t_R FILLER_210_178 ();
 DECAPx10_ASAP7_75t_R FILLER_210_200 ();
 DECAPx10_ASAP7_75t_R FILLER_210_222 ();
 DECAPx10_ASAP7_75t_R FILLER_210_244 ();
 DECAPx10_ASAP7_75t_R FILLER_210_266 ();
 DECAPx2_ASAP7_75t_R FILLER_210_288 ();
 FILLER_ASAP7_75t_R FILLER_210_294 ();
 FILLER_ASAP7_75t_R FILLER_210_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_304 ();
 FILLER_ASAP7_75t_R FILLER_210_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_318 ();
 FILLER_ASAP7_75t_R FILLER_210_328 ();
 DECAPx4_ASAP7_75t_R FILLER_210_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_369 ();
 DECAPx6_ASAP7_75t_R FILLER_210_406 ();
 FILLER_ASAP7_75t_R FILLER_210_420 ();
 DECAPx2_ASAP7_75t_R FILLER_210_442 ();
 FILLER_ASAP7_75t_R FILLER_210_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_450 ();
 DECAPx1_ASAP7_75t_R FILLER_210_458 ();
 DECAPx10_ASAP7_75t_R FILLER_210_464 ();
 DECAPx6_ASAP7_75t_R FILLER_210_486 ();
 FILLER_ASAP7_75t_R FILLER_210_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_502 ();
 DECAPx2_ASAP7_75t_R FILLER_210_509 ();
 DECAPx10_ASAP7_75t_R FILLER_210_526 ();
 DECAPx6_ASAP7_75t_R FILLER_210_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_562 ();
 DECAPx4_ASAP7_75t_R FILLER_210_569 ();
 FILLER_ASAP7_75t_R FILLER_210_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_581 ();
 DECAPx4_ASAP7_75t_R FILLER_210_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_631 ();
 FILLER_ASAP7_75t_R FILLER_210_653 ();
 FILLER_ASAP7_75t_R FILLER_210_675 ();
 DECAPx10_ASAP7_75t_R FILLER_210_701 ();
 DECAPx1_ASAP7_75t_R FILLER_210_723 ();
 FILLER_ASAP7_75t_R FILLER_210_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_751 ();
 DECAPx6_ASAP7_75t_R FILLER_210_758 ();
 FILLER_ASAP7_75t_R FILLER_210_772 ();
 FILLER_ASAP7_75t_R FILLER_210_794 ();
 DECAPx4_ASAP7_75t_R FILLER_210_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_839 ();
 DECAPx10_ASAP7_75t_R FILLER_210_843 ();
 DECAPx4_ASAP7_75t_R FILLER_210_865 ();
 FILLER_ASAP7_75t_R FILLER_210_875 ();
 DECAPx1_ASAP7_75t_R FILLER_210_880 ();
 DECAPx2_ASAP7_75t_R FILLER_210_888 ();
 FILLER_ASAP7_75t_R FILLER_210_894 ();
 DECAPx4_ASAP7_75t_R FILLER_210_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_912 ();
 DECAPx1_ASAP7_75t_R FILLER_210_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_943 ();
 DECAPx1_ASAP7_75t_R FILLER_210_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_968 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1213 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_211_2 ();
 DECAPx10_ASAP7_75t_R FILLER_211_24 ();
 DECAPx10_ASAP7_75t_R FILLER_211_46 ();
 DECAPx10_ASAP7_75t_R FILLER_211_68 ();
 DECAPx10_ASAP7_75t_R FILLER_211_90 ();
 DECAPx10_ASAP7_75t_R FILLER_211_112 ();
 DECAPx10_ASAP7_75t_R FILLER_211_134 ();
 DECAPx10_ASAP7_75t_R FILLER_211_156 ();
 DECAPx10_ASAP7_75t_R FILLER_211_178 ();
 DECAPx10_ASAP7_75t_R FILLER_211_200 ();
 DECAPx10_ASAP7_75t_R FILLER_211_222 ();
 DECAPx10_ASAP7_75t_R FILLER_211_244 ();
 DECAPx10_ASAP7_75t_R FILLER_211_266 ();
 DECAPx1_ASAP7_75t_R FILLER_211_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_292 ();
 FILLER_ASAP7_75t_R FILLER_211_315 ();
 FILLER_ASAP7_75t_R FILLER_211_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_326 ();
 FILLER_ASAP7_75t_R FILLER_211_359 ();
 DECAPx4_ASAP7_75t_R FILLER_211_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_399 ();
 DECAPx6_ASAP7_75t_R FILLER_211_411 ();
 FILLER_ASAP7_75t_R FILLER_211_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_427 ();
 DECAPx2_ASAP7_75t_R FILLER_211_445 ();
 FILLER_ASAP7_75t_R FILLER_211_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_461 ();
 DECAPx4_ASAP7_75t_R FILLER_211_468 ();
 DECAPx6_ASAP7_75t_R FILLER_211_500 ();
 DECAPx2_ASAP7_75t_R FILLER_211_514 ();
 DECAPx10_ASAP7_75t_R FILLER_211_542 ();
 DECAPx6_ASAP7_75t_R FILLER_211_564 ();
 FILLER_ASAP7_75t_R FILLER_211_578 ();
 DECAPx10_ASAP7_75t_R FILLER_211_616 ();
 DECAPx4_ASAP7_75t_R FILLER_211_677 ();
 DECAPx4_ASAP7_75t_R FILLER_211_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_721 ();
 DECAPx2_ASAP7_75t_R FILLER_211_744 ();
 FILLER_ASAP7_75t_R FILLER_211_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_752 ();
 FILLER_ASAP7_75t_R FILLER_211_773 ();
 DECAPx6_ASAP7_75t_R FILLER_211_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_795 ();
 DECAPx2_ASAP7_75t_R FILLER_211_802 ();
 FILLER_ASAP7_75t_R FILLER_211_808 ();
 DECAPx4_ASAP7_75t_R FILLER_211_818 ();
 FILLER_ASAP7_75t_R FILLER_211_828 ();
 DECAPx10_ASAP7_75t_R FILLER_211_850 ();
 DECAPx4_ASAP7_75t_R FILLER_211_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_882 ();
 FILLER_ASAP7_75t_R FILLER_211_893 ();
 DECAPx2_ASAP7_75t_R FILLER_211_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_923 ();
 DECAPx2_ASAP7_75t_R FILLER_211_926 ();
 FILLER_ASAP7_75t_R FILLER_211_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_934 ();
 DECAPx6_ASAP7_75t_R FILLER_211_941 ();
 DECAPx1_ASAP7_75t_R FILLER_211_955 ();
 DECAPx6_ASAP7_75t_R FILLER_211_967 ();
 FILLER_ASAP7_75t_R FILLER_211_996 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1005 ();
 FILLER_ASAP7_75t_R FILLER_211_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1202 ();
 FILLER_ASAP7_75t_R FILLER_211_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_212_2 ();
 DECAPx10_ASAP7_75t_R FILLER_212_24 ();
 DECAPx10_ASAP7_75t_R FILLER_212_46 ();
 DECAPx10_ASAP7_75t_R FILLER_212_68 ();
 DECAPx10_ASAP7_75t_R FILLER_212_90 ();
 DECAPx10_ASAP7_75t_R FILLER_212_112 ();
 DECAPx10_ASAP7_75t_R FILLER_212_134 ();
 DECAPx10_ASAP7_75t_R FILLER_212_156 ();
 DECAPx10_ASAP7_75t_R FILLER_212_178 ();
 DECAPx10_ASAP7_75t_R FILLER_212_200 ();
 DECAPx10_ASAP7_75t_R FILLER_212_222 ();
 DECAPx10_ASAP7_75t_R FILLER_212_244 ();
 DECAPx10_ASAP7_75t_R FILLER_212_266 ();
 DECAPx10_ASAP7_75t_R FILLER_212_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_310 ();
 DECAPx6_ASAP7_75t_R FILLER_212_335 ();
 FILLER_ASAP7_75t_R FILLER_212_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_351 ();
 DECAPx6_ASAP7_75t_R FILLER_212_362 ();
 DECAPx2_ASAP7_75t_R FILLER_212_376 ();
 DECAPx4_ASAP7_75t_R FILLER_212_392 ();
 FILLER_ASAP7_75t_R FILLER_212_402 ();
 DECAPx6_ASAP7_75t_R FILLER_212_410 ();
 DECAPx1_ASAP7_75t_R FILLER_212_424 ();
 FILLER_ASAP7_75t_R FILLER_212_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_436 ();
 DECAPx2_ASAP7_75t_R FILLER_212_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_461 ();
 FILLER_ASAP7_75t_R FILLER_212_464 ();
 DECAPx4_ASAP7_75t_R FILLER_212_483 ();
 FILLER_ASAP7_75t_R FILLER_212_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_495 ();
 DECAPx1_ASAP7_75t_R FILLER_212_518 ();
 DECAPx10_ASAP7_75t_R FILLER_212_528 ();
 FILLER_ASAP7_75t_R FILLER_212_550 ();
 DECAPx10_ASAP7_75t_R FILLER_212_558 ();
 DECAPx10_ASAP7_75t_R FILLER_212_580 ();
 DECAPx6_ASAP7_75t_R FILLER_212_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_639 ();
 DECAPx10_ASAP7_75t_R FILLER_212_652 ();
 DECAPx4_ASAP7_75t_R FILLER_212_674 ();
 DECAPx4_ASAP7_75t_R FILLER_212_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_752 ();
 DECAPx4_ASAP7_75t_R FILLER_212_759 ();
 FILLER_ASAP7_75t_R FILLER_212_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_771 ();
 DECAPx2_ASAP7_75t_R FILLER_212_778 ();
 FILLER_ASAP7_75t_R FILLER_212_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_786 ();
 DECAPx2_ASAP7_75t_R FILLER_212_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_818 ();
 DECAPx10_ASAP7_75t_R FILLER_212_839 ();
 DECAPx10_ASAP7_75t_R FILLER_212_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_883 ();
 DECAPx4_ASAP7_75t_R FILLER_212_894 ();
 FILLER_ASAP7_75t_R FILLER_212_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_906 ();
 DECAPx1_ASAP7_75t_R FILLER_212_919 ();
 DECAPx2_ASAP7_75t_R FILLER_212_930 ();
 DECAPx10_ASAP7_75t_R FILLER_212_958 ();
 DECAPx2_ASAP7_75t_R FILLER_212_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_986 ();
 DECAPx2_ASAP7_75t_R FILLER_212_994 ();
 FILLER_ASAP7_75t_R FILLER_212_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1171 ();
 DECAPx4_ASAP7_75t_R FILLER_212_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1214 ();
 FILLER_ASAP7_75t_R FILLER_212_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_213_2 ();
 DECAPx10_ASAP7_75t_R FILLER_213_24 ();
 DECAPx10_ASAP7_75t_R FILLER_213_46 ();
 DECAPx10_ASAP7_75t_R FILLER_213_68 ();
 DECAPx10_ASAP7_75t_R FILLER_213_90 ();
 DECAPx10_ASAP7_75t_R FILLER_213_112 ();
 DECAPx10_ASAP7_75t_R FILLER_213_134 ();
 DECAPx10_ASAP7_75t_R FILLER_213_156 ();
 DECAPx10_ASAP7_75t_R FILLER_213_178 ();
 DECAPx10_ASAP7_75t_R FILLER_213_200 ();
 DECAPx10_ASAP7_75t_R FILLER_213_222 ();
 DECAPx10_ASAP7_75t_R FILLER_213_244 ();
 DECAPx10_ASAP7_75t_R FILLER_213_266 ();
 DECAPx10_ASAP7_75t_R FILLER_213_288 ();
 DECAPx10_ASAP7_75t_R FILLER_213_310 ();
 DECAPx10_ASAP7_75t_R FILLER_213_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_354 ();
 DECAPx1_ASAP7_75t_R FILLER_213_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_446 ();
 DECAPx2_ASAP7_75t_R FILLER_213_455 ();
 DECAPx10_ASAP7_75t_R FILLER_213_478 ();
 DECAPx4_ASAP7_75t_R FILLER_213_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_516 ();
 DECAPx1_ASAP7_75t_R FILLER_213_568 ();
 DECAPx6_ASAP7_75t_R FILLER_213_594 ();
 FILLER_ASAP7_75t_R FILLER_213_608 ();
 DECAPx6_ASAP7_75t_R FILLER_213_622 ();
 DECAPx1_ASAP7_75t_R FILLER_213_636 ();
 DECAPx2_ASAP7_75t_R FILLER_213_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_675 ();
 DECAPx10_ASAP7_75t_R FILLER_213_696 ();
 DECAPx10_ASAP7_75t_R FILLER_213_718 ();
 FILLER_ASAP7_75t_R FILLER_213_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_742 ();
 FILLER_ASAP7_75t_R FILLER_213_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_751 ();
 FILLER_ASAP7_75t_R FILLER_213_772 ();
 FILLER_ASAP7_75t_R FILLER_213_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_798 ();
 DECAPx6_ASAP7_75t_R FILLER_213_819 ();
 FILLER_ASAP7_75t_R FILLER_213_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_835 ();
 DECAPx4_ASAP7_75t_R FILLER_213_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_849 ();
 FILLER_ASAP7_75t_R FILLER_213_853 ();
 DECAPx2_ASAP7_75t_R FILLER_213_891 ();
 FILLER_ASAP7_75t_R FILLER_213_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_899 ();
 DECAPx2_ASAP7_75t_R FILLER_213_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_912 ();
 DECAPx1_ASAP7_75t_R FILLER_213_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_923 ();
 DECAPx6_ASAP7_75t_R FILLER_213_933 ();
 FILLER_ASAP7_75t_R FILLER_213_947 ();
 DECAPx1_ASAP7_75t_R FILLER_213_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_989 ();
 DECAPx2_ASAP7_75t_R FILLER_213_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1075 ();
 DECAPx6_ASAP7_75t_R FILLER_213_1097 ();
 DECAPx1_ASAP7_75t_R FILLER_213_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_213_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1211 ();
 FILLER_ASAP7_75t_R FILLER_213_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_214_2 ();
 DECAPx10_ASAP7_75t_R FILLER_214_24 ();
 DECAPx10_ASAP7_75t_R FILLER_214_46 ();
 DECAPx10_ASAP7_75t_R FILLER_214_68 ();
 DECAPx10_ASAP7_75t_R FILLER_214_90 ();
 DECAPx10_ASAP7_75t_R FILLER_214_112 ();
 DECAPx10_ASAP7_75t_R FILLER_214_134 ();
 DECAPx10_ASAP7_75t_R FILLER_214_156 ();
 DECAPx10_ASAP7_75t_R FILLER_214_178 ();
 DECAPx10_ASAP7_75t_R FILLER_214_200 ();
 DECAPx10_ASAP7_75t_R FILLER_214_222 ();
 DECAPx10_ASAP7_75t_R FILLER_214_244 ();
 DECAPx10_ASAP7_75t_R FILLER_214_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_288 ();
 FILLER_ASAP7_75t_R FILLER_214_295 ();
 FILLER_ASAP7_75t_R FILLER_214_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_310 ();
 FILLER_ASAP7_75t_R FILLER_214_319 ();
 DECAPx1_ASAP7_75t_R FILLER_214_327 ();
 DECAPx2_ASAP7_75t_R FILLER_214_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_346 ();
 DECAPx2_ASAP7_75t_R FILLER_214_375 ();
 DECAPx10_ASAP7_75t_R FILLER_214_418 ();
 FILLER_ASAP7_75t_R FILLER_214_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_442 ();
 DECAPx2_ASAP7_75t_R FILLER_214_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_461 ();
 DECAPx2_ASAP7_75t_R FILLER_214_464 ();
 FILLER_ASAP7_75t_R FILLER_214_470 ();
 DECAPx4_ASAP7_75t_R FILLER_214_494 ();
 FILLER_ASAP7_75t_R FILLER_214_504 ();
 DECAPx10_ASAP7_75t_R FILLER_214_512 ();
 DECAPx6_ASAP7_75t_R FILLER_214_534 ();
 FILLER_ASAP7_75t_R FILLER_214_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_571 ();
 DECAPx6_ASAP7_75t_R FILLER_214_578 ();
 DECAPx1_ASAP7_75t_R FILLER_214_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_596 ();
 DECAPx1_ASAP7_75t_R FILLER_214_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_621 ();
 DECAPx10_ASAP7_75t_R FILLER_214_642 ();
 DECAPx2_ASAP7_75t_R FILLER_214_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_692 ();
 DECAPx10_ASAP7_75t_R FILLER_214_697 ();
 DECAPx1_ASAP7_75t_R FILLER_214_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_723 ();
 FILLER_ASAP7_75t_R FILLER_214_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_751 ();
 DECAPx4_ASAP7_75t_R FILLER_214_764 ();
 DECAPx10_ASAP7_75t_R FILLER_214_780 ();
 DECAPx6_ASAP7_75t_R FILLER_214_802 ();
 DECAPx1_ASAP7_75t_R FILLER_214_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_820 ();
 FILLER_ASAP7_75t_R FILLER_214_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_836 ();
 DECAPx6_ASAP7_75t_R FILLER_214_860 ();
 DECAPx1_ASAP7_75t_R FILLER_214_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_878 ();
 DECAPx1_ASAP7_75t_R FILLER_214_890 ();
 DECAPx2_ASAP7_75t_R FILLER_214_908 ();
 DECAPx6_ASAP7_75t_R FILLER_214_934 ();
 FILLER_ASAP7_75t_R FILLER_214_948 ();
 DECAPx6_ASAP7_75t_R FILLER_214_956 ();
 FILLER_ASAP7_75t_R FILLER_214_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_972 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_214_1187 ();
 FILLER_ASAP7_75t_R FILLER_214_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1209 ();
 FILLER_ASAP7_75t_R FILLER_214_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_215_2 ();
 DECAPx10_ASAP7_75t_R FILLER_215_24 ();
 DECAPx10_ASAP7_75t_R FILLER_215_46 ();
 DECAPx10_ASAP7_75t_R FILLER_215_68 ();
 DECAPx10_ASAP7_75t_R FILLER_215_90 ();
 DECAPx10_ASAP7_75t_R FILLER_215_112 ();
 DECAPx10_ASAP7_75t_R FILLER_215_134 ();
 DECAPx10_ASAP7_75t_R FILLER_215_156 ();
 DECAPx10_ASAP7_75t_R FILLER_215_178 ();
 DECAPx10_ASAP7_75t_R FILLER_215_200 ();
 DECAPx10_ASAP7_75t_R FILLER_215_222 ();
 DECAPx10_ASAP7_75t_R FILLER_215_244 ();
 DECAPx6_ASAP7_75t_R FILLER_215_266 ();
 FILLER_ASAP7_75t_R FILLER_215_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_325 ();
 DECAPx1_ASAP7_75t_R FILLER_215_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_344 ();
 DECAPx4_ASAP7_75t_R FILLER_215_351 ();
 FILLER_ASAP7_75t_R FILLER_215_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_363 ();
 DECAPx6_ASAP7_75t_R FILLER_215_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_392 ();
 DECAPx10_ASAP7_75t_R FILLER_215_421 ();
 FILLER_ASAP7_75t_R FILLER_215_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_445 ();
 FILLER_ASAP7_75t_R FILLER_215_468 ();
 FILLER_ASAP7_75t_R FILLER_215_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_488 ();
 DECAPx1_ASAP7_75t_R FILLER_215_523 ();
 DECAPx2_ASAP7_75t_R FILLER_215_537 ();
 FILLER_ASAP7_75t_R FILLER_215_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_545 ();
 DECAPx2_ASAP7_75t_R FILLER_215_555 ();
 DECAPx1_ASAP7_75t_R FILLER_215_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_571 ();
 DECAPx2_ASAP7_75t_R FILLER_215_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_600 ();
 FILLER_ASAP7_75t_R FILLER_215_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_639 ();
 DECAPx2_ASAP7_75t_R FILLER_215_643 ();
 FILLER_ASAP7_75t_R FILLER_215_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_677 ();
 DECAPx10_ASAP7_75t_R FILLER_215_699 ();
 DECAPx1_ASAP7_75t_R FILLER_215_721 ();
 DECAPx2_ASAP7_75t_R FILLER_215_747 ();
 FILLER_ASAP7_75t_R FILLER_215_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_755 ();
 FILLER_ASAP7_75t_R FILLER_215_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_764 ();
 FILLER_ASAP7_75t_R FILLER_215_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_817 ();
 FILLER_ASAP7_75t_R FILLER_215_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_823 ();
 DECAPx10_ASAP7_75t_R FILLER_215_848 ();
 DECAPx1_ASAP7_75t_R FILLER_215_870 ();
 DECAPx2_ASAP7_75t_R FILLER_215_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_926 ();
 DECAPx6_ASAP7_75t_R FILLER_215_955 ();
 FILLER_ASAP7_75t_R FILLER_215_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_971 ();
 DECAPx4_ASAP7_75t_R FILLER_215_979 ();
 FILLER_ASAP7_75t_R FILLER_215_989 ();
 DECAPx1_ASAP7_75t_R FILLER_215_997 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1150 ();
 DECAPx6_ASAP7_75t_R FILLER_215_1172 ();
 DECAPx1_ASAP7_75t_R FILLER_215_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1190 ();
 FILLER_ASAP7_75t_R FILLER_215_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1196 ();
 DECAPx4_ASAP7_75t_R FILLER_215_1202 ();
 DECAPx1_ASAP7_75t_R FILLER_215_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_216_2 ();
 DECAPx10_ASAP7_75t_R FILLER_216_24 ();
 DECAPx10_ASAP7_75t_R FILLER_216_46 ();
 DECAPx10_ASAP7_75t_R FILLER_216_68 ();
 DECAPx10_ASAP7_75t_R FILLER_216_90 ();
 DECAPx10_ASAP7_75t_R FILLER_216_112 ();
 DECAPx10_ASAP7_75t_R FILLER_216_134 ();
 DECAPx10_ASAP7_75t_R FILLER_216_156 ();
 DECAPx10_ASAP7_75t_R FILLER_216_178 ();
 DECAPx10_ASAP7_75t_R FILLER_216_200 ();
 DECAPx10_ASAP7_75t_R FILLER_216_222 ();
 DECAPx10_ASAP7_75t_R FILLER_216_244 ();
 DECAPx10_ASAP7_75t_R FILLER_216_266 ();
 DECAPx6_ASAP7_75t_R FILLER_216_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_308 ();
 DECAPx2_ASAP7_75t_R FILLER_216_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_327 ();
 DECAPx10_ASAP7_75t_R FILLER_216_346 ();
 DECAPx4_ASAP7_75t_R FILLER_216_368 ();
 DECAPx6_ASAP7_75t_R FILLER_216_384 ();
 FILLER_ASAP7_75t_R FILLER_216_398 ();
 DECAPx6_ASAP7_75t_R FILLER_216_414 ();
 FILLER_ASAP7_75t_R FILLER_216_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_430 ();
 DECAPx6_ASAP7_75t_R FILLER_216_448 ();
 DECAPx4_ASAP7_75t_R FILLER_216_464 ();
 FILLER_ASAP7_75t_R FILLER_216_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_499 ();
 DECAPx6_ASAP7_75t_R FILLER_216_512 ();
 DECAPx2_ASAP7_75t_R FILLER_216_526 ();
 DECAPx1_ASAP7_75t_R FILLER_216_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_558 ();
 DECAPx10_ASAP7_75t_R FILLER_216_582 ();
 DECAPx10_ASAP7_75t_R FILLER_216_604 ();
 DECAPx1_ASAP7_75t_R FILLER_216_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_630 ();
 DECAPx4_ASAP7_75t_R FILLER_216_653 ();
 FILLER_ASAP7_75t_R FILLER_216_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_665 ();
 DECAPx2_ASAP7_75t_R FILLER_216_695 ();
 DECAPx10_ASAP7_75t_R FILLER_216_724 ();
 DECAPx10_ASAP7_75t_R FILLER_216_746 ();
 DECAPx2_ASAP7_75t_R FILLER_216_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_781 ();
 DECAPx1_ASAP7_75t_R FILLER_216_842 ();
 DECAPx10_ASAP7_75t_R FILLER_216_876 ();
 DECAPx4_ASAP7_75t_R FILLER_216_898 ();
 DECAPx6_ASAP7_75t_R FILLER_216_936 ();
 FILLER_ASAP7_75t_R FILLER_216_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_960 ();
 DECAPx1_ASAP7_75t_R FILLER_216_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_973 ();
 FILLER_ASAP7_75t_R FILLER_216_981 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1030 ();
 DECAPx6_ASAP7_75t_R FILLER_216_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1146 ();
 DECAPx4_ASAP7_75t_R FILLER_216_1155 ();
 FILLER_ASAP7_75t_R FILLER_216_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1170 ();
 FILLER_ASAP7_75t_R FILLER_216_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_217_2 ();
 DECAPx10_ASAP7_75t_R FILLER_217_24 ();
 DECAPx10_ASAP7_75t_R FILLER_217_46 ();
 DECAPx10_ASAP7_75t_R FILLER_217_68 ();
 DECAPx10_ASAP7_75t_R FILLER_217_90 ();
 DECAPx10_ASAP7_75t_R FILLER_217_112 ();
 DECAPx10_ASAP7_75t_R FILLER_217_134 ();
 DECAPx10_ASAP7_75t_R FILLER_217_156 ();
 DECAPx10_ASAP7_75t_R FILLER_217_178 ();
 DECAPx10_ASAP7_75t_R FILLER_217_200 ();
 DECAPx10_ASAP7_75t_R FILLER_217_222 ();
 DECAPx10_ASAP7_75t_R FILLER_217_244 ();
 DECAPx10_ASAP7_75t_R FILLER_217_266 ();
 DECAPx10_ASAP7_75t_R FILLER_217_288 ();
 DECAPx6_ASAP7_75t_R FILLER_217_310 ();
 FILLER_ASAP7_75t_R FILLER_217_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_333 ();
 FILLER_ASAP7_75t_R FILLER_217_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_342 ();
 DECAPx2_ASAP7_75t_R FILLER_217_354 ();
 FILLER_ASAP7_75t_R FILLER_217_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_376 ();
 DECAPx1_ASAP7_75t_R FILLER_217_399 ();
 DECAPx6_ASAP7_75t_R FILLER_217_409 ();
 DECAPx1_ASAP7_75t_R FILLER_217_423 ();
 DECAPx10_ASAP7_75t_R FILLER_217_449 ();
 DECAPx10_ASAP7_75t_R FILLER_217_471 ();
 FILLER_ASAP7_75t_R FILLER_217_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_495 ();
 DECAPx10_ASAP7_75t_R FILLER_217_511 ();
 DECAPx10_ASAP7_75t_R FILLER_217_533 ();
 DECAPx1_ASAP7_75t_R FILLER_217_555 ();
 DECAPx1_ASAP7_75t_R FILLER_217_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_579 ();
 DECAPx10_ASAP7_75t_R FILLER_217_586 ();
 DECAPx1_ASAP7_75t_R FILLER_217_608 ();
 FILLER_ASAP7_75t_R FILLER_217_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_620 ();
 DECAPx6_ASAP7_75t_R FILLER_217_649 ();
 FILLER_ASAP7_75t_R FILLER_217_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_665 ();
 DECAPx10_ASAP7_75t_R FILLER_217_672 ();
 DECAPx10_ASAP7_75t_R FILLER_217_694 ();
 FILLER_ASAP7_75t_R FILLER_217_716 ();
 DECAPx1_ASAP7_75t_R FILLER_217_724 ();
 FILLER_ASAP7_75t_R FILLER_217_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_750 ();
 DECAPx2_ASAP7_75t_R FILLER_217_771 ();
 DECAPx6_ASAP7_75t_R FILLER_217_783 ();
 DECAPx1_ASAP7_75t_R FILLER_217_797 ();
 DECAPx6_ASAP7_75t_R FILLER_217_807 ();
 DECAPx6_ASAP7_75t_R FILLER_217_841 ();
 FILLER_ASAP7_75t_R FILLER_217_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_857 ();
 DECAPx10_ASAP7_75t_R FILLER_217_864 ();
 DECAPx6_ASAP7_75t_R FILLER_217_886 ();
 DECAPx1_ASAP7_75t_R FILLER_217_900 ();
 FILLER_ASAP7_75t_R FILLER_217_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_923 ();
 DECAPx4_ASAP7_75t_R FILLER_217_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_943 ();
 FILLER_ASAP7_75t_R FILLER_217_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_964 ();
 DECAPx6_ASAP7_75t_R FILLER_217_974 ();
 FILLER_ASAP7_75t_R FILLER_217_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_990 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_217_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1159 ();
 DECAPx6_ASAP7_75t_R FILLER_217_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1204 ();
 FILLER_ASAP7_75t_R FILLER_217_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_218_2 ();
 DECAPx10_ASAP7_75t_R FILLER_218_24 ();
 DECAPx10_ASAP7_75t_R FILLER_218_46 ();
 DECAPx10_ASAP7_75t_R FILLER_218_68 ();
 DECAPx10_ASAP7_75t_R FILLER_218_90 ();
 DECAPx10_ASAP7_75t_R FILLER_218_112 ();
 DECAPx10_ASAP7_75t_R FILLER_218_134 ();
 DECAPx10_ASAP7_75t_R FILLER_218_156 ();
 DECAPx10_ASAP7_75t_R FILLER_218_178 ();
 DECAPx10_ASAP7_75t_R FILLER_218_200 ();
 DECAPx10_ASAP7_75t_R FILLER_218_222 ();
 DECAPx10_ASAP7_75t_R FILLER_218_244 ();
 DECAPx10_ASAP7_75t_R FILLER_218_266 ();
 DECAPx4_ASAP7_75t_R FILLER_218_288 ();
 FILLER_ASAP7_75t_R FILLER_218_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_300 ();
 DECAPx4_ASAP7_75t_R FILLER_218_312 ();
 FILLER_ASAP7_75t_R FILLER_218_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_324 ();
 DECAPx2_ASAP7_75t_R FILLER_218_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_345 ();
 DECAPx6_ASAP7_75t_R FILLER_218_379 ();
 FILLER_ASAP7_75t_R FILLER_218_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_395 ();
 DECAPx1_ASAP7_75t_R FILLER_218_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_407 ();
 DECAPx4_ASAP7_75t_R FILLER_218_430 ();
 FILLER_ASAP7_75t_R FILLER_218_440 ();
 FILLER_ASAP7_75t_R FILLER_218_464 ();
 DECAPx6_ASAP7_75t_R FILLER_218_472 ();
 FILLER_ASAP7_75t_R FILLER_218_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_501 ();
 DECAPx6_ASAP7_75t_R FILLER_218_519 ();
 FILLER_ASAP7_75t_R FILLER_218_533 ();
 DECAPx1_ASAP7_75t_R FILLER_218_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_561 ();
 DECAPx6_ASAP7_75t_R FILLER_218_584 ();
 FILLER_ASAP7_75t_R FILLER_218_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_600 ();
 DECAPx6_ASAP7_75t_R FILLER_218_627 ();
 FILLER_ASAP7_75t_R FILLER_218_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_689 ();
 FILLER_ASAP7_75t_R FILLER_218_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_715 ();
 DECAPx10_ASAP7_75t_R FILLER_218_744 ();
 DECAPx4_ASAP7_75t_R FILLER_218_766 ();
 DECAPx6_ASAP7_75t_R FILLER_218_798 ();
 DECAPx1_ASAP7_75t_R FILLER_218_812 ();
 DECAPx1_ASAP7_75t_R FILLER_218_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_823 ();
 DECAPx1_ASAP7_75t_R FILLER_218_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_834 ();
 DECAPx4_ASAP7_75t_R FILLER_218_838 ();
 FILLER_ASAP7_75t_R FILLER_218_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_861 ();
 DECAPx1_ASAP7_75t_R FILLER_218_868 ();
 DECAPx10_ASAP7_75t_R FILLER_218_889 ();
 DECAPx10_ASAP7_75t_R FILLER_218_911 ();
 FILLER_ASAP7_75t_R FILLER_218_933 ();
 DECAPx10_ASAP7_75t_R FILLER_218_982 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1114 ();
 FILLER_ASAP7_75t_R FILLER_218_1120 ();
 FILLER_ASAP7_75t_R FILLER_218_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1133 ();
 FILLER_ASAP7_75t_R FILLER_218_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1158 ();
 DECAPx4_ASAP7_75t_R FILLER_218_1180 ();
 FILLER_ASAP7_75t_R FILLER_218_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1192 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1196 ();
 FILLER_ASAP7_75t_R FILLER_218_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1212 ();
 FILLER_ASAP7_75t_R FILLER_218_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_219_2 ();
 DECAPx10_ASAP7_75t_R FILLER_219_24 ();
 DECAPx10_ASAP7_75t_R FILLER_219_46 ();
 DECAPx10_ASAP7_75t_R FILLER_219_68 ();
 DECAPx10_ASAP7_75t_R FILLER_219_90 ();
 DECAPx10_ASAP7_75t_R FILLER_219_112 ();
 DECAPx10_ASAP7_75t_R FILLER_219_134 ();
 DECAPx10_ASAP7_75t_R FILLER_219_156 ();
 DECAPx10_ASAP7_75t_R FILLER_219_178 ();
 DECAPx10_ASAP7_75t_R FILLER_219_200 ();
 DECAPx10_ASAP7_75t_R FILLER_219_222 ();
 DECAPx10_ASAP7_75t_R FILLER_219_244 ();
 DECAPx10_ASAP7_75t_R FILLER_219_266 ();
 DECAPx4_ASAP7_75t_R FILLER_219_288 ();
 DECAPx4_ASAP7_75t_R FILLER_219_340 ();
 DECAPx2_ASAP7_75t_R FILLER_219_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_362 ();
 DECAPx6_ASAP7_75t_R FILLER_219_377 ();
 DECAPx10_ASAP7_75t_R FILLER_219_414 ();
 DECAPx2_ASAP7_75t_R FILLER_219_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_442 ();
 DECAPx1_ASAP7_75t_R FILLER_219_472 ();
 DECAPx1_ASAP7_75t_R FILLER_219_487 ();
 DECAPx1_ASAP7_75t_R FILLER_219_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_501 ();
 DECAPx1_ASAP7_75t_R FILLER_219_509 ();
 DECAPx1_ASAP7_75t_R FILLER_219_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_539 ();
 DECAPx6_ASAP7_75t_R FILLER_219_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_560 ();
 DECAPx4_ASAP7_75t_R FILLER_219_567 ();
 DECAPx6_ASAP7_75t_R FILLER_219_594 ();
 FILLER_ASAP7_75t_R FILLER_219_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_610 ();
 DECAPx6_ASAP7_75t_R FILLER_219_617 ();
 DECAPx2_ASAP7_75t_R FILLER_219_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_637 ();
 DECAPx10_ASAP7_75t_R FILLER_219_661 ();
 DECAPx6_ASAP7_75t_R FILLER_219_683 ();
 FILLER_ASAP7_75t_R FILLER_219_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_699 ();
 DECAPx10_ASAP7_75t_R FILLER_219_703 ();
 DECAPx4_ASAP7_75t_R FILLER_219_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_735 ();
 DECAPx2_ASAP7_75t_R FILLER_219_748 ();
 FILLER_ASAP7_75t_R FILLER_219_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_756 ();
 DECAPx2_ASAP7_75t_R FILLER_219_777 ();
 FILLER_ASAP7_75t_R FILLER_219_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_791 ();
 DECAPx10_ASAP7_75t_R FILLER_219_832 ();
 DECAPx1_ASAP7_75t_R FILLER_219_854 ();
 DECAPx6_ASAP7_75t_R FILLER_219_906 ();
 DECAPx1_ASAP7_75t_R FILLER_219_920 ();
 DECAPx10_ASAP7_75t_R FILLER_219_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_948 ();
 DECAPx6_ASAP7_75t_R FILLER_219_955 ();
 DECAPx2_ASAP7_75t_R FILLER_219_969 ();
 DECAPx10_ASAP7_75t_R FILLER_219_997 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_219_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_220_2 ();
 DECAPx10_ASAP7_75t_R FILLER_220_24 ();
 DECAPx10_ASAP7_75t_R FILLER_220_46 ();
 DECAPx10_ASAP7_75t_R FILLER_220_68 ();
 DECAPx10_ASAP7_75t_R FILLER_220_90 ();
 DECAPx10_ASAP7_75t_R FILLER_220_112 ();
 DECAPx10_ASAP7_75t_R FILLER_220_134 ();
 DECAPx10_ASAP7_75t_R FILLER_220_156 ();
 DECAPx10_ASAP7_75t_R FILLER_220_178 ();
 DECAPx10_ASAP7_75t_R FILLER_220_200 ();
 DECAPx10_ASAP7_75t_R FILLER_220_222 ();
 DECAPx10_ASAP7_75t_R FILLER_220_244 ();
 DECAPx10_ASAP7_75t_R FILLER_220_266 ();
 DECAPx6_ASAP7_75t_R FILLER_220_288 ();
 DECAPx2_ASAP7_75t_R FILLER_220_302 ();
 DECAPx10_ASAP7_75t_R FILLER_220_314 ();
 DECAPx4_ASAP7_75t_R FILLER_220_336 ();
 FILLER_ASAP7_75t_R FILLER_220_346 ();
 DECAPx4_ASAP7_75t_R FILLER_220_354 ();
 FILLER_ASAP7_75t_R FILLER_220_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_366 ();
 FILLER_ASAP7_75t_R FILLER_220_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_377 ();
 DECAPx2_ASAP7_75t_R FILLER_220_386 ();
 FILLER_ASAP7_75t_R FILLER_220_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_394 ();
 DECAPx10_ASAP7_75t_R FILLER_220_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_437 ();
 DECAPx1_ASAP7_75t_R FILLER_220_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_464 ();
 DECAPx10_ASAP7_75t_R FILLER_220_509 ();
 DECAPx2_ASAP7_75t_R FILLER_220_531 ();
 FILLER_ASAP7_75t_R FILLER_220_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_539 ();
 DECAPx4_ASAP7_75t_R FILLER_220_551 ();
 DECAPx6_ASAP7_75t_R FILLER_220_567 ();
 DECAPx1_ASAP7_75t_R FILLER_220_581 ();
 DECAPx4_ASAP7_75t_R FILLER_220_627 ();
 FILLER_ASAP7_75t_R FILLER_220_637 ();
 DECAPx6_ASAP7_75t_R FILLER_220_645 ();
 DECAPx2_ASAP7_75t_R FILLER_220_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_687 ();
 DECAPx1_ASAP7_75t_R FILLER_220_708 ();
 DECAPx10_ASAP7_75t_R FILLER_220_715 ();
 FILLER_ASAP7_75t_R FILLER_220_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_739 ();
 DECAPx10_ASAP7_75t_R FILLER_220_743 ();
 DECAPx10_ASAP7_75t_R FILLER_220_765 ();
 DECAPx10_ASAP7_75t_R FILLER_220_787 ();
 FILLER_ASAP7_75t_R FILLER_220_809 ();
 DECAPx6_ASAP7_75t_R FILLER_220_814 ();
 FILLER_ASAP7_75t_R FILLER_220_828 ();
 DECAPx10_ASAP7_75t_R FILLER_220_833 ();
 DECAPx6_ASAP7_75t_R FILLER_220_855 ();
 FILLER_ASAP7_75t_R FILLER_220_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_877 ();
 DECAPx4_ASAP7_75t_R FILLER_220_887 ();
 FILLER_ASAP7_75t_R FILLER_220_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_899 ();
 FILLER_ASAP7_75t_R FILLER_220_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_924 ();
 DECAPx2_ASAP7_75t_R FILLER_220_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_937 ();
 DECAPx10_ASAP7_75t_R FILLER_220_960 ();
 DECAPx10_ASAP7_75t_R FILLER_220_982 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1140 ();
 FILLER_ASAP7_75t_R FILLER_220_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_220_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1176 ();
 DECAPx6_ASAP7_75t_R FILLER_220_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_221_2 ();
 DECAPx10_ASAP7_75t_R FILLER_221_24 ();
 DECAPx10_ASAP7_75t_R FILLER_221_46 ();
 DECAPx10_ASAP7_75t_R FILLER_221_68 ();
 DECAPx10_ASAP7_75t_R FILLER_221_90 ();
 DECAPx10_ASAP7_75t_R FILLER_221_112 ();
 DECAPx10_ASAP7_75t_R FILLER_221_134 ();
 DECAPx10_ASAP7_75t_R FILLER_221_156 ();
 DECAPx10_ASAP7_75t_R FILLER_221_178 ();
 DECAPx10_ASAP7_75t_R FILLER_221_200 ();
 DECAPx10_ASAP7_75t_R FILLER_221_222 ();
 DECAPx10_ASAP7_75t_R FILLER_221_244 ();
 DECAPx6_ASAP7_75t_R FILLER_221_266 ();
 DECAPx1_ASAP7_75t_R FILLER_221_280 ();
 FILLER_ASAP7_75t_R FILLER_221_306 ();
 DECAPx6_ASAP7_75t_R FILLER_221_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_335 ();
 DECAPx1_ASAP7_75t_R FILLER_221_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_362 ();
 DECAPx1_ASAP7_75t_R FILLER_221_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_396 ();
 DECAPx6_ASAP7_75t_R FILLER_221_414 ();
 FILLER_ASAP7_75t_R FILLER_221_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_430 ();
 DECAPx1_ASAP7_75t_R FILLER_221_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_457 ();
 FILLER_ASAP7_75t_R FILLER_221_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_472 ();
 DECAPx1_ASAP7_75t_R FILLER_221_486 ();
 DECAPx4_ASAP7_75t_R FILLER_221_502 ();
 FILLER_ASAP7_75t_R FILLER_221_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_514 ();
 FILLER_ASAP7_75t_R FILLER_221_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_527 ();
 FILLER_ASAP7_75t_R FILLER_221_545 ();
 DECAPx1_ASAP7_75t_R FILLER_221_555 ();
 DECAPx6_ASAP7_75t_R FILLER_221_576 ();
 FILLER_ASAP7_75t_R FILLER_221_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_614 ();
 FILLER_ASAP7_75t_R FILLER_221_661 ();
 DECAPx4_ASAP7_75t_R FILLER_221_669 ();
 FILLER_ASAP7_75t_R FILLER_221_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_681 ();
 DECAPx2_ASAP7_75t_R FILLER_221_705 ();
 FILLER_ASAP7_75t_R FILLER_221_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_713 ();
 FILLER_ASAP7_75t_R FILLER_221_748 ();
 DECAPx1_ASAP7_75t_R FILLER_221_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_771 ();
 DECAPx2_ASAP7_75t_R FILLER_221_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_828 ();
 DECAPx2_ASAP7_75t_R FILLER_221_849 ();
 DECAPx1_ASAP7_75t_R FILLER_221_909 ();
 DECAPx1_ASAP7_75t_R FILLER_221_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_952 ();
 DECAPx10_ASAP7_75t_R FILLER_221_975 ();
 DECAPx10_ASAP7_75t_R FILLER_221_997 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1113 ();
 DECAPx4_ASAP7_75t_R FILLER_221_1122 ();
 FILLER_ASAP7_75t_R FILLER_221_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_221_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1210 ();
 FILLER_ASAP7_75t_R FILLER_221_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_222_2 ();
 DECAPx10_ASAP7_75t_R FILLER_222_24 ();
 DECAPx10_ASAP7_75t_R FILLER_222_46 ();
 DECAPx10_ASAP7_75t_R FILLER_222_68 ();
 DECAPx10_ASAP7_75t_R FILLER_222_90 ();
 DECAPx10_ASAP7_75t_R FILLER_222_112 ();
 DECAPx10_ASAP7_75t_R FILLER_222_134 ();
 DECAPx10_ASAP7_75t_R FILLER_222_156 ();
 DECAPx10_ASAP7_75t_R FILLER_222_178 ();
 DECAPx10_ASAP7_75t_R FILLER_222_200 ();
 DECAPx10_ASAP7_75t_R FILLER_222_222 ();
 DECAPx10_ASAP7_75t_R FILLER_222_244 ();
 DECAPx10_ASAP7_75t_R FILLER_222_266 ();
 DECAPx2_ASAP7_75t_R FILLER_222_305 ();
 DECAPx6_ASAP7_75t_R FILLER_222_325 ();
 DECAPx1_ASAP7_75t_R FILLER_222_339 ();
 DECAPx4_ASAP7_75t_R FILLER_222_357 ();
 FILLER_ASAP7_75t_R FILLER_222_367 ();
 DECAPx10_ASAP7_75t_R FILLER_222_375 ();
 DECAPx2_ASAP7_75t_R FILLER_222_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_426 ();
 FILLER_ASAP7_75t_R FILLER_222_433 ();
 FILLER_ASAP7_75t_R FILLER_222_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_450 ();
 DECAPx1_ASAP7_75t_R FILLER_222_458 ();
 DECAPx2_ASAP7_75t_R FILLER_222_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_492 ();
 DECAPx6_ASAP7_75t_R FILLER_222_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_515 ();
 FILLER_ASAP7_75t_R FILLER_222_588 ();
 DECAPx10_ASAP7_75t_R FILLER_222_598 ();
 DECAPx1_ASAP7_75t_R FILLER_222_620 ();
 DECAPx1_ASAP7_75t_R FILLER_222_630 ();
 DECAPx6_ASAP7_75t_R FILLER_222_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_664 ();
 DECAPx6_ASAP7_75t_R FILLER_222_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_704 ();
 DECAPx2_ASAP7_75t_R FILLER_222_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_733 ();
 DECAPx1_ASAP7_75t_R FILLER_222_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_759 ();
 DECAPx4_ASAP7_75t_R FILLER_222_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_792 ();
 DECAPx1_ASAP7_75t_R FILLER_222_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_817 ();
 DECAPx6_ASAP7_75t_R FILLER_222_821 ();
 DECAPx2_ASAP7_75t_R FILLER_222_835 ();
 DECAPx4_ASAP7_75t_R FILLER_222_850 ();
 DECAPx2_ASAP7_75t_R FILLER_222_866 ();
 FILLER_ASAP7_75t_R FILLER_222_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_874 ();
 DECAPx10_ASAP7_75t_R FILLER_222_909 ();
 DECAPx6_ASAP7_75t_R FILLER_222_931 ();
 FILLER_ASAP7_75t_R FILLER_222_945 ();
 DECAPx4_ASAP7_75t_R FILLER_222_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_969 ();
 DECAPx10_ASAP7_75t_R FILLER_222_976 ();
 DECAPx10_ASAP7_75t_R FILLER_222_998 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1020 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_222_1130 ();
 FILLER_ASAP7_75t_R FILLER_222_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_223_2 ();
 DECAPx10_ASAP7_75t_R FILLER_223_24 ();
 DECAPx10_ASAP7_75t_R FILLER_223_46 ();
 DECAPx10_ASAP7_75t_R FILLER_223_68 ();
 DECAPx10_ASAP7_75t_R FILLER_223_90 ();
 DECAPx10_ASAP7_75t_R FILLER_223_112 ();
 DECAPx10_ASAP7_75t_R FILLER_223_134 ();
 DECAPx10_ASAP7_75t_R FILLER_223_156 ();
 DECAPx10_ASAP7_75t_R FILLER_223_178 ();
 DECAPx10_ASAP7_75t_R FILLER_223_200 ();
 DECAPx10_ASAP7_75t_R FILLER_223_222 ();
 DECAPx10_ASAP7_75t_R FILLER_223_244 ();
 DECAPx10_ASAP7_75t_R FILLER_223_266 ();
 DECAPx1_ASAP7_75t_R FILLER_223_288 ();
 DECAPx4_ASAP7_75t_R FILLER_223_327 ();
 FILLER_ASAP7_75t_R FILLER_223_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_339 ();
 DECAPx6_ASAP7_75t_R FILLER_223_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_368 ();
 DECAPx10_ASAP7_75t_R FILLER_223_377 ();
 DECAPx10_ASAP7_75t_R FILLER_223_399 ();
 FILLER_ASAP7_75t_R FILLER_223_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_445 ();
 DECAPx6_ASAP7_75t_R FILLER_223_476 ();
 DECAPx10_ASAP7_75t_R FILLER_223_502 ();
 DECAPx4_ASAP7_75t_R FILLER_223_524 ();
 FILLER_ASAP7_75t_R FILLER_223_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_543 ();
 DECAPx4_ASAP7_75t_R FILLER_223_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_598 ();
 DECAPx6_ASAP7_75t_R FILLER_223_605 ();
 DECAPx2_ASAP7_75t_R FILLER_223_619 ();
 FILLER_ASAP7_75t_R FILLER_223_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_667 ();
 DECAPx10_ASAP7_75t_R FILLER_223_674 ();
 DECAPx2_ASAP7_75t_R FILLER_223_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_712 ();
 DECAPx2_ASAP7_75t_R FILLER_223_724 ();
 FILLER_ASAP7_75t_R FILLER_223_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_732 ();
 DECAPx10_ASAP7_75t_R FILLER_223_752 ();
 DECAPx6_ASAP7_75t_R FILLER_223_774 ();
 FILLER_ASAP7_75t_R FILLER_223_788 ();
 DECAPx6_ASAP7_75t_R FILLER_223_800 ();
 FILLER_ASAP7_75t_R FILLER_223_814 ();
 DECAPx6_ASAP7_75t_R FILLER_223_836 ();
 DECAPx1_ASAP7_75t_R FILLER_223_850 ();
 DECAPx2_ASAP7_75t_R FILLER_223_901 ();
 FILLER_ASAP7_75t_R FILLER_223_907 ();
 DECAPx2_ASAP7_75t_R FILLER_223_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_923 ();
 DECAPx2_ASAP7_75t_R FILLER_223_926 ();
 FILLER_ASAP7_75t_R FILLER_223_932 ();
 DECAPx4_ASAP7_75t_R FILLER_223_940 ();
 FILLER_ASAP7_75t_R FILLER_223_950 ();
 DECAPx10_ASAP7_75t_R FILLER_223_972 ();
 DECAPx10_ASAP7_75t_R FILLER_223_994 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_223_1192 ();
 FILLER_ASAP7_75t_R FILLER_223_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1208 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1212 ();
 FILLER_ASAP7_75t_R FILLER_223_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_224_2 ();
 DECAPx10_ASAP7_75t_R FILLER_224_24 ();
 DECAPx10_ASAP7_75t_R FILLER_224_46 ();
 DECAPx10_ASAP7_75t_R FILLER_224_68 ();
 DECAPx10_ASAP7_75t_R FILLER_224_90 ();
 DECAPx10_ASAP7_75t_R FILLER_224_112 ();
 DECAPx10_ASAP7_75t_R FILLER_224_134 ();
 DECAPx10_ASAP7_75t_R FILLER_224_156 ();
 DECAPx10_ASAP7_75t_R FILLER_224_178 ();
 DECAPx10_ASAP7_75t_R FILLER_224_200 ();
 DECAPx10_ASAP7_75t_R FILLER_224_222 ();
 DECAPx10_ASAP7_75t_R FILLER_224_244 ();
 DECAPx10_ASAP7_75t_R FILLER_224_266 ();
 DECAPx6_ASAP7_75t_R FILLER_224_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_302 ();
 DECAPx4_ASAP7_75t_R FILLER_224_314 ();
 FILLER_ASAP7_75t_R FILLER_224_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_346 ();
 DECAPx2_ASAP7_75t_R FILLER_224_353 ();
 FILLER_ASAP7_75t_R FILLER_224_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_361 ();
 FILLER_ASAP7_75t_R FILLER_224_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_379 ();
 DECAPx10_ASAP7_75t_R FILLER_224_410 ();
 DECAPx1_ASAP7_75t_R FILLER_224_432 ();
 FILLER_ASAP7_75t_R FILLER_224_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_452 ();
 FILLER_ASAP7_75t_R FILLER_224_460 ();
 DECAPx2_ASAP7_75t_R FILLER_224_470 ();
 FILLER_ASAP7_75t_R FILLER_224_476 ();
 DECAPx1_ASAP7_75t_R FILLER_224_491 ();
 DECAPx6_ASAP7_75t_R FILLER_224_517 ();
 FILLER_ASAP7_75t_R FILLER_224_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_533 ();
 DECAPx1_ASAP7_75t_R FILLER_224_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_546 ();
 DECAPx1_ASAP7_75t_R FILLER_224_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_558 ();
 DECAPx6_ASAP7_75t_R FILLER_224_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_599 ();
 DECAPx10_ASAP7_75t_R FILLER_224_611 ();
 DECAPx6_ASAP7_75t_R FILLER_224_633 ();
 DECAPx2_ASAP7_75t_R FILLER_224_675 ();
 DECAPx10_ASAP7_75t_R FILLER_224_684 ();
 DECAPx6_ASAP7_75t_R FILLER_224_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_720 ();
 DECAPx10_ASAP7_75t_R FILLER_224_754 ();
 DECAPx10_ASAP7_75t_R FILLER_224_776 ();
 DECAPx10_ASAP7_75t_R FILLER_224_798 ();
 DECAPx2_ASAP7_75t_R FILLER_224_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_826 ();
 FILLER_ASAP7_75t_R FILLER_224_862 ();
 DECAPx2_ASAP7_75t_R FILLER_224_867 ();
 FILLER_ASAP7_75t_R FILLER_224_873 ();
 DECAPx2_ASAP7_75t_R FILLER_224_881 ();
 DECAPx2_ASAP7_75t_R FILLER_224_897 ();
 FILLER_ASAP7_75t_R FILLER_224_903 ();
 DECAPx10_ASAP7_75t_R FILLER_224_961 ();
 DECAPx10_ASAP7_75t_R FILLER_224_983 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_224_1121 ();
 FILLER_ASAP7_75t_R FILLER_224_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1133 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1165 ();
 DECAPx4_ASAP7_75t_R FILLER_224_1187 ();
 FILLER_ASAP7_75t_R FILLER_224_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_225_2 ();
 DECAPx10_ASAP7_75t_R FILLER_225_24 ();
 DECAPx10_ASAP7_75t_R FILLER_225_46 ();
 DECAPx10_ASAP7_75t_R FILLER_225_68 ();
 DECAPx10_ASAP7_75t_R FILLER_225_90 ();
 DECAPx10_ASAP7_75t_R FILLER_225_112 ();
 DECAPx10_ASAP7_75t_R FILLER_225_134 ();
 DECAPx10_ASAP7_75t_R FILLER_225_156 ();
 DECAPx10_ASAP7_75t_R FILLER_225_178 ();
 DECAPx10_ASAP7_75t_R FILLER_225_200 ();
 DECAPx10_ASAP7_75t_R FILLER_225_222 ();
 DECAPx10_ASAP7_75t_R FILLER_225_244 ();
 DECAPx10_ASAP7_75t_R FILLER_225_266 ();
 DECAPx6_ASAP7_75t_R FILLER_225_288 ();
 DECAPx2_ASAP7_75t_R FILLER_225_302 ();
 DECAPx2_ASAP7_75t_R FILLER_225_325 ();
 DECAPx6_ASAP7_75t_R FILLER_225_350 ();
 FILLER_ASAP7_75t_R FILLER_225_364 ();
 DECAPx4_ASAP7_75t_R FILLER_225_394 ();
 FILLER_ASAP7_75t_R FILLER_225_404 ();
 DECAPx1_ASAP7_75t_R FILLER_225_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_416 ();
 DECAPx1_ASAP7_75t_R FILLER_225_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_477 ();
 DECAPx6_ASAP7_75t_R FILLER_225_489 ();
 DECAPx1_ASAP7_75t_R FILLER_225_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_507 ();
 DECAPx2_ASAP7_75t_R FILLER_225_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_517 ();
 DECAPx2_ASAP7_75t_R FILLER_225_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_573 ();
 DECAPx2_ASAP7_75t_R FILLER_225_607 ();
 DECAPx1_ASAP7_75t_R FILLER_225_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_641 ();
 DECAPx10_ASAP7_75t_R FILLER_225_645 ();
 DECAPx4_ASAP7_75t_R FILLER_225_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_677 ();
 DECAPx1_ASAP7_75t_R FILLER_225_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_702 ();
 FILLER_ASAP7_75t_R FILLER_225_732 ();
 DECAPx1_ASAP7_75t_R FILLER_225_742 ();
 DECAPx2_ASAP7_75t_R FILLER_225_774 ();
 FILLER_ASAP7_75t_R FILLER_225_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_788 ();
 FILLER_ASAP7_75t_R FILLER_225_810 ();
 FILLER_ASAP7_75t_R FILLER_225_817 ();
 DECAPx4_ASAP7_75t_R FILLER_225_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_840 ();
 DECAPx2_ASAP7_75t_R FILLER_225_846 ();
 FILLER_ASAP7_75t_R FILLER_225_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_854 ();
 DECAPx1_ASAP7_75t_R FILLER_225_863 ();
 DECAPx2_ASAP7_75t_R FILLER_225_875 ();
 FILLER_ASAP7_75t_R FILLER_225_881 ();
 DECAPx4_ASAP7_75t_R FILLER_225_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_911 ();
 DECAPx6_ASAP7_75t_R FILLER_225_937 ();
 FILLER_ASAP7_75t_R FILLER_225_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_953 ();
 DECAPx10_ASAP7_75t_R FILLER_225_974 ();
 DECAPx10_ASAP7_75t_R FILLER_225_996 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1128 ();
 DECAPx6_ASAP7_75t_R FILLER_225_1150 ();
 FILLER_ASAP7_75t_R FILLER_225_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_225_1191 ();
 FILLER_ASAP7_75t_R FILLER_225_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1208 ();
 FILLER_ASAP7_75t_R FILLER_225_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_226_2 ();
 DECAPx10_ASAP7_75t_R FILLER_226_24 ();
 DECAPx10_ASAP7_75t_R FILLER_226_46 ();
 DECAPx10_ASAP7_75t_R FILLER_226_68 ();
 DECAPx10_ASAP7_75t_R FILLER_226_90 ();
 DECAPx10_ASAP7_75t_R FILLER_226_112 ();
 DECAPx10_ASAP7_75t_R FILLER_226_134 ();
 DECAPx10_ASAP7_75t_R FILLER_226_156 ();
 DECAPx10_ASAP7_75t_R FILLER_226_178 ();
 DECAPx10_ASAP7_75t_R FILLER_226_200 ();
 DECAPx10_ASAP7_75t_R FILLER_226_222 ();
 DECAPx10_ASAP7_75t_R FILLER_226_244 ();
 DECAPx6_ASAP7_75t_R FILLER_226_266 ();
 DECAPx2_ASAP7_75t_R FILLER_226_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_315 ();
 DECAPx4_ASAP7_75t_R FILLER_226_322 ();
 FILLER_ASAP7_75t_R FILLER_226_332 ();
 DECAPx2_ASAP7_75t_R FILLER_226_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_362 ();
 FILLER_ASAP7_75t_R FILLER_226_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_372 ();
 DECAPx2_ASAP7_75t_R FILLER_226_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_401 ();
 FILLER_ASAP7_75t_R FILLER_226_428 ();
 DECAPx6_ASAP7_75t_R FILLER_226_436 ();
 DECAPx1_ASAP7_75t_R FILLER_226_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_461 ();
 DECAPx6_ASAP7_75t_R FILLER_226_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_478 ();
 DECAPx10_ASAP7_75t_R FILLER_226_485 ();
 DECAPx10_ASAP7_75t_R FILLER_226_507 ();
 DECAPx1_ASAP7_75t_R FILLER_226_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_533 ();
 DECAPx6_ASAP7_75t_R FILLER_226_540 ();
 DECAPx4_ASAP7_75t_R FILLER_226_560 ();
 FILLER_ASAP7_75t_R FILLER_226_570 ();
 DECAPx4_ASAP7_75t_R FILLER_226_600 ();
 FILLER_ASAP7_75t_R FILLER_226_610 ();
 DECAPx10_ASAP7_75t_R FILLER_226_639 ();
 DECAPx6_ASAP7_75t_R FILLER_226_661 ();
 DECAPx2_ASAP7_75t_R FILLER_226_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_681 ();
 DECAPx4_ASAP7_75t_R FILLER_226_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_698 ();
 DECAPx1_ASAP7_75t_R FILLER_226_710 ();
 DECAPx1_ASAP7_75t_R FILLER_226_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_724 ();
 DECAPx2_ASAP7_75t_R FILLER_226_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_744 ();
 DECAPx10_ASAP7_75t_R FILLER_226_751 ();
 DECAPx1_ASAP7_75t_R FILLER_226_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_777 ();
 DECAPx10_ASAP7_75t_R FILLER_226_800 ();
 DECAPx1_ASAP7_75t_R FILLER_226_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_838 ();
 DECAPx1_ASAP7_75t_R FILLER_226_850 ();
 DECAPx2_ASAP7_75t_R FILLER_226_860 ();
 FILLER_ASAP7_75t_R FILLER_226_866 ();
 DECAPx2_ASAP7_75t_R FILLER_226_902 ();
 FILLER_ASAP7_75t_R FILLER_226_908 ();
 DECAPx10_ASAP7_75t_R FILLER_226_924 ();
 DECAPx6_ASAP7_75t_R FILLER_226_946 ();
 FILLER_ASAP7_75t_R FILLER_226_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_962 ();
 DECAPx10_ASAP7_75t_R FILLER_226_993 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_226_1037 ();
 FILLER_ASAP7_75t_R FILLER_226_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1145 ();
 DECAPx4_ASAP7_75t_R FILLER_226_1172 ();
 FILLER_ASAP7_75t_R FILLER_226_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1188 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_227_2 ();
 DECAPx10_ASAP7_75t_R FILLER_227_24 ();
 DECAPx10_ASAP7_75t_R FILLER_227_46 ();
 DECAPx10_ASAP7_75t_R FILLER_227_68 ();
 DECAPx10_ASAP7_75t_R FILLER_227_90 ();
 DECAPx10_ASAP7_75t_R FILLER_227_112 ();
 DECAPx10_ASAP7_75t_R FILLER_227_134 ();
 DECAPx10_ASAP7_75t_R FILLER_227_156 ();
 DECAPx10_ASAP7_75t_R FILLER_227_178 ();
 DECAPx10_ASAP7_75t_R FILLER_227_200 ();
 DECAPx10_ASAP7_75t_R FILLER_227_222 ();
 DECAPx10_ASAP7_75t_R FILLER_227_244 ();
 DECAPx10_ASAP7_75t_R FILLER_227_266 ();
 FILLER_ASAP7_75t_R FILLER_227_288 ();
 FILLER_ASAP7_75t_R FILLER_227_296 ();
 DECAPx1_ASAP7_75t_R FILLER_227_316 ();
 DECAPx10_ASAP7_75t_R FILLER_227_334 ();
 DECAPx2_ASAP7_75t_R FILLER_227_356 ();
 DECAPx10_ASAP7_75t_R FILLER_227_387 ();
 DECAPx6_ASAP7_75t_R FILLER_227_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_423 ();
 DECAPx6_ASAP7_75t_R FILLER_227_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_452 ();
 DECAPx4_ASAP7_75t_R FILLER_227_461 ();
 FILLER_ASAP7_75t_R FILLER_227_471 ();
 DECAPx4_ASAP7_75t_R FILLER_227_495 ();
 FILLER_ASAP7_75t_R FILLER_227_505 ();
 DECAPx6_ASAP7_75t_R FILLER_227_527 ();
 FILLER_ASAP7_75t_R FILLER_227_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_554 ();
 DECAPx2_ASAP7_75t_R FILLER_227_577 ();
 FILLER_ASAP7_75t_R FILLER_227_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_585 ();
 DECAPx1_ASAP7_75t_R FILLER_227_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_596 ();
 DECAPx2_ASAP7_75t_R FILLER_227_623 ();
 FILLER_ASAP7_75t_R FILLER_227_629 ();
 DECAPx1_ASAP7_75t_R FILLER_227_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_643 ();
 DECAPx6_ASAP7_75t_R FILLER_227_656 ();
 DECAPx2_ASAP7_75t_R FILLER_227_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_676 ();
 DECAPx4_ASAP7_75t_R FILLER_227_716 ();
 DECAPx6_ASAP7_75t_R FILLER_227_759 ();
 DECAPx10_ASAP7_75t_R FILLER_227_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_857 ();
 DECAPx4_ASAP7_75t_R FILLER_227_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_882 ();
 DECAPx6_ASAP7_75t_R FILLER_227_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_904 ();
 DECAPx2_ASAP7_75t_R FILLER_227_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_923 ();
 DECAPx6_ASAP7_75t_R FILLER_227_926 ();
 DECAPx2_ASAP7_75t_R FILLER_227_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_946 ();
 DECAPx1_ASAP7_75t_R FILLER_227_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_962 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1089 ();
 DECAPx4_ASAP7_75t_R FILLER_227_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_227_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1188 ();
 DECAPx6_ASAP7_75t_R FILLER_227_1194 ();
 FILLER_ASAP7_75t_R FILLER_227_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_228_2 ();
 DECAPx10_ASAP7_75t_R FILLER_228_24 ();
 DECAPx10_ASAP7_75t_R FILLER_228_46 ();
 DECAPx10_ASAP7_75t_R FILLER_228_68 ();
 DECAPx10_ASAP7_75t_R FILLER_228_90 ();
 DECAPx10_ASAP7_75t_R FILLER_228_112 ();
 DECAPx10_ASAP7_75t_R FILLER_228_134 ();
 DECAPx10_ASAP7_75t_R FILLER_228_156 ();
 DECAPx10_ASAP7_75t_R FILLER_228_178 ();
 DECAPx10_ASAP7_75t_R FILLER_228_200 ();
 DECAPx10_ASAP7_75t_R FILLER_228_222 ();
 DECAPx10_ASAP7_75t_R FILLER_228_244 ();
 DECAPx6_ASAP7_75t_R FILLER_228_266 ();
 DECAPx2_ASAP7_75t_R FILLER_228_280 ();
 FILLER_ASAP7_75t_R FILLER_228_308 ();
 DECAPx1_ASAP7_75t_R FILLER_228_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_354 ();
 FILLER_ASAP7_75t_R FILLER_228_366 ();
 DECAPx6_ASAP7_75t_R FILLER_228_374 ();
 DECAPx4_ASAP7_75t_R FILLER_228_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_408 ();
 DECAPx1_ASAP7_75t_R FILLER_228_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_419 ();
 DECAPx4_ASAP7_75t_R FILLER_228_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_441 ();
 FILLER_ASAP7_75t_R FILLER_228_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_452 ();
 FILLER_ASAP7_75t_R FILLER_228_460 ();
 FILLER_ASAP7_75t_R FILLER_228_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_466 ();
 DECAPx6_ASAP7_75t_R FILLER_228_495 ();
 DECAPx1_ASAP7_75t_R FILLER_228_509 ();
 FILLER_ASAP7_75t_R FILLER_228_529 ();
 FILLER_ASAP7_75t_R FILLER_228_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_551 ();
 FILLER_ASAP7_75t_R FILLER_228_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_562 ();
 FILLER_ASAP7_75t_R FILLER_228_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_587 ();
 FILLER_ASAP7_75t_R FILLER_228_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_596 ();
 DECAPx1_ASAP7_75t_R FILLER_228_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_609 ();
 FILLER_ASAP7_75t_R FILLER_228_621 ();
 FILLER_ASAP7_75t_R FILLER_228_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_651 ();
 DECAPx10_ASAP7_75t_R FILLER_228_676 ();
 FILLER_ASAP7_75t_R FILLER_228_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_706 ();
 FILLER_ASAP7_75t_R FILLER_228_714 ();
 DECAPx1_ASAP7_75t_R FILLER_228_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_733 ();
 FILLER_ASAP7_75t_R FILLER_228_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_743 ();
 DECAPx10_ASAP7_75t_R FILLER_228_761 ();
 DECAPx2_ASAP7_75t_R FILLER_228_783 ();
 FILLER_ASAP7_75t_R FILLER_228_795 ();
 DECAPx10_ASAP7_75t_R FILLER_228_819 ();
 DECAPx4_ASAP7_75t_R FILLER_228_841 ();
 FILLER_ASAP7_75t_R FILLER_228_857 ();
 DECAPx10_ASAP7_75t_R FILLER_228_868 ();
 DECAPx6_ASAP7_75t_R FILLER_228_890 ();
 DECAPx1_ASAP7_75t_R FILLER_228_904 ();
 FILLER_ASAP7_75t_R FILLER_228_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_932 ();
 FILLER_ASAP7_75t_R FILLER_228_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_943 ();
 DECAPx4_ASAP7_75t_R FILLER_228_961 ();
 FILLER_ASAP7_75t_R FILLER_228_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_973 ();
 DECAPx10_ASAP7_75t_R FILLER_228_991 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1101 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1141 ();
 FILLER_ASAP7_75t_R FILLER_228_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1152 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1174 ();
 DECAPx2_ASAP7_75t_R FILLER_228_1196 ();
 FILLER_ASAP7_75t_R FILLER_228_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1212 ();
 FILLER_ASAP7_75t_R FILLER_228_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_229_2 ();
 DECAPx10_ASAP7_75t_R FILLER_229_24 ();
 DECAPx10_ASAP7_75t_R FILLER_229_46 ();
 DECAPx10_ASAP7_75t_R FILLER_229_68 ();
 DECAPx10_ASAP7_75t_R FILLER_229_90 ();
 DECAPx10_ASAP7_75t_R FILLER_229_112 ();
 DECAPx10_ASAP7_75t_R FILLER_229_134 ();
 DECAPx10_ASAP7_75t_R FILLER_229_156 ();
 DECAPx10_ASAP7_75t_R FILLER_229_178 ();
 DECAPx10_ASAP7_75t_R FILLER_229_200 ();
 DECAPx10_ASAP7_75t_R FILLER_229_222 ();
 DECAPx10_ASAP7_75t_R FILLER_229_244 ();
 DECAPx10_ASAP7_75t_R FILLER_229_266 ();
 DECAPx4_ASAP7_75t_R FILLER_229_288 ();
 FILLER_ASAP7_75t_R FILLER_229_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_322 ();
 DECAPx1_ASAP7_75t_R FILLER_229_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_369 ();
 DECAPx2_ASAP7_75t_R FILLER_229_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_440 ();
 DECAPx1_ASAP7_75t_R FILLER_229_450 ();
 DECAPx6_ASAP7_75t_R FILLER_229_461 ();
 FILLER_ASAP7_75t_R FILLER_229_475 ();
 FILLER_ASAP7_75t_R FILLER_229_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_519 ();
 FILLER_ASAP7_75t_R FILLER_229_542 ();
 FILLER_ASAP7_75t_R FILLER_229_550 ();
 FILLER_ASAP7_75t_R FILLER_229_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_563 ();
 DECAPx6_ASAP7_75t_R FILLER_229_581 ();
 DECAPx2_ASAP7_75t_R FILLER_229_595 ();
 DECAPx4_ASAP7_75t_R FILLER_229_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_621 ();
 FILLER_ASAP7_75t_R FILLER_229_625 ();
 DECAPx6_ASAP7_75t_R FILLER_229_650 ();
 FILLER_ASAP7_75t_R FILLER_229_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_666 ();
 FILLER_ASAP7_75t_R FILLER_229_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_674 ();
 FILLER_ASAP7_75t_R FILLER_229_681 ();
 DECAPx2_ASAP7_75t_R FILLER_229_691 ();
 FILLER_ASAP7_75t_R FILLER_229_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_699 ();
 DECAPx2_ASAP7_75t_R FILLER_229_713 ();
 DECAPx1_ASAP7_75t_R FILLER_229_750 ();
 DECAPx1_ASAP7_75t_R FILLER_229_776 ();
 DECAPx1_ASAP7_75t_R FILLER_229_795 ();
 DECAPx6_ASAP7_75t_R FILLER_229_816 ();
 DECAPx2_ASAP7_75t_R FILLER_229_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_836 ();
 FILLER_ASAP7_75t_R FILLER_229_843 ();
 DECAPx1_ASAP7_75t_R FILLER_229_856 ();
 DECAPx1_ASAP7_75t_R FILLER_229_867 ();
 DECAPx1_ASAP7_75t_R FILLER_229_877 ();
 DECAPx2_ASAP7_75t_R FILLER_229_918 ();
 DECAPx2_ASAP7_75t_R FILLER_229_926 ();
 FILLER_ASAP7_75t_R FILLER_229_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_934 ();
 DECAPx10_ASAP7_75t_R FILLER_229_999 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1153 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1182 ();
 FILLER_ASAP7_75t_R FILLER_229_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1190 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1210 ();
 FILLER_ASAP7_75t_R FILLER_229_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_230_2 ();
 DECAPx10_ASAP7_75t_R FILLER_230_24 ();
 DECAPx10_ASAP7_75t_R FILLER_230_46 ();
 DECAPx10_ASAP7_75t_R FILLER_230_68 ();
 DECAPx10_ASAP7_75t_R FILLER_230_90 ();
 DECAPx10_ASAP7_75t_R FILLER_230_112 ();
 DECAPx10_ASAP7_75t_R FILLER_230_134 ();
 DECAPx10_ASAP7_75t_R FILLER_230_156 ();
 DECAPx10_ASAP7_75t_R FILLER_230_178 ();
 DECAPx10_ASAP7_75t_R FILLER_230_200 ();
 DECAPx10_ASAP7_75t_R FILLER_230_222 ();
 DECAPx10_ASAP7_75t_R FILLER_230_244 ();
 DECAPx10_ASAP7_75t_R FILLER_230_266 ();
 DECAPx4_ASAP7_75t_R FILLER_230_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_298 ();
 DECAPx4_ASAP7_75t_R FILLER_230_316 ();
 DECAPx1_ASAP7_75t_R FILLER_230_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_347 ();
 DECAPx2_ASAP7_75t_R FILLER_230_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_360 ();
 DECAPx10_ASAP7_75t_R FILLER_230_372 ();
 DECAPx10_ASAP7_75t_R FILLER_230_394 ();
 DECAPx2_ASAP7_75t_R FILLER_230_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_422 ();
 DECAPx10_ASAP7_75t_R FILLER_230_440 ();
 DECAPx6_ASAP7_75t_R FILLER_230_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_478 ();
 DECAPx1_ASAP7_75t_R FILLER_230_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_500 ();
 DECAPx6_ASAP7_75t_R FILLER_230_523 ();
 FILLER_ASAP7_75t_R FILLER_230_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_539 ();
 DECAPx4_ASAP7_75t_R FILLER_230_553 ();
 DECAPx4_ASAP7_75t_R FILLER_230_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_593 ();
 DECAPx10_ASAP7_75t_R FILLER_230_614 ();
 DECAPx2_ASAP7_75t_R FILLER_230_636 ();
 FILLER_ASAP7_75t_R FILLER_230_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_644 ();
 FILLER_ASAP7_75t_R FILLER_230_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_670 ();
 DECAPx6_ASAP7_75t_R FILLER_230_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_729 ();
 DECAPx1_ASAP7_75t_R FILLER_230_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_762 ();
 FILLER_ASAP7_75t_R FILLER_230_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_791 ();
 DECAPx10_ASAP7_75t_R FILLER_230_799 ();
 DECAPx6_ASAP7_75t_R FILLER_230_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_835 ();
 FILLER_ASAP7_75t_R FILLER_230_858 ();
 DECAPx1_ASAP7_75t_R FILLER_230_866 ();
 DECAPx1_ASAP7_75t_R FILLER_230_881 ();
 DECAPx1_ASAP7_75t_R FILLER_230_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_897 ();
 DECAPx6_ASAP7_75t_R FILLER_230_904 ();
 DECAPx1_ASAP7_75t_R FILLER_230_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_922 ();
 DECAPx1_ASAP7_75t_R FILLER_230_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_949 ();
 FILLER_ASAP7_75t_R FILLER_230_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_969 ();
 DECAPx10_ASAP7_75t_R FILLER_230_987 ();
 DECAPx4_ASAP7_75t_R FILLER_230_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_230_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1098 ();
 FILLER_ASAP7_75t_R FILLER_230_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_230_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1157 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1166 ();
 FILLER_ASAP7_75t_R FILLER_230_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1183 ();
 FILLER_ASAP7_75t_R FILLER_230_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1216 ();
 FILLER_ASAP7_75t_R FILLER_230_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_231_2 ();
 DECAPx10_ASAP7_75t_R FILLER_231_24 ();
 DECAPx10_ASAP7_75t_R FILLER_231_46 ();
 DECAPx10_ASAP7_75t_R FILLER_231_68 ();
 DECAPx10_ASAP7_75t_R FILLER_231_90 ();
 DECAPx10_ASAP7_75t_R FILLER_231_112 ();
 DECAPx10_ASAP7_75t_R FILLER_231_134 ();
 DECAPx10_ASAP7_75t_R FILLER_231_156 ();
 DECAPx10_ASAP7_75t_R FILLER_231_178 ();
 DECAPx10_ASAP7_75t_R FILLER_231_200 ();
 DECAPx10_ASAP7_75t_R FILLER_231_222 ();
 DECAPx10_ASAP7_75t_R FILLER_231_244 ();
 DECAPx10_ASAP7_75t_R FILLER_231_266 ();
 DECAPx10_ASAP7_75t_R FILLER_231_288 ();
 DECAPx2_ASAP7_75t_R FILLER_231_310 ();
 DECAPx10_ASAP7_75t_R FILLER_231_327 ();
 DECAPx4_ASAP7_75t_R FILLER_231_349 ();
 FILLER_ASAP7_75t_R FILLER_231_359 ();
 DECAPx10_ASAP7_75t_R FILLER_231_389 ();
 DECAPx2_ASAP7_75t_R FILLER_231_411 ();
 FILLER_ASAP7_75t_R FILLER_231_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_419 ();
 DECAPx2_ASAP7_75t_R FILLER_231_431 ();
 DECAPx2_ASAP7_75t_R FILLER_231_443 ();
 DECAPx6_ASAP7_75t_R FILLER_231_488 ();
 FILLER_ASAP7_75t_R FILLER_231_502 ();
 DECAPx10_ASAP7_75t_R FILLER_231_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_532 ();
 DECAPx4_ASAP7_75t_R FILLER_231_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_565 ();
 DECAPx4_ASAP7_75t_R FILLER_231_573 ();
 FILLER_ASAP7_75t_R FILLER_231_583 ();
 DECAPx1_ASAP7_75t_R FILLER_231_607 ();
 FILLER_ASAP7_75t_R FILLER_231_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_641 ();
 DECAPx2_ASAP7_75t_R FILLER_231_648 ();
 FILLER_ASAP7_75t_R FILLER_231_654 ();
 DECAPx10_ASAP7_75t_R FILLER_231_660 ();
 FILLER_ASAP7_75t_R FILLER_231_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_684 ();
 DECAPx4_ASAP7_75t_R FILLER_231_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_701 ();
 DECAPx10_ASAP7_75t_R FILLER_231_715 ();
 DECAPx10_ASAP7_75t_R FILLER_231_737 ();
 FILLER_ASAP7_75t_R FILLER_231_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_779 ();
 DECAPx6_ASAP7_75t_R FILLER_231_817 ();
 DECAPx1_ASAP7_75t_R FILLER_231_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_835 ();
 DECAPx4_ASAP7_75t_R FILLER_231_839 ();
 FILLER_ASAP7_75t_R FILLER_231_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_856 ();
 DECAPx2_ASAP7_75t_R FILLER_231_879 ();
 FILLER_ASAP7_75t_R FILLER_231_885 ();
 DECAPx2_ASAP7_75t_R FILLER_231_900 ();
 DECAPx2_ASAP7_75t_R FILLER_231_916 ();
 FILLER_ASAP7_75t_R FILLER_231_922 ();
 DECAPx2_ASAP7_75t_R FILLER_231_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_938 ();
 FILLER_ASAP7_75t_R FILLER_231_982 ();
 DECAPx6_ASAP7_75t_R FILLER_231_990 ();
 DECAPx1_ASAP7_75t_R FILLER_231_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1020 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1064 ();
 DECAPx6_ASAP7_75t_R FILLER_231_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1136 ();
 DECAPx6_ASAP7_75t_R FILLER_231_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1171 ();
 DECAPx4_ASAP7_75t_R FILLER_231_1193 ();
 FILLER_ASAP7_75t_R FILLER_231_1203 ();
 FILLER_ASAP7_75t_R FILLER_231_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1216 ();
 FILLER_ASAP7_75t_R FILLER_231_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_232_2 ();
 DECAPx10_ASAP7_75t_R FILLER_232_24 ();
 DECAPx10_ASAP7_75t_R FILLER_232_46 ();
 DECAPx10_ASAP7_75t_R FILLER_232_68 ();
 DECAPx10_ASAP7_75t_R FILLER_232_90 ();
 DECAPx10_ASAP7_75t_R FILLER_232_112 ();
 DECAPx10_ASAP7_75t_R FILLER_232_134 ();
 DECAPx10_ASAP7_75t_R FILLER_232_156 ();
 DECAPx10_ASAP7_75t_R FILLER_232_178 ();
 DECAPx10_ASAP7_75t_R FILLER_232_200 ();
 DECAPx10_ASAP7_75t_R FILLER_232_222 ();
 DECAPx10_ASAP7_75t_R FILLER_232_244 ();
 DECAPx10_ASAP7_75t_R FILLER_232_266 ();
 DECAPx10_ASAP7_75t_R FILLER_232_288 ();
 DECAPx10_ASAP7_75t_R FILLER_232_310 ();
 DECAPx10_ASAP7_75t_R FILLER_232_332 ();
 DECAPx10_ASAP7_75t_R FILLER_232_354 ();
 DECAPx10_ASAP7_75t_R FILLER_232_376 ();
 DECAPx4_ASAP7_75t_R FILLER_232_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_408 ();
 FILLER_ASAP7_75t_R FILLER_232_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_461 ();
 DECAPx10_ASAP7_75t_R FILLER_232_464 ();
 DECAPx4_ASAP7_75t_R FILLER_232_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_496 ();
 DECAPx10_ASAP7_75t_R FILLER_232_508 ();
 DECAPx2_ASAP7_75t_R FILLER_232_530 ();
 DECAPx10_ASAP7_75t_R FILLER_232_542 ();
 FILLER_ASAP7_75t_R FILLER_232_564 ();
 DECAPx6_ASAP7_75t_R FILLER_232_591 ();
 DECAPx2_ASAP7_75t_R FILLER_232_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_611 ();
 FILLER_ASAP7_75t_R FILLER_232_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_628 ();
 DECAPx1_ASAP7_75t_R FILLER_232_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_639 ();
 DECAPx6_ASAP7_75t_R FILLER_232_646 ();
 DECAPx10_ASAP7_75t_R FILLER_232_668 ();
 DECAPx10_ASAP7_75t_R FILLER_232_690 ();
 DECAPx10_ASAP7_75t_R FILLER_232_734 ();
 DECAPx4_ASAP7_75t_R FILLER_232_756 ();
 FILLER_ASAP7_75t_R FILLER_232_766 ();
 DECAPx2_ASAP7_75t_R FILLER_232_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_782 ();
 DECAPx1_ASAP7_75t_R FILLER_232_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_810 ();
 DECAPx6_ASAP7_75t_R FILLER_232_833 ();
 FILLER_ASAP7_75t_R FILLER_232_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_849 ();
 DECAPx4_ASAP7_75t_R FILLER_232_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_874 ();
 DECAPx2_ASAP7_75t_R FILLER_232_886 ();
 DECAPx2_ASAP7_75t_R FILLER_232_912 ();
 FILLER_ASAP7_75t_R FILLER_232_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_932 ();
 DECAPx1_ASAP7_75t_R FILLER_232_940 ();
 DECAPx10_ASAP7_75t_R FILLER_232_958 ();
 FILLER_ASAP7_75t_R FILLER_232_980 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1016 ();
 FILLER_ASAP7_75t_R FILLER_232_1022 ();
 DECAPx4_ASAP7_75t_R FILLER_232_1027 ();
 FILLER_ASAP7_75t_R FILLER_232_1037 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1042 ();
 FILLER_ASAP7_75t_R FILLER_232_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_232_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_232_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1208 ();
 FILLER_ASAP7_75t_R FILLER_232_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_233_2 ();
 DECAPx10_ASAP7_75t_R FILLER_233_24 ();
 DECAPx10_ASAP7_75t_R FILLER_233_46 ();
 DECAPx10_ASAP7_75t_R FILLER_233_68 ();
 DECAPx10_ASAP7_75t_R FILLER_233_90 ();
 DECAPx10_ASAP7_75t_R FILLER_233_112 ();
 DECAPx10_ASAP7_75t_R FILLER_233_134 ();
 DECAPx10_ASAP7_75t_R FILLER_233_156 ();
 DECAPx10_ASAP7_75t_R FILLER_233_178 ();
 DECAPx10_ASAP7_75t_R FILLER_233_200 ();
 DECAPx10_ASAP7_75t_R FILLER_233_222 ();
 DECAPx10_ASAP7_75t_R FILLER_233_244 ();
 DECAPx10_ASAP7_75t_R FILLER_233_266 ();
 DECAPx10_ASAP7_75t_R FILLER_233_288 ();
 DECAPx10_ASAP7_75t_R FILLER_233_310 ();
 DECAPx4_ASAP7_75t_R FILLER_233_332 ();
 FILLER_ASAP7_75t_R FILLER_233_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_344 ();
 FILLER_ASAP7_75t_R FILLER_233_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_367 ();
 DECAPx10_ASAP7_75t_R FILLER_233_371 ();
 DECAPx10_ASAP7_75t_R FILLER_233_393 ();
 DECAPx10_ASAP7_75t_R FILLER_233_415 ();
 DECAPx6_ASAP7_75t_R FILLER_233_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_451 ();
 DECAPx6_ASAP7_75t_R FILLER_233_458 ();
 DECAPx1_ASAP7_75t_R FILLER_233_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_485 ();
 DECAPx4_ASAP7_75t_R FILLER_233_492 ();
 DECAPx1_ASAP7_75t_R FILLER_233_509 ();
 DECAPx6_ASAP7_75t_R FILLER_233_530 ();
 FILLER_ASAP7_75t_R FILLER_233_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_546 ();
 FILLER_ASAP7_75t_R FILLER_233_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_555 ();
 FILLER_ASAP7_75t_R FILLER_233_567 ();
 DECAPx10_ASAP7_75t_R FILLER_233_578 ();
 DECAPx1_ASAP7_75t_R FILLER_233_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_604 ();
 FILLER_ASAP7_75t_R FILLER_233_619 ();
 DECAPx2_ASAP7_75t_R FILLER_233_632 ();
 FILLER_ASAP7_75t_R FILLER_233_638 ();
 FILLER_ASAP7_75t_R FILLER_233_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_650 ();
 DECAPx6_ASAP7_75t_R FILLER_233_657 ();
 FILLER_ASAP7_75t_R FILLER_233_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_673 ();
 FILLER_ASAP7_75t_R FILLER_233_677 ();
 FILLER_ASAP7_75t_R FILLER_233_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_693 ();
 DECAPx2_ASAP7_75t_R FILLER_233_711 ();
 DECAPx2_ASAP7_75t_R FILLER_233_725 ();
 FILLER_ASAP7_75t_R FILLER_233_731 ();
 DECAPx10_ASAP7_75t_R FILLER_233_755 ();
 DECAPx4_ASAP7_75t_R FILLER_233_777 ();
 FILLER_ASAP7_75t_R FILLER_233_787 ();
 DECAPx10_ASAP7_75t_R FILLER_233_809 ();
 DECAPx2_ASAP7_75t_R FILLER_233_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_837 ();
 DECAPx2_ASAP7_75t_R FILLER_233_841 ();
 FILLER_ASAP7_75t_R FILLER_233_855 ();
 DECAPx10_ASAP7_75t_R FILLER_233_879 ();
 DECAPx10_ASAP7_75t_R FILLER_233_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_923 ();
 FILLER_ASAP7_75t_R FILLER_233_926 ();
 DECAPx2_ASAP7_75t_R FILLER_233_935 ();
 FILLER_ASAP7_75t_R FILLER_233_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_943 ();
 DECAPx2_ASAP7_75t_R FILLER_233_958 ();
 DECAPx1_ASAP7_75t_R FILLER_233_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_985 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1109 ();
 DECAPx6_ASAP7_75t_R FILLER_233_1131 ();
 FILLER_ASAP7_75t_R FILLER_233_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1156 ();
 FILLER_ASAP7_75t_R FILLER_233_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1164 ();
 DECAPx4_ASAP7_75t_R FILLER_233_1173 ();
 FILLER_ASAP7_75t_R FILLER_233_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1192 ();
 DECAPx4_ASAP7_75t_R FILLER_233_1198 ();
 FILLER_ASAP7_75t_R FILLER_233_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_234_2 ();
 DECAPx10_ASAP7_75t_R FILLER_234_24 ();
 DECAPx10_ASAP7_75t_R FILLER_234_46 ();
 DECAPx10_ASAP7_75t_R FILLER_234_68 ();
 DECAPx10_ASAP7_75t_R FILLER_234_90 ();
 DECAPx10_ASAP7_75t_R FILLER_234_112 ();
 DECAPx10_ASAP7_75t_R FILLER_234_134 ();
 DECAPx10_ASAP7_75t_R FILLER_234_156 ();
 DECAPx10_ASAP7_75t_R FILLER_234_178 ();
 DECAPx10_ASAP7_75t_R FILLER_234_200 ();
 DECAPx10_ASAP7_75t_R FILLER_234_222 ();
 DECAPx10_ASAP7_75t_R FILLER_234_244 ();
 DECAPx10_ASAP7_75t_R FILLER_234_266 ();
 DECAPx10_ASAP7_75t_R FILLER_234_288 ();
 DECAPx10_ASAP7_75t_R FILLER_234_310 ();
 DECAPx10_ASAP7_75t_R FILLER_234_332 ();
 DECAPx10_ASAP7_75t_R FILLER_234_354 ();
 DECAPx10_ASAP7_75t_R FILLER_234_376 ();
 DECAPx10_ASAP7_75t_R FILLER_234_398 ();
 DECAPx10_ASAP7_75t_R FILLER_234_420 ();
 DECAPx4_ASAP7_75t_R FILLER_234_442 ();
 FILLER_ASAP7_75t_R FILLER_234_460 ();
 DECAPx1_ASAP7_75t_R FILLER_234_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_511 ();
 DECAPx1_ASAP7_75t_R FILLER_234_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_522 ();
 DECAPx1_ASAP7_75t_R FILLER_234_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_571 ();
 DECAPx1_ASAP7_75t_R FILLER_234_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_595 ();
 DECAPx1_ASAP7_75t_R FILLER_234_603 ();
 FILLER_ASAP7_75t_R FILLER_234_622 ();
 DECAPx1_ASAP7_75t_R FILLER_234_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_650 ();
 DECAPx2_ASAP7_75t_R FILLER_234_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_669 ();
 FILLER_ASAP7_75t_R FILLER_234_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_724 ();
 FILLER_ASAP7_75t_R FILLER_234_733 ();
 FILLER_ASAP7_75t_R FILLER_234_741 ();
 FILLER_ASAP7_75t_R FILLER_234_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_765 ();
 DECAPx6_ASAP7_75t_R FILLER_234_773 ();
 DECAPx1_ASAP7_75t_R FILLER_234_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_791 ();
 DECAPx2_ASAP7_75t_R FILLER_234_814 ();
 FILLER_ASAP7_75t_R FILLER_234_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_826 ();
 FILLER_ASAP7_75t_R FILLER_234_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_856 ();
 DECAPx1_ASAP7_75t_R FILLER_234_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_891 ();
 DECAPx1_ASAP7_75t_R FILLER_234_920 ();
 DECAPx4_ASAP7_75t_R FILLER_234_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_942 ();
 DECAPx2_ASAP7_75t_R FILLER_234_957 ();
 FILLER_ASAP7_75t_R FILLER_234_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_965 ();
 DECAPx2_ASAP7_75t_R FILLER_234_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_983 ();
 DECAPx10_ASAP7_75t_R FILLER_234_990 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_234_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1123 ();
 FILLER_ASAP7_75t_R FILLER_234_1133 ();
 DECAPx6_ASAP7_75t_R FILLER_234_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_234_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1176 ();
 DECAPx6_ASAP7_75t_R FILLER_234_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_235_2 ();
 DECAPx10_ASAP7_75t_R FILLER_235_24 ();
 DECAPx10_ASAP7_75t_R FILLER_235_46 ();
 DECAPx10_ASAP7_75t_R FILLER_235_68 ();
 DECAPx10_ASAP7_75t_R FILLER_235_90 ();
 DECAPx10_ASAP7_75t_R FILLER_235_112 ();
 DECAPx10_ASAP7_75t_R FILLER_235_134 ();
 DECAPx10_ASAP7_75t_R FILLER_235_156 ();
 DECAPx10_ASAP7_75t_R FILLER_235_178 ();
 DECAPx10_ASAP7_75t_R FILLER_235_200 ();
 DECAPx10_ASAP7_75t_R FILLER_235_222 ();
 DECAPx10_ASAP7_75t_R FILLER_235_244 ();
 DECAPx10_ASAP7_75t_R FILLER_235_266 ();
 DECAPx10_ASAP7_75t_R FILLER_235_288 ();
 DECAPx10_ASAP7_75t_R FILLER_235_310 ();
 DECAPx10_ASAP7_75t_R FILLER_235_332 ();
 DECAPx10_ASAP7_75t_R FILLER_235_354 ();
 DECAPx10_ASAP7_75t_R FILLER_235_376 ();
 DECAPx10_ASAP7_75t_R FILLER_235_398 ();
 DECAPx4_ASAP7_75t_R FILLER_235_420 ();
 FILLER_ASAP7_75t_R FILLER_235_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_432 ();
 DECAPx1_ASAP7_75t_R FILLER_235_461 ();
 DECAPx4_ASAP7_75t_R FILLER_235_486 ();
 FILLER_ASAP7_75t_R FILLER_235_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_498 ();
 DECAPx1_ASAP7_75t_R FILLER_235_506 ();
 DECAPx1_ASAP7_75t_R FILLER_235_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_542 ();
 DECAPx1_ASAP7_75t_R FILLER_235_554 ();
 DECAPx4_ASAP7_75t_R FILLER_235_564 ();
 FILLER_ASAP7_75t_R FILLER_235_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_576 ();
 FILLER_ASAP7_75t_R FILLER_235_584 ();
 DECAPx10_ASAP7_75t_R FILLER_235_592 ();
 DECAPx1_ASAP7_75t_R FILLER_235_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_643 ();
 FILLER_ASAP7_75t_R FILLER_235_649 ();
 FILLER_ASAP7_75t_R FILLER_235_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_658 ();
 FILLER_ASAP7_75t_R FILLER_235_662 ();
 DECAPx2_ASAP7_75t_R FILLER_235_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_678 ();
 DECAPx10_ASAP7_75t_R FILLER_235_692 ();
 FILLER_ASAP7_75t_R FILLER_235_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_716 ();
 DECAPx1_ASAP7_75t_R FILLER_235_726 ();
 DECAPx10_ASAP7_75t_R FILLER_235_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_765 ();
 DECAPx1_ASAP7_75t_R FILLER_235_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_792 ();
 DECAPx6_ASAP7_75t_R FILLER_235_800 ();
 FILLER_ASAP7_75t_R FILLER_235_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_828 ();
 DECAPx4_ASAP7_75t_R FILLER_235_834 ();
 FILLER_ASAP7_75t_R FILLER_235_844 ();
 FILLER_ASAP7_75t_R FILLER_235_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_856 ();
 DECAPx4_ASAP7_75t_R FILLER_235_863 ();
 FILLER_ASAP7_75t_R FILLER_235_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_875 ();
 DECAPx2_ASAP7_75t_R FILLER_235_887 ();
 FILLER_ASAP7_75t_R FILLER_235_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_901 ();
 FILLER_ASAP7_75t_R FILLER_235_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_912 ();
 FILLER_ASAP7_75t_R FILLER_235_922 ();
 DECAPx1_ASAP7_75t_R FILLER_235_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_971 ();
 DECAPx6_ASAP7_75t_R FILLER_235_978 ();
 FILLER_ASAP7_75t_R FILLER_235_992 ();
 DECAPx2_ASAP7_75t_R FILLER_235_997 ();
 FILLER_ASAP7_75t_R FILLER_235_1003 ();
 FILLER_ASAP7_75t_R FILLER_235_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1010 ();
 FILLER_ASAP7_75t_R FILLER_235_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1016 ();
 DECAPx6_ASAP7_75t_R FILLER_235_1022 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1081 ();
 FILLER_ASAP7_75t_R FILLER_235_1103 ();
 FILLER_ASAP7_75t_R FILLER_235_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1110 ();
 DECAPx4_ASAP7_75t_R FILLER_235_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1161 ();
 DECAPx6_ASAP7_75t_R FILLER_235_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1205 ();
 DECAPx4_ASAP7_75t_R FILLER_235_1211 ();
 FILLER_ASAP7_75t_R FILLER_235_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_236_2 ();
 DECAPx10_ASAP7_75t_R FILLER_236_24 ();
 DECAPx10_ASAP7_75t_R FILLER_236_46 ();
 DECAPx10_ASAP7_75t_R FILLER_236_68 ();
 DECAPx10_ASAP7_75t_R FILLER_236_90 ();
 DECAPx10_ASAP7_75t_R FILLER_236_112 ();
 DECAPx10_ASAP7_75t_R FILLER_236_134 ();
 DECAPx10_ASAP7_75t_R FILLER_236_156 ();
 DECAPx10_ASAP7_75t_R FILLER_236_178 ();
 DECAPx10_ASAP7_75t_R FILLER_236_200 ();
 DECAPx10_ASAP7_75t_R FILLER_236_222 ();
 DECAPx10_ASAP7_75t_R FILLER_236_244 ();
 DECAPx10_ASAP7_75t_R FILLER_236_266 ();
 DECAPx10_ASAP7_75t_R FILLER_236_288 ();
 DECAPx10_ASAP7_75t_R FILLER_236_310 ();
 DECAPx10_ASAP7_75t_R FILLER_236_332 ();
 DECAPx10_ASAP7_75t_R FILLER_236_354 ();
 DECAPx10_ASAP7_75t_R FILLER_236_376 ();
 DECAPx10_ASAP7_75t_R FILLER_236_398 ();
 DECAPx10_ASAP7_75t_R FILLER_236_420 ();
 DECAPx6_ASAP7_75t_R FILLER_236_442 ();
 DECAPx2_ASAP7_75t_R FILLER_236_456 ();
 DECAPx2_ASAP7_75t_R FILLER_236_481 ();
 DECAPx2_ASAP7_75t_R FILLER_236_494 ();
 FILLER_ASAP7_75t_R FILLER_236_500 ();
 FILLER_ASAP7_75t_R FILLER_236_514 ();
 DECAPx1_ASAP7_75t_R FILLER_236_524 ();
 FILLER_ASAP7_75t_R FILLER_236_572 ();
 DECAPx1_ASAP7_75t_R FILLER_236_604 ();
 DECAPx6_ASAP7_75t_R FILLER_236_633 ();
 FILLER_ASAP7_75t_R FILLER_236_647 ();
 FILLER_ASAP7_75t_R FILLER_236_652 ();
 DECAPx1_ASAP7_75t_R FILLER_236_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_674 ();
 DECAPx4_ASAP7_75t_R FILLER_236_683 ();
 FILLER_ASAP7_75t_R FILLER_236_693 ();
 FILLER_ASAP7_75t_R FILLER_236_703 ();
 DECAPx4_ASAP7_75t_R FILLER_236_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_729 ();
 DECAPx1_ASAP7_75t_R FILLER_236_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_741 ();
 DECAPx4_ASAP7_75t_R FILLER_236_750 ();
 FILLER_ASAP7_75t_R FILLER_236_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_762 ();
 DECAPx2_ASAP7_75t_R FILLER_236_778 ();
 FILLER_ASAP7_75t_R FILLER_236_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_795 ();
 DECAPx1_ASAP7_75t_R FILLER_236_802 ();
 DECAPx1_ASAP7_75t_R FILLER_236_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_848 ();
 DECAPx6_ASAP7_75t_R FILLER_236_869 ();
 DECAPx2_ASAP7_75t_R FILLER_236_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_889 ();
 DECAPx2_ASAP7_75t_R FILLER_236_903 ();
 FILLER_ASAP7_75t_R FILLER_236_909 ();
 DECAPx2_ASAP7_75t_R FILLER_236_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_925 ();
 FILLER_ASAP7_75t_R FILLER_236_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_950 ();
 DECAPx2_ASAP7_75t_R FILLER_236_954 ();
 FILLER_ASAP7_75t_R FILLER_236_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_962 ();
 DECAPx1_ASAP7_75t_R FILLER_236_993 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1025 ();
 FILLER_ASAP7_75t_R FILLER_236_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1040 ();
 FILLER_ASAP7_75t_R FILLER_236_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1052 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1070 ();
 FILLER_ASAP7_75t_R FILLER_236_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1166 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1188 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_237_2 ();
 DECAPx10_ASAP7_75t_R FILLER_237_24 ();
 DECAPx10_ASAP7_75t_R FILLER_237_46 ();
 DECAPx10_ASAP7_75t_R FILLER_237_68 ();
 DECAPx10_ASAP7_75t_R FILLER_237_90 ();
 DECAPx10_ASAP7_75t_R FILLER_237_112 ();
 DECAPx10_ASAP7_75t_R FILLER_237_134 ();
 DECAPx10_ASAP7_75t_R FILLER_237_156 ();
 DECAPx10_ASAP7_75t_R FILLER_237_178 ();
 DECAPx10_ASAP7_75t_R FILLER_237_200 ();
 DECAPx10_ASAP7_75t_R FILLER_237_222 ();
 DECAPx10_ASAP7_75t_R FILLER_237_244 ();
 DECAPx10_ASAP7_75t_R FILLER_237_266 ();
 DECAPx10_ASAP7_75t_R FILLER_237_288 ();
 DECAPx10_ASAP7_75t_R FILLER_237_310 ();
 DECAPx10_ASAP7_75t_R FILLER_237_332 ();
 DECAPx10_ASAP7_75t_R FILLER_237_354 ();
 DECAPx10_ASAP7_75t_R FILLER_237_376 ();
 DECAPx10_ASAP7_75t_R FILLER_237_398 ();
 DECAPx10_ASAP7_75t_R FILLER_237_420 ();
 DECAPx10_ASAP7_75t_R FILLER_237_442 ();
 FILLER_ASAP7_75t_R FILLER_237_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_466 ();
 DECAPx10_ASAP7_75t_R FILLER_237_505 ();
 DECAPx10_ASAP7_75t_R FILLER_237_527 ();
 DECAPx4_ASAP7_75t_R FILLER_237_549 ();
 FILLER_ASAP7_75t_R FILLER_237_559 ();
 FILLER_ASAP7_75t_R FILLER_237_570 ();
 DECAPx6_ASAP7_75t_R FILLER_237_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_592 ();
 DECAPx6_ASAP7_75t_R FILLER_237_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_628 ();
 DECAPx2_ASAP7_75t_R FILLER_237_632 ();
 FILLER_ASAP7_75t_R FILLER_237_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_673 ();
 DECAPx2_ASAP7_75t_R FILLER_237_679 ();
 FILLER_ASAP7_75t_R FILLER_237_685 ();
 FILLER_ASAP7_75t_R FILLER_237_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_695 ();
 DECAPx2_ASAP7_75t_R FILLER_237_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_713 ();
 DECAPx2_ASAP7_75t_R FILLER_237_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_737 ();
 DECAPx2_ASAP7_75t_R FILLER_237_750 ();
 FILLER_ASAP7_75t_R FILLER_237_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_758 ();
 DECAPx6_ASAP7_75t_R FILLER_237_772 ();
 DECAPx6_ASAP7_75t_R FILLER_237_818 ();
 FILLER_ASAP7_75t_R FILLER_237_835 ();
 DECAPx4_ASAP7_75t_R FILLER_237_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_855 ();
 FILLER_ASAP7_75t_R FILLER_237_859 ();
 DECAPx4_ASAP7_75t_R FILLER_237_901 ();
 FILLER_ASAP7_75t_R FILLER_237_911 ();
 DECAPx10_ASAP7_75t_R FILLER_237_926 ();
 FILLER_ASAP7_75t_R FILLER_237_948 ();
 DECAPx1_ASAP7_75t_R FILLER_237_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_978 ();
 DECAPx1_ASAP7_75t_R FILLER_237_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_237_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1041 ();
 FILLER_ASAP7_75t_R FILLER_237_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1062 ();
 FILLER_ASAP7_75t_R FILLER_237_1072 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1077 ();
 FILLER_ASAP7_75t_R FILLER_237_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1095 ();
 FILLER_ASAP7_75t_R FILLER_237_1101 ();
 FILLER_ASAP7_75t_R FILLER_237_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_237_1125 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1142 ();
 FILLER_ASAP7_75t_R FILLER_237_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_237_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_237_1176 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_238_2 ();
 DECAPx10_ASAP7_75t_R FILLER_238_24 ();
 DECAPx10_ASAP7_75t_R FILLER_238_46 ();
 DECAPx10_ASAP7_75t_R FILLER_238_68 ();
 DECAPx10_ASAP7_75t_R FILLER_238_90 ();
 DECAPx10_ASAP7_75t_R FILLER_238_112 ();
 DECAPx10_ASAP7_75t_R FILLER_238_134 ();
 DECAPx10_ASAP7_75t_R FILLER_238_156 ();
 DECAPx10_ASAP7_75t_R FILLER_238_178 ();
 DECAPx10_ASAP7_75t_R FILLER_238_200 ();
 DECAPx10_ASAP7_75t_R FILLER_238_222 ();
 DECAPx10_ASAP7_75t_R FILLER_238_244 ();
 DECAPx10_ASAP7_75t_R FILLER_238_266 ();
 DECAPx10_ASAP7_75t_R FILLER_238_288 ();
 DECAPx10_ASAP7_75t_R FILLER_238_310 ();
 DECAPx10_ASAP7_75t_R FILLER_238_332 ();
 DECAPx10_ASAP7_75t_R FILLER_238_354 ();
 DECAPx10_ASAP7_75t_R FILLER_238_376 ();
 DECAPx10_ASAP7_75t_R FILLER_238_398 ();
 DECAPx10_ASAP7_75t_R FILLER_238_420 ();
 DECAPx6_ASAP7_75t_R FILLER_238_442 ();
 DECAPx2_ASAP7_75t_R FILLER_238_456 ();
 DECAPx6_ASAP7_75t_R FILLER_238_475 ();
 FILLER_ASAP7_75t_R FILLER_238_495 ();
 DECAPx10_ASAP7_75t_R FILLER_238_503 ();
 FILLER_ASAP7_75t_R FILLER_238_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_527 ();
 DECAPx10_ASAP7_75t_R FILLER_238_531 ();
 DECAPx2_ASAP7_75t_R FILLER_238_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_634 ();
 FILLER_ASAP7_75t_R FILLER_238_659 ();
 FILLER_ASAP7_75t_R FILLER_238_677 ();
 FILLER_ASAP7_75t_R FILLER_238_709 ();
 FILLER_ASAP7_75t_R FILLER_238_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_722 ();
 DECAPx4_ASAP7_75t_R FILLER_238_778 ();
 DECAPx2_ASAP7_75t_R FILLER_238_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_827 ();
 DECAPx2_ASAP7_75t_R FILLER_238_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_846 ();
 FILLER_ASAP7_75t_R FILLER_238_852 ();
 DECAPx2_ASAP7_75t_R FILLER_238_862 ();
 DECAPx10_ASAP7_75t_R FILLER_238_871 ();
 FILLER_ASAP7_75t_R FILLER_238_893 ();
 DECAPx1_ASAP7_75t_R FILLER_238_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_921 ();
 DECAPx1_ASAP7_75t_R FILLER_238_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_954 ();
 DECAPx2_ASAP7_75t_R FILLER_238_963 ();
 DECAPx2_ASAP7_75t_R FILLER_238_975 ();
 FILLER_ASAP7_75t_R FILLER_238_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_992 ();
 DECAPx1_ASAP7_75t_R FILLER_238_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1015 ();
 FILLER_ASAP7_75t_R FILLER_238_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1028 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_238_1043 ();
 FILLER_ASAP7_75t_R FILLER_238_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1064 ();
 FILLER_ASAP7_75t_R FILLER_238_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1075 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1081 ();
 FILLER_ASAP7_75t_R FILLER_238_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1115 ();
 DECAPx6_ASAP7_75t_R FILLER_238_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1151 ();
 DECAPx4_ASAP7_75t_R FILLER_238_1158 ();
 FILLER_ASAP7_75t_R FILLER_238_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1174 ();
 FILLER_ASAP7_75t_R FILLER_238_1178 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1203 ();
 FILLER_ASAP7_75t_R FILLER_238_1212 ();
 FILLER_ASAP7_75t_R FILLER_238_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_239_2 ();
 DECAPx10_ASAP7_75t_R FILLER_239_24 ();
 DECAPx10_ASAP7_75t_R FILLER_239_46 ();
 DECAPx10_ASAP7_75t_R FILLER_239_68 ();
 DECAPx10_ASAP7_75t_R FILLER_239_90 ();
 DECAPx10_ASAP7_75t_R FILLER_239_112 ();
 DECAPx10_ASAP7_75t_R FILLER_239_134 ();
 DECAPx10_ASAP7_75t_R FILLER_239_156 ();
 DECAPx10_ASAP7_75t_R FILLER_239_178 ();
 DECAPx10_ASAP7_75t_R FILLER_239_200 ();
 DECAPx10_ASAP7_75t_R FILLER_239_222 ();
 DECAPx10_ASAP7_75t_R FILLER_239_244 ();
 DECAPx10_ASAP7_75t_R FILLER_239_266 ();
 DECAPx10_ASAP7_75t_R FILLER_239_288 ();
 DECAPx10_ASAP7_75t_R FILLER_239_310 ();
 DECAPx10_ASAP7_75t_R FILLER_239_332 ();
 DECAPx10_ASAP7_75t_R FILLER_239_354 ();
 DECAPx10_ASAP7_75t_R FILLER_239_376 ();
 DECAPx10_ASAP7_75t_R FILLER_239_398 ();
 DECAPx10_ASAP7_75t_R FILLER_239_420 ();
 DECAPx10_ASAP7_75t_R FILLER_239_442 ();
 DECAPx1_ASAP7_75t_R FILLER_239_493 ();
 DECAPx1_ASAP7_75t_R FILLER_239_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_507 ();
 FILLER_ASAP7_75t_R FILLER_239_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_543 ();
 DECAPx1_ASAP7_75t_R FILLER_239_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_573 ();
 FILLER_ASAP7_75t_R FILLER_239_602 ();
 DECAPx1_ASAP7_75t_R FILLER_239_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_620 ();
 FILLER_ASAP7_75t_R FILLER_239_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_670 ();
 FILLER_ASAP7_75t_R FILLER_239_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_676 ();
 FILLER_ASAP7_75t_R FILLER_239_686 ();
 FILLER_ASAP7_75t_R FILLER_239_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_699 ();
 DECAPx1_ASAP7_75t_R FILLER_239_714 ();
 DECAPx2_ASAP7_75t_R FILLER_239_730 ();
 FILLER_ASAP7_75t_R FILLER_239_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_756 ();
 FILLER_ASAP7_75t_R FILLER_239_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_771 ();
 FILLER_ASAP7_75t_R FILLER_239_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_796 ();
 DECAPx4_ASAP7_75t_R FILLER_239_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_841 ();
 DECAPx4_ASAP7_75t_R FILLER_239_850 ();
 FILLER_ASAP7_75t_R FILLER_239_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_865 ();
 DECAPx2_ASAP7_75t_R FILLER_239_871 ();
 FILLER_ASAP7_75t_R FILLER_239_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_887 ();
 DECAPx6_ASAP7_75t_R FILLER_239_908 ();
 FILLER_ASAP7_75t_R FILLER_239_922 ();
 DECAPx1_ASAP7_75t_R FILLER_239_926 ();
 DECAPx4_ASAP7_75t_R FILLER_239_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_946 ();
 FILLER_ASAP7_75t_R FILLER_239_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_954 ();
 DECAPx10_ASAP7_75t_R FILLER_239_958 ();
 DECAPx6_ASAP7_75t_R FILLER_239_980 ();
 FILLER_ASAP7_75t_R FILLER_239_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_996 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_239_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1034 ();
 FILLER_ASAP7_75t_R FILLER_239_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1066 ();
 FILLER_ASAP7_75t_R FILLER_239_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_239_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1162 ();
 DECAPx1_ASAP7_75t_R FILLER_239_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1175 ();
 FILLER_ASAP7_75t_R FILLER_239_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_240_2 ();
 DECAPx10_ASAP7_75t_R FILLER_240_24 ();
 DECAPx10_ASAP7_75t_R FILLER_240_46 ();
 DECAPx10_ASAP7_75t_R FILLER_240_68 ();
 DECAPx10_ASAP7_75t_R FILLER_240_90 ();
 DECAPx10_ASAP7_75t_R FILLER_240_112 ();
 DECAPx10_ASAP7_75t_R FILLER_240_134 ();
 DECAPx10_ASAP7_75t_R FILLER_240_156 ();
 DECAPx10_ASAP7_75t_R FILLER_240_178 ();
 DECAPx10_ASAP7_75t_R FILLER_240_200 ();
 DECAPx10_ASAP7_75t_R FILLER_240_222 ();
 DECAPx10_ASAP7_75t_R FILLER_240_244 ();
 DECAPx10_ASAP7_75t_R FILLER_240_266 ();
 DECAPx10_ASAP7_75t_R FILLER_240_288 ();
 DECAPx10_ASAP7_75t_R FILLER_240_310 ();
 DECAPx10_ASAP7_75t_R FILLER_240_332 ();
 DECAPx10_ASAP7_75t_R FILLER_240_354 ();
 DECAPx10_ASAP7_75t_R FILLER_240_376 ();
 DECAPx10_ASAP7_75t_R FILLER_240_398 ();
 DECAPx10_ASAP7_75t_R FILLER_240_420 ();
 DECAPx6_ASAP7_75t_R FILLER_240_442 ();
 DECAPx2_ASAP7_75t_R FILLER_240_456 ();
 DECAPx2_ASAP7_75t_R FILLER_240_464 ();
 FILLER_ASAP7_75t_R FILLER_240_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_472 ();
 DECAPx1_ASAP7_75t_R FILLER_240_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_483 ();
 FILLER_ASAP7_75t_R FILLER_240_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_576 ();
 DECAPx2_ASAP7_75t_R FILLER_240_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_603 ();
 DECAPx1_ASAP7_75t_R FILLER_240_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_625 ();
 FILLER_ASAP7_75t_R FILLER_240_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_749 ();
 FILLER_ASAP7_75t_R FILLER_240_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_760 ();
 FILLER_ASAP7_75t_R FILLER_240_772 ();
 DECAPx6_ASAP7_75t_R FILLER_240_780 ();
 DECAPx1_ASAP7_75t_R FILLER_240_794 ();
 DECAPx2_ASAP7_75t_R FILLER_240_801 ();
 FILLER_ASAP7_75t_R FILLER_240_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_809 ();
 FILLER_ASAP7_75t_R FILLER_240_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_856 ();
 DECAPx6_ASAP7_75t_R FILLER_240_865 ();
 DECAPx2_ASAP7_75t_R FILLER_240_879 ();
 DECAPx4_ASAP7_75t_R FILLER_240_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_930 ();
 DECAPx4_ASAP7_75t_R FILLER_240_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_946 ();
 FILLER_ASAP7_75t_R FILLER_240_955 ();
 FILLER_ASAP7_75t_R FILLER_240_973 ();
 DECAPx6_ASAP7_75t_R FILLER_240_980 ();
 DECAPx4_ASAP7_75t_R FILLER_240_997 ();
 FILLER_ASAP7_75t_R FILLER_240_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_240_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1059 ();
 FILLER_ASAP7_75t_R FILLER_240_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1079 ();
 FILLER_ASAP7_75t_R FILLER_240_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1106 ();
 FILLER_ASAP7_75t_R FILLER_240_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_240_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1175 ();
 FILLER_ASAP7_75t_R FILLER_240_1184 ();
 FILLER_ASAP7_75t_R FILLER_240_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1193 ();
 FILLER_ASAP7_75t_R FILLER_240_1197 ();
 DECAPx4_ASAP7_75t_R FILLER_240_1212 ();
 FILLER_ASAP7_75t_R FILLER_240_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_241_2 ();
 DECAPx10_ASAP7_75t_R FILLER_241_24 ();
 DECAPx10_ASAP7_75t_R FILLER_241_46 ();
 DECAPx10_ASAP7_75t_R FILLER_241_68 ();
 DECAPx10_ASAP7_75t_R FILLER_241_90 ();
 DECAPx10_ASAP7_75t_R FILLER_241_112 ();
 DECAPx10_ASAP7_75t_R FILLER_241_134 ();
 DECAPx10_ASAP7_75t_R FILLER_241_156 ();
 DECAPx10_ASAP7_75t_R FILLER_241_178 ();
 DECAPx10_ASAP7_75t_R FILLER_241_200 ();
 DECAPx10_ASAP7_75t_R FILLER_241_222 ();
 DECAPx10_ASAP7_75t_R FILLER_241_244 ();
 DECAPx10_ASAP7_75t_R FILLER_241_266 ();
 DECAPx10_ASAP7_75t_R FILLER_241_288 ();
 DECAPx10_ASAP7_75t_R FILLER_241_310 ();
 DECAPx10_ASAP7_75t_R FILLER_241_332 ();
 DECAPx10_ASAP7_75t_R FILLER_241_354 ();
 DECAPx10_ASAP7_75t_R FILLER_241_376 ();
 DECAPx10_ASAP7_75t_R FILLER_241_398 ();
 DECAPx10_ASAP7_75t_R FILLER_241_420 ();
 DECAPx10_ASAP7_75t_R FILLER_241_442 ();
 DECAPx4_ASAP7_75t_R FILLER_241_464 ();
 FILLER_ASAP7_75t_R FILLER_241_513 ();
 FILLER_ASAP7_75t_R FILLER_241_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_547 ();
 FILLER_ASAP7_75t_R FILLER_241_580 ();
 DECAPx1_ASAP7_75t_R FILLER_241_587 ();
 FILLER_ASAP7_75t_R FILLER_241_597 ();
 FILLER_ASAP7_75t_R FILLER_241_609 ();
 DECAPx2_ASAP7_75t_R FILLER_241_617 ();
 FILLER_ASAP7_75t_R FILLER_241_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_707 ();
 DECAPx1_ASAP7_75t_R FILLER_241_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_787 ();
 FILLER_ASAP7_75t_R FILLER_241_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_861 ();
 FILLER_ASAP7_75t_R FILLER_241_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_867 ();
 DECAPx1_ASAP7_75t_R FILLER_241_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_917 ();
 DECAPx1_ASAP7_75t_R FILLER_241_931 ();
 DECAPx2_ASAP7_75t_R FILLER_241_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_946 ();
 DECAPx2_ASAP7_75t_R FILLER_241_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_964 ();
 DECAPx6_ASAP7_75t_R FILLER_241_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_987 ();
 DECAPx2_ASAP7_75t_R FILLER_241_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_241_1046 ();
 FILLER_ASAP7_75t_R FILLER_241_1060 ();
 FILLER_ASAP7_75t_R FILLER_241_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_241_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1078 ();
 FILLER_ASAP7_75t_R FILLER_241_1082 ();
 FILLER_ASAP7_75t_R FILLER_241_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_241_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_241_1134 ();
 FILLER_ASAP7_75t_R FILLER_241_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_241_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1178 ();
 FILLER_ASAP7_75t_R FILLER_241_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1189 ();
 FILLER_ASAP7_75t_R FILLER_241_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1204 ();
 FILLER_ASAP7_75t_R FILLER_241_1210 ();
 FILLER_ASAP7_75t_R FILLER_241_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_242_2 ();
 DECAPx10_ASAP7_75t_R FILLER_242_24 ();
 DECAPx10_ASAP7_75t_R FILLER_242_46 ();
 DECAPx10_ASAP7_75t_R FILLER_242_68 ();
 DECAPx10_ASAP7_75t_R FILLER_242_90 ();
 DECAPx10_ASAP7_75t_R FILLER_242_112 ();
 DECAPx10_ASAP7_75t_R FILLER_242_134 ();
 DECAPx10_ASAP7_75t_R FILLER_242_156 ();
 DECAPx10_ASAP7_75t_R FILLER_242_178 ();
 DECAPx10_ASAP7_75t_R FILLER_242_200 ();
 DECAPx10_ASAP7_75t_R FILLER_242_222 ();
 DECAPx10_ASAP7_75t_R FILLER_242_244 ();
 DECAPx10_ASAP7_75t_R FILLER_242_266 ();
 DECAPx10_ASAP7_75t_R FILLER_242_288 ();
 DECAPx10_ASAP7_75t_R FILLER_242_310 ();
 DECAPx6_ASAP7_75t_R FILLER_242_332 ();
 DECAPx2_ASAP7_75t_R FILLER_242_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_352 ();
 DECAPx6_ASAP7_75t_R FILLER_242_359 ();
 DECAPx2_ASAP7_75t_R FILLER_242_373 ();
 DECAPx2_ASAP7_75t_R FILLER_242_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_391 ();
 DECAPx10_ASAP7_75t_R FILLER_242_398 ();
 FILLER_ASAP7_75t_R FILLER_242_420 ();
 DECAPx10_ASAP7_75t_R FILLER_242_428 ();
 DECAPx4_ASAP7_75t_R FILLER_242_450 ();
 FILLER_ASAP7_75t_R FILLER_242_460 ();
 DECAPx10_ASAP7_75t_R FILLER_242_464 ();
 FILLER_ASAP7_75t_R FILLER_242_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_529 ();
 DECAPx2_ASAP7_75t_R FILLER_242_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_548 ();
 FILLER_ASAP7_75t_R FILLER_242_559 ();
 DECAPx1_ASAP7_75t_R FILLER_242_579 ();
 FILLER_ASAP7_75t_R FILLER_242_603 ();
 FILLER_ASAP7_75t_R FILLER_242_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_736 ();
 FILLER_ASAP7_75t_R FILLER_242_757 ();
 FILLER_ASAP7_75t_R FILLER_242_764 ();
 FILLER_ASAP7_75t_R FILLER_242_806 ();
 FILLER_ASAP7_75t_R FILLER_242_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_862 ();
 DECAPx1_ASAP7_75t_R FILLER_242_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_893 ();
 FILLER_ASAP7_75t_R FILLER_242_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_968 ();
 DECAPx1_ASAP7_75t_R FILLER_242_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_987 ();
 FILLER_ASAP7_75t_R FILLER_242_993 ();
 FILLER_ASAP7_75t_R FILLER_242_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_242_1011 ();
 FILLER_ASAP7_75t_R FILLER_242_1028 ();
 FILLER_ASAP7_75t_R FILLER_242_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1070 ();
 FILLER_ASAP7_75t_R FILLER_242_1084 ();
 FILLER_ASAP7_75t_R FILLER_242_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_242_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1120 ();
 DECAPx4_ASAP7_75t_R FILLER_242_1124 ();
 FILLER_ASAP7_75t_R FILLER_242_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_242_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_242_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1210 ();
 DECAPx1_ASAP7_75t_R FILLER_242_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1218 ();
 FILLER_ASAP7_75t_R FILLER_242_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_243_2 ();
 DECAPx10_ASAP7_75t_R FILLER_243_24 ();
 DECAPx10_ASAP7_75t_R FILLER_243_46 ();
 DECAPx10_ASAP7_75t_R FILLER_243_68 ();
 DECAPx10_ASAP7_75t_R FILLER_243_90 ();
 DECAPx10_ASAP7_75t_R FILLER_243_112 ();
 DECAPx10_ASAP7_75t_R FILLER_243_134 ();
 DECAPx10_ASAP7_75t_R FILLER_243_156 ();
 DECAPx10_ASAP7_75t_R FILLER_243_178 ();
 DECAPx10_ASAP7_75t_R FILLER_243_200 ();
 DECAPx10_ASAP7_75t_R FILLER_243_222 ();
 DECAPx10_ASAP7_75t_R FILLER_243_244 ();
 DECAPx10_ASAP7_75t_R FILLER_243_266 ();
 DECAPx10_ASAP7_75t_R FILLER_243_288 ();
 DECAPx10_ASAP7_75t_R FILLER_243_310 ();
 DECAPx4_ASAP7_75t_R FILLER_243_344 ();
 FILLER_ASAP7_75t_R FILLER_243_354 ();
 DECAPx6_ASAP7_75t_R FILLER_243_362 ();
 DECAPx2_ASAP7_75t_R FILLER_243_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_382 ();
 DECAPx6_ASAP7_75t_R FILLER_243_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_403 ();
 DECAPx1_ASAP7_75t_R FILLER_243_416 ();
 DECAPx10_ASAP7_75t_R FILLER_243_432 ();
 DECAPx2_ASAP7_75t_R FILLER_243_454 ();
 FILLER_ASAP7_75t_R FILLER_243_460 ();
 DECAPx2_ASAP7_75t_R FILLER_243_464 ();
 FILLER_ASAP7_75t_R FILLER_243_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_566 ();
 FILLER_ASAP7_75t_R FILLER_243_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_661 ();
 FILLER_ASAP7_75t_R FILLER_243_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_827 ();
 FILLER_ASAP7_75t_R FILLER_243_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_918 ();
 DECAPx4_ASAP7_75t_R FILLER_243_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_944 ();
 FILLER_ASAP7_75t_R FILLER_243_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_986 ();
 FILLER_ASAP7_75t_R FILLER_243_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1075 ();
 FILLER_ASAP7_75t_R FILLER_243_1084 ();
 DECAPx1_ASAP7_75t_R FILLER_243_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1095 ();
 FILLER_ASAP7_75t_R FILLER_243_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1132 ();
 FILLER_ASAP7_75t_R FILLER_243_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1148 ();
 FILLER_ASAP7_75t_R FILLER_243_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_243_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1214 ();
 FILLER_ASAP7_75t_R FILLER_243_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1223 ();
endmodule
